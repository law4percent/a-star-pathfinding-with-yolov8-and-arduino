PK   �>�X*M��l  ��     cirkitFile.json�][o۸�+��jޙ���s�}�m���CS�D5:��9��n��?C9qdǲ��Nw�h���p����Q�d����rٺ�G׮��";1�.l[}�ëd�]5�Y��}h��Ev��ϻ�W./��W˅[t3^��e�;�伲U��\2RÙ�f$;{�OXe�l�rKk�˵S2W��R
*]�g&{?y��32e1CS:B��X�G��*�`*�V�S��Bj�CU�$�*�"n�(�:j�ƀ42=�������JCJ��0@sn�vm)�@�
 �k��#�(BÖ:N�ŉ�8q'.��U���L`b����M��$�j�
�Vefghijk�#�Md������c;c ��z�R���#QO#QO#QO#QO#QO#Q�"Q�"Q�b��x��u#��V
/s�(
s�sSK�+Y���Bc{e �:l�8*�uSr�����,9��uM����c��@E�"B�Z����Z�e/�Ӯ�Q��wCk��3
���U"B$�%͌��th��@�H�E&Ѣ�h�I��c\\$0Ҡ����� � �@�`ҀL����4Q�Ƕ������\H��T�4(�iPLӠ��A1K�b��,�8��Cˑ�+�<�h�����v.��/�u��y$Տ�B�haǴS�x-G�L�j	���Z��(���k9���T?^�H�E&Ѣ�h�I��4�K�4�4��4��4 �4�4�4�4 �4(�iPL��4(�iPLӠ��A1M�b��4�i�4(fiP�Q��(�����R�[-H���n}O�Tfg@&٧�u����UͰX��k��w{� X�����Ζ�s[�\�B#m�(�#@R��+aA��+NH�%��h4�X�Le*-
�?�x��#g*�F���cnq�S�9���ޑ�Z��P��ƭ�%��K�֬���豽#Y=��A#���A#��s	�+}w�*,�V�V@��p**!����9f�rl��6��x7 �N� ���g%�%�g���9�f�	�x�)b'ɟ��'@X�)���*P��$T14�#��y��Zw���$�.�}|����H�{?x���-ހH
w2�f��<��7 ��6�	�]��,�OB�Z�$��d��1�,��'�@(<�B�`o���7��G���]�1y�1 0��5 pI`��������K��.��I_L����a�8��5��X��O�����[�F&ԑC��8AF�2���?�M��|/���mu�,6'�6ߗu�m�s]7U�a.���C|�kG�H�>�5�<صc��>ᵣNE�
�}𙯰���Qu�y|)���ȳHy)/"�e�����i�e��~�+fz�O�(�"b!
��X�B,J��[Q
Ll��E"�Δ{6��m*��Vئ~n+j��8��8��8��8��8e�8e�8e�[���|�*��º���$�S�T�������!�������~��_�B�Q(ĥ�G�d���5�/�|��+\�;��ໂ��3��ໃ�^ �����%���^�z	�%���^�z	�%��`�9�����r�'��[e /�)KG
Rڛ�)T��p���0�%��uU�4����y�C�(Ѳ�sV�sPuV:/kn�1���%e��� �<���e�յ�]u�.���; lә
�*n���%Z[�S*�P]s��ߧ�ػ^Cn�:���ڲ{<.�덞�`�}���GOr���v���c\�7����D�캟Rӿ��)n��c�O��m��>&�c���^x�݇w�D�7��&u�I�4��M䦩ߥ�|>+Zg�bi[�^��ͪ[���'V���'�/��7��ʵ]��V��p�j��E�����J����b�%S{����;��3#�tW���0�͙֕�F�Ԙ���%�ݾS�N2�k;�(׊�v�I�l�b��f�W^wӖsw3C�SS1� �O����/rآo[��*�h���u�,7f0eS��?�5`�5"%GwI��93p���jpUY�&'VT9Ή��X@.d�sJ�-����+�g��h�j�f���G��x��{�;�W��K4���}��W]�,>��{����d���_�����_K�z�hP<ßZ���u襮�v�J�m�t��7�6�Wn�t�uu���z�V\eg�����@�T��իە{Ӕ�7�ś�ؽZS����zQ��}�ύQw������˺�����+[n�|� ��6��A�>I��~�:��&�T[/���/�W�q�����F5L{���i_��>2o'��6S���Z`�b�M���\Hb����&��T���WP��,��jk9S��zo��n܇���q�dA��+]����^������9V�c�Ic#tJ)��VE�	P9�L`K��[N�A��ibu�
�j�&�K1�zʑʡ#nH�p�%�\�Ν�kArM��(QTTDXAS*���)���I�f�9�	3��g��4wn�ǋDJE����5�`�R�-���
"�A�B�@�KBV�&S! 7�5��%���(��Ė3�d�@$���r���zbniI�c�~g�b"�.W�30��\xo�g����"��	땻B��M8g����aE׷�u��&ۓ\���.�w��¯�F�T����11�x�M�5�&#rLB��w�+�)���Hl)�m��u�a�d�6��d~~}�u�]���R
�d`4i9U)6h2����p�w�x�D���N�Z$�J��E�!ʆ-���P����m;��Q�W��h�/�]�.��{f��L��U��*�b�"���41�#�d�|��\�4Ea�#��QQ���sh>��S���#$(����S��3�4�ARHI�8Ml=���W���������))o�9B�j.�����RL��MzZ��!�F��!�嘐|�������K�b=#I(�SSu^�
��/^��Å�֟��sG��r�Ŗ��n��M���o������v����yֿ��<;;�}_�y69�ta[��U���G׽6���
{�ޫj�ImC��Ng�ղ��e��^ח����?�}]��o�$��W����w��۪�}�I�Ȱ��F����Vu�m� �=�=Ͼ"�Q�~]t �+�(��B8�`[ �b�CQ�?���_��n��G<��}L��M{Bx�t�Љ����C?:��I
[��B�m��K��,�Do@:��C�����U��N7�G�P���M��nI�<D��!�8��y�<.1����)A����n�y�A�x�ϒ�!H��L�<��C���A����nL��jN�-4��D ����A-�xm8�`Z �`���?Q�&ۛ�������Kv���,�L��K��J�!��kl����f>]�h;�6v���<
V���/W�h�v�����]���_A�\������ޭʶ����}�?PK   l�X,qJ؏� �� /   images/278ed6c5-ad12-4b42-b098-da68003ec988.png�zeSL�5��ww�ŝE���Ⲹ��ݝ����ު��3S3�a��z����1j*��HDHPPP��rRPP�|����N.�=��@�k�J@�ΐ�AAQ@�K�ky�\�<':����>�������w�«P0~�o���b���F��a9�5E�5�P���H�B�V�Z 
"D2�[��B��^:M�r]��/6߶:�Ӧ��a���X�9�lz޸0���W��L5HƴSʹ߯��l��4d���}[%�7u�[����;;KW[��1̈́��0�7��0 �LN�c����UP�ǒH'�13���1���#��Y{�Y�"[Bźq�kL��ʾ<�p��������#G��	��Ṧ�aj\��L��T�6���)e�矌v��������P�a\�4��Ԭ����ŐyA�^�pMZ.GZ�)V�:�S�J��		�t�¿E��!�Ӗ��}��}s7~!�t��(t<H�У�H&�K������e���qҭ�%&�8�R�c~ꉑQO��DE3'��t���k�{`��>�'.�
�1_,B6��<-�� ���m��1*���s*�{�YuK��^�w�B@z�R��&ed`?{�J��q��L��e��P�U��v8p����a'Af�N-��O>`��t`zi#������ap1�Ę'�pB$�,Qܜݥ ��ՠ�����K����H��������l��t2}�*����>ZM����u��=�~>�Վ��ih���!�y�tt2������дd���>�kL�E�W�X`_O��N	�w��3�V��ݧ�}/�-aDX;ڢ�{�Y.f�/�����>�
2����!���(1��H0/��D����(����yA�w��Op�׶b����(QQ��O��Ó��������
��|�5��a�a�<jUMBLp��R�1��	$~�������:\@qj_X��М�7��ɟ��PL��58��_��A/]j��R�RcG\�e{�ljS�?�H�+�[�$lz��X���i�:0����}����C�y��33�]`:sd�] )Ã૞6CTE����6I���֪�I���vr��;��P#�]�P�[���,2m[N�Ay�JL��4�!$&�b�2�HE�DŊ8�TVI�Ǽ�K�W�s%��5�gz�(��j��晎����O�A�8�/,4�ح���H�p*z%�Xa��p���]$�M7��8l�[�c���ӗjt���Q�������V��G�F����[�7�4���InM��A�;&��0�[&�ޘ&���(y�DT>�x���iN&�hTw�$M[hb��:�{�[<�F���_zf�FB*���Q���=�0���Y���.��\%7�h����#P��n��PmUҬ|��n�O>�{�5���4/J=J`��� ��f,���<H���n��*�������U�*
ć�#!y#�1�6!ӧ��R9��y�3)fH7��2�����Z|�c�����}7���t�u�`&Ԋ���p`mG�l+���O�|�,W��R<���o������lV?�ʈ.�� �犣��6=<���_��153�3=l�ѵ!�:/�[:n����@k�����zhygm9�҈Vd��O/�m��R�+�7���U��m�v*V�8�e�v��G��p�5Zr- Be�|N��,M�	re��ҝ,��s��7���C���8�(�jY��>y�Py�%;���"�u)�hq'}p��'��N!U����֐��$�Paˈ��&���?��(:�{i���2��e\( 6�>��%'�g��� ��C//��\��U+��Med�C�g1�.I�v0�n��5��'�â�F*�f�J�CqIcyKJf��C��%|�ڵ�r�w7&c�o���|y%%N��Rႆc`��f�P�g�X��~�[3�;�����"��2�>E��2���Hu Gcab0�k�UG�ӑ��2SHAQ���!:�}�Ӣ�c�}��<A�O��Naz�T�kB�:��Z�HV�j�I��9i�2;d�=*��48�:Ρ��g��ҭ~���#�^W ~'�T�������p��Я2����U�Ĳh|�q�`קJ�b|�D`b��g���'��fZt`��%���c��bȬ���n�B�!|���Ma���H���"Rc[������N�7�I���C�M�q�gY�bh.g��88�2G�w�(s�:��X���9��$�eM�.�\��)�9���03܌�2�m��9B�ƫ{X�%�vhe����u�z�3i��!f"E�L�-G��XL��RFE�����\^Z�kUy�B�w�-V�V��%[�������:~���/9����X���ұ�ef;d�w�����O����ݧ�e�s�1u�g ��
��.�
a
7���D��[E$%̬,��R��p�I�bȏ;����aP�lJ-*����h9�-E�Z�H�!*է�/����~�e��[@�"v����9.����:4d��w����5L���K�˴
���a5���Y��M~��9����f����*�Z��X�n�u8Vd��C����I�.��e��|����q{`Y
�eRJ]mW���K)����������c3�Qu�����w֟l����T��B�;���^,�m�[��`������~��"�$f���euÄ�";�Ƴ���`J��7]WU>b��Љ��>�(���qf	����\]ܪ��ԣ8x�fk�h^=�rN���B�WK�8��ɰ��.`Y	�#����������b�_����-/R��cdiS#Rd�n�Ǆtq�i�nQL���S�!0��n���^5�s�󕫙�6�{�q������S9�g���Jl�wu�|�]<IݎL�{j���[ 1��p˪ҏ��  ��3`�3�ײ���1�݊>w��Ȩ4��D{�.�|9*�
"��8$�-�j�$f�"zH�����!�,�^,Q��x����K�]%g��Ǒi�j��d���j����莁�f}�t尿�-�����_�@>���5G�x+�P�_�,u�:�Ao��
 f�!S��k
�x��$�c�Kt>1�Is�ؾ�*I3�Dhpf�8��0� t �Ķ��)LH(y42�9sbZ��<��*�u�%W��R�Km.�����f��7���\��Уc
����1��S��e �:�3�'t�VqT!�7�us�a�^^a%�3v��d<����S��Ub�G�x��{gg-,���6��!�r����������Q��a�"��6�Y���R�����J�5b�kP��k[����4�:[�&�2d&�]�h���58f�w��$�]�g�h�R�!OU)�����D����x/<��{�je߱~��3�%�gmZ��'K<�@��*��N,s_�u����F��S�K�`q�U1���?1릂��MC1u�bDj���F�	!7���߅=0{P�H5;[����r��e!�}EM�jqT�1�$WS_�,N�ǁ�B#0q���wfh<GK]_=�;s��I��m}Y%�jG@E_Zo(�R �3�2Cl�]��IN�u�;���"1�M� �C��"�Ը�W���h_�+%2�Ѿ�*��43�4�1�-�(�}D�W�-ڸ�E�rS��3����U�Q�'6.��H���; m�"=.�m_���^0z�F�������@魈5U��� �u���a�g ��[�Q4돿�DXg!*��~�� ���kL[��>0�`j"�ߙ��b�X���j�9�� j�#s��M��r#��`����n
��oUt,�b��/o|}�)*6p�c����0�G%�����?�{��>�wRK�I��)���E�K�ze2�@?��+ͅ�@��/�,�"8k-�U�SU��t��Gd��Zr��)�ޛ�臆w�(��t-��m8��[F�]��?��gGnH'1� R܇0)5�j�F�X#��bCl?��H�Z��T�nh��]��#mO�=8�����[�$>,��5)���Yb��H�z��]���*�����u8ߪ6��LV���[�r�)-�b=����Mǖ�*+�����5��,��$_�u����"��Ăa_��Dj/փ��{(�yE�ܓe���G�����ť�i.�j;P$�%��;Rx0e��Ss��d��u ���)�XF�t��K\�?���;6�2�I^}����P
J�b�J �F|�M�&��K�M0>)�����P��6����|�J�\����YC��)��]V���ÏLS�[���h�Ȭ9�Q��#M�Cӳ��~�3/�ஔ E>~�_�]0{Q�ϔ|�����ǋ �	���O�/��h���k��?���g���|ɕҜ2�w�i
N+�o7d�G�z.�2)G<�eޓ��-�L�ʳ�g
��fq
K�#&��34��O�� �$�H�2�>d��p�W�r�_�on��YlU�a��,j���)����<e�CWٰ(C]'��5�M���;;���Y���f��G0�.4	�63�	��:�bT	<Ys���BЌ�c��H��>��Pz�-j�
?�10�T����e~ȳO�>����r��]�É�-����'�oX����1W]�=~[����aZ����f}A�d�n��V�S��h1ʢ��+��lq.����>'�ʴ,(�Q���V�:{PynolNa$�f���;�352���2�	��.PPB��UζGUǪ7��$a���=ll��Q:NZ��v�zַ<&�1�'�(�v���`o[��2�b�:��v5��:��𚧰D���Ï�á��@�M����5i��d�<Q*8ci�K���p.L^��u�z�VWv>v顜��K�>=�/��!�`|jV:�E��!;� ��pAx�U�.
��9��񣄞m,��P
Y�1��xґ�x�Mz{_mOM��Q;m&[8�Nq��W��H�-m~[�y@H�i�'��!��p��O�&�P, ���A�T$'�T<ݝ~�`��&��yY�F���S�?�Q(��C�+�);��d1n�8��^.L��Y#��W;�]�V�T�V��..�Ջ��}6�VF�C�t���,������m�׉��*�q� 6D�@��7�{�ő�@���V��J�t��ƅ��� utI ���ڂZrw���)�\'N��s�#��.y:���'�3T�-�����&5�><$f)R��s�M�p[}���F��F��X붣�$���%��XtCCF�m#���5O�^�+���e�~���t��c�umYȘ�}=����sk�R�c�<�����3\�� Q79�3�~��XP%�rb�RǦ<ɐ�#"�q�PKw�x����h(1����!8�S]�˱s�ӵW�m����K�$Db�>���oy�rA<�Q�(��#�>�5B���u^���m��&f��E�4#�E�7�6��+šR�0$pLPAX"
��8&�h:�D=��-��&-!�����]�l�܌�!n��Y�ڀA����j�,m��FrQ�X�92,V�TF�x(�l�v��X���G�%a������\'J�+�>�"F}�y��
�k@�7#aJ������:@�їK��>|�%�: �\ª�	����`2`��޵T9q������vʿ���Nyq���o�����dhS�ȕ��}D�]e��@	 =2(�?k�n�eA�8�5�:��L��;!>��p�SO�[�}Y�_7��4�`��/�� 4�,�/��lMd�'>O�`������xk�����g��a���
�x�sd��5�㟕��6��[���k,k'N�16�{�X�БF�K���?2&�	����N�[�	�҆ �}��)k{r3#� eg�l�-���RH�{?2W�w�Q��ڡ-|�h����]���@grS��k���Ԇ�^7���8Lp	c$kZ���F�y�6����"���hBry�j	C0��4��+�DoG<�]7�#DBe, pcߕ,9�`k�e�\:��ΝN�� �Uv$áD�I����p�9�,���M.��s�S!��p|��R^�M�t����8��u������^��j`ð~*?��� �4F�XY��M�ǿ�b#���ic�?�P
���VlL,"�pw��6l ���U�(�L���cZC8`#�N/�,�y&b�Ջ�`��S�p8�1�qRϠ(��aAF����=}�UR�.k��i8�����W	o�E��g�|�6�$�}3|NY�ӞIST�=�����Ѭ�w�[�`�r�:I�Օ������^&ͺ�'�[�(�06Fa����������6��j@.�����v��A?��e�/{�s�}�i1�[?�W�g�v���R�EEG���QM��ң�ux�Mb,َ+�8S~6 mFy	GUS�`#=�?�8�>�9�'�)����T'����!�(L ��DHp�{�m|�����2��<
}�����i#7%� ���+J�Wv`k$3
� `�� d���S�m�ϡ~�؆"�*:��4��F@p����ɦ�	&���x��yD��O�IH(���vo]�}���5i�Z�{�v�{v�|J�[bQ��`#�Qd��r��fȶg��B�A��U.h��A-I�jki��	>���|e��rm(#�V���:!.<�����	���o�	����:��p.� ����vX
�[RE����� C��?��T���(g��߮[#9�8f�&qz�����uc����Y���	y�[7�瞟�sFqxՆi2�{J�f���0e�!">��nF�*y��E�[&)R��F�sR��D:گS������l�m�ibh1��ā��xo1L�`�PG��;ZhSh���ֈ5Ƒ�כ΁r�A�[�3Գ�s=^������������p	�3�/eX��������{���#k��,����Lo�P�),����|�AAe�J'�,��R�E���u_�ͤ��	/FjN}x`�/���]�_��%_QN�;����*�f�������N?�L������ ���W��'��|�F�f��Ws�;A<-���H���$�9��]	x�լ�=�/z.D�XRK�(\�N�ᓖ!%gP�q��b��鮣C���N�&,����"2�vCCIxh�)#����~�zU�#�}NY�X��t������R4Fd��"�	@�e�ǢD5Tm	JC�5c�p�Y���g�?BX���)���^���9�J �O�w��˛D߱n�P�3?j[����3��tϞ�B�(�N�����- ����>@7йe�lߛL���TO҅X�C4��&g&�k(��Nm�2�}�-��Vg��ʂ�<�1�RA�L�s,=C* �q��`�p���-L��k��~�WO��C���HI`�]�����$�Y�����Ƭ���W�+b���&I^��`���aKT���Ǘ�<$��YW_���8�fAҟu�w��$bo62��������Y��x����{͉6'�����'�\���s��a��J���ݔ(��_vI^Yх���4���I�hP^�&h`[��u��,QZL�r�����a�T	A(-Ee���	�W��gà�����ݞ�^��A��D�����>!z�[���e����z�Z����'�k�-����HS�/Ew��)c�= ��+[��!Q�[��H�����bmI��U�{~�ϡ��:���^�, Z�M	)���.�~`��s
$ܧ/8,��O�3�P�>%w��m�W#P�)z|.ܵ:�g��+'������Ǖ�fÑ��@M됺�����ŀ�uE��.�Mza�E�X����ҏ��Wc~3{��!&�V����՛�&��r��N�VM_�Gi.���8ޗ�J@s!S�4P[:]��O�n��R1.eܨjX��P��
y*�,$���;kn(�Á��ո�@Ʀ"�z��|�e�}���~_�JKH����
�e��-9�G�4'��U�煮z%��|W7P��""�NG��u6w�l͙O�3T���ޛq{���������*�k��wxIP���	]ՂaGR�	{���}�#���9��9:ʟv5"�'�S��%5�x�&\e'5FI4ƾ~�_/ ��G���g`�43A�C�ߪ:�|r�x������/�746��-�s%��JwbyN��H܌or����v4�ّ`�#�g6t�ҏE�W^L��]f�g�r��sh�v'�p2�;�}�w��T��c�wA*KbٵޤX�<��6�mm�WS��4e��R�i�&MD��x��R�+��	�҈���0d�6�/A�fS��f���� ��Ń�g��ܐi	X�Ÿ�m���`Ċ�ǑM�75�O֤9�A.����}��~p@f�/�����:O�E�MG��9hGB��p�����i(�]Z��b��	7����-Ɩ�6��U��8��?���|/$��bSlձ�:Q�a���E��Ö�	��G=�+�
z��#
P��H;�����]���y��e���ρ4݉��S�9᲌�i,��QJ$�y����~\N�P����$؈ ��G|��qs�������N�ȣ���o����Q�(�xYj%��\ACb�=ew=E��G�Ţ���'_[}OC�O6�kG��y�?x�KɆK�=�ܥ玎I<�B��ަ�e�lԜ�5@��D��O������������r�S�=�� �� ��KYbD����RKhMq������e4Ҙ�憮(���rMJ�<դ{tR�&�P�~gx�>̫�lS$p�Kp��	\Wa����]�U�*~\����I0**!�B��}�-��|z�����f�T��+iד����A��l�r�
{k�"��b��Z�ZP�4b��������'��#��S�v	6���A�d��_1.bz�uGp��݇���d��g�g4��I���%佰3��ɉ,8�@�.&���ed�S	�d��*�/�$�Ҧ�mJHf��0��Gq7���#u��=�9�d-J8P���K�븻4�[}��6�FԘ��gbU- {MG�V)�<�:<�����3�5&՚���"�IE����*��ߵ��B�؂J��M�fH���2��b6d�R̃]��e�!��s�B�`@��mR-�,�|ʳV+]�_�F�1�|����.݂z*'�չ�~�i�W���-#PN&dS��n����hW ~"�EŠ$w������:��"bn���ߗ��*��j666UN��Þ�:϶V�N���HXv0:�?9�����p;��d�|5�e�M4CN�)D��&�����=�A�r�U^9���#-���3�u@[p��`����ҟK�6ϧ|�q���.`+,&XV*���v�Q�|*cU�-]���C`��L�;e�ўvt�Hs�3� ��ըe-�m�� �J�ƵȒ�`}"��ĵ�U�^dzL�y]l���4�I�E����=}�p��z�+���b��r�T�rD�y؅V��ٵ4���]�G��|TY�h�V�����n�ƭу>y%!���UXl�AioP3p&9�ݪ�~�2�G�ԵV�9�ӏ�Q��N�Bs%�m&���(w�h���2&�=��j��zK͘;f&D�ߐ�>N	KR&gO
�ʋ�B�y�@y�Dۮ�����Siw��Xj��ƾy�vJ�DQ�Cu������B��u�����2qjR֥�9��?�?D�!eT]�%�L����y������9P�=*��S��s�X.����55�*�q#b#[O��~|�l�Ӣ_+���J�D�ea�e��lvn��n��R�.tR�Հ6�`�4I�f𛳧��p]Ҥ�(\Ԣ�ϣ�խ~�Ⱥ�^��nu��r�� �Ξ�h�
EӮ�k�\��ҟ��d�F�����q�Xٍ��L� O�<��������7u����cOl�_���-�8��4e��zZ�����.ggI#����
��'�bRܓ${���E��OY�ѹϐ& ��pC�076d����,���^|��A~��5l+�j�?5���h���˳���؎�b�R�蘆�8(��/�g��H��f�Dퟕ֚�Tжs~�,]���}�w�
���y>ݞ���:����������;8pDGZ��]<��
��pʬ�޸Ҽn�x���謚.l\�#n�q&�q��7{�w���n��	4y/�6��zbB�B6�;�3���DJ�3�g,�M4(<� ��S'[=iϊw�c���ѴPY,��n��&�m Hb{@���䕴JN'��H��Z��=k7�50�!�s��@<n/�3�~�D�s%��!���Mپ�#��S�+N˿�Ke��ւEM�  �5/�?��
���R%��FP���8c,����	v�!!Q]p�iRP{�|GS&�FA[#���޹r;�`���N�]h=�& �8�1�nP�2#}�)c���OYnkʚo(J���h��^����g$K���m�br�ո���e���M��M^��k�J���S=E��%@�^�oVѢ#��)�[�6����s���M��}y@p��'������-0�<�2�L)_�ԻB@�ګ��%�΢f���`tV�b��4����xj= *�k:���	Nyܓ�+~�Qo����*��H(�I�b�©�PG��tH��=�Q'dʆK>�!o����Ysʃm<!D�S[@���eֻ�����	�y����y[b�y�e�D�d����SE�6/Urt�g�SѠ�Вu��E��T��ZL���H`ɀux�[葮��Ǒ�T���$��z�4T��K"�V�<")|UppԞ�\���MI�����^�{fn'n�-���zHұ˯���%`L�Q�p�W_(����~�AlW�ԝh��{]
���J�xe�1\����Ñ#v��'��<�$��j�����?��3��ߪ/[԰�.O�"J�z E>f�)���F{6�%���y�u*��;��)�I���ImĐ"15r�1��-)!�Y���`o:��Ǥ��Ь�F��)����/��ì9^y$�)Q�'�ƨm�t��V�����.�3�>J*����K�R?�i��9Lca���vdz��3FB���-���tU�ib��6�kP̉'_E�:G�I=���$r`mZ�mR��OC>M�����<"�͢�m�	�ߛ���F���,�g�5E�$�����ߦ%�D ��Ύz����A����"�0B�������_}�z�;�"��m4BSR���J:8�2�?�d2��8�|[��yҢm�Qo�zd�W7<mP�mc-��n	�T�����E��#I�[�^!�X�Z��<#}�>��&
h���0�TYjsſ�x���\�;o3}K}Y�O���}x��
�	�:���۠�_�Z�֑]}�G�^sjm0q*!\Q_ą��/��g�c@��˻0������/j�n0XKz�������_.����t�
��_/�(�&��v�yG�<��䤦��aW.�"��.�!�8�j�D��K�R��4��RG�������Դ�t�}0�
�K�j�����hm-�[�z��#�t�Wo��փ���D5}`�@��κ2L���XA)\r���J�#� �+9a��z��N�bL�e�Fp#�!�:�QO3��l=�I����=��[Ðf�閄~�\{R��
*�J���P�\+ts�O�j==��iqh6y�����F�)�`R(�Ǎ�1��b��t��Ϯ�H��fQ����}��pp�P�f���c�2�[�{CM�5��J2�����&���(�O�-ۙ<e��g��)RO�wA'nԡy/�����ޞ�co��k��N)�Y�܅�\��s�zcjtTn��#�UL��KR�UV�ne�@�a)���C�Y�sg��`�������T��4�7Md�v���1��df��L
�L����忐�3��	��=^��j��x}�cP2*����A��͜h"�m�y$�8�q
�q�����`�w��	�T��=ȆL0胛�w���)V������i�J�9�f�r�)t�rB=X̧�m���Z$_E����2�U��,̷�����)n��h���o9ʀ�")�06�|�y���qi��?^)gG�N�^�#l|��h�����7��Q3YH���:M�<��駒�e�b�%g�#V�\(L��Ǫq�n��?jw��$�̭w��n�.�~�͝{���JX�����+PXY�������}58CYzare�z��eI|�H���
��a�8��-n�V�C$\"������-<�X�Mf�{�L�(�R�}D����/+z&���Tl��4�[����nw6d@%�;��\Ke����ie��a
�qr�t*�OVՎFp$�i�G��{r��l0��"�~��}ؒyۘ尢�G[T�WH����b��<D�y�6Y��Y�x��B�O�Y	�����qԈ�|��m-N�U�g��S��Ë��;Q7����IKi�|�!	2�qK��~�������YG1��v5�ONT����9��$�ö����l�����G���Զ�H��zvP@`ȸ-�u��h��"���Q���:L6���Ov�A�	e��P%	�6M[M��df>�|+�Y��n�������)�w?:{��6�˅��ף���?ώͧ����Aɤ��p�%��*!������kve�aվ��Öx��I,0d��)҉p�#/&��B
��]`|�L�.����i��W۩x|���~�z��Ԇaw��x�Ȣ����>��v�?����g��}��nQ(}�fl^�3�b��"�Ġ��Gwr�7�j�c����yH�E$���Y[驭"F�َ��@���_�eb,#?�Z*�Yi����Fboh)�r�W<��k�h�Ƒ�؈��$X6��<c�ה�h|�c�Ƀ��o���:�!D=Q�#�b��X�"0�@S����%�uT{�̽��BQ`�\&Q���U����]%�N�z���jQ�M��<��b�*�M�g�](/�ڹ��Hg .)itԴM��Q����(�<ơk��Ü��\ٴ��Cw��T���:g>9��?��g��/%���^��u�<�y���J��E[��-�ķ]:_���IuF.��]mIi�,�}�F�ݯ/�b3<R�{�/^�"���'��U�Г����KB�%��*#�Hh�)���V�#�+:d֗c�g�hg�#�����巸H�����|\@�5%�����o?x�pߖ@��[Hwn�h�Y����:�SA	P�{�X����E��j,ݻ�mh�we���n*����d㥊_�	�;�L9�%���u��������0B�&�n�
!��K�Y�3�T�{��>̔z9C�m�=�1�J�9��������������)��hm���05�-����p`'+~���������v�:��&բ�g�tũ�Tz0�%���,p<?�ڢ"-yڲR�c,K[�p������=4���yo�^1�c{�ƛ[�ᴴqʝ��)> �a����;a��=��p��ZB��B��<�C�u&G&05���� ��N�͞U�zȝ��@Ra�%�` Q���&т+�=��t�Q�!	��FE>�H)Q���mg媜!���q.̏��%��UWs=���+{;R��w�ԫ���v�&o>�&J�uF�s`�GF��,j2=Ƙ���ՆF��4W�	�
�V�1�D���)�Zd$��G	珃����+����y�ZN�q87���LvO����˩��l�$�=]+b��-l[ �K�K:(���MD�l�'�}��}Ps0	��1*���Սz����|����8 :ls��f�³��S�t	⁨�Ih) N�3RYS�!C�o��C�.����;×�����y�m�P��Ϝ��C�d�s�Z�LـV�a�N�!:�1�����/�'��Y�c�9eA�DπJ(����YU޶�#��7Ag�3/4��.��7�����aw�|��Y7�� J�+3�$��ܣŶ��1Ms�b��G}�tm~\��Ƽ�^3[�G"rL�dO�w�zc�����[xcO��4���ZM�ea��z���������T\�
~�#ϒ�S����}�c�U������w�������؅�����V�ʆ�����!y������xg�"����Ӿ�{x��V����i&*pN$DƓ���5fp�=�V���2%5��ؤ���w[�N޼�`�M������풚.�6��T|���t&`�O����R��eK۬+/�Y��5z$�JJI��][Ӽm�A���Ɓ���(!���P0&q"���!�1Y�����`�p3�"ʛ��KY�t����_!�,�k���G�~}�?���������Y����$?f�A��aa=���:,-"�"�|�����.I
��>��hmcc��^��_���~��O����!�h�����^�9��mw �]�+O�?��;>�X���dŶ`��>ȫc���6��Y1��b�����3(O�47�@6�U���o�),$�� ��Ŀ����e�|2d)��Jј[J����X���J�/M�����-�����G�D�����<��Z����C�b���hCK��%E(c�d)7�$�ٓ�l�NR�\��dHl�-��/d=�K+<�+�7�;Ɵ+."�e7g�O]ooB��q����AW,�Z�	�Y����H�p@�[�k�_�>3�r"�r���%~"v��c��a}%�MQ����ZM�mK����� �X#Ų2��6X�)7�����c�h��y*�u��7�_���{3q�謻�$�B�Z�]9O�oL�?_ĺ��}_v�:��[	 6�-�H���� �L�+8��d�˯��mm�1�v#t�c�vN1�h,��h"i�JVW
1%
}�;�g�Cc-�Df�\3Gߤa9�t=���qB0�� �&a�ɳ�ce�♼D��U˙m�rf�?چ>������\�S��-7�s���~�x4o��)=6�Pv�	[���N�0G-l*�<�D&����/��(ntb5�dB����,le˄�^Ka��]?�^��=��T;��q,���X7����������9���`�`V��bpD�5�`J�:Su%�s��vpO-�S�ؖ7�������$�K�L,�eP(��hjB�6�c�ĝ��v��f��T���`��w9���ܷ��=�,6:���EN{���Y�XE�=v���`���>z���~�G��������2��~�`��J�&����x�7Mꑷ�1�B��|�i���W3x���Z(A�6��.7[�a��(�*w�g��mz�mm!�.��w[���]!\�`��[Gk�t���v��\(�\��²:w���#e`��
#ʥ�}p��������5�A��S�8y}�~x=�Շ=g�:8�O&³��e1Z:�9f/R�6&�W��}��'�D0g�����N�{�6f���jc�C��&��It�=����_�r9�k�!�-�[�C[��V�e{�F��l&��AK�|�:�e�1�a.8�D̑��M!�WKo��T��_���G"��
���j�����0�D��e-��H[�{�h��A�{mkcV�~��ؠ���7��7�K_�k��&qNE��x�� ����x�L�m#�r@F*��F߼ no�өA3}-�������زej�$��
���'st����z2�t<cz
}s��9��Ҕ���js"��r��EĢ�t���T��;�y��ة�,n��*N��D��;[z��e�4�f93�D>=�'��`�*I�L��K�ʌ
���v�5H͕�+J��������O�aQq_q�7�	��1n^�J҅1����}��W�7���נ���V��Օ�<�v!�u�uiuU������^$r�H�d���ŝ�/ǋ���z��`��;��M�Ŷ�Ah��>�
��hmx�$��h�Ãnњ=]%ah�`g�_pDRI��[j�Z'��`��-��+���þ�+�5p'�KJVB�3Y+�m]���]���ʢ���HB��QZ����>�P����V��+�#��{���|w^㵳��1��F����U��S��p`����=�
�����;�a{"O`
����"�:��/��/RS�vQ�~�*���u#���0�yW����֥�pR���=�4R��� �齔�N�.��[
�:��^�$��&y�M�wy���p�*��f]v�A�n��w??L�w��T��7��rף$l�~)��$�S�3�e����=��}��m���M1��9�lL?X�w�@ eP����� �'��o+��Xs�TV���RY_l���)p03�ҳI^]�<C���I.�������3O�Gb��+w��C��~S;��F@�|I:Y�����"�ӵf۬������}��Dz���� 1@ο�;=�1`����c���T�i�˄��r`�y��Oe�ܕ��]yH��:����Y�2-+��p}���dݙ��kJ��nwZ]IV�;�
w��3ߑӚ�h���L��\4�5�:�jq��y�������cL�q��IS��O���;��10鏥e�k��X۸�R,���SI�	�cW��6�[����&�,����#�����i�!s���'�h�䐦�������P3;I+�X��R�{&��J��=R�-��-P�R�̽G����x�y�h��s\��#t|ԛ-8��Mְ#�k[��vĨޞ]!� �E����}�L���Tp��p�b�T�4`}x.�@��J��oon}�o>�S_�����õ���9���u��/F�8p�lm��s(_#hT4Cd�q���>i�L���vsʎ�˲���M´|6��ux����Qw_ߺ/��茦v����p:�Q���ˡ)81�8Y-����Ǜ�b�����^����q�\�<U)*���w�Z�«���C�L���{�5�����������}Vl���s�ŽWi�ￎ�J[v��ѵ��LlPo���:w7w���)�V�]_\b<��jʟ0��|z���3\\_����ɿ��`��E�ՕҞ��%��}I�sAt�]���g�$;Z<(B�v����u2$�����4q#� ��*b!��aW�5�J�*e��?>x���P̙�1qb2�.]Wy~u6>���L�,ӞU���,��N�|("���q�eXJp3@���il˶ly�T-� l�z��T�҈a�	ERp�)�Y�zP�1�-�b�p|�z�%̍�� �1v���^�`�ݒ	�޴�h�����d����	k������h1���)N���f����l�[�U�à.a<��W/0M�X����ÚWǃ�=���2K�]���D�t?1��PVJ�����l�KX�L�p�3��H��������&�G��]��R�5T�X�D�i4�ۃ��M�sDi�rc��PG$����0��pq�Τ����MRAg�M ����_�����z�_��M����A�rt������h�x9���p�qL��j��:p��&'�)�hbx��ܑl;|�.�̊�ƀ̀�'V�����������a�ޕ��/�p1b�/�9\&�)%�T��1��H���=��w{����x8�˃}|z�/  GȉfS���MT���/�1B?��Fc�j���yI��/�p��g�n6����ob��$����O^��WR�J@統�[����AMy]]KW��Z���kaTϏ��1���v��Z�7�=�rZ������-�7�k��{��3���c	c�fx�H;����߽�Z���/�^�r0��Ύ4R�V��67k:ЉR�V^�""5�J�z��'8��2AT�1;��ϥ���kzy�F�RYa�ͫ�	�l��{|F�[����Ķ��c�h�L�ڞ��b#O��x���s�h�ݰ*QA�	��n���S_3 ͳ
WI4Ro6%�?q�N��l�-Ƹ��5~�J����6�[4��<=�x0�>��Z^�.�F��$L���֠sN��k1osc������&�-���z���|"YҌeMܘ�|��0>�4A U	�)AcG_�_�$c���p����Q)4��1��K�_�7��H���U&�V)�0[�$�qisʁ0!�y����]1�S$��}`B
i���J�
�＾��k���@��?|��s=���U�[�Ѹ�jr���Ø�o�wK��&�6�[y���Ow4�T1j(O@,%�fI���T�Fû0-PI�������lW��,��#a]l�2Չ�/X�u}�I��	,��'9�v�xsW ��x)pqy���H:,������D�w�����XX��ݵM�t7��X�8����?>|.m�x��.���oJ�i.��� ��G�/ğD��kACt��;w�t̯Lf��ȫW塿��S|J=lp-�D�erf��&��k�wP�*�__b8H��n�%M?S�����������:�T%Tz�{�����OO�N�B�.M���S\�_���L���������T�'WG����^�₭�L��dΘ!c+w۲�Z��x�s�^�4F,����!��w���b�Up�Nג�-$\��5��d2�P�]����dcUa�`����D�	��U����Q.�	�&@<7�͂��f�NN��p<���'#aml�?*9��T�fҊ���Zn ��8�?D�^ܭ?Py"ِ��N*�%��}���5����f�c� ��:��"��o��qӋ��W�)C�A���C��l^J�լ@1#��N�W�HB��ͻ�5̮G�'3�L��.�FM����I��<�YE�y��$�x��D����5y=-H��G��U��V��[�0����Vm���_�������s��'�4ϣ�o�����.���h$]Ab%�=�s���
7Z,t*]�3��Y�i���a�L�&���� R#�2���*����6�����z���V�q�	�;}!��S�Bmw�k�{�6��Z]�@�:�d&�d����Q/� ��:��h ;�﹒�����쵷Џ&x9���t�����0m0-'�^��O?z��bd���x�է¢Th2W�qy/l_�ؕ�P��>��j��NS
����T:�0��f���0��{xc�.*:������P;��z��[��g����ở��Q�/F�x{�~j�ZA��d���K����ְ��`~�Gc/�quy)!qX���֑��o4�j˳h,����pM0��Enϣ`(X���]J�2�g7������Oi���Y{�(��2��C��$������[��ye	�8��sL��Hv�`������P�\.F��ߨ!hTE�=�>�񠏓�DZuIa8=��t�H���X����i���K8r(��cs�l��D�o3m>G�f6�~����Igvz��E$�iN��YY��<7c�Ô�zF���Ȕ��3.7a��p!�$K��2ֈ�����P���N�0:�����]ӛ-���D�	=�7�&�(�q�	�9"�!���f<���A������I�BZ�qO0p��8���Z�ƃj�{o��~����������ӿ�pˣ����/Ώcා��:
�--\�r0��B�V]2�L&�NA�����s��lG�m,�V&�b�2i(�l"#�R� 4��^[��z�s�I;��1N^��Sn��7/��:!z^U��vg����Rq�3���Z]����O�H2a(�������m�6q���/�߿���ev���|��t�:h˽L��ы����sb����1y�>�l졃��k9��o��@T����3<�:���J�X)�w�]���|l���E��5�om"��G��>� ���]����:�n���}����s�fS�}9���@vJ�l1�K]���Sn>C��ss�FH���!~����j6Ģbz󱽻l[&EgCH�tT
����N��nle�?�����˹e5��	���U �tE�tK��*yFn����sY9∿���an�4\Ut}ScJ�$��N��LF8�8�97wCI@�<�z�38�0yX8u79LYk�+����34�r
�#�,P�d��4ղ�9��}�{��\$�ȩT���I2;N2���27nӲ���(�۶Gc/I��<J���<�?�3�Ј43]�<۪u�̑�� ���@P�ʜ,
�nJ�:�o�T/�@Hd��}�><�Ǆ��f��WE����$qƤkg��To�ۿ��'�s{���vpv�+�@���dc|����B!R�ML�����v�NK:10����RGl�����#�1F�p�t��N.a)e�y*��{Ua7d^���*\��q����L��~xy��Mۛ>I��w}O�{eVem]��t�,wB���	k�`��+G8º�[������1B��_����$+l�Ax����vO����^�U���9'+����^�2뗿�9�y��OMv���L�⣮��VE��Vn�)��)~��@H�+�S�����D��vqqa��u��vQ^�W�����kO?��o���(������w�^\����ݳ�����x�l2/$k���=�i�+%��"@?9ۗ�	=5�+���׮ʜ��-۫W����+�B�w�X��jG������������ V	�oo\��Rզ�����dz]��E �OE��:F��4??�P�B��b:��G�/>������3�n��C���u>w���r$��5M}Vz6�-c�x�	��QjI[o81� ��?�4�5�뒨\��XkKN`�Kv�a���·޷ʠ%[�Z&+��A�X�8����5���M¨��H���N�AcG|�`i%��Ap@�ՠ�̶#�,����mP��2+<�A��]�𺰰k�E�4��!/��c4�*6�H�T�y(�M�͓v%[��+u�QY�� ��J�T_QO� A�(:q��`�SY��V�V�>}j��<�l����t�wϔ�|A-+&���ۍ��>�������g��O=s����������d���~s�y��^�έ;w�y�[o�,�l!c�U�[M|j�nt�
J��dxp�q���,HNL�=����
l�z�����;�h�Q��ΦC;���"nx3���3�����^��H�Z�� �1a�B�r-`� ��o���О0�8mX��B}W7�m�\Ӵ�i�̾�졝t[
nd�uTPJ5���>oEN��Hgt�軹AKZ|[�{;7�V��������$����S����ީ$dFc��_ߵ��	�e{���<)|��6��t>��?������m�<�[:��I���+7e�c��u��1e]�VmhCWn�����MJ%V���������o��Ak��Y9aX̭Æ�Oh0���iPџl��d��PI�g�OM����s6��X@�&��h�qoT�z�"��&>����eϣ��t�r�50O��1�����oF@�֏|.ZR�AO?�k�QA�e�6��j�a�8D�m�����q��A.w.(j�~��)���w��P��paZ*���2]O*C~�L��6�-3�-c�3O�V�l��������	WJV�V<H%��P�ɢ2y+�+V\�h_7N��G���g6Ȧm�����frj��s��K���An�V￻u�K?}�O��zp�gO��{���ͤ��~�y�5�[g��07"�rp��^�UEX�/�I⡹1�#����E~���,�zR������jlr�w�m���Sۿ8����ڙ�d�Q�e�6�d��B4���l�*��&������^�r��k���i�JY8���MdO���M�zi������d�u5٪��j�~���Y5U4���L����}���eN=��Q(~g��X��?�e�ESYJa�j�R��zf=��.-@  �~v�����c+��={�����P�v��u�n�[����g��}|O�[]BA%��[������,��<7l��ܘ�0�w�qq���;L��i��V^����e��ũ���nO{���ՃŌ�'�S�q
��u�e�W��(��}�����k�od��bQ\`�)+d�xӦ(Ie���Unl�ː_"�QZKG/@QD�p&�,AO\�\��(�����b�F�9�H���̡lf�M�ƿ�B��C{���y�;�$�-{�FO�נ0�Z>d��T�
;}���y y�$&z�*cCEC���U�O��&3K�'�c���X(&V������N~�nml�SU��Rъż&��*�N\\6�/H�%0>1���S���c���Sq�KW����	¾�7U��ٜ��i�,�޻S���O���۽{��O�����J�7�݋ݧ���`���[6ҍ˅��R�����.L�bp�E��4��|�Eo�((K�	MJ˳��O	lL<1�`6;m�֓��mHi�^��|b���f賱֧L�
l7�v�&��vW��F�a�~_�
)��o�����Ll��'/����v|rfk���]�ز���(g���}�����q���@�ҫ���;�Y-[�Q0�x��=y�J�}ʴZ�lw���[ۻ������R������Ǉ���?=֔�MF�d�٭���E{�쑽x�L85L{�67%�������s`�
L�����[��C����ྮ��m�V��������za�^_�\*+��׼�K���i������٣��53��2*����W2$zNP��b��4ذ�u�V�xz����R�0H[�T������,��+�R&EO�^Q>#%W�����oJ��yp�8JWB��rm4�0f��V� ai��I-�x�S��w�d�l�R��^�zMݮ~Ǭm��l	n��y1�&�%���+��D��x���!1p�%��iT>��彾�_|#܇`8MR�?9�BH�3��Ԭ:q����۩���E��	u�\��C�D3�ǃ�`2���3���S{L�m8�Y!#�n���rI'���2����M&�y|�\��nm�K_}����O?s�������W����׻��%��ſ�x�1��APɠ�&S��M�de�@pSO@^wE"�qr�`" qL9y{s��"�e���xO�W�4�dl�6���Fт���~�n�7m=Y�).��;9>8�����5[��5�F�����>}bGG'��n�\U��^��h6�����)��������Vϖ� � j���H'��Ų��sU�Z��|6�fk
�B}�Rٜ����Sp��� �+HO��۪�Y:���/۳gϴЮ_�f�[[6��=�{�^�L&+H�J�h[Ud���yt�v�B��T��jkO�����v��#a�nE�@3E{��]�{����gO������n['�����i% ��L�Z��J$>�>_�̺��:}e��|��u}���q�Z�l��ғ1U�X2��D!�jp�3.�E#9D�n�����x��Z!��4��u���V�L� �����Lf(�Cp��*��+���\A)������#��Ȭ4h	 �f%���Ւ��Tt�O����WN���1�I�t���?�}�<�kZ<n�lr޴d���2IZ%�l�ꅲ��ܱjP��������:�/ټ��};l��G/���TA��%�9�U��!1Bb��bN��Ap0l+���V�Fe�����/���w?������T����L����ō筦��ܰ���0����b�}��nH��|=�QJ$�+��o���YR��Cn$YN5U�	(�G�/���A�&����k������,�tO*m��M��@DO�
K����4}%�^2��/m���:���nn����j�DN���2���틆Đ�ښ��{�n�6�bN�o�)�r�"`ϛ++V.�,��Xo2�������)���Y>�e"ŏ��P�L�X4��kkV�0��������+Q���^�,�un�g'jēa0��	p�HRYk�έqv&���ښe�EM�����/�X[�)J%M�߿q�޻yW|�.��sj��ߴǭS�ȑ�QZ��+��+��6lw��G��hHB�Lm��ٸ7P BuT>
�Y�5��P�W8-�\
K����[i�b�M(P9�sPjP�e/Y�ܭ�
{���	�����<0��~�28d�N��;�E��RY(e�P���:���b��(���C	�ó� ��lC0|=�-0�� �~7��|T-�I��n��$�LiE��n�L��,5���i��Ya4��$a��D�P%A�i�ه�`�*JIe;����ϥ� -�y1o�H�!��Z���abn��2|�����5�Q�}t�����៽��V����%���o�x�n��~�H��Ʉr�Ӌ�V��� iKӀE�i��.�n<dw�* )-i$��go728hX�7���_��fv>�ڣƞ=9޷꧅�����C�%�Sy�-⟺&���̊\�糱�_@\��-&F}I�<}�\e�c׮�fm�J��Ok����m������?�ݏ�    IDAT��sl�J��ԯ�-h9�Z�t�"�Bl��ן�ub���E�ey�U�^]��8hm�"e������p>g�L\�n��P�7��ڵ�i�M��Хs�?�MK����tfG�"ts0mno
��9�o<{$h,2#d�y������Z>Q���oOG�}��|2�pS�1=���tz��Ï�sq.!�ב˦��_�T������Lq4������C�P�W��]��jYN�(�LȄ2>���v������ԱoHt�}��s��ÓЮ#(RƓ�!N�)^�yώ�}|]�t��J<�%KE�D��dT4��De-��A����Ofn��]�{��NY��>j1�ʜ;`�U=��)j�d���C��T��׭� "��T\o����W�x��4�T��0DR�A�)�6ۓ�u����!x=~f!o�\�0iF��B%��'?����n�
�땕��������Sn��<�����c�L�_�.n��l�}a�	^��/UA
ٌ�֪��Y����An2+�d�7�w���ɪ��������}k�nW���@ے��Ɂt���oQڅ��I8 �����.��k�_��$J�q�X�f«�5/���L�X�Z�nׯ]��lA=	&���Oͬ9٣��;x.&��tz-SP�x��%����"�U>��vl�qb/����Œ�^�ت��	�x�;Q�΅2B��{~�g���
n7�w����0I�@j=ܤ����z�H/^>a͹+׮Z���W�3���'��t3.Pɖ$���7߳��!�ԜtD���G��`�u�|$��Eo�`�h���葍�=�����T�o�խʐ�P�����lw��j�a��g~A9��)n�Zm{��Lw�~�ǰ5$�*���%,]n����)<w)X?W�|��=k������ީo��E^����gM����#�L2�%G{�w�A��Pp���7����1y�l�WXܖ��(O5H&<��
HX���.�LPP�-"�y2�`���K�!�%�0��O���O�����I% ���AS*4�TJ��3Tq��1�1��@6��DJ�T��G�*�_�Ͼ��o&���o�H39���^��^�#O�J�����V��hj'�>
4��k�d�*�5 \w��E�^A	Z	�D&���d�:�<���t(�Dq��hel���/��&�.2L@��¬#��J�
��[��&z����Sm(��L�0�EE[�'�*ɤ��=;���e�e��;t��f����)��nyU<�Z��^*g��g~�{a/ώm�����<s��U��^Y���8�lzרp4�62f�"���A��:L�,a��]�o�ݝ�V�3ov̗6�F%f��ؚÞ=|�XN�4�77������.4����Q������œ��ݱ��{j�����u2�� �K
)�h�ƅuON��՞%F#e�������BS:���-�iB�S�X�B�6g͖Tn���MA6��ٹs�j�����n���VP�V����{�ܔV"�226���0(�@�n�Q�COL_�G��9�/ q��;8�����h���@;tR{ 6�+ý-�0�~n��T3��ϋA5NKcp������ z�ʋ���	{Gz{�Sw�S��h1�E��Nl��I �i�7�~�).8�f�Q��}�eQ(j�,!Ӕ�$��)2ⅼt���[=7�U�&��zꗯ�3V�aT�~�������7Q�����o|���$��{��p�z��� j���~!��hܳ� �ɎgpLK@C���ݟ ��H�i�G�"糺Qh\1ES�����w+�R2�DF�*�Z�s�k��d�V���d,��y6kyyZ&5�d�X!���r�j����K��p��˗�PNE`�k��Bߧ���w�۔we��%�̔{h��ȕm�P%R�N�����u�a�D9����K+ꉬ�V�m˄�Y�.t�Fۿ8���c�L�j�۸��,��߲'�׽��I_��b��7k��Ǝ���=;;�
�^iqA 'S��y2����u�N�w~n�t�6V���ή� .Wl6������yOFS������<?��GGҽ;��P�P��c�[[V�ٲ����x�(�eJ�``�,)8�)HE3ᐹѻ�ِd�B��|��2��@$��`���ܔu���Hg(Cxb-BB����xZ�
As����yp#�� H�L+LV�{��Kp��P�W����i�Q^^[�v��s��Kug�G��#R��rF3A���0��{e)�B��L�:��2�e<��]!yz���~�A�T%��u�KYe��+���v�˿����(pC~�޷��Nj���������u��r�W+�� nk+��q�����2�މ^�2�FzZ�|	��TdH�x��oJQP�G-�&�0`c�'��T#nzy<���3����66���@L��~r��5<�,d��JZ>�����{�C�a8��2�$�
,Ӊ#�	n(w�n(�rȣ5��  ��@��8 ��L�k�^D��Jq����h�R�g3N�W_$���k/Ϗ�=�^�R֡�x��=�C
W��ȏ�RE��R� jپn�Q �d��d�������3k��x��a7vw�R�u}���uϛ6도�ÿ��X��ֆ%�Ee�4�_�ۣ�Wv�n[�����6��t�R��U�.��^2؊�3��d�72M2y`M\=3c={y��Xֆ�&m��8s�5��k�ܖKWk���I��-�����Ջ JR��pp��\V������G���U��n����<���Y�� �i�hm�Z�
��0����� ���o�#����w��dқ�h�(��͞ڠ�'jGUk�čj���\���_x��?}(�7?����~�e�y�aK��[n���s�,
�fD�+.4q�H��X�R�B��)� �Ç�3��^� S��&��FV7�4F+q
��2=�I��_��-���E��wx_N�Мv��Ь���4��-k@�%<|6�Rz�B���gs�;�=�$q��']�&��	)��:��)1�ZY~\_6�.V#�	ƈrj0=6�g�ڔۀ�O9_�s�2;g�%�&�Z`�Z�)�`�l澱i��E!�3wK�.�������l&S]�ܺGG��+؝k���R��Ǣ������u.Z6���͇C����2+�n�k2��'��ϟڋ�#9���5۸q�ҫU7���ܝ�����x��~$�
G����0\����^!�$�*�G�wKJ���bƶ�u�;ۢZ����2�͗�c���<^�p�XJ
<#�%��⥠� χ�����%r�t糀!T�($#*i��cȒ�x�#����k����q����=R���F@=I̠ӱa���G��dҮW�>����_��|3�ۯ���/v��_��]����B�Gdn7�C0�-fnL�(����J��dL�K��ƓџNtJ��)�D	��Z9��]�	��[Ӊ,�Z�!��I��L|�s�@�`��Ef&g��Z��6����sH  ���V5�q�m�Wx�HQ�l�z�f�f��.�fZ�L��o$YXj�R�4Α���u����5�p��YRT3Q��($�+2�.�c�ϝ��]�$��Dod�Sl�&�5�;��p/��aZ	r_���c|?�#�����=4�l�Z��ߺmwn�Tߓ���ɹｲ	�2n5����v���=�1�~m��v�,��"���<�{/�˻��vc׊����C�g�M)W�5n���j. ������æ���e�8�:�| ��O�F����9�ָ^����/��9k��q���!��Ep#��L�$*�D.i���n��Czi�����we�P2(���Qr������8T�SoK�"�����4��W�!#%�-2lwl�i�`��YM��Z���W�����O�}�Z)��{��w^t[�*�!�Eb}n�<P�� ��` �x	ntAbp��wHi;'�Y������.C�s9e�}T:��S_dA?�HTQ�i��W��O��C/#��c@^%��F't������ד]�A�Q���U�?\�g�	���� ���"��h���G$�+�I�~y����d��?�e��+����Fb3@Y�u��@�Jd�D%yVp��F�fP�:�>|a��~�k��N�}ї������ū��ڼݲ��U�»o�{o�U�ot��b'��3d*c����3�Cύ�v��;��{E��?��=x �YP�U�^q�s�bz;��=�������p8����r%��:MNAHA��Cv�9_�VA0��ŀ(���I����q�iMj����������	*�B� %�IL�إ_���:��X�k�-`	Z� �yJ�4cŢ�F���a=����ٯ�=#��C��"X=&&aD��̍�k%dn�g��9�Q]���捯�������_�˙���+�ɇ_���<�+����^��
n@/<t0_��Fp�8_�VZ����$*b�R"�SvG��G�o4�U`�M\�%��ZɾI�pSq�̐����দ/Z�����m��ZY��!��g'=3~&:Zj�� �R>�Ұ�>���1�]Dk���`B�h]'}pH���zM����QFb���UpKӌG���1��鋦�I�.�!��ӐԀ�ޤ֦�_E(�b�/��S��������(��͊������O���9�Q��]���;�{�>s�m��v�����O�uz��-س���4�����{�_\���Ͽo7߽+�>����c�F��%��l���k6+ᰞ�YƁ����:���+٥?L}�\�E�_��$<p�W�3A�c��Ob�X���=�p�}�z��kn���Y����t�	Ϫ"4�@�,�Ḟb�KҸ~����D=f^�1������E��bJ��g>'TD��M=D�<Z4��q7Ț�������� @J��;b�$Q����e�vce�[�n_���}ǟ��B������{���^b������}8��t���̓��J�H�U�ג�� ���Ybp�&�nP��\.�7dqN1��`/$��θj�^%�[�)J�59���P`�3e)S��ēe�+�����\jƬ��C�CH�lU�y)�����]�pJ�ᩅCp�e0!��P���R���F��oi����%����7| r*�ۚ�G"��r��@��B�w�l̠������"���e��n�l��{B�^�Au�`3 �V�����疄r�HM���[��}|f탖��ֿhJ߂�`L�g
n�Q"[>ew���v�;޳f�o�|���{��>>8��0�p�nZ�Z�I&�iZ,K_�ܔ	�m�33��,(
4 mRpx�@�*��R�y^�F��$��	�6�qd��� ����$s
%�4J���*�r`:�gnq»Ȭ�����%ʕ�WC����дN���!H�
K٧$�F�T�x��v�&Ke��h�-��AIK����&��	l�V�R7��<s�ƻ�׾�s_��O߷��k|�[�ѯ�L����x�m��L��<d�p�_��m�Z�M��-�iʨ��S,N�����!�r����!4d/�� ��wA"�=��d���,0n:7�gt��4�r.�u�	�`Z�Ҩ}���E��҄*�I@��CEj�9_.\JB�GS& B�M��W�en�#����1�dqp2ҬE���{�R)����c W�����%�@��Y�&��ܖ�Zn�Ә<���3��b�0n\��6<:�D�k;+5�������Z�ٵ����:j�Fß��i�!5�'�:J�6ϧ���������Q��۷�?������֚]}�m��G�D�@1\h\�&�y��X�A�<$��kǽ'���t>�L%��k�S7!v�m�U��*�82]Jϩ̓���#~ͳ/O�o�<�t[C@���|=sM2���J�޸gD�Z�u�����]�{���� =�X[�[�5Fd�.������!�ܘAƌR�W����8�dճ�S�X��LY|��l��Z���ۛ[_�����O�����[��}����Ѵ�|K���2����� }<�X.����U+=zI]�r ��8�Ԋ�B��>=��s.8�+>��&�JЃ#������#HH�؅����b��喔fy��3#"��x����M��Ұ��׬�b�.'��bZ��`�MP"0�>���K�.e�Bb^�e
� �G���H;\�C���Ү�e�%;Yn�<�&�9��X�Bh�G(L,a�����=ٜ?`�0M���wtj�W{6i6�F�n��}Ǿ��w�]?;����5�N�(l}7hq#�c�O�jEKW
���[v��M;h6��)���;�V�n���6�&m�v5�jy����o*�tA��I���I��Jls0��7������u�� �5� ��*'�����F�~j(���m�����O�/��ƀ�վ�ղ c
<"ԇ����1X^քQ!��!�\�f��&��7z�E|Ո��d*C��+�b�Z�A�x�$�!3��j-���B���T�
���z]�6/�yrf��Ȫ��frv�����/������܆��h��.��^�i]���c!�fc��V)[?�lF����m,����JY[8U"R:��:pCV��6������ƿ��}E9�M?b����22�%h(��5fz��U^��Q:�9c�L�\��3N�������Q�,F��!��{t���S�#��N�O�`�e�^3?���"�����`1�)&�l�2�� 	�u�^N�dY�Cb��)�H���3;y���ggv�Z��o߲Ͻ��U�%kv�l��Nl�ș��6)�MFC�������m^ߵ�kW,S-۫�c��o߷��{`���77l��V��!�xA��@��b�L~U��J��~�2���A�L`�`4�X�`4�π���0���9�B4�t<�y�sܴ�CSeY�S]�1�����(�,0�����U!�����4�X�4�����Fp#�f�E�a�}	ؼ�>$>�Jh���Gց��� �X�|�2x���Y��N�VRܣ}��J�$�?�ҽN���;?<�$�-��5n_kc�K�{~��bL����c��~���<������'��=s�M�Q����6�v|�\�Z�l�\F���c)�pbVG�Q�o��4(�ˆ)���nUl �������e�8�W��IF�b
�I�.!{�Âۢ���~C�;�|D@�� P��AZY��`26��K�4)�1�d}���O�FD�{҃���
��g�u<4�cpW�ʧ�-���侄���_|*K	`�ȜC�\_f8�a��Ξ�s;��b���\�woݲ��mˌ��:���k���l8����ӱ�77�Ɲ�v��Y�\��;<������gr��_�j�wo�����d�Mh������~D��&��HO�� �}�@bK"f~����ʠw�����L���<���±�&{�)��*��Z��B_VW�G��<_>�MH����߅��⿝����f���2�K�9�����2Xv>m��Ot�f��>��=��c���.g������&>1�9z����8�����p�W�{����;�������}3=��ѷ��|6�GG��_v��-���7Ce���JE�~��Cp������N'A�8��P�."�aI�A,��5}2��p_ �f� ����6�����GMl���&����"f.ң���� F�C��c�B���+B�zk���%6�>`n8=J��5Ђ�LB�t��K�j�ZBp�%8��{!�r-*��n�\��Q��3��%f�.�,�2S������Ȧ�d>mw��Ş��,?��nm���ݵw�߲�|UM}TB����8�a�e=)��Vm{{ۮݺi�ׯʆ���P���������Œmߺn[�oX?�SdD?)�����a&�9���#鵮��'�g�{�ed�� {aヰ�����M
��F�GhDI�0�Jk��t�z�/+o�h@�:	�i$�+P�Q��奷`B��:�?�1\�(Gcv.�Q�;�|��L����^c&���{�o%�0�    IDAT�����NK�{9���h������Cѹ�gg�r��{�������o�n��������{(p���Ϟـ���	n��u��I.WH�sٔm��(���(K!ד�)[�	��A�a��a�-���&%�/)�.�C-��K�-D '@ؿ!_ȱ���S� ��)�`.��ʽ�3#��ǣ>��7�`x�8���<FJG��E\�M�gL`�Ld��fR���?�l%��)f�
�K�����׵�	-���i��M���/�P0/�9.��Ѩ3hv2�~ߺ۸ѰJ6k�k����v��!-~�A�ٔ9����t�v��X}}�Vjk6��%��t�Ց�?}n'Ñ6�m��v3	����y�h p�`E���@�0��x#��ǀY�1.�4
&h�+k_�*p�5qV�^��K஫����{�漃�cOX�����cЦ
tSX)����k �F��dv���,��'�'y"L��^����ơ������A������TZ3_2��ts����)�����р�ZK���45�~���؍���wW�_�����o�~�k�}�b<���Q�Ͼ�6l���_\s$�|S�ꕊ�d�M (�5�Iצ�*24a
��%���rOA�gR������)C����?i|\\��
���@]���E�QX�(��M@�c�"��8�
��¦���E���A�}ye�d�Jz�V�-�A�����M����cQ��]Y����(=�ˁ��#JZ/eǱ$�����6�g�p�����	���+���*1g����u�ʒ��D޾~�n�^�+�V@�+�p��WKTB�=���Ɖ=y�Ҟ�|a��^�)x�\֪�;�~u�*�����1cc�C*� b����db/�R�B
o�>��a��u "���C�i�(���p�	�(V�}f�����KߌCl�8Pp�wy@ꀉ�~i4ٙL�Ճ-�R�Bo�C1��lKx���ˈk�ZY�f�,�c���"k�~ z9���	h��%^&�6
b�>:�+R\"Y}N��CA�2Y�����L��@n�^[�����?���������[�?|�1������;g�n0�D7��V[)_���
�i�0(����?�=7q�B�_g,CC� �:=�������U��ei��2��9u*������,��!����v,P Y�g�B�1@N"�1�;h���Yc��_���L��Q4�q�� �Tt��8���-�/���%a�*�z����m\_���w	ЌX<�v³
�zra
F�IT��u��:x� �*n*���e���H���kW��΍[��Yw叄����|��O�2T����e�DS�\����v���* os<vK���������+�'����c���$�"BVM��Nc���B�`Ʉ�ҍ2k��.�l��=F�o*%��{�\B��D<�*h �a)�r���_)[�a��Q�(`��P��e���
�:^z3�->�����Q�Őt�Oh������~	�!�f1N�I
�풵��!������oPia>�
�M��Z�xxgm������O_ύE�;��9w~e����dn����g��T�e���)[-�4-U㑑5zN�U�%�E+bc�o�(f��i�J���ͣ�E?�Er�CRf�Be1޴es������2�t�f�hQ9�xh�E��)�xH��<<(ʘ$���(A�D���IY
�)p27Jt�^�Q ұ.], B���o�,�`�E�/ �������^���q�
�}�����̘Ž��-�"�/��>�\��+���<8�&�Ε-�zu��[u�y��|�8�B����� $O���
n��"PY�ش��W-�|�4H��/O���A��z�[>��p��t$�F�����@.�������@b�r�e�@BPQiK=�el���d��9������D�_@�s��S�Lʮ+���P�v�-���C
�D�)E���?������C\!��+"�ju��ʩ�3�P�K�zAǋ�"���}�kI�+��̞ܒ��K���A����2әU�YqKo���nm}�o}�_�_�H������t�?�4�E�̎�7�S.xhBͧ��V�Vv(���s}��-l�� P�<��c��ʦ:C/B=2nZ֋�<�U��K�?��MҠ����4��o� ��G�
F�yd�L�u.�� �%�SS���=�X������&%HJ�M"�$�,�4��zw(���*$�45������Ri�����&z>����������eE�/���@#�$��0��f�a��D�)�W�Ҥ�#k�:��}\�mkc��;�
n�ٳ��m�t��B��	���	����{2�)Wk���mk�ۈzO7eγ*�����F�G�CF�+}�{dݐ��y��L�1F���Ñ�;=yAH�k�'FP����L/���V,S*Xf�$@1$��̤�t(-�]��׀&LK�n6���Z��p іp�\ē��Q��^Zڃ��X�Z�	�'��Ik���8���
�A|�6�7V´��oCG�Cܜ�+ /\�%U����vvp�~-&�8�ߨ�������������F��o?|x�h���G�������-�*p�/�a�$E �����Ven������
S;�T!��iq��)W����jn���.M>PXj�Ƒ:�(o�_^�sC�� ��Ù��*K������~hDx�rI
�\n>����F�q�$T W��=E�m�'P�h�r?������o�qPKe!�z`���J�B�/e�
1j���@A�1�8ڏ�M���;Rsh�Ee4�%�8��xb�k�ڳ�鹭����ΆK���1��yhzc��Ȗ��e�Ik���CM�ʵU[�޲����Ҧ))�6�٫����.p���ۚ����2����[��o�??�n�-E�v�S�YHbǁ��v���:_]�L�h�k;
�����R �\����?�.l�D�/�}Ե����b���5��o����Q�\88�r�>��W�QkE ��¡�8ߏK��װ��W��F��Rp������M��w�C �g �Of6���Xx��t�Ꙝݨ�?����տ��~�y#���ݻ�O~���ꠇo�X8#` d����WVl�Zu�����P	�-"��8ʝ����F��Z�,����zhQ�%6a_n1P�����ˆ��X� ����Ұش耬�H���}�:pbȀ��p�7�-�0����3M<#��ņ
��"Ǿ���=Ì �8Q^d`l�n����M`��?���D�����g�1���U|G��,0�ܦXz����liY����a�d.E޳����׬vu�V��,���X�i�&>,Io�Xd~�_�:я_�۰;���U77�0͂��*�q�(�QZ.ʦ��E&g�E&�x"N��G6j��}xj��@" �R��Ŋ�rY���F�<Me�ݮ7έC�/�KbN`+��Q:C��3�	YSQ������ x������Q��eq��!�8���� ��$��}R;�"��z�6&���3��5&Z�A�P�6еbO�nB�Z'\���I��?�,�m��׳���g&[�zV������_��?���LY�����i$���p��K��~�Zӑ���8�K"e��x�R��ZUcp��h�3�rnd�u�s����}7��!���[���B�%BA�C��=f���s(Y���r��l��*���k��ظ��)�B��
%�f�����Z0Xp�鿂CP��2;�0��>c��Bv'��^hRD5Y@T�K�-�L�,s<�x�%W<r�Or[�=�@M�����W�.��@�D���Ԕφ��pz<��ށ��ط�鹭��ٴ��
�6v$-2?�9���RM�X�4e�/����+���kV�r�V6�%�I9:I���\��5�C�>`D�sh�3�
�9I�2;�6[�?���E�*�]��Y�#6�J�ads6�~^%�Ս�䘎��i���Cy�V�r�Z٬�N�=�M�6Ce;����5�eb<��S�����A�
Ce��{lj�Kn�:Y��L6-�2�x��h���M�.�z�ڇ<�@	n�PՒ�[ƃ(,���{&�A��&M�#�8B�&&�1�����-i����9�����z����?y������K�������IDs5�������p�y=��܉�R��O�tc�2��SϘ�)Sa���?(���zm����Η�S� ��uOJ���QElZ�6�~e�z"�`�d�X(�;�t����R�$ʀ���XP�6�`��l
T�s���)���*>i9�LEb��P�ohH��B�F�r1��\:�JT~٥z9NK�i]
�Ll\]�8:�+��:?��:��ۿx�o�W689���u+�lXi�&��<�� ��l���,� w���"��Zmc�6�]�1�����i��Z& �#OWc;z>��32�.��	 �V׆gM�^�,��J2m�\�n�����3o�ֺ�} \�C:m��TϹ?�E�k����<:�g���G�3K�3�R�&]msݲ���������鵅��Ӷ��NS�̸�
���v	�mM�CpS��χz�J2����r���r	�F�A�.ZHA��&�|�c� �s���N�@�t�2OhX?�|Ђ��oY)���b�j���V>ڭ���/��~3=��x�����ˇ��?��рi�gn���R�EP[�,����	���N��1�ի�ORGb�Z>"�'��h�bAh��S(��R�`�� B �T����A�~ɴV�HȌ�Y.#g"1���-�Tl"p���K.�3u��c�8���>b(9�A��AC�u�Ӝ?E
���)�i����ؗQ9A��~��	�JV� �� �d�:����52 �P��4i �,*Sڵ�������d�\��e%�S6e#�N3�	�Y7qh<�0KI����+;z��f��hY��+�ו�����9=����F��
Su�D4�կ;/�ٸѴi�mU��J5{o����ڶ;W��Z����#��Ƴ�@���T8��hl����N��H������;���V

n��U��Lz�Ҕu�lH��x���I �j��
 @Č���s ؾ����d�RY�a�Y8��쇣��9T�s}3��K$9Tj����e�� t��1�p�D��PYiR�e�T �N��TZ*̳nOmx�7d�7�����������)K�ɇ�lLz�`o����s;v�5C7ߧ����s�9<7����@-Z��ďL�d�@�2D�X�.��1Ê�S�(<Xŉ���Xp��/�'����,�.U_��
��4�tr�ƭ �.�G0Ҵ��	���|J��r<�%ϕ�e�(A�`Z�97�1%���2UpY��ʢ��	JQ�
3����d�;��C'M�Y!���7�?k�/��w��.prl!(3\
n���in2��љ�2�<8����ֺzf��Fi7�v�L�Ge)rn�T���徂��ƺ[%��dI�vc��)�L��B�h|2:a���ڴѲ�i�2���Y߲/ܾk_��m�**M�Aw���1�\�q���NXG��L���v����\��t��V���+�ʖ)��3�\�,�a�x;��]���שHS�@u
�X�&��M�B�_�a6���-�G�3jé�;�"bq8�Cm��co8������Ak��3���Xդ%������2۴ӵA��Vsy��NӒ��/��̗~�ߏ~���,�ߺ��ab�K����?G�wam��S��T����JE�W\�[=9�S��A�#B���=�%hT���b����z���e<c�iX�����H�^V��Ȳ"4%Ja�}B���??����)fNy�|rm* �����$I����"#y�e`�$|�[�f?|�@�T)�˩O���BiA�jv���:�^�/���Opk�����H��<�Q���b.�kl��Ȇ�9.�b�dqjf���	�g�Ⱥd��{ʝx<��e��a��{��?�B�j����qmG� �	Ls�!3Ar6��,���utj���*��eW+���!��>��A��L�ik��hOe.�M�
�������Ƕ>I�F*g�s�=���>oo�\�N�a�'�"�c�S-����6K�,�8
�ٜ%s9ktZ�vf��_��q��:���
��5���-_)�Ӕ��S5�=�:�.(�(�
Su��z��!N��^������UAɇG(�q�k�Ԙ`�׀y��uE�b��>���UV8�n%g���Hi9y>t'��`J ��2��*8:Ɠk\H��Wf�<	轒��F>o�d�6s���j[_����!���x������G��_~�:M�.��*ͽ����W�@A���F�*��D|�Ȳ\~%�2�i]q/	$�`O��+�[�j����7?]P*N�TN�t:���?@%� '��q�������G����
�|κ��BbH�=����^*���.��b�J�L����^6'�9����ﹼ7�{7��:�����r,�EIr(%�5=v �C��(e�_j�E���BH���R�'1�u�O�}�PZ]��+��DPp�i��+�4��+&�)�}h�Mgv�w`G�r5���Z�VR�n�NY75�)P�� P���(���>��t&Չ�Y˦'��~�gW�Y���i����ݾ���}v|b���ey2i���]ͦs��RE�Чٌ{��X<����+;k^��yÚݦ�Ĭ��H;]��?��#�w�f��R�2{�#!���uf���P������epsO�~K9̄��[R �h�) �������e������89ȓ�%�%�����P���H�����I�o�ߠ�i@�KF�"=P�z�yBÄ�L֮���lm}�?���pK	n�I��mn�skL�b,7��
UP���b�!�6)���H�W�'�1c�1��x�pɿ�ZZ��%B|��8-�O�F�F�߇<�N�y��(���P!�#H�?�pX�|&�y	�T$l"��`�K��OT���>�.��y�g�k��ط�e��L��B/��X΋?�p!�8e����-�=zn���[d1뙰p�Y�K�v\8$��-�Q�Nj���3���9�Ȟ���-9[���N_�[���V�׭~m���Rh&��q���+������+k� Y��-�ZR�6�g�#��gY�:����U������5W��8���6<8��q��*��w^}˾��_�d(�c��Tr<ku���U�%�� ���7�������zސ�j�Ӳ�V�F@D�vS`"�T�l;�SPbMh��l2R�«����	�XC��$��f�^��0�CBa#��΄��(xQ�J��ɡ%aWS��6����:�AȪ2��9Ӹ�J�
�@�8H���5�ւ�:������j�w^�θ��}t"�[<K7��^Y{����/}���|x���x���'��st܂�rd�s�ep��k�m��O{Mb\)+����=�8���2`�t
���O-��?z�"q\�`�;�%�W�b�*M6���6��1��2D�J�(�%ˠR�dAfH}7�SL'ɘ�
n9>I;S�^��<
	��V��[�u�qC�q�<c��:Qf7��l0)� �� ���x�r���` � ggS�>*�i�Nl2�R\d� �$!àI���@��Rޫ$��R�A�)L�
�Ol�^��[�mmg���senP���2 �Iijbv�����S�y}}�*����n�(�i~��9���<q٪����/Isx�`l�Fӆ{��k��ݱ/�y�n�n���vzt(sh̎��u��Vk5����� �ƕ�S���	i^���hbpb��s�6Ì{D�S.m�lJ"	4�a�`|L�C����5�]*�� VI0+b�]�I9���*�a�Y*�-����?�ˈ�J;��M��1��d�>Y��<�l����S���tgؚ�̥mF�W%��Fc���$ ccVD?ήS�!ӛ���[!ܷ��xF9��&����,3�[�U(�
��������Ko�����ݻ�N�����1sk�'2~��Q�s�Y[]�y�-��1�ɍ�q �^�~�i�ȶ��E��d���    IDAT%xǲzO�� ��zX����ô���\��c�M<�CL��,�2B
���(�޴e�'CM��Wd��I+��V�:O�L2$k��7���m0���)䊖�h �@RtO�D�ol�^�� &�W:m�NV,b�H�ޥC�(H&�7�1љ���h� ���NF֙e�,S�ࡊ�=R?�}�;28�%�pe�A�]��Pr��,㩥(�)�jk  έ��e�+���4��Ҭ#{�xi��uq������Փg�B�W�l}g[�3�M@�rz���ax�b27�	��KYy4��ѩu_Y�ٳ��;�{���` �/^���
E��*2/��Z�^�r��y�����Z�߷��3�h�����:���_<?����G����+d�V)t�&���3�W����1�D%�Br�(�*��e� �^)�J��k*�
zO����rYK峡A��A%a�t�JlKkvX;kw�9Zk4�TK ;���ƛ��)��V?.���E�MK����Oң��d5!�9�١D�C�	�OC��Pb��T�6�y������ͭ/�ܛ����\k���h���g�$���t��dgSvk����rU�8� ��pWS4�2T�@�K��EI��[/27o]F�c�fC�z��^B:�z�8X����(2< L�q�,�����H�f��mVj�^�Z1���ƹ�5,X��������U�y+���X6�'�	��U�z`����0�$X���W�E��8��TFY�;H�3)L�7,\�F�N�6�m6�>�w�5H���ײX�"oN���o:�b����^�&v:D|�&��@��o��L-75����N41,l��ʕϸ�t �$�x�"�Ϭbi+'2v�乽|�D���zݶ��X�ʦ�)� %A
J}'-G"����L���y�f�A�p��Ƈ�V�������}~��T����.έ�R�r��u])�ʹ�����JyŚ����G�������ҧ��6�ӒL�8��e23+p8%R6L�6�J\Z�U�>0��T�I��g*m�l�j47�**V+���Rԟ�H�3����>���;�Ǹ�&�@�&Rf��#�h��E��Z�ױ�f�·I��(6���l�d�BQC�d�ȇ�VM>�����Hj�)�L�>�We�ʰ�=k@���
ȋl�n�k��޺��?�?-��ڿ.������ÇW�����p��+O�'��fc��Ƨ���e*�mu5dn��Ud+D��PS���� UM�X܁�A�Z.G՛����g�IQ��
u<�x�OqA�5$�p$�lz��1�!��܂?!x�:I��ɰpߞά`�8i��n��������t58`�II�� 뢔�4NuE*��RK �	��M�f!�������dp��"�^(��ZD:��\N�R# �� ���U>4�=���"���:ӑ�㛣�����K�u�r�E���>��ٱ��^�����\���əӯN�mkk��;u��3��R����#��k<��<��~�8��m�붵�c��d*K���:��IFJ]�#��;����a�f�vr��Ʈ]-�X���c�i�T��b!��<��gtk'�����8<<�o~�=/��A+K�Dq#��M'*,M�!�a�+clCx�T �=)PAd,K��y+���5uK!�V�K�J1g����V�V)��R��Z�'��"��[�=�K��!zod����Zdn����{v����E�Z����c�M�Z((�3��\xm�B����K9�W*6�g܍\$��p������x��`s�������QI����;�W���ߏ����7���ۯ?x�s��݃A�=i�������d���y�):BA(���D���U
�B)�K\3*�/�@���ר��k�ޫ�}9y�����8/w��.�
$��r���q�Jl�ғ�{�f�.*H�3��%s�C�TɲVN�l5Y���v��i9zOé{]��V�笐-H6�EE��:�FQ斤w�ʦRҠ������[��ݨ�SsU
�tk2E0�8���.U���tt�P�AV�i��:}.��%ď���=ꫴ �#���q
����M�Y�1�zt>P���s���Ȅi'F������i{w�j�V�׬G��7��9�!��:[afVIe���{�̭����k
���\����\_Ӿ�=&���6h�1�[�շ�q����Yݲ+�T(�J�C'������+��ʦt��
`�����h4v�޽�lA�
%2�R�P?�Ih�Q�F㞳HT҈�f�8GW�����w�r\-8ZD����I%Xo��Y����r�V�˥�V.�m�\�|!+s9t�J$�� 6����l�T��L�?��2�s̳[=�����`]�J��%2�w^�-W.�k�P)Y>���}1c��$?�i�ܚ6�f>#C�$�t�`zhhTL�ܮ��>{o��O����;Ϟ]9�������?m���_�X/��Q�T���b榆�z5#97qCT݇M�8�����Ş�ņ�ӯ�\x/���JQ�6� қr�4'�z"t�u�?���(y:;��f����P�w��A��6�aݞ��
��md*rU�(T����x8=���ɸ��	��Kf@#f�����E�o�S����*��	�v�c�aϱB2�ť�UW�`^6w�\QpC��+&xm�,F�ܒv
υ	+Y���Tk:��^�.�;"�9�1zR���Lσ�I�c��
a~<��{��5U�n޸*U��q�� �{n���wcZ:���v���5�Ҁ�˧um�9�x��:%�M��sj����gM+��v��j���3�.U$���u��m�� ����D��jY�?�~x�fggg�p�`U�#ę���LlZ8��Mq�
�|��)9������AL�)w:z��E�O4�LNY�?�Y9�}��N{O�TT+D�R�9�N����1���|no� �m8i_��3�&����	fꕩ�
A�
@��Y	\��
���W�V�	��r�晜��A>m�b��oy�yd0�8<9V�Cp[Ie�����w6�����27�������Y�,��uf�\J��(%�Z[�Z���$��G?aJRN���WI/%R��r/����R�P��!��`d~%-$�����@�9�>���d��h|�r�)�ԕ)��POe�Lp��,��m�PUp[�V��
�4��P��B��B:��Nw6*��� �ٍ�OK9�CZ\h�y��E#�0�0�M�~O��6Q�(�v�-�� ɩ����\AGc����c#��U&�	)n�w�-�Q�A��sa��s��۔����`�MPSF��")���������Z���a�wm�����LuY'i/-ūM�\(r8մ�a���g�o��-]�@��B�Z�0�lR)��	|M��T����<�v�捖�[�NV���&��Pxr���g ��G@��Y�^�oϞ���Ź&� �ONN���H?�P sJ�{}�ӱnD�=5�(p�="ecJ^����5���pZ��%���(q�)5RR^AV*�z�E�4aʹ���B 0�eq�6��G�Ɓd	�ѝͬ��e*7��G(� �r��5�	V�j/ŁP&���z��ڊUkkVZ�Z��f�"�(yW
�^�[;�� �I����*a���!�|%������ln����s���HY�;��_9���Ѹ��=�4�7܆4f��i:�(�M8ͧ|��IJ�IK\�e��,8v �#�	u��]["�������\��$��Z�Vx�8�2 ��)e �G0%ԟa�`&ʈ��
ɤSi+�3*S����T�6
%����V�E+1k��jڠ��b���ɺ�x�M/D�;���S��dVx7M@�Ы	�5-L��Y��O��& /(\ɤ�2a�8[�����$=<7l�8�.����R����%5��N��6$S/��un�A׎�m`%�i��2D>��k@��3ff��#M;;Ƕ��i;��Պ���kM�
n��s��GSKC����=}n�fG�m��U��^�Y)��8J��1?S(zzX�樯�ĝ����Z=��]�V�mm���D����&���� �wi!PV��C��N��N�N���T����3!��Y�wB��A84��L:'�Jyɿ�%x	b	��1<�&�Pt�R�ϓ��lb��X�nR6�-QR����2���O�h*��dB�}�h%3xg{ON4�OV;jED�<�IK��N��0��?�ڪ�VQE�X�T��j�:�������u��n|ur�-�TƊɤ]�֟��y�������	n��v<��$��ʎdf���
�`�ŀPe��j�:w�#�WC��4�4n���X�JF����B�Ʀ	�:�Z�'%W��0S�9i�Y9����\4]��jジ>Gb��BY���z@��np~�PZ-���m=[�j:oID�#AB8uz:��EeN2���H.W��i���F�֌r6��
��z!���@!(��^�0���GV@��W�^�i���ܸo�L(��NOtP�*�E��|еT�h���m޼���������Y޽�y�s�]�]�}�����&G��(��Hd	%�%(����A�3E�8XQ� E"���>>=5�y^�<D�����E�#�J�]�5���Z����s?���l���0������S.R0�)$bJp:����l
oNCq\\i{oO�z����݋������7A���z^�x�܅���:y�R��Į"���v�*�̓��
�����`}�V�H~����*��\�uF~�r�^�B���(��=�&�O�4�M��<�^_^s�[��P��7��PI>C�>�&)V��`Z:�8��d� �`s�����<�p��7�R�r��v�f�̦.�\����+[��ёZ���p�:Y��{�7tmKMaF�	�/�d
�عqbF��;��0=1*CU���A����*�*��U�J��m׵h��F͓Y�hp��a7XE��v��z�l�|����������ڊ[7����ɿ�|p�{޻��2(�mx�6��j�N�|��Y���]��z�����M��"i4�j��p�$ܴ�.9�eY#s�p��_���V2U�Ug�<^B�l�����ڬ{5}�����ZW���>�����tl\ J��+h�^�v��������C��b�?�I̅�Q��ظA*�ڧ�ډ���Id:������֖�{8����gKG�2;��Eȅ-R-$`�aC�!����t��	#�ƹ�T�����/]�V����T�ZE�J�7���+s���1f S��>(e£�/Ի���ޞS�_��+f ��S-T $��@��G�>���4M�
���j���m�c��q�ύ�ր<b�hWo^#N!��
k6����F˫�r����E�Sym��&��~��E�G�F�l�.�8���Wn��'�l��0nbĽYKՊv���l�+���$�K~��w�M.r�-8�u:�D'G�;�h=+5��D�����ۡI`�Yi>[j�h<Y�uq[�5烿�I+vN�o�A�����*`n���.eyy	����FGq��)U�ʗ�~��V�ZE����2��&��^�z:�������(2���v���_����^[q륗�j��e�p1U����0��e������Vf�pAc��ѧ�`���J|���IcĴ�zt{��W�A���En:68Q�:���v���U�蠒�2�r>�Z��� ����N{]�&#��b����%��FL�- %�wXRg�-����5rZy��PI��+Z��-�`#�H�8���8l�ӯ�$"� �=_B#�> � Q�5�E��[0�LrF��j�>@uԍF}0ٔ�].FnF�ӫ'cwc�N˧7d�|��q���aj�>�ijm��@����/��g���w���:���˃R=�͚�:(��ʭ�>�?}����p��Ζ���U��xc�g�.��U�ͻ!�d�����%�':���n ˫[=�������խf��F��8@������+`h�����y��&���á�D��w6���JV�%U!��h��3p���]��[2<����<䵔Z��Ȓ�b�k��ťJ4b���ឤpZ�J�Ɣ5���Қ���.t<1y�bF�-7.����@��:D1X"�hOVِ�ˢ�[᜛�r��<&%6��RU"�'WT�VѢZQ�U�׼���/&���OM����REq{g����O������������/]-ǿ���&�7��G
��V��v�鋂Ԧ�r�غ4�(p�Y�=����Qqta�0;ڸ$x۝� �~�A01��\^;����5��E�kt��T`�Z�� ��[��GR<��n��3b���*W�,��кQ@5�i�)�\�)"A7Ͳ!gAζ��r��~�:�~6�o{�h�c��>�К��Y<��d>t:�R�H�D����8�-y��DF�]���7B�"a�1GFQ��c3��sC���M�6�az���)�kTUh54-�u3��z1V�Q>R3��=��]�������7���k������G�a:��r�m2:����3M�5�;��s��>0��^Ӳ4�Ʊ��sc�DT�&���B�ۑ&'z\mbi��٥�X�.������L�9�6�n'>W/s80���!z챽�/���;+WJ��:2N���*��>&PQ�x^���!�N�HG/����`L8�z��z	��-}H碸��c�kF��,5c<��Mo���=d��`2�-����xj#�2˥��5��i��,�iV�J�R�r��^,�SQ��P��ЪTR���fM�jN�ӡ^n������\*���[{�?�K�k,��~��Y�������٣Q�{��۟��Z��{��߁��'#�z�&v��
c�#��Ŀ��]\�J���YT/�	s����c�LN��*�ݯ4�](i+_1�ݝ�O��bͳY- })pZ�r8�y�F���E	�M�RQ=_��75��H�r����֬2�2 n9#"xl��.DAYh<�߂��tgA�:.F�N|:`:4�4ِy���b��*!�Y�<��{�h�����I�T��
�i��E�S��l9�6��Y20n%Pr'�{nl}�]���U�}�r�nS]�z���b]��:�D��������Q��5vw��l�A�ơ��J I"�7�N)�J�����?�[�ၚ��%h�Vt�ɖ=)�v�g�ǸeHJ��lb��?����딚��zG'�2JӜ�G!�L-YJ0��&v��H?_�ͺ;�`Mŵ�8F��QrV��$ �֖_S��9U+Gbfh���	�3F�ȕ�����ɩZ`A��s�Bv�N�Q�8}�QU�VU�k\1�l��	��L:{:���lK�T��ӹƣ��l����nG�w�'S4�ge��p�Ԙ	�,�5ꏔ�t�)�0*��ރ|��r��FkK��m�;��mwpjT4�t4��]��L>mX�A�u����?��~�����ҹ�_Ϟ�],F�l��/{W92�٥G Z u�Ro���o����)"�î�ݜ�lt�.�}fcd�ZG�[�K�CmtԵ�<NQ�n�*�]���	=t`�P�꛴�rE=,V�����ZÂ�'I�[�������`���9ԟL����M��`n� �v��ra�{�j�|1�1_	��kLg5��5����bv�c`W�DN�E�|��Ä��p��V6@a�׆�M�����8�1�-["]�5�;:�@0E� ���.2.��*-��M����K>��nW71S�f�\�> |��U1����7C:1�/�ya����y��;�L��g\������# 8*���Ͽ��O�i9�������=s��)��V�E3��\踾�S2=�������L�5��ղ7�Ÿ��fk��c�{}�Y��2���<װ�2]'檺�`KUx��
����h������?�	<�K���F�������a^ʶ�XP��P���|�W)�R�XT�V�v���V]�FU��}A�$��~p�裯8|����58��-M�g�������uM��bn������ڑ��l    IDATF�"J|逧����?�tV�JE�ZSͭmU)p�;ʴ[�4*�I�t��ߜ��g+���A�����?���_�B�+n�K����`0���d��rz��#}��;z�sߣ���J���Y�R���c)]���7KqC��
��@�����3&Z��d���+A -@ҿ�+�l0��9�z�.�q��7[=����3��y����JZ�rʔ�.Bto4p��؆���-�%��M|�&!�^ �}7��=���0bXL��~���;�&H:�``ƚ�1=������I�����1�9P��xQ����r!��^GRM��_��ō��OA��KW���GV�t��hc&r�,#W���6KI��T���]�h:s�JaoK��{.h��"�����y��lC���?fm�f4u����c�<�7!�m�ӳ��c��i<�|���=a��]oiq}�Yw���3s���~�".(�������7���h�1hD<�¡���c`n	$k��֒�3c8�l:�c���q@��8�nX�Q ���e|L(����N�ZȩY.��@~Usq+�r��&t'�$�$4�����B�w�ZR\Wv�@z�Ot~���`�.�\n�!ov<���;�2�U�PpJ��1���bŤ�r��ڃ�Ju�4j�Z��r6ԗ�+����&:�j:�����o����?���������<�p�?_����{W9��n��0�ֹH����7����t���<���ӗzys��:\��>��ƺ�\�w�M1s� 9+踈��r���l�s�Jg�\����Kzow_O�����g����u=c$I�r����{*�R*0A�J�	��[MK["�|o�6E|�l����ڄ9�bЏ�Ǥ�xs�!��j�yW� �˅#��+?�ո(_�e�l,ls2����()PIԠ��c;7��d�0���K<��P�
L&�cC�焦�c�A��v��Py���I½�X�RI�3�f���k�Ƨjݬ�~ת��rD�����[�� 8{
��J�������}�˘ ����g��
���֎���e4���鋗�^�h=�X�����Z�nW�����$7���VK�rm/��z>h<��Α�gջ�j6�c�@�� V
5�����pp'Uc����c ����F���+��Vn 9&M<�1Ai�
�ze=�b�DA�{t
}��������S���kCbd0��f8��hh�m4v�c�H\��(���̏�ժ�/�1)[zOV1p����մn5���5+u���x5ыލo/�g�Z�f��>{gg������3�' &tnÿ@q{ٽ�!�eC�xӢ;����Է�xG��ﹸ_��ӓC��44��W+���nE%����\���~Ҫ�5�BB���Y-U#iF��Z��X��T�s}���wp_�Zm˟� ]�\��������hn����VgW�J%H�,�N���w�7>ӨVT�x�Mr�kE|���B �JRX�� v��J
Z2f�q%`j�r#��IW�/r��E�%9�걐M�#� tfI������<G2�&l}^Gr��_���ⷵS�F�Z��	��4vt�`q<�_@��kA:�	|����ty���;;ʳ���tzu�'G���H%���Z�r�NRK�,��l��^@ОK�TV��sg(�/����5=x�P�vǣ)#1 P�U0qOGR7W�Z0��mo���\]���X�^�]ܬ7�0i���4����ļI����ӥ4�)�G���ҹ��d�Í�<�]��|�@���c�ό�yl��l�Mc�� *,�q����J��bZ��m�h��l�����j6�v�0�bI�R�m��Dn��|�$�dþ*5Вe*����R��ܘ�xc<��q���a�����X�UJ��˪�.U)U�u.V���r$�U*��j���f���B7����}=�:�l=W��|^�Z[�?������w�����:��l�ߝ�{?KqC��O-�s���]T7Y}����;��ή/��ٱNz�v��T�I�)��	7Ϡ�I",�hml���R�����s�W�&3en��]u�����w���������N|�F]�2����֞Z�m�<4{z�e�+,���}�U6j�^,`-��bθX����@����P��Ů�R����4t|�ڇ�#vmM"}#)R���(����tݠ=Ei�S$/�~�CGyVI��8��������L�����}k2ICφ��߅�i23&�g7��m�4��(�אׄi"��*͖N.�����=���(��Ъ�����Zj �L4�i��S8��ip~���S�&#����uv�T�j��,g֨�!ڹ"ʮl"�
��V��F��W:z8j&�Nf\�j>�����D~͔%c�����ȃL
���ʊ�
EJ6��x	}���U.��NGc����{i�
�M�n*��B�d��riOh��ڊ ��1�d�3�p�I٤�A5��� �/C��>&���Ɓ�������R4��MQ�~�.�I0���s�\�wqkTk~��"��-�ku��U�ke�y�汈�.7K���P/n�5[�U�e�*�fk�˷ۻ?�'~�5Y�ڳ����/_��?�t���ōu�f23���{o�?Փ�{������ͥI���(<fF�$E�i<�,�,���t���W&dR�36SԠ�..�*N�J]w��KUGs��h��ֶ�:���f�I���?PFӝ�=x����0��`4x�U46��ɘ��(�CM�x�$87��X��z}�dDD�tHN-�~���b"��T�X߸�=���9O"k��%J�d4E�̩o���yͯ����������!�x�y�&�󛍱3
�����Ύ�!3���Bm�fП�tj����J�m���������~�}o�N��,��ɬ���5˦5�nt��z����1w�lr�R%��zcO�I��W(��lwt��C8��7�IG�cU�l��BH����5��5#p����|� �E�%�D��TL��ύbu��./(T�Kc{�l5[�J����ت'���hhY�5���e��v���-��#��%�Ю&,�ت��Ce��B�5�T���*[�<�==�6��>�1o�����
to�[��w�+��o	Gk �JDu]\>�.<�K�[�Q�ĢzE�fE�zI�RQ���b���AWG�+�5�v)nO�[/�lm��?�S?�������ۻg��_����{�;u5X�ܞ�=� ��3zo�~��z��К7nH��*lĒ�����#���ѹ��6��,6�$�--��׃[]z�F�S
��S�ϯ4q������E=h4l?��l�La���0[.k�࡚�]�M��hn�Cwn�z�ap�4?����<��nGc�s�(�l�f�E��[.��ᱬ3�R����=,-��,���'�Q/��K��k-��K�/����)�ɲ�K�W2(�-�/�c�r�m�郅_|O�	�^���sP]0Q�2�#�Ya��tg�5�N�wp��i�qoV:[N4���^���A���R�rA�4��Aci��������Z�>���0�	v��w��B��T�� ��C����^:��*���;�9 �|ecz�pӺ7Rf8Ѫ7r"=KH�[��c��[p���z��X09�w�`S(Df����8
��j5z�N;o-,�S򙅭o��� �5CNi����\N\A(l��J��`G@$�is�-�|�/e�L�B ������^�!�R=A/��*��m�뀶2o��_D_����r��u��i��u�)5�I-u��{��B��	��X���:z�����������T���WT�������=�-���l���{����F��/�Ҥ����@?��;z��c�q-�e��Pɉ�/��s��e��4^�|rY�Mڔ�u�#]���ɱ.��*u�JsZA�=9���Z������u�6�z��ox�|����*S���h�Xj<�9��+���;8[����1V8S4��#_$�����H
P�o��q#|����8.��Hw(jh)l��S�3H�d��$�.~�}���2�*�@x��MC4��8%��0Ʒ0tG����t�`s���Ł�āģm�T������p���z�@b�x�0ª(�����r���@]���e��p�l���7���R%l�zC��c]�!��J�j���*;m+$�����U(+�0y,��[�� �@�	dcwX�N(v���e�%vG��,���-��w��י�8-�
�����3�'$<���ó���l�M��茭Q$P��9%rQ��=�-����b��&���vqmA=�^r� �V�Yc}	�F13�ď.oΩ�2H�fPB��0�A �.n���A��?ds���E.�A�sN.��;7����F�m��ۺXҬ^Ԧ�T��P7���z�/{W����zt�X,�U��?�;�����|'�����������?߹Z���t��F�Fq��EØ�-��/����y�T_��D��o���a^.� �gDp)0��	a|r1����R���PSߜ���K��\��WSj�P�;��g_h~t���0��t���O���k���㲂o6�~�ӵ:v�GO�&��*�u�2��-�� >��"vW��k�"T(6�67[��?�Se���G� �
�ы�+6�����B�+>�ŝN��pS�����{IA��%��p�Z%_��X��4���W� ؊Nq��Ԧ���Es��;�1d�G���/d��P=�Qe��ϼVŬ�thٴ� ���n�={�j4�g�)M�����/��h��ənN�4���q)ת�vZ�<<�y妔�.��l�c��q��ª
67��%利fd�x"�l��d��n�ZGZb�>���G\�S2j��0U�{�剢6�Y��^S�2NL��9�
�
K�H�t�k�4��&��mf�E-�$cuT�a����1��<��'zf��b��j2��'`
��@Dk�f�MG�h����Q�!Q.���&m#όm�J����m�q���j�a�:���6,��zE�v]g�>���G�ϴ̬�f��eQ]<����[����?���!\������>�l�������;�^��&���u I7�xX������<�� @i1�_�tc��� �So\�����8|��ֈ7��*��"��k��}�w�S��z������ҷC�+��].������R��<�X�YA�]p��r���(7lFwL4�Kiwxr0����6�[Ŭl2�V
@�al���΍��{4&���������w	7�3п�)���[�h��td��DRВ�3[_-l��	�W��е���\���x�����	��L�W�S� v�z�8����|V3���;���H���Y��C5B�y�tǛ���,ŀt������۞���CYf��P�����a��J�M��o;���`w��) ы`I��r������,��S�qAM4�,�bhIW���avN+�`X
��Z�v���bWb��k��RC��t��;�9���+4)��Ì�b�U	|-�W��W��S�\��x���򵢱�D[
�G�Yg��s����"�ko��x��|��􏉺�,����C�����(L�w���^����{��r��j�������FM�zY�뙾�]����6Q��R��tPk\>�t��{�_=��o}���8=�K���xy{YDh�-�Q$Q����A	A��F�{m��Ajn[jˮ 6cn)w��>k#�7��\��1Fq���V�Qr�������ˮ*��Z`e��;���_���}O�zCk����n,L0���a,�y�_�S�qf��Y���^W��(tM����F�i�:
��{l��Q��5L�>��oouqqf﯄�pВ�l�n\锂CE � ��p���d�`�H��ݛ�?jU������H���5�iB@�k�:#:���d!�Z���sH�8�1&�ᠡ�Q�y'*uW�:�5(���uC~Cj�ʇ�R�x����*d�<���-��g�}��/���`d�o�L����c:�c �/~́��ҹ���(�rQ���᪍f.v�Ñ�˩?_;Ҙ*���7,��roh20B�lp[�h"ާ��l�������j�iJ��=��3�&�|64e�1f��p���U��U/�\�y-[J�J^�r�!1Iqs�ÂhJ�H�՜��+��#쾗�&&���X�Џ"�1��&����v�!���]�S��أ3�"���To������ֶ��\��U��I����D��W����f��� ��h]����g^[q��}Թ�.�|6��7eS;�S� �%й�����O��Goy]Nh�秇vq��e�f�4xe�(���i�CL|��HK�2a��^�%-:��լ�{~�Ï>��gϔ�,���l�v�����?�o����?O��\�:(fr��^^��Mۛ��-�����o��ڧ�j��j�;>��╅���$:3(wY���=��Ҩ��$�h��%2.�W��牄�d�LT�٫]X��%�c�����k_��l�L��_R�X��"�U�Rqq�d�rw�PI����	�hS!�*_��������T�B�4:�g�k�,'�hU�?61��l��>P���щ~�{�����ڽwO��U�M�ջp m�9`��ۮ�h�+`G����ޗ4?{YD1������2�K�!D��1q t��[t��B����8�T�9`�tp`p��]e��#�|�1,��85'��m�����3ˮ*�%*� �jֵլ�ި(_�/p�L1g:� ϳqiK.�J�cvC�^1{�/�Ď��h��e���K����N�����<��%
��8���،�tr��
�����w����SikK�vM�RA/��?<~��z�%����ɛ{��{[����2��o/��/R���d��=���b5�%ǘA��9O�����׏������-U�}q�\��L�~��]�&[2&�;�m2=-j��`,0&��-��h�L��x�������O-vN���lC�E'�{o����}_O�~[y�+���~�-h4#L()M^��泰����m7#�H���8V�E��2tT�W+�H`i5p5�0r���J���J�		fFwh�-$�h�H����#� y��Dݤ�s�-�(��	��;�o4�L�IGI}��O�����5V��1��C�e:f��A�;M�.{p�TJ7}�W/5;�V��zI�\��|>��l��אd��_n�O�˰����=}��'�<;�뢓�wZ���S�QW�^����,>y�B���4 w�t��F��FM�̘�G^0��U���X�P����6K�$�
I�E#�28�еQ��7-����1���{�	���Nӯa~*�K�)U�� ��UԮ�`(�L�U�U6�-�3E!��#5c�
#j�)'hgIU�� ��r ���MOW�������y[��p�I�M��d-�Q�#��N���ƥ۪w��8�S��ֺ^Q�����Оn���2���I:�4x�����z�����Z���{��y9��٤���^V�I�F2ov�G�J��=pq{���UЧG_跟}��IO�RZ�R�Ft\��⚢�q���5��ؕ��m`��0��+��L���g��Ï4���f�g���o4��O����ꝷ���+�e ��}�q���N
�
''p&�k%2䖲H������ُB�`J�tN�������P����^Rm�zr:�񥢰:�D#J�Kp7~?�����$I#Od`����4)`�vo�ޫ�Ɗ��������dc��P�.�D�.2����6@��b��.3���KEq@n\2JŊ��nOǗ��ϗ*tZ�=�����~��P狉����X�[,�E�;Ś��[V��}}�ɧ���t�;?=�V�����6�luڦ������G�ܵǑ�s���r�h�iB�TQ]�2�(1Ju��zc�@��#�n{Zv�>�+dI�g�Z(A(�ټf( ï�WN69X.�m�pnf����2�2��bN5�9/� �Z��1���	Da�\�v��"�RȻ$b���7��x�;�E�� �c�4��    IDAT���ʤ���Q�8�-��7�Y{����*��J5���
�ͤt��t6���s�s�F��v��>y��������^Kq�_?���[�{6�����u�bе�^T��v��o�����޹�X�lA_>���>�ɴ�~I�`�1��-�R:0&H[�����A+�� �J[��Z��N?�\�~�Cm����NVf�?���O����Otppp7�����k�w�؍AFğ��#t�nW�� �-Q��8�moo����9�3�\j��[{�������<,\La���vwQ���Q��C"q���L�����e�n�dW�.�:D'&E7K�d,�
�'e1�ş�������p���N�+�c�c�h��@�i��b����e��=�ז�l��u��l��4�ZJ�l�s��9p�B����YK�V#]Ri�sdos�V�	�7痾��q��tT�5c���I&8�B6�e�+��\m6�l���q��LNE����.~��_�V��6�ㅖ�}��W��q����L��+�G	q I�J�`��m�A�dܣ��қ��U �B�&(.�*!mib*H���R�=�a�`��Wo>�UY�@�K[���v8v��{u��f1�k���=����%�8ԓJ��%y�lKk��-ձ��a[�j�̮\P?�	ҫ�D�ӑ^�^(U��j&�{������_�����[o�O���������?��F�d�����u�i6������>j�����zzp����#}v�R˱zi�[k�	�+d�<�(�-7�v8aA�.�?��U
%��ʺ��.?}�����!]�
�������ӧ���w���Ύ�Y����\�S��|��0��	"twM$_��hŖ(��|F���vvw]�z���Ł!�n -����ΎOt����s|�e5Aj�?�1o���K˘Ƅ0O���M�L��#'�P��X���y̤�s]�]��%�*��9������<�&K�N���.���1
���)\����c$�H�ܕZ`�sB��@����d�/-�F�=����hXH�6�Q/�Ҡ ��Y�
���Kn�V�{N�1$ܥ.^���\���!��
T��;8�����gG�{6�P ���t��v!�Ȧ�&���Ik�#�9qK/7gifC�6<�Pz4U~�R��t�!.d@P��b0�D��c|�/���ɇ�5A)��İ���F7��J\���l�j��q��0�<@��ۗBO�dk��,�L�
�s2�j֨6���R0� ��zc����#�o`fe��4�Mכ�Z�_�J��f$��2����#��by�.`�sqۯ��5�~�O��|�&����*n�������NF���tp۸�Ldy�t�ff����Vs�θt3K�.�:�hQ"jYH�$P�eNH\<l)PX���Ʉ�8�|�l�q�ⰻ��ku�U�婞���6�T�^p|󇾥�}��ڿw�r�$���e2a�*U*�:H�n]0�\G�zw�$��J����5Z-尿����6���/R�٠W�>ݬt���w���}�e�7k~Mv� >R)��� �r�o�rqF#Ov
�/H��0�X�Hh IK��$y<^a��(~e��~����rH����P(��^7V:5n�5���WW, 许б��:"��񁣾���s-W����V������ 2��!k!X-q��a)�c��ճ#�|`[�ɂ�6�ፆ��T)�`��G�0�,qg�d�W����w 6[w�-�,W�LC�&���ŭ�N+7[h~�Uj4Qi�Q��r���|�4{�>���V�p�r��s�����M�d�e���'Yta��gB�K!�R^K���RU����Z��>�N$�B��8v^�{��+j�Ӗv7�	
�� �=8�.c�����iTH{�y'��Xi:H�q��-���3ثow���4)���gu<����OϏLq<`!��j��qs�����o���{�#�\��������Ϝ�z��I��A�F�!����k���dzTn��WoX��Rޱp_�����K�x�h9���^a�����^(��/{�/g���-&���^Y�k)����f�.z:�͏4>�v�ս{��#?��z��wT�C0�j��+���dK'���:i����D����/2n���]����/4
r�V
ܵ~�4��� ȧ���`()V,k�$۱\-�����YJ�v�ؒ��qNqK
O�0m�����1�C�p�
��D�����h'��i	�`R���u�J�z�`�t��F2�ɽ���U�n|t��������鉾��-�y��U��[�~v�nz���.1ĕ�����$<�Їݻ��
mi�`�x�]���h��`�Pk{��ܑ6O,�Zt�����D�yP�E��.R�o���,��]�(;�'7WeMVjJ�ye��R��e<u0\C��ȯ\G��!��c�/��Q��Uŭ�ƞ�^��]B�x8�M��Es��j��̒�F���\��D�=�p�S�R� e���ب �_�P�a5�=�ڬ��\Y�z��tPL��4���-m�닧��C=޺F�)��E���G��_��{��������_U�~���������l:�#Gݛ6��Z�goO�]��ʖ����������3���T4�J]=�/�Tw�EsF�T��<�Im՛z��V=S0?�"6ã�\��T�Ӂ�N̧XZ�i�ګ��'�]*7_��������i��?��
ޕl��Q�L;��c�#u�7�uG	��/������f�����h81�vtt��SwM�hE�Q
�q�h��s�$f����O1*͛�u�Q
�eЦ��d�H��7j1�4��(&��d�}�2�HJ�+LQ�!��D�ղ t-Iq�s�!��Y�S�/��KF�����cz{�F��9�W{��R�n��ř�o�4$��]ӺQѤ�W//�JY[���6Z�mOn���q ��#�#u��J3����m��`[�jI�|�n9��/�	K����.����;��$�����_Bx�ղ�wq�{�&uJ���`�D痎��.Z���?,4�];��Z���.�u�;q�|
)��ݚzKo,�H�r�+�p}��ȼ,
���8����Ƙ�]�
ml�m���B?r(��c']�W�\A(l�z�|;�~��fp�:�n�4oT���烣gN��aQrPi��~�k�_�K?���R��I�����N&�����z��6Z�"7�g�����M��>Ճ�m��rI\m����М7V�ncWi�:z����F[�ٚ�f�8�V�h�����r��7�:�8Sw>4�:�~��Ŗv�%�F+��D�Y�Tv�7�0�2\L0ݓNd4�G|����qyy�8�*��A>$q���#�T$?����/���ёo��p`�Ð��7s�����P]��E�4�}�������y��}G;$㆐z#13)^�jƂȯ��-�����Tc8�,�Ϲ�[��mޓ▼t��a9�+X"%��ɜlǢ��l��?�xmй��3��l(W-;�_80Y�o��\]p݃���ԺY�4���[#Qp~�R&�J
�5��o�&ҿ������z��R�e|�_?����3�Yi�w��-�48����y(n\�n_��cۖo�l���U$��g�эy����YQ�����;1��@���,���PR�y��p�otm�D_�ˍ��P6�k+�7#Ɋ��;lK��D]J3�F���\Т�o3�=�:%x-�y�H)����FC�f��+e_���2����n��{���������!�\}jA{���q���<�����tn��g�ɤ���'�?qԻݹ�������(���s��}���������b',no�tL�F��zc�l�i+6�Nf���J�����pt��Wg~��QO�vM�rE��ިoiGe��ym�Zfx�Z�
ax��!���P.�<c'c	���7�&��n�[������8k{��@���>��s�v��7���"x�S>D
_�$���"�P?���J�ם�̿�$r��y���Z�L-)��"!�N�.0�~�Z��^�x%<Bw^_�B'����Cka]���wˌp$�b`��LG����(Ij*U|�����U�������JG����O�|���w5�t<��z=��;bD��}B�����A�Y'�^���L�[wb����ڻ��S��Fl�����k� g���h6"������!e�d���irq��x��V
���p�y�4�Q��� �װ�ʓR�`W�ɒ�`�C"��#z��|�bF��Q-�	�R���B�X'2(�_E6�!��l8�2üJ���h27�c<��;�d�r�s�[\�m�{�7aDu��+.Ҏd� ܄N��2�b|1��O�RS��R��вY׹fz1욢3����n�z�����_{��_{]��Uj�G�'�?y���]L{vgl3�(a��X��/���o��5���>__�{�%Ņq�~}[Oh��QUy�gc�i��tZ���fC�TF7끎n.���ݞ��,�U.k/S֣rK����o��v��3�
Ix�O7����m$���jc|����b\D.1��V���y!W��l��p����|yd.+�V��L������,��s�8$��o�8V�k��#�ω��)�B�)v�ȅ�(���y��7��$��XD|.)��P��r�H�L刅#,@��ՉY�`�V�1/ ��+R/nڤ({\�}�ƛ���I-����M�;�@��F7ݾ��=���	�kP��:5� ��0O�B���0r%����?~f�gP2gW�==� �������Mj"��ǁ3H��| ���ƞ������M��$��y]�t�LU��TZn�r�M���8�yȾD�1��v#�AO�cg�,�vݡ4t��v��VB����N�j�?7�/є�����mW�΍�/�����2���\�R.���A�p��h6�AD<� [��̖d���k�t�`� �2!�|���x�,�eh8�Dj����-�M����Uwn���5U��
����f��}���lK��=��N�����p>����� ����4'E�|���SՋu]�ouһ�gG���$�um�*zP�����,�|2]�������w�մ������ŪH?=�>�g'����L�:'^Y�ي���_lj�X�������F'�b4��7�':��0hV����d3�jm��֬�BH4[!I7�]�<��.���&L(�S�͍&][�j5��%cb���c�e�Mtqa�x�H�m~��!q��[ut�H6m���V2�&E3����\���3죏�R�ڂ�67+�ƌ����`���7v�����Q@:�7��� 1�6��b��Ⱦ|��yҳb���(�m�6N��f6�N�yͪy�8F���"�N��β��<��
�{�K���]_^���\�r9l��U�UN�]�,��(���E�)��N���y��@M��ܵ�+ՕV-��r��8�<�-'6�t�&��{�EB�@��3���M�|�V��T)�Li�)l5��_�1���V�@_�����_���l�$�G\��fs;�4�,tqE��L��D���ս�X���9
���X\�'�1�v�>�G\����-��l����b��L��y����X��7�����/��^�~�����o�=��Mz����C���/���o�c-�!�bv�Wq��R���~G_{�m�r%wk�/O�ԟ�_+�U�T՛���ߛ��x��G:���E��.��oכz�w��֎G͓ޅ���lp�t��dkSнbCo�v�_iɆ�(�؂�
�f�\�C�����u�_\[�\��]��kkkG�;�N��������ű>��S�����^t<7=�Uz7��W�[�S���q�HK��0O,r�� �ޝ\�O�����+�J������_uTu�n��'ʳ�	DL,8���+�!���P݂]�}�Mi���(����hOH�8$}\'zX�~�4�������þ��ך,&vW�8�y�b�<E�X*�M�-KN�]Sz�-ujYT˚D����Zr�ڎ�#�	!̮S�e��tu{y��/_
S��v�v�i�o7�*�Ѕ�*�O��Q���>���+n`�
͵��OTFK����vUWJ�UZY��p���J�.Q4*eg�X^�(��ǜ�I��|0�Z���̻Q`�E[��hh�Y�V� ������Jhzc�# &sL� j��а�*厎�6�R�7ֈ�h8U�������1����]��]�#W�:3�(����K{���쨰���v88ڏ�F�;�{�\�~�q���o?}�W_d�٤~��s'��u9�?`�\!)|г���jm}��z��[*�����C^����Ʋ����zw�������(���g��q��T��FGo?zCD]��������vM�RQ����5��.�]���@;�÷D�x�A��!�BZ䋳s�|���#6� ���ڍ�	�bYy8{|�7��胏���%"`|�4r�Y��;{n>d��|�Q*Y�Sd`޳�� =E#qqg�
��U*]Q���j��d�M4�t��t�
\N��~�qp���Gx,��n������
y��Q�pǻK�􊭦�$J����X�1���`ID2�M	`�� *wXu&��I_�jQ�VY6��ZԊʴ���Z��RNW�&􍆹&�B<�
Ǽ;9Ҩp��>�P��J����+��ν]���q%��3�ǘ>;h8!~���$�r�2���rE��zo��6�=-�z�^�3嵌no���U�CJǖ;؏���-�Yb�:v!��ou�WD�0�oT��m� �U�N��B�+��W%8B��e3�t�,��6E�EN,��ڮ 䂀���0Y����p:3�D�c�0f���1�� �����xX�d}	nK����w봕uni]�˹��s��/����J�������'��_���������A����?t>���t���9Ql���v���.n�x�-����*eK:�k;?����	�x��C}}���-u6�����^�6u5����k����������L�חjn�ԩ5���t��V��z��5{( �d|����`�l!�4�1��'���8�s���%�xN�D`\!t����V�/]�e���A���y����XY���&PF�D�%
�UJ�Z��)����`����\��[�L:E�/���BĝY����E�Ɣ��m5�O��,��`n��.�}�~��>)`�N^��"���3qݏ��p9���l9�p>��#NqC2�g�K:����ۤ��]�ϵ�����(f5���s�M��{ ^!�2�d���F���,E� �L���5�DP0L6+[�$&�YT���ܝ���\�TA�lAovv�����j����Z��z@?�FǶ�.n]�����c�	 ��e	4@&M
@�.�Q��W%O��[���Z5X�'�kV�0:	э��sc:��M'K0��p��:��g焳�]pLR�(\ȥx���[�H����p^[u�_1a��Zבat4[~u4�x�ӊ~hF.nolu~�����_��7~�|2���t��!�,O�q;{���7�zG_�������gzvq��>. ��O��˺������^�\�EP���H��O:�z���B.k?���c]^_��n������V���r�\��l�X���?��R'b.���Cu��5��Tr��s!T�5mmm����ay��P�}��P���[��9j� ��EA�CoaD4X�
(�I�ȟ'r�d�c�t�p��\0�aH�2^���<����$���A$'�J	6�=[�+>�G^��M���sb�!K:R(%.��O�\��+���"ctpV��q�15���JW7��Jz��ͫ^����q����0��.t�Kk\ʪ|o[�-��Es)-K9M��(�өo���q����6r����c�O/5%dh�V�QSc���N+���}!5D5=V12X.�.�7<�������Rñ����
%e�ý�k|�� _
�-V�K������T
o%)p�_��F@�6�`Zɵ�IdVV%�N(��֮B!�+�Dp;��Yz��`�0	��ʄ���    IDAT�
*�� �r������ [��k;�ch �Y�q8j���]��`��s������	���u<�h�Ӧ "������v���~�o������?�C���;���c��c�d�$��Zڮ���O�ѷ�{_�tIW�=?;����8^�����z�H�U���^t�����M���n @�ǥ�����t�������K�u�w:�&}��Uӗ0��Ѕ$`�Y���[~�r�5Gӑ>��ͧ!Aޜ�(�bM�:͖G).���}��'����ܶ�<��[���&
]B����N�[�դ��+�|�W�T�p���QCC�b#�����|H�ӄ8;CF+�r�q��L6��o��P,-�>5)�Sr1_���D'�?�u��^=�?�荆�:Q2��F�J2r���ե.�/D6j����ٜ�>���K�u���ӓ�D�J^�ݶ�vmQ��(�[�`�l~��6mj���ar����R��KM�nMf���j���mO8�8�ߡɍ�'�'t��z6k�ک�eB�m��H���������s�\�h��c#��ϝ�F����~0�'�ӂ��c),&( ��R��® A~���FvA6e���k޹���QXO%v�l�і����Z�x�	��%M&��\
�X�!�<
(�h�E,�"M�
�q��ܸ)p���jEi�>:-[usi��Mt8�鋫sͳa��o�~��}����|}��}���ݳa��N��'��e+v/����R�����7��
�(T4�Muty�����=s\ܻ�{�{���V8|vu�_~L	7!���-���X��Σ��n��� G���H�~O����mݫuT����n2/@��[�/��V�j
�3ONO]l�)��ku�+����y�ŲG�g������q��ݱ�<`ٔ�`���������������ǘ[�B�h6#/�c���r�_&��to�L�*�E.Q�X�n/bx��J<��o"�O�E:7~@E�"#ʯ?.���X�$#h� 1�]\���¿cLj�0r@��{kD�W��6��y�����^p��F�Fٌz빋��z�T����]���jY�k�������/��ϸn�s��I�k��.���?���~�&�>Ák�l)SB�\1`��=O�W&/��!d�"��̕�TYnTZ�l��tŔ3Y�Y�I��`b�zm�A� ��R��C��lP22��K�������[!�*9
tS�WD��Y�a�~Lt���̽��	u�U*�Nm��"{��T,lA����֋��"9u�j��,RX,d�^�X[��nH�K����Jm��j�t��[[�Y%�R/�������7���ײP�����Ϝz��Q�����H�	�G� �r%}��[��w��f�j<knNf�� ����Һ]���ő>:yxs���W�BE����Zz���J���zj7\4�\P[Œ�I��5UBFmRe��������\&\:^�L4��� �;�����5�m�Tno���}���Ӌs�i�DU���8�Q2&kp3�k� ��D*��.zQC�����Q/(���O����ȷb�㒷^�st{\J�me�-M����<*
f*�"�.ql�����Yx�r�P�(TIg��P$M)!�/�H�2��� 2�,rmE��h0T�wk�����`��x��� `;�Ԩ���bb�ԺVT�7<�����=sc�D:Ǻ�=6�m�i"i�o����i|��ʅ'�t�f]�z�txp�c[�uʃ���VN�V&��K��>�5�Ψ�ߐ<E�.ט���	Zah+�B������ �l.����fГ��*�[>�
Z]�5^t/�s�������#<O(�tmx�7r��2B��є�҂z��!�ti�sH�2�I�63f���DR˱~%uu��0�T��3������֦�Pj����ʮ ��"(�M�#ݩ�{�������,n���o����w�.#d>�ϧ4�m%˯�q��~��wlM�.f�9`U:��O��z��O���W8�R3S�v���������Z�(�٤Ɵ_]Z�D�q���n���JC%��%���r*��,���|���]�����j�R�������b��be�7~�Y�5�M��4�� ���2,-^-l�(<'��wQ��t`,)ҩ�K1�>���F¸�kyU��1ۤL���p����Sch�"J�B^u�M�.��،�ѡ"Y2����1��[D�J
���a�Qn����	ō�J�|�D�%㷥N��hҽ�������B�Q������@�|F�RN��]bI��y��j���45ɧ4!u�0o�� }C�y��Xa��8ʂM�U��oo8�S��6��r!8��8�f��݌��%�fq{å����Mם":U������㑱/˪Џ"�*�Ł�ӵ0��k������rB0K��3�������C�!ۉ:��&��#��K�dJ79��	�+SF(flK�P�"��1Y������uNݴ�H�@9��Âz��Ǔ{��L������.R{��Ɨ�i��;]ה�Z����֟}���dyě���wN���E����㾉�����$ c�Q3���v8�ꍝ����E�(s���p5����>��|6��}6�ڈr�T׻����u�I����f��Ǉ��*�����ÁQ���"!;{L��!#7*�2�`e��_�\k�Bt����ԏ�ֶo��vG�j� 4��>�P���ߺ�Ar�Q��:1Z�E�{�2$rٸy�0� �z˩Z��K+Hw��ţ���0So�-�A�0M�1�X>�����Մ{����(9���p��$E�]&�tx�;z��6
<�}�T�6v涱x��ű�x�>������Z)V	�8)h�2#�ɛfA����ω"g��@�B�ωi��涧��Z^��o��_ε��C/�;�;5��5��C��I�Tİ�s�	j�`�B��l�X>�D����g�.���/{8#�΍���8��0_�����Ԁ�ҙ�ۻ�jԔY�տ�	�;�r�k+�Y��lh����"���]�j!e|P�o���1�t�f)�ؘ"�r����eJ�f���)v��ٴr��J����l�.�� /�U�a�W
p:ez�BX.���_�US��b�/ju�kU���U&倠����'֢��Uk׏�;�'�����y�;�(��>����dy��7���9�����I���ӁW�"XN�(YY��_�����4����}ߗ�׭�����d�B`P"�	J,�$2QP��(Dٔ����xc1�e<��Q"G����鞞����Z�sϾ����<ϭ2Q4�sZ��:���9���<����R�6v�p�Ne2�d��x���zԷ'�g�Q��rp��r����S�+��:6�u�wӲ�h$}��m+_�jl��Z�'Kf26;8���N����XQ��ɠveɨ�V
E���67HH�W� ����O}&0D,>9wc�����>cIg\0��5X����V$]��Ӗ:5}�_��g$D_�Zn<O����~�	��^�7YS�(�G�247��@�#k�kM?i�Sʠ�������4�H�t2���a���3u�:�%�&�TT�`��xj3t� `���M��?Pp#��D~�i{�ݩ�l{���fncۘ�SQ�mTm���,���v�v^{h�zI|dR@��lZdpd~8�S�� #�
�j����]v;�B9c�T��0'���7�:>�b:���i⓰���۷j!(�F�����n��N�b�a�F��LY
��M	�i��W�7a� �Br-b|FA�����+V��sJ����YKf����D��5�����ʍWSF&��no`����S'$���7˼��6��2�:#��\��w������v���	�J��躕˖*U-U�����nZ?�g�����c�/pn�J�+7w���������sᖲ@������y���'��C����ዩ�(�R�؇��=h��v���4�@2.�3Y
����s�.jɨH�x0�#)�Wݲ�BY6�u�\��5��HL� ��ۖ\Ω��WAd0���'GjD�����E<��	��\(X�RB�� pqv�����;Η�w���V<P��^��,nT� �q�\+?��(�F27��z�UQ�2imlAO�� ƽ�/841"�O���`�Pv==2Ѵ��#�}��V $�3��m$��� RD����P�������Y�>+��F!�:Z��-4��3*�s<P�zx��^))��6�T��۱!�$,U���n�0�nl�J��|b��Y�Y����������2��揉_,���{��21\ s�_t�wݨݷ�uK��Z�&��*Ns�9S�G�u�n2!�0�wK�e�"\F����S���D�y4TP!��P��,�g�j�0C����+�P��4��d���Y�\�ݭ�~��{!M�#���1~��i�A[9�ͅ�S¤�I�
�����0VfKk��r������|as�T�½��ʹ��J
q��%u�P8ᾎN>˕r��Vq�<6;;�l6��سN����O�3X��XE��*�Νj��=[o������|2�o��[_��v�y6��lҗz)�(z%�\�x�U�2��d�0v@��E��9�`���-m��ˁ�M6��f2g��B�m3u��A�m�d�Uc��ʶ���>}�T�fЁ|��$Q�ղ�nGVb8\s���8�{sJq�"ΆD�nc��f5��>�&��%�2��ra�����¦fJE&��e�W�����Y���Ea����<��M�����r���X��W����W�4}p���w=��E�X7�*	n���[\�(����Q=�TJ�O�V����%p/J̾4��!j�Y�n,L{�C T=�pa#�����9X�6;?�
.*㶵u`d��\�b֏��E�eW��Y>m5��v,Y)ؚM�K���T9?�dt�`���)���/��ou��;=k]^Y��R��8hax��������rt2���/�U��+�-�B�l�� Ѐ�8�� ��̉\F�M9�� �u���8��IQ��RߪU�R̫���� w�"�`&��y7��� ޥlȌ�ED�m8YX��W���l@o�S�y��B�|���E��S��e���cM�0���eMY$W�����[)��b>����ɑ�l.�����Z{�\��~h��k�[Y�7���_<���y2��0����(���|��޷�틇��-(0��>��^[k!����$8�雌h�@fDZ_Kfm+[҄i3��x2��zi�2���h��֎�y��t�٤��N[��)(k����K���l��Д�l��D���c�o������W�j�8�$���i�Ԯ����R?*��@��'/{h��J�0Y�V	����L��E�L����}m|�P��EWf��J��ZCώ�@��A2�٠���1d� ��vvd���u�p}�?����h�d\E���g�`�C�V\�]: ��=E>�2>LH '�R]�'��X	ٌzm8�u�����&��Rي[u��4-Q�Y�\��&���� �1ML靑�ჀrG�)YV2-	����}��c���.�J�H =<&��d#�z.o�v�l��۪�w���F
&�ʅ%��Y}8�2�d�3��`r8�_'�3�7N��;#�Y&���{!��d�R	(MBJTO�b�2٬Z��M���՜ �Z%��Q������<.�g���Z�L�d�D��|^	U?���K�M�g���L�U*c�J�"���b1{1��k��׶��$D�JF�Y,_�)W���9���?��G~�b�s{��.�o�w����g��J�0���x��썭}��݇���+Z��:����3á���+�C�A�X#zzSѕNS�>5za�,���#-�҈����]�AL�Z5���Ɩ�����N�eن�X*����s��i�n��=Fؖr���]����B:::������p1� Ǎ�-g.��Cp�W�[P�ı\�ޖxv�D��l<��	48>*� �?��󿔉y��Y3�A)G0`S��-<I���4�����pL�9vo�	�aHA0�Z�"����mepH��`C�kt�� oN��SU1+|��)`n �	nj�{1�cm��LA� ɿ�P���$?�L�I����A�`��弱.?=?��C��ֶ��坦���C����Q���b2��Q4�Ԑ)Z��i���Nߎ?�u�-7�@L�RE\��S�N�z�wG�g��@���w3����,M���
C/!�Zs�%�a9�ش?�!>��W:H.�1�P��֖���~2�)AN�N/N���~����g*U�o0�A<�	9{6j+a��¹q� ρe������$��*�F�������^:��*�/[�X�E*i��ʞ��v:�K�r	�`��kJW����_|�k��W��ȿ��w<P��o���'�������T8w|�� �����r��^�:�3Dwܯ���.;������`=��㫠RL�sqD��L<aL�91gk�r�F��ի5ȄX��W��Ռ����M��f�n�8�]�����{��#�
�����������L5 -:��!}Ʊr�.�߼�$��-��+$�mOm�T\�@�Y��R��O3.,ж@Q�}�]S�

V�"��zo��2���[��J��M��z�Y����L Β�Z�R�&�%m��V(C.�NC��-�:!��`%t�7�	eo�7�s̅��T�+U�d�ָdm��*u�c�r�������
��ked�|����m��*�!H)cp�����;\̧�\�OPA .IiJF�}pݵ��u�Z�'F�PB�:����52���V �S����` h�T|��]7�֯W߃w.�pf�`GP�`��tc'֜ӨB����CB��n�3�g��u�&:pŦq����0�R�������j!�"�߶���>\�/��nJJ�[����gN[��2Zne˗���[,�*��a,jgө����I�¦�V�I��Q*]=����#_����?EP��ޏ�qp��{x>�������<t������-�Ca�~�/ڗ��ai[�����>�8�S��l�p:��OE��9����~��2&�3'��\6��BĬ8YYe����,=]�j4��vlӘ,�8OOυu������ �?5�K�s�������7������5��Jx8�Ar#��4�S����&����K>�J@�>S�D������D��(�F-X�M��ƢTs����||�������W� �%.s
���)AC�[�s�ET�(F��v87]{.����?��j�)�C�H���@�!�����&�D�ގ2�xRSm���9O�����t���t��LFmH�Q���vB6i����;-;���n��&y2���V�v���ۤ֞�l�,���'�����D�07ܯЂ#`�n�/����&��t��~.�VS�a��gҨ�t��t����wa��H���b�'�h�**9=m�����
,Zb8_�Ĭ�^v�`ހy��#aT/$��/!ɻT)�����:�/M�y��T� �ޗ�p��|a�
��*�ד⇞��g:�>�&�U����ɣm�A
��筛���|l����j���&��f�r�hw�O��_�c'��3�>88�����A����c"1sR%�6k�����{���Ν{�[j����{f�/��Űm��X��q<�����gr���E�e���s�'�R�PI��Z.���ba��¶#);�嬴�۴�Q�+v����J��Ϗu��˫�kg <q�n��D
������
pdP�>z��@��K���( �.�d�E���#���3&���w4�ہ�?܄�B�Q�|^����,N^��A$��[��?��|TC�Wq٘�W�Ρ���`�%��,��q%�+eC?���/�����sLO$Ž�H��g�|6�`S	Ǽ`��#7%E�F>A�ҋ�L���^�un?o2*��M�`�zA�-Z/�*��k���;���A:UL��G�t��b����Ώ�����_=G0eж��%2�b�>��x����f`��XA����=m%�rф�2��    IDATE�lNmvӱEo x���dl�9���OU�8<Z���u�(I���zr�mlVn��̸�A�-�+��S������P
�$�$�$9+GsT+o3�;ŧ��� �J��t"�����']?����\
��-S�$��R��ժM�C;�gǆ^d>�Mdi�R�����^��?�w>���o?~o����g�ֿu>��;�;A�l�S�Z�~��/)s�+7�����=�<�O�Nm]ix@Yz��o�jVʔ�3���Ҟ��(ZS*��s���mD��-�V��mk�{ي��Ul�Z*�1�Ҕ^7���T}�H4�$]nBH��*�4m%˒�j,mo���Q�R�~�����ٙz>�F*��XF��Sݫ�B��	��T���Ŧlϋ<�s�W`���ml>�-�k�j����F��ŦN����-h{57l�^�;,���o���y���W*>kp��`�V,޾?����{:BE�&�k�K�p)�8A� Ep��у���E T��q(��e� t��*Gc	w}}7��`���xdn���Ewj�\�36�G��B5��Lk4�D$n����wI���1=��	������O]/��"������LC���6�jۨձ�hl�t�*���bq����;=����E�b� *��P`������<M���A���=5¡�^�"�����gРl�;�		�M�]L3ɮb.x��J֩���e���������t��S�x�V//dz	z���%�ί�{l��%-���k�H�i�"��m��V�����G�v�k�p1�h"j�R�ug��_��?����E��D�~�3����wwO�_x�k���i?��E��B:V?��;����+�ܕt�n_��i�l�1��;[����VJ��f6�������qd)uI��6���,;_Xy���h�^+6�n�!h�U�Ʌ\�����~	�v��IY ˍ6	'/���E�
lp^�^�=9?sY��i�66��Ғ̍2���Gh���PI E�֌�5���5��A��%S9z�BA�Gld`;&z�4���K��/8�H�pm77�Kޫ~���2Q�E�
A�N���ß�9� !��F� ��,�������+��j ��6��ե=?>���S�9�iO���ݗf���&��-��fŢ[e[2��4����Z���3T9%�mig[�4�E{Ӂܯ���B�FS���5�Ɯ�0˝b.�����HԷ�����b2i�D�
@K�Au�6���b0tަ0衑7�	����}.F�7:��{8h9:�i �JγF^������̷�`^Pr��:���M^��E(T��r�808�������^�r4���)���y���H�E���L$��H'�g����2fɴ-�s�l�f�֥�}|uj'����}K�c�U-��i4������?~�ѣ�gZ��k�b����֏�O��q��A� ���V�=�w��ڝ�΄�q��?��g�6KFlIp[����{{�d�ړ�]�;���X����H�@ NF-Kv6�[a���d�^�n۽r����Ŵ����ܮ�a�~ry���C��&�{���0�eJZ(�ɓ'��.<#!d\�J��˾`EGXt�&5i������G@�,HD�MO�($�����R�Њ fU`�p �94CC���tb�!{
��@���9G�"$�C�r���=O��2�Ϝ�/ב�n�R����֕�������S�K��\*P�%U�ִ���n'g�������]���V@ �����ỚJ�,��鲒��NEr��T���G66Mկ�]˜����X�[mwK���r*��R�$����>�}��=3�v�tI�Nm��X�������WL$�Li�L+��5���|4�,�ܫ�*WZ�r��ʩiHM�ݴt�?`4���;��s#_�^>�T�Q���ڧs�����˗�8�(��8�����
)���]>�b���p$vˢ�J�g� ����*K�ڊ[�	n
l ��E�[&Cpk�U
���Ԟ�/���$l�V�����������7��O�_L������^��I�g���b�?�M��?���}p����$Qt3�iZ����mjn6���C���-I�堭�/���$��El-�~�������}�wD�"s㴄H���g���'�Y�.�ɉ���hø^��./.��T�&b:�ܻ�,�Ӈ))�!�UФ��=(q�����u�,��a���8��'�O�/�\�98�dn�z3�P�9��T��0]�6�[��e����'8�RE��I\p �X�Δ�r���C��w�2b�q�-�tW��f�6�uht�|�O�1d��\*[6��T6�qW�kk���a���١�9�=��_2|[3)�%�։,l�v�n��Ld&���/�U��yK}0|䈕J˴$��E.�R�v��C {�I5��9.��3A(��!a4����n�.m9��u���iej��-�	�x(#��)E��+*��\i� �[�\`*ԫB	\�˃�=�{T.�u���)��WbF���k	�/[A������j�u���E�3����.��b1q[��6�HXaȞ�(����
E��R��G�'vҹ��T*�z��٭T�ܗj�����W�߫$����R���x���F�?v9r�� �S��[4m_���
w�{�����=�:���6�Om��@$jo?|ݾt�5�ǲv5h����=~�\n���Z K�2.�Yz���%�~�n��l�\�
�m�+vrt"�U�Z���	�P�����7��k��dtϦ��F�4�L��Ө�b�T�7�)B0P�a�t�� ���j�)Љ�#GX��2
@��X�e�t&^���Y�%o��k��C&#d}�+���kP�x-���J@�g(C�=�t]�_���e^@+�	��hԭ�l*P�g2z�XrpU�`��^������j����~8T`�W����r�)S~"�5N��8��>��A���u�-��h���~���d�rI������Z|�a��m[T�ց���x&�r�H�i#U�b<e�O��u��ViT�P�2��P,��8=�%�N�{�g"@���̦2�a]�dКJ���A��/�!���´9̣�9r���1׫|���ޙI��0��)*c��J�%��{���T�����\�@租��<u*JT����Ap���\
L�/��d*��F�rE��߳Q�F+VЕ*�䢆	�xn2�5o�L�"��-�y[����ՙl��a�*�w+���ˍ��_pe�~�G/���N('-N�ˍzn���M����,��倅���|�o޷��}+$2֚�}mO	��8���T�1��SpmS�%����m���P?##���g��]j�K�����$���,(�����l�F�n_�җ���ߟ�8��pF�d���u# �,0�� 6�w�
婀�c��t&��zC��l6���Y��d)d{dq,�S�p�'�1�:Yq���dN�FCY(?#[�%h=6*�!]`��kJ0Q%�Z׳����-(�p]d_Loy�)����t恚y�ˢ]��J&d�g}#���|��3��!�#s�����ե4��1U�N��/�R�ar�x߫Y�ޞ-�$"bm	������1k����ĬzeOb��k+�*�تk�Ջ%��201�#A@0qa�l�>Pq.�wٿu}m�vO0o�!���Z�:�5�}EV �)S܅lG@^����2���0�N^⧝r�b:�Wc��*�F٩Jx��������|L�e����y8qs�wK�q�(��W��-��Y�Z�c�#� 7XD�(��^����hlY!_�������u�e�6�n죓#�v�/�g�^,�6�?�}_|�7?7�J
'��_yֿ�w.���<b�nӥ��q��G_�w����nlgг�jj������JͶr%KŒ6�N���
�KSW=7�U�.qJ�Ƕ������a�nw����/�x8P��A��̛!C|���4����EHp����-������Cׯ����:a���T���L� 0B�C��1xZԊ�i��?�	�� #������P�����0�$������̕�Ng���������xq*F �k��g�,`q������=�����O�/4�Ĳ�Mv]f�g)�ᡌ�9$�5g6W ����Ж㑂e�2�)z~N而H��΍�[��i��t2 T������XF"�_�l���f�dv�m�Fή���V�I&<�	�7��Zr����S;}v$�GTw�w��`wϚ(0��N6n�H���]�7Y	�.%`Z�gݞ�kf>u
)��$H����X�
P�e@����!��� *��|�ҕ�xCޗ���d�n=M��t{��a p�i� 
���� �q7�z�O	P���Ry�[(W^S��?�eq=�;mNdCe	,+
`�J��+֛�u�Um����bf<bW�����G�Q,��j?��[o��?��/�	��x���R2�����[
n��j�ӛ�-��ڿ��M{��C;��6P<��L�}S�� D�(�.-�ƺ����w���p��4v	�1zݾM�o,1[X#�mUda5�A��Rv|tbg/N��%�������l�7����f�j�Z�n�dE,`~��M�zX��`�H�zD`����j±�N� 	�ґwٍ(�Q�o�Y_Uv��	 <�(���FH��L��R�g�T�iR;���I<������� ��-��ŋv���>$z^�qTc�R���4X�����5tzm{��ȎON�g�
���w�	C�Sؔ�;��O��p�Ab"�9��T�sܗn��h�\�'���]�[����π�D,��H"i���Ʃ�-�9[�Tm\�۠��NteK�Zә!���o���Z�=���S���| )�v����tG�m\�,�����2?1�����P� rM]7�	ĔmXJ��#�y�<��$�2����~z���R�g��@���%$�i��h~��a�������)�L�cC�Wի��R�[ghc���T�ك� 	S0�[��O�dX��9��_E1�O[<��J�V@͚�ָϬX��fi�[o>�(Z���U��~��?ߝ�_����W]�w;������u��h��#��8����)`�Z"oo޷w�n���s��ϻ��j��#L���s�����*����ق��jKFf�RXӔ����XL9;7�����)���ڧ/����BZh`���6��%����(�I�~c1�Ak��*�L��g����Aa�C��SaB�
dr~N�c�Vdqd���L�Y��|1� W�P�ך~�}���ٱl6��Wvqq�@F��)LwC���ޅCZ���C�%�c�������������Y�B=�ة�B͉[�����B�ٺn�,�g3�8��3��%LJ��Ю�/����i�aj�L9A�����(�E1m��M�9k��6��lI�Ak0n5KZv���uߞ|�}K̖V�'��������m�k6�4`�	Ԩ��z1���[⩛r���k�\u� ���٥* ����P\W�1�QɊ3X̩�Y[��7��O�����T��k}�DҐ s��#� �OBU�z)�p���u��~��.�T("�a ��l%_�2Le~���{Qma^����WX���E�/M�)��lZ�`�2�[2 ��%V���zO�{�����ݭ��<����
l���E���s���{{G��7N7����+���r�N�����}��vj�W(��K)x�i�;m@e;�@E�G���g���l�;}�F���x�"��4�a>�ۧ�?�^�	K5�>R�����h
��F���հ��ݤ��y h�C�<�7��M�Z-7�L'��s�� \բƪ�/@�|��'�O��t��zi����J�^Oٍ�>"�L/C�zk5g�Kkb������B���w�VF��s�:h\��`�b^A�V���u$3�=���K����v<re�+S>iZ�7=$l�zCφ�>�n\y��&��Yz�6�67C���n��$��p�G>'0�b�֙���Ӷn�m\I[�����+]���IZ�R��,����O-6�H:�+o�i�4Áj�ZX-$��*M������s���i�OA�'�Q�{6t����(ŏO^X�۵�V[�A����%o���Q���Y&8A~�i'{$���?����,o{r�Ӕ���� _�/�[TJ�EC�C�p�~M8\�2=@�7��]N��_�	�DNId��$�45d�S��+%ySd�In�e3ME�M���H9Q��r�����Ӈ��o|n��>�'���7N��i-Ƒ��~MT�W�~2�5�U��ܶj���F��w�|p���ρۑ�lā��47i���B��ئ;��j#g���m�8���da(7?��6��(*զ�j�SpO�v}y�`���W�@��w����`&<��6��$�VR�p�o�6�A�Jwt&��Τ-,$2T����\斛Ҷ�rN9�ѯ��Lo�pa�J ����n:A�R��g?��qQ]�ǵqݠ�]��	��#P������������gx�L���[9�&=A4�5=�'tm���N�����`��;�'�'|����87�g47���F��n]����Q�&0n�9HȢ��u�d�jں���QC(Gmf��*n�������i�,�2z���6	k �zG�[{vq|b���;z��M��jV�n�9Nv�Z��s����x�����s;����S�`���0��#�O��*�|>�6A�|��@�j��TX��|��$s�U��.�0��m������$��eb�� �K�sCG�ww=n��z���ɾ��%P�a��RknY�Z�\�b�R֬P�5#.x������Bix�����{ۿ��Kp�Z�"����E�0�Yln��ԋe'/N�D��Mk���&�N �HU�ZY7-C5U�xl[�=�n�w�j��8�%x����>��RJ�bV�m);��J��Ln��n)��;]7$���;�w�i��z����G>_G��qC�,�ƽw��N���,e)7UYf����r
`281TR:���T��L^���h\�tB�M�"�qw0��dl7��;u}D�0 H����ce	x?��w�
lP��l�20�W�Dx�J�Z�9<xR�
��5
{FII-��>�Mݤ��?��\�}����R:4���E�[f��.elQ�۠��n>a�LD��2j����7K&vP��!ex�b�Ѹ�	�_�p��={�D���L�M��=�F��npL��4���J��׷����~1��E�wH�;lG���	U1�_e��fl���6���{
�W�U�"�:���&J�Jʗ�А�w���I仩�˾�G�rkL8<���m��M��[Ω�Z@��(�u�{dx��Uv�,W�Jl��YZg1���X2��R��4���r��޸s��kp;��~�Š��/��X/2s�$�x6"�HZ5_��FIm��jt2p���>H�њ_.e��29��K'��:��hn���V���]{��e#q�A�^-���������Ǝ�:�^��� ���H�o�L��ww���������Wp��*l�\��Q���q��`�6e��䄍ʍ��Υ=�&x�{X!Ɍ{�I^��3@9B���%�O�/L��d196ߖpf��X�'Fps H����)�7�{}/���:�MS�v��9g�L�Hp㥅�t}X�4�ᙼU�׷DD��m��CL0�k�ˡc��r��	n��LF�����E�hkJ�\�ƅ�u3��6�&l�{2��En��9�Xr8�u�;��~�f��Le��VS"�~�����l��~s�޽g{{;�)fe��w5�G�5�=�	��o�3�8?��d*�	���L�X�6���o�:#w��h}��Lg�P*�p��	��{b�[�I}��n~���	~�CG^��ԃc=C��d�{��Kk<�zkd^@S���l`J�����k��Pg���^��F�/���	i�b9�M+ժNg�^�x!'E��̮&��ΈGT�����n��ފtH    IDAT�w�/���k��������l�K�7?r1$����-�;�2��|p�|�BQQ7��lF��1Bk-���iÃ���	 T#��L�72��N��T���v��%*�$�$�p�������::S�������9�{������Fc�h��Ν}�x���N���v�F�M����p�-���:� )@ֿ[���#� r��������;4e6^���*�W��ټ{�+\�=2��ύJ�< *5-T�S*���l�TxCf@�R9�r8��7�!k�9L�0 �P�0(�}�Bo�ϱ��[@D	2ڝ=�{���ɑ�rM8Z�!��;}Eޗ��mPϛ�7�����P���Dٿ9f�%[gS6��l��['�Qp��6��-��myٱ��kˎ�Zc�޹��1�_���j��>�������u{��}��/�_{Ce*�3T� H%�Ě�l��|4�����=y�L=ڭ�]p�B��Y�Q+��'k�@��f��
D�E��C}���֎zr(`�2`p��K(���~�����\r��6�&�$�z��Z��H)�� ]��e	__��%���B=�����l�T�9����0k��ڨ[�[�Jc�6���6+iC�"�YN�z4t��F��J23�-������_�k�ߖ����w<P 
�b������=��S��Zzn��n�K5~�(�2f&;�����9t����	��E*|�R��t�$)��K�����n�h���<"1�����B���{_J��'	�ٔ���ĺ�����)C ��������v7b�24��*7R�i)X���I�g�>�/{Z�<o���ܮ>�
��:Zv^M#�l�����U��E��Щರd�V,�`5qP
�L �JZ����J��L��%�IZ�/q�*v����D��<�}O�՛C�����l�f$����6}0��Π:��^����ޙ��zn����X��<
�l1o�B�ɸMRQ��6�%��=7ݏU�fg-�][n���ܻo_y���q��e��Bm1�_�{߾����Q�7��G�v˙�kggK����Y�<��S{��MN�1�ؘ�k�!~� v�h�-m>�+���mT������i�k�6���B��\�G��_(I_-[�A(�c� �8��9��;Bp+��A�E����d� �����-�|!k{�������*G�.eֱ�zk����\���s���m�H�f)E�j*;�)������y����l�̮~�Y���N�i.���6"<��bIz�jh�%FB���}5�I(W	۬��3,�g/����ʡ�Y�%{cc�Z�$m;���> ,P�����T+Ȥn�~�q��f
n'/^81ß��&l7�NAןZ��ܸq�h�z79B8�T>8&P��]:m%zB^W�M!]x��[�l�����%8�`���	?+���bїq�̅̒�H��;��
��+��笪�5w�pNTz�+ZR�����^�?l� `2gwʛ�>*8�^ϕ�6�ͦS���tؐ�����s�'�q�ahA��u���h�e)��	�eЖ@v��I�0�O�lU�ۼ��~!m�\\e)Gm|ze��WV�o�^�~��VffӉ-���{��������Af�����Y���}�W�"Ƀ��L�6���ũ==�-G�iz`2���)���fe��������)�J�%���r��N82�4x�)��tN5�m����<��ՃJٛ����P-�A���(Z5E�+u�ʊ�?�bZ�V~�AB	H�c�0� 0IR��������_��i���<֞=2XT]6k��"��t�S���Xv��E5��J?�����/����	����}�q9k�������M�~��������l�@�˼��Ce�����R�as���Ur%-��|��}��3�h���|m���v0���l+��J*k�lN����f�裏l�s�(���C�٩����t�.�&HHON�5W������P"�/�	&�VS�����v�S��E>�P���ES�l�v2ɟ�lZ���4���&���|g��h�J!�a@�����1�P�qF/��^���h��B��#��&��t�(r����K�pz�\����O�N@�����`�?��-��Qו��is��	���z@���^���Ip?xM/����L�"��Ev�6,e���(�q_b����y�R����o����W�7�`��Ȟ�؎&o\�%l\'>�ֵ�����=�۱�Z�JY<6�N-�3�<��/����ߘ�)SQ���z]��Ǐ�gO���!�%R��q�C�<�q�p8#��A�0nz?^����sCI��=��|)X�=&�"䣃�����P��l�HA��!��ޙ Œ)����U���穐���+�������ﳽ�}[m"֛��ӵ	��hD#���'�wG��Uӹ��z�'^���K_�ϧ,%�]�o���A�O\L�Yx{dn¾�ˈؤr�N&��
��c_��K$�є�i��N�n�BE'�GOۧGO]�٬-��|<��Xڪ����
V��-�`$j��]S��\�T��Ɔ"��&�FB������B�׺���Wn�7�إx�<��̚�D�=�t�������1�Д��Z������dw(��+����#�a�x�a��{�	$[>�dC�R�(U�D!�@���|!�����,Np,f�F�6�Qj�i/��f�������
A~h����o�4����b�� ��x2;�?���b#	:�i;���[hF+=66Cn�J�6�UR6��nqn���fm[��-5���d�<|dwww�I�=;��/�s	r��
���{�}c��ؒэmWk�Ň�m���8P��%WQ�LW־l�B8=�PomN�������&���J�S�?�Ğ={.�X�%ZnN�ٙ��w�6sL�s.�K��Ȱe��!�Ttc�u}6(T��\�Bp�(��}qN=�C�ee��x�Lydp���ܓ\<�@�\�㮮����s)�7v��Cۻs ^H������6��,nb�`���$j*�dj�_)���������P��w�m<��~�h�����0C�Mp�i@p��P<E��`,�[�܄�����&n��m�klY�\ї�ѧ�ؓ���j�<ܶ�ikD3�W*K��-){DQ�I���%�-� N).ݱ����iZ�7%�c�s{�e`�ʅޕ�llF�U�v�f$H\�_(H2���sYAй��v5�y��jKi�6M�P2M�n�N	�-2�.�x����AHʏS�Uʮ��wF�l���υr2�p���^�^���]en|v2�00!�i2�t��u�`��@'�L�L2Y�"���%��>� �O8�{(H ,��)�ӔoD��[ωk2�%��3�G})��f��l�V��-����e6���,mrֲ�iK���ۻk��v����֍��m���A^Y>R網�h`3��ԛ��7�v!�^]li��B5]ڰ;���k;~qbWP�`Z$c�FJ�6����
Œ�^�}a���i2ϡ
^��$�����K	���2M��k�6���p>s����E�$	yR������Q��}_Ϸ,���xB�#�1` �OP��aP��{V���MD���s¢/&��=��ߵr�a�|�:���ш��&�V�k�ݲx��J��p�T�������������<�~�h���.��T	..L����B���t�ܸ���&'��J22p��ܖ+{�٧���XAI�y��G3�I�l/]��JM=��l�J4�&ˍ=��3m66J*��s27���5n�e%W�57�A\��#�'��B1���f��U�@\�,L˕���ä)��,���1B�L(*X� ��y8���L!0���^����zd9L՟�M��R"������R9J��FS�O���s7��l��(i�,P��Qzp4��Tw�$��V���ǹ��(��ʣ���P�K��)�:O8Oԑ�i2Psb>�ޠ�̄)$��V�ز��y5k�R��ٸ�Q�H&܆�W6;���pno4w�Ѵz�`�,Qo w*�\=**��@t��|�)�Y�~�fo?�k;Ŕ�f��_ll��4?NdNsѾ�.���ʲՒ�51��[Ph)���na7ܴa3\k��M�R��v%r�j�i�%쏡}�7dX�hVLs��W�n�E���;�ظ!����0+4\[P�%�q_Q�m�x�dmrd37��5������s���߱���Je�gR��A<�h�Ƒ� !���Q��dT5��K�����ʏ~�����{<~��ҿ��?�:��x��:�M=7en!@.��ː�]34�"  σyP��V�v���Ϟڳ�c5^���sPdv�y;,��N�&���x�&����9>��Cѯ��r%m@n,���t�e�/��2��mW^zV�}H�
P���$�w�fA��jn ��gQ�p��2��� �f�\Z╞O���{w����F!{�uh�kQ%^J�/����^��`�{��gϞ��`3)S�t�I�R@ǔ����n�� ;{���㲳���#�+��N��)�D-�p�K�a��L�ɷ|X��}�46~5sӵb$�G�x.4�ɔ���d<t��`<���M���f,V-Hf|R�ج^�>����M�6>o���-�bͶ�#\ʚ��\[ji�U���ՙu�M��B$�+5{��53Q畀��bc�����Mg+�hݸ�6���\W�Z�g$cK&��4�s �%��OJ��汋� .����RM}�$I<��3��Ø�%1C56�����	G/ύ���]��`�M����������e-�A��L�R�c�m�S)!�?|���2r����ƪ��D�&���)5��¼nֈe�*տ����_������
l*��E���s^	n�r>�v#K�W����&��6\Q����$��L�U�$$:y��k�jM��gG�����`��/�������*b-,�S�^.��l����\�贪V�j������u�eW����:O��͕��nT�=I|�^���Bp��c���A8<A��&��὜v[V=��ė
��6S��� 2,Q�������y�|27�k�\Y(�|�P�D��!��_K5ڝ��{8}6��{%K�O���(�>x:��
b�L��vO��_�s��>s�PS�W�������<�j��M�Cd�oZ.�����pՙ��	[4K
n������m�����m���j�$���
Ʒ�Ym,�Z%�@�5u�����[OgVJ��~s�޺�k�����f+Kn�[El9[Y�ӷc&���M	홴շ�\p+�o��:f��P%'A��l%����\�*�sa��Dw2i��Ӈ���s�~����՚�=�^�7�a0����%;�p�]�{_����&/��	`�dUI.s�tڽ>�7�mwܷ�	
��d/��f �q��"( �� �:��V�8�S���;��?���~���ngn�x������g�G��lǖ�I�����W�JV,��t�/� ������e3���B��o��v��&-OO�t�G��ܹq�j����.�^�l) ���U�r��ط��-��jic��۷��A�/�?&��~lo۩U�������b}j�n�a��k[@	Sj�2�0�r���tJқ���N�����d�xu��:��smxk<5*&�޹'�l �cҌGj.�����(в�o�obx��h�j䀔ay=��W#�{0����ʰH��H����@��:םN�}�F4DxE��o7aVO�;f����y���ZE��E�B�����i�e��t{}-f�m�U�
n�B�换��)�h�Hb�Ӗ��;���m�T��Ib���bey�Z3[�Z��k8>;��ֹ��7�Ϭ��Pc�4�VM.-��¬��a=c��О=?���/�sc�D�2�������#Y����s���BQ�"��<C��+GA�s��K��#�r]��g��V�UU�^u:vvu�w:w�`�����@YL�����VM��	eў����.�d�X
*�4Mw�=�mHa�.�ʶ��e�{{V��l�^�u2�)A�6�T\�iw5�� ��w�X=_��˿�Ɲ�?�'��������27
ǋ�O�n���b�oG�6&���
�2�7�j���8�	�2fҋ�m%r�W(��ƾ�V*�n��I�
aB��[#��f*o;���y�j���g+{��w��h�=�L�.Ps���4���r*:�� ��LU�A�����$A@ ��e����#����bE	?Zt��-�4��|*�YaS���\�ç9�)�lj��0��)����Z�E���7� �2>::r�
802Vk4�����#��H�KYQ������:�O�Ot��QfP���M���/\��p�S�\�Ec�,�O�^�h�)��ۀL�M���R�-�����;���h���7�,Z��$�Rp[6�6)�l��Iq&��hn�k[\v,;_Y9��/�1+Y�
����d(�\\_ؠ߱�fi�墆Z;��5�Q���j���%˦�vuֲ�>zl�=ngX��	n;x���/�L��S�'vqղ�̉5�ۃp�Z�0_P�Ɵ9(����G�8'kʧsb^KT1��&�W�-;>?�˫+iJU$@<�L��tJ�,mJCz������Fɮ5ϯmwh;� �s��؉ftg�!i$�d\����F����\���!��	��ŜE�9�6ֆ+���o�u(�esӝB�y���?��ל$��v���?������Ǐ�7����D�6$ݕ*-kKF�V��:uS����H*�W��D-��Xb���&a��5{�~`{���W��=��ϏU�R>�ᖞ̭h�C�Er��Ҩ�ԝ�Dnח������*�̟��|��N�������@F�)#�
��<h����@q�B����&JvLX���!�S���]L+�ޗC���>���P2�	$��SO|NF�>����WGL�1��OJb&o�뫖vĝ@��޾�u�9���s7�έ$�2�[��!PFr�`enїB��@���i�su}a�N�#d��%7Y��?�y�>�K��Px��D��l�������-C��K;���X1g�b�f����[nUm^��*��5U��ڛ��[m�tG������J�b	+D�VHe$k��`g���|ҷ�|b�r�v�+�W���X.�=p�8�#�~m��{����p��Jp�P���H��Z*Z���&���{3;:>����t�P�j�V���ҥJ�
��	/^���'j��G�f�j0�*U+�����/�4�����Ӄç"��Y�V�;w��hj�����u�0 {3���@O��.�p���ٕz؈UdE���"��D��&FJ���{S.#B��
LXs��%�[�26���V���3LtK�Id���R�_(�~��_�׮�W`������w�a�d:�sG��?u2�ۑ��s�bC���O�%#�)����"+='	Ek���*"(��R�ި��v�b���>x�}x~dXfs�O7�[�����^�jە���i��C@��߱��ʗR��2.r�KdS�AD�A�ߵ�&���Ʊ���z������t�&bpĂ
U.VD#�A�(�X��Y𹬌����c�I�J@���s*�����
�,�M�Wf܂��/i��DK3���d���x��o8p4.J 5�;=7]����\O ��=�%�N�	[8���1��� ������Ȕ��i媾��95��ǹ�v��o;ͦu;7vyղ�n�RՒm*�Vr�Nml�(۲�7�gԓ����Vݡͮn,=Y	$^\�U"IH�V.��}Hy���۰k���ꅴ�+Y�F����Y%����]�� ��|qn���}�;�`8W�|�L���s�o�jŦ}|X�ֺ��ӣ�R��U9�C�v$��C2�V�e�/���gOl=�8�DF/~�X)�VsG�S������%kS���)����={��@�(#Av~%W��֪�鴮�Zs���*"��hj��+�n\��G!o��{�-8������\b\�|�lN��B�bI������)D��rà�7Oc    IDAT`2\�r*m[���~�����~��>���������l�g�����ٴ_�F�6��4*p0�1�晰��fF��t@�eS�7
n�M�rˈ=(7��ځm+6�L��OۇgG⬊��\[~�4������+$3�;"���'�ڋ'�uܘ!̴��٬l8!��#�:
nLC���j�����P�Y��,�xD��5@9x^�x�`%l���N�!�p���5�cASXi����A��?�=�ks2��'�%�gđ�Q�e�p^a�R�@�؟��~��� O~�);��Ӛs�)>K�*Y��[�.~�j>�x���z��4���]Mpen�LƷ���T|o�+���!�i�t⮹Z��?i�1LX3���W�ۨ��U=o7TK6b;��E�3�\jj��V~����V�l���K�+~lԷE�c���ŴU�	K�g��nU����,�<=���~l�|��Mf��"j��{
�[��m��7���}����:-Χ��5�[v�@�TQ�Xw��]�\I���gO��Eb�J�ԏ�pSokgO�	2B�2%�N�Y�,�ϋ)��k�)�~��j��ŕ���l�ͦ&��%��+WJV���aT$�8ln���J��Ҩ���_S���G�۱��3�����g1�X&c�|ֲ�ެ:vM2)��M.c�d�z빝q("�n+&�VO�w��_y����쫟SY������������Ӌٰ�pc[ђ^m�Ɗr @�U|cs���R����E,��*��Tv�Ɓm�k6�M��O?��^i�Y,-M0��-�cSp;�6d�ֹ�R �����S�裏��ʤ�Պ\�,�t4(�Z-ѵ����ց����y����ɡ�l.(*"d8wbaӆ>��&��sٖ���`(���:��H<'�){�'�t (����n�?�Q��	���N�,��
}5��)���z�ۉn&�ԇo�����
�2L5��ޠ:��D��4%�����l�u��� ���^�	�n���� �)!s�q��Ԡ!�u$a�b�����kW�R������=�`aTz���ڦW�����ږ�m'S��J�*���4|�ߵͰo���j٘��	�F�_I��N�v�u��{��O��ob�?}n�9��S;8�#��^s˘�#z���O�ً�L�K&dPs���v�ܐ(�b��Z"�JБcb�I��Y��5�4)������ى�8;� ,� �&�7~��ݽsW?�`6K�;�>�]���T!tJR2���wM�'/����ɳ#'�P�[s{K�)�r����T�6�����z���:1ThhkR����Rn�G��_/�׶(�1Q�t4�rrX�~���O����?���_����x�n��/����z>�r.��7�cqy�[��hb� pJ1hM~�����ʶ��u`;��S�����'6�,%Yǈe8��p�2�N�n�պ��̗2x����޷������M�lx�9��W�◂"�v:����(M���9J��uR�]�ߩ�乐!��
�q���n�_���d��3B�{����\�8H���B�w��ɭ
�4H��6;�<��s�+��k6�
B����8j���-9�/��!���8=7u�I�krY���Ʃx��ʌ���CBd�3sL��p�zMJ{=��\�������s��l��ڸ��a)i�r�F��M�I����6qa��ӕ�N�l����É�F��h5pP/&S[�f���Vsk$cVME��NX)mvo�dw��P����᷿kG=�ӧ�]E5Y��LÄ;w�؝�}KD#�&8\�؇�}f/.�Ĵ�^���;*IU����'o����ե=;V�n�XY��V*9t��Zò���C{qun��-u��m�w���$�@�Mj�Z��e��,M���_~��Ւ�-��Dy0m��u[]�89Uն��m͝m˕�6���؁�
�)��_��UO�AUU6W��`]��ØY��8�؋�kqpS�cq�e��[�_x����}nP�����-���?s2����rV����+���fI7�Ht)���(K,T��	�,�ִ���
n��-m��O>���?��r.��xb���b�7m��+Y�߇}*眫n�ط{�gvf�\��oLZ�-��`ʆl���W�-�$�]�J -��6�֒Z�N��ps���N�S��|��Ӣz�;htϽ��N��9��	�)�l������_���M�S���������SW�t
�t��J��xRM�3ї2!|����IT�ʴg��&CvJ=ƽ2�T��&��[$Ϻ[S&,�M
�e��A]��g��m��_���>W+t���z�ʭ$���2	n�1�<Om9u�K} ��n0Z�RQVx��g+�	8�]V�U9��ߢ�ݒ�ib1W�p���f��&��}���ׁ��k1�{�E���<y[1�N<6-�b�c�*KBg+节��`*�d�#��,�4���p0�7�Ä]� bb�V�mv�B�t��)b�.&�\ӆ=[`�X `�Q
�p�J��#��㰖��QCl�	���7����#&�� V���2��?8���s-�n�����XWq�����K�k��6B�h�������u�&�{NĤ�V�G
�hS�Bg<B��dJ����1�O���	�!���h2E�7����˵H�H�&�=}�T�y����L�M�?$���`*][�ZE�QE*����z�{�e���AOrHYr� ��JIf�pca�6.�����#LqN�""�Y��ҏ�{��Á
W��o���o��n���j�#����0r���v�
gB�����	�+�u�
��b�K�pZn`�T)�Wo���%�+;ާ� �XJ[��AF�~%��)t%�}1��^�y��(hO'���F�y�L6�]L�J�nWtkj��@(�ـ�,��U�7H��;y?ȼ�b�$+�J��#�|�6zK�ZT57����B�P�Hy,oC�W����S�s���ƪR�м���* nP��ל������H�S�2�j,JR�w��Pɧ�mu��c���x.s5_k0�}�AY�&�@�W++7��6�ع �Y#�@�5n���c.�Eɝ w@y�QSLƐ��aF|J0��`��`�h+�
3eJ1��2V�5]<t�dK�s����L2|���l��v��d�D�T�\O�j8>ك/��y��~��CX����	������=4�MDb1t:]�_���odʪ��^{�*���T�{�J�����{�Z]�RJ'3ȤHr��e���?�����Z�$-�RF��l�����a@�P�+�Vg�:��5E�i���cd�I��)`R�Ֆ��`���i:��ViTG����3�������C�߅�X���7
��v�f����/o.�[�Ꮔ����b�~���ώN?�Bᇟ��Rǚ���5�[㵛X���f|�X����|'�V����X-Ŏ��y�N�c�|0��/�F$��b�rU@�����\����9�H�"�
�T���e�F�)m������W����LV�lK9{��Q�@$�� �@�Օm�h4�u���S����ܤ��Oޝ���G��W<�m�m���������M�)	
z�`r�o'���s�2%%B���VJ�̤&
�5���ؓq��Y@S�l*B�T�v˱����� ��(�g��_�����|~7�تVµ��x�<���U�����*�1xVH���X�Tv���[�`�5�յj�W2O�Ĵh�BN��-d�*1G!#�a#�u�zB�x|�G���|�bxu���D#��~�!f���r8v���f4��t��4�>zZ���#��	��Q���~�3ؽ)�s~�Cj)
���s�ud�Iѿ{���^~�
���W�^-��Y�V�*;��H%���[��>b4�!��#�N!�߉Y&�$� q���	�3���� *�a�h�g�X��P]�M�:�R����SÒל���r�4b̧��}�yg�Ώ~��Y���F��R+c�`O��������]�����������L2�|��8��ri� S)���%�cLH�FQȤ��J�N�{?����+F[���i��^��5���m��@X��q�K5� �wŐ�X<"�`ZS+ƨ.!
nw���b��3xV;D�P�^�^�M��D[G�hvs�����{�qu��
ܹ���K|?�����f�X	�юœIq�O?~&�?��a2Q�l�O��(�rӤO6�^;�X� �[<�E���Ubn޼A,ť̾s�P�jaU5�~�ؔ���5M�ǣ��`D%@���}J�hة+��o��HkM�fi����ñ��%o&���e��eR�-�E֕���2X�Ұr�"�=���ǒ�V]̨��r�k��y��htr�%�&"SB���7Ǳ��ce͍Oh�X���a��c[j��nF6*��xD�$!sĶ4�M�����br׆9��j�\=��ra�]ȹ�f<�f&�g�<9��v��":C�������b;��5�]˦>Q*�����6�e2�h�����.�^���(@�JFł�R+ɒ����j+������]��H��nq�G9�DnV^3�.p���!S*I�%־{5J"T�=����5�\¡!)�4�yrH9_b��
[_H�'���*p��2�X.�Z����j���ܷڸ��E�ے�����6�xF��r�LV,��o��� �F|���Ԣ��������������}7����_[[�����Y�~���͞eČd��TyR=�"ORa*)_g��M���(-i��6 ����!�GO��m`�<\���5���N�р�?Ö7lK���~��r[ӑ�/��|s�[�����yY�tJ�dV�hQ.E�yn��	hf[�gBg�׫�&'��[K"��\��e��=!8Of��1fR��|�K��s/��M,�d�N|�IT����;G������S*J���y�,���:"@��_�	8*���܊@��Q�/��jH�+Fu�j�/%�8��T"�i0`V���.�v������7ź��?�7.dKJ��mԽz�-_/37{�R�^�o'S�8������0`D VG�R&���06ܪR<��'�"}� �V���C�n�D\f�ܴK�I��)�B��m��N��a��2{5��#�.���/���b.��	�V�^��'/�٫ßN�������7�x��Ũו�A2E��<J{�5�/�$xڱW�����N�^T��-��0��;�����]o%�fLW��
!�[2i����),H^/rq%u��-|��lC%�
��dDfd���B���-��CGX7͇c5��UH�~rE����R�x2T��lJ��O��t1��baLC~�-���7f¡K%��z&���~�?�`�GJ8?����-1s7p������խ����1pƚW��|�(����D=�Ó�#ԳU,��Y���wbIM��-�~�B�ݢ����O�q��?��d&�A�<��B>���E2�A�W4�r}e��6��h�+DV[G��x�����<�(��
�� L^�<�@jV9xM*�.{����R����N�m��m^���:����rPe�F�vʐ��j���V뜁(�T��-9<feŴ&���)��R��;�� �)&<NE?Q�YM��q�qDv�T�'���tP�J�ƓFod�����=@g�J�TPc�~����r�&��+�vi��d�tD�y<�E��r2	ر���V2�M)'�:�T�;V&|ɱ܆�uG=�1�tEKE@�\P�;w��c#eۨ�W�[&�B~e���d{�"j�"8�ݷ�>����g�8�B��\,�C�h���@�V�/�z�C����W����c6�H'�� S̢v����	��"|�\/l\_\�����6��1\�D��A�f��:r��T��y2�#�@C��z[O�
��1�`�9�M��\c�d8!U�蟷+��ŜpV��S�ș�a���0cw;YT��)�0P�@�euH*û�9�{�j��b!#m5�!��),c��� ����1z�\���Xl^��胂��s[���9�����\���pc�a`�E4��q������6pyU�����;�i�+��T^$[�A��������Ybg;�6�/F�K����'�PJrH:@��A�f<	X���m)y7��ڂ������s��Gn�(�b.?o������Q,d�k̔�y�2[3 ��!݅'�^�D�*=?����~陘���x�E�P[O�<�6R��`
��3w�{qz��0�<�LF���&��)�J���5]fǲ�#�C��0�dO�����T*�"��I���v�~�n�]T�c@�S��T%$��7�z�A�2a�/ �����Vg:���%���c���l_,�0�l����hw�+���&�JE$_�'��ĭ6R��7~$`��c���l�C8E*�E�T����a�FڲPv]�9�� �r�޳�ky��yl�%��h��B����N��}$�Op���H��&��}�ޛto�M���E�)�P?=���H�� G�9.�\���5:�eso.��+�Ѩ`��HZO����nuP�C�(���'�*{5�E2����Dq���pvlk]V��\��w�@�^��s�K0g)r-V��x&�R1+��b���F��w~��:�)A?E��8ܫ	����U�Xf��Y8�E$��v�{s�������X�,g���O��o��ʇiK�P,�ߺ7G�I�2�O>n�v+	�l6H�CxR��ZG�!'���ib�Y
��4�����@:Fx듊j����aÓ|H־�b�0�ꏑ���K�O���@1�Ĵ7D��^�ٮV�G���R!�Ѹ���Ɍ�I%S���dއ�{q���J�\6-	�|^�Z��J��E̽_E	��9�m��ig]5S�{�RP�֕�T���y����T�u+�8�X:��e�ɡ��\K "�M�H�'	���Ȝ����e�\��g�E����C��^[Ma>��u{���c���'P{bj��Tg�w3=!��ӝ_�̡%����㸂�nPsER4�mi*���uD�ʚ�T�h��c� ��J���'�d��%����S����7P��Hl�H���>�}k8@(���)^ʩ��� b[H�&*�%
�9�#a</��=A��BqV3�;<�:Ǣ=k|V���A�^B��?y�d�Ds3�|6�y@����GL#�����7��=?�����bQ��p��[ܼ�@����h�M���<����g���g�"Y������Zw����2g$͉���AC���T.�s�T���r�ٜ�GRw"��[ݫ�x��ӲŪ��^�|8��jE��hׯ�9��|0L��w���|8�o��ϊQ,-�|����>`�7l�`-�!���W��U�f�᳽����-��gZl�˿{g�Ӷe�����%�;*������?A�'�r���
��+s:�I� ` �v�JbF@����s/w- ��pzC$�5>)5�����E��x$WJ��ZR�I���-RVtl�dV�;�ʒ���R�9�C%�f|�P%�t�M_O���.����ݐ�7Ot�(�tVGlG5�iՂ&��6:]�?SvG�ws7�iT�(3)O�O�Ἃ�R��a��/��\��en(���`��V:Q؊�����'+=����0൪��Ǫ���7�8���i"���_Iˢ���	7JR��ǿ�=��(�y-��ও$fI*gBUH��J�m� 䌹
���3�;��^qj��siK�Ɉ��l�	��9�98�ֱ �A��	nhB@h@��"��w}���-��1<�����n��4�t�3,T��O�|\*�ϞH�B��52�����W��-���[c�!�(����?B,W�a:I`ty���T�n��d�(5Q}q���c��M���q��\�<��%3c����8|v��/>F�� �Y��޼���뷸9��b4�]�N��8�nMȾ�i	o��a:��'�
s�MJy�dJ��,X�1�jj(p����i9�j�Z���|��~Z6/P#�ۛ�g�B�UPȤ����֏)Z��`�)�-E��f.�q�93L��b:��g���7>�������wg��e&��O�R6��T�I���)~��r�$f���T��k��b��ʕD�d��d    IDATmd'�}��)'_���	���s��<N.��D���pǙB�9]V.2�tq(�ZA�. s�B"�F2�FR��i5CJ������=����i?���#Vd���$8�!X���I��M&��^X�^�YϤ6[U��/]�iN�xhy�	��7-�"��+�#M�U��\G��R0�*-q��Ԕ����Z��[i���
h� @����� �w4IX7�OޗV/����^�-�~>�D�{���y�@ͯ��'�R�=:�r��&1P�5n<~/S�y��[[���L:p���I��+��-g�+g������S�\���_lO�vS#nK}�\[���\�lR�c�o�u�3-U��'�4�S)�3��rI�T�[#ܿ���+��8�b�]"�l���c�<�`*�}�l���k���0����[��*���	JO��?l��ˊ�����kܽ�0�C���
�N������@,�W�/p���o/`��HE�==~���=d�%�r�-[4���R�0]B�6�8l�!W�0����4�j�e��n�D�M�l�V��AC��l�n��^������Q4+%�3Id�1D��������ho�n���!2GKN9�����?��&��̭eM���z�Z��@�X��^y��n�Z"���໴��$G�*�����d��a���9\�%nв��Y~����R N�{	9d3�.�s�up�/�&��C!����4C�B3!�FIDś+-+�d:#�����"���^K%`���񀹌g��<��﷜Rq������ �[G�6�����2@��&��>�f���<.=S�le{I�#������ ��s�\��R%�VR�*���T��RY*<[R�sxU��u;�]~y����F$�r�J:��&���fWm�U�P^�ⵉ�hY��a���\�PdY�T*4�y?t�LS8��l�TD	�BkVo������%��]p�E���`571oa��X�$�����ā#���ʥ���Bz�@nj�f[���ǧ�
����XT6���6��9���5��lW[�d����>�`��z��ͫ��_����4��WA�g(�!IZ/P�5����~�����c��5������Z�ı��q��
�o.�24�c$S	�Jy|t�R��d���X�)eTCtzC��3�j�Я�QC��D&�����/)V����5�*2�JbHY����Z����fs�������sD�;�J6�Œt��_��g;`
a���[�֘��^bKR"���?��������~��k�������v̈J��2;��
�h�k{xRo�ImO,�C��Ba�vЙq���q6@?`a��"WR�sI��B�֎��4��l���D�Y!��!��!?���N������:���e��u87�:�r9������իW�I�Ғ�e$�L�q��]����=�S|3�r��.X]�:ANoP	���7��*�B|���d�dK�������e�w߬�p��3Co�~U���@�����}�<OJji�c�������BF�y1"@�L��uo|j�C��[&��b��4E��G^��� n��S��|1�6�{�{;df+f@�QX�(�d�l�ı���.Ϲf�na����B��h�|�bV*�Z���i �� 1���,Q�,|R,⳽^4ȳ�]Xx��K\�>Ǹ;@�V�z<Gu����c�=9�]l�h���������)����P>�C��T>y.�3�|�&_����9��7X���'�(�h<=F��a�4�~�GZ/�0�~����|�p*�\��Ƴdke$H����g	��;=��3�3��T�TD��P,�≄8�0ǖ��w���E��H�e�ptr(��k���`>�����hЁ1�¿Y	�U%��y$S11�\�ic�Nc��εqg[�3_!(��e)��g�}��������/Ҹ_N������m��lKiR�M�j��r�l ��|��n��#��"�(�7���o]���6��lmI�a@?)JP���3��k�;�_���O�B��~�$b�
QZ�/׈�H��B7`�#z��@ҁ��2��{F(�b� ��ъ�s7:�L��>�'��g��+�g�#ٍ$*�Y�'��z�}mv�!�nE�}�c,Oz�R�{G���W Y�{�&�"/Toa��PR�s9�tZ����
����E���o>�<��&�f�}�
Lxna%w�kEp�~�l�*�']���ˆ6��HQ#xQ~R	!1�4��J"��4-���.l�ʇ�V��W����	&�9� ��v�$�h��2QlRQ���*��a�2YY��]��`�~�ppG��A��C(�>�~z�-�ȸk$�&r���i�Y>����𢹇|,k2��?��g�������d��}�?9F�� ��$�����o0�~`��p܂1?OOP}~�ҳSD2 �-�_��sv���-���]x�h*�j����2�GЅ����/�0�}���2�����WQv�T��h&��d����rAa��;�О�	n۹x�e�R��6��~l���]Z�Ϧ(�r(�S8x����#Y⹮���h0���F�6��^�};�*�22�����h1y,��4ƽ��~��s@��e)���������7>���_��^o9���9�w:�"hl�f�@� ��?�dF� �\�T�t^ldA���1�X,�8<�=S�6>�P4&�O	��p�fIٿY��ϱ����OJ�Gl鸻�"-����=�a�^��X���A��9)��eɊ��&���U�\F�Q�Ko^�n�N��

����QY��R�̼��s���R�DUV)�~\�4��JOX	��7�F�=��<l�\/�2����9u�W�ɤ�X�rK7�������R��\1����
Vfo^��<gRM5��2�K~��FҸ��$>��J�y(䗙�mbm/��,ȟ��65ĴΙs1���e�bidp�V�"X�`C`�SP.�>?����h&�tV�II#a7S�!��c�gZ�
;���0k��2Waj k۲Xx���{��p���^���粡$_��+�*��e�i<yz" Whԁpk��˗oк��AM�҅��������G� $ˇ(0�q���2��tZbC����%pp����R�� 7��
��
��G�y^-M$*�}t�t�e���qʙ����G:�F�Ԍ-DF���[*�p$��r�Ao���;<�<`<�4f�V��6�nTU�H�8�k,�y�}��a���d �]�ry4M���H�pv.Lw���v8�I8�G�\�i��kozY�g��'O��-~��ͮ=��wF��u�Eh����1�X�a#�V�� e!;?��,�+��E��Ƞ��	n{��k���Zyj���ٗON:�ă��j���5ͅ��&�HЋ}�ia���l��1���:;	N�IE�Md��E*OvΏؚ^��U~=#��r�уJ�/�Ei�;\�����H�w��+�����Hd���]2$��ύW�uU���V�7�
z�-<& �	�����Y�`x$c-��n�X0L���ȹ���T�x��XL
��.��]���2ó�
T��A��&�+_P��E���_N�v�3�i�b����'�^^�䞌��	�`Q_�#Z+`�I*2H9b@J��]���Qo��`8�&��?&mdj e/M��(�>+W�Ǉx~p��k��������h?t`-LY>�݃r�b1��^<C�B��H+!���k��X��1��)�0N����}�	n�lMp�g_`pw/\��f� �4���v��D� �氚��]?�����x�`� ��
�����d� _:#�qk��}��D����������"$^Gb�,��7��w��)���z%�R%��~�JY
��a1ui�4�w1��Ǯ����♘(�掋�vF0�y(��f��z�>�i�Eg�n����ǧ/~�7>T����3�����kcZn��W��R
��[�Yz��H�B��ɇ�8(װ�� Ð�@![T��Xy=�i/��?��?��c��?���-<\\��$7��#K �D&Z`��� ��(����ᐛ�x��]x�����l<A�w{����!ĺɫ�x�2D��ƪPY�+�%���1W��o[2%�"�H��ȹp��w�M����բz�e������"�*����6���c��9>Z�{m�n5D�W:�Z�r�S-o��Ĵr��' �ce�X]�I����{���ڊ\���CW���Z����<3~p:��m)bֆ?(�\(|��wn���*���xD�2n�"��b؆����l��k���ᷖyV�2�Z�x��.6*0D3�-B�"s	�B�;Dzn��t�i������^��L����s!J���Wr#� ��(^|�\fQea7>��]�Wv{�(���nOE�ѧ/�
Bpds�2몃��3L[=X�1�[�L�z	��Q?�G���Jc�����|�G���P؏�A���l`�~3��
��!.�0��:�\�S�T��b	�JE쎸��9+�;n���4�]M��B��A�VD�ԕ`Ғ�^�`�QU�c�E�R���[&I�6/�=�1G �`��m�E��H�#	�V*��/�|��~��ү�|�q9���|�k]c6]u�c;���(������)�1׏\0*�vP�K�JYή��R,�Ew�#�c�VE��0Of1;?�m�p��%n^��
��"�YrE���n-aNXb��8��o[b���FגD��<E�j[�����Ź����H��9`0(rn	���Cً���j�J=sS
���[Q
�y	��RVn٬���څ�'���%������,����MD�������������#��0Y���z��K�N%����RTZ���0B��Rn7��^=���i�<�MW�J��$j|���f�RM1I^�z��M�����/jZ= ���$m�&��X@�/�y���� � 1jO��"s7r�)QsKQz.��{���q���'[i�d�."I�B�7F�\����;�^T�h��2{y}�/�x)���RG��
���G��|���Z�����_}����r�H󃨟���'�P;�G�`�L��ww��'��f�i-�ݹ��WP���������nm_�a3] �#�|\G�YAn�&9`n���ઃ��;�:��ͨ?:�T�5�kud�e��q!�W���Ad`l�iG��ֳ�A�V@��6�� ��C��G�.&�.Lc��������#Ԛ{�R���M|ss���0:�-��B3Ä'��[.��;��󃵥����L��v����9�+䫑U�senf�N:�|"�t ��j���Ar�G#WƓZ�bqnE�t
���N��7b������]�;�������9����9;�raJ�Z�PF��%g%65"��m������"m�"r:�s�)�+��	���/_��ؒJ�iX"���A}�"V:2{����OҢuCrO=p{��%��`0G�{|��15x�g�xdګM��tK*6GA����Kp�-��f�䴆���)+ts���4�|6'���\���MR��>{��Iɼ?��T�ތQ܋=�^�?M*?i=]Y(��Z����r��}4���g��<*]���\�@���_�HQ���\`����FR:d,�H��D�b�R�L>nX���a�v�l�O�5Q���&��&(�.��^�8�P�e�+`>�7/_IR���h�"7�y4�ѓI����8;;ǛoΥ�g7��
�HH��O���yr���p�F�.�\��?�\>��m�\��i����ST������py���ߠ{v	��"E�U2��i���u�B$���F���g��n=-q�ϭQC�^k�*|�� �='_�^2T���3��a�zYL1i"�kt�uz��X�3l6�T��j���ͺ�/mt�3|qq��6 #A�Cw�b�[cKC�Lz].���֏��F����w}�.���b��w�ydF&6���=^$��T
Yr�躻� �	�K��-��/��. �|R��|i���e�g�(��XD�a����"��׷x���?��x�b<�R*+�Yl�7�%37j�ș���h>ň!�k�B�u�
�IKGyOR�to߾��� O�D�հ�N��NƔV��+=���j� �u��7��p	n��R^�~�Xy�*�rC+x���n�Ҷ{���
����t���'��剜M���\u5x�6�?#�Q��� �cd��L�m�!����-eӤ�y���3������d �W��[��hM��ۮ��9k��|��e8����lS@��`&������'HW��.&����E��eT��@<*j�B�"�K��8�~~�>v �׬���r�4V�,�ܲEg�Sz�e�(�R�N&x�tqvv!x��7^��!?��%�+E<9<@�T�M���K\�_	��[bΓ3��4N�����2�Ak�7�����L�+[�"�B����}|��J<_n���K��|+ˇ/^�S1�=�G頎��X��X��]�pw~c>����w���ZU��T��!��n�>�����۵�h�7+�;i�\�H)��V�]*/����t�Y!����l��CXX6�c|~v���3��;tyQe���)�]�ҙ��t���w>T@̏_��ڛ�f����9��w�g;����&D��+�����p��*��1D�FX�w�掅�c�^��>��Y�Ц�n����#3c.&�wW���#h,�DQ�&��
~J
3TE��e���v��6�L�漉@E�B2�N.��^O�!RdS�S��liEs�N=�n�z��\ϩ��&����&S��~���x��X�l9�"�B'��xz�o�G��Ĳ��*7]jAJ�j���d	�zs���ya�ǣ�C�������d�_]]���n�y\\H[I�;{Tϒ]��Tk^���}�b��)yl�מ�$AY�+�K��h���t�p�a��^�d��.�ٚ�� �M�|x$�6[���0%�+Y���"!1P`F&�5I`�̎f{�����G׋%w���Fz�"�d����h����~"�&�.t�5l<�������E��o �l�2N�MĂQ�Y�}}�G.�%��+�pZ��5�t���>N\羍���x��[�R��l��*>��9�K�ŏ���9�XE�M�>ca�A4�`��1������u��M=z�s�8
t��ŭZUr1��<;�j�����P`'����}�(�b��n`�V<t1�,o>�Ҟ2�d�z��C�
14`(�]o��.o��G�`�ݠKL��4E�Ī�+���������}�PfZ��G�s���Ͷ���}~�l#Wl1|�6��+�GH���f�8�5P�����d�qE�p�x��d��VʺgG/(���_ڞ�C�pL�I6���o�#��"��µ>B�$H6%�ML��R����@�z���-�_ɟb'��[���������`iøE�]����S�w�&�7�w�K�<[TO,/���2���)�c	�Q,*��J�@(�U��yL�_�|?ӄ�����荨v'���u���Ǎ1�!%;cx��q����H��[t}U�I�kh���%r� ƞQrU�����E ��!���K�q&H��ͷjҁ�s,O5H��h���B�VA�ԍH@��h!���IiQ-�Ffr!ʯ����@���!usvg��8�J���`���Ep�"�b���?�"�)"����x帲�6Zd����IW��-	���~��v���c���@�7�.��J�u6F.�ē�C<9=���G@8���+�˟��.�BK�PЇx"�J5��}���L�%�����뷒��J��P?j���H�8�[�^ߣ{5��Ӈe�drN�:����z��D�.�]�aJ�x���Zvȕs�4k(��+��,:W0C���+���l�F�f�lЛLq���G���[o���!� o0fW��I�����(�zX��n1����L��PAn!��W[Y�7�E���׭�ɡFo~��j�3c{��I����"j��i    IDAT�C��.?��落�]���J.��4��W�u&�OM$w429�QI��썃a��d(Qj9�x[�:r����V0&��6lIy2__\���* ���)a}
1`z'�v����⼽�y9�Z1�r��ß���#�����T\<<�q�{���[q��ykZQ��j�x�"C�u˸�[��
��=x�r���1%��gn�JЏO�߭I�%�_匒*"����}^�F���N ��G#16pL/�j�4�JvG�ӠlJ�z�m�N@jAw߀O��ù�d]:!�x
�{���Ÿ����V���,�q+�,Z@����5VKl�����Y����"=_#ҟ қ�ov�C���<��z���V�����S�L����h��j�J��
W痸8��|nʅ���X,�T4 �����x����n}���|��7h�wT�R:���n�t&��|�����'r8?������Q:�\R�*{���(��J%L��܎0��,�;a�ͥ�R���X���,,�!�NI
^�e��&<�E��C�YA�恛�¸3���p��9�� �� Q� ר#S���L���?��Co�BJ����]/ѧ��	&ާ�V%���'����?�k�w[����k;������J{e��1�:��0#a!��P2����'[��rO�PNgP�䐌%�1���s��ctfCt�	�[>����#,ɝ��zY�&{���*[=x��K��.6�)B��T�\9k��x?��d�'x�ӕA.Txo�8bT.D#R���C�*~���<����@N���i	���c*�NW3"#y���S_���=��~���"{�w�6�^,o��� ��k/ס�?�6��I�ע�V*�J�ƽ����f*�զd�z��PPU�z�(8�����W���d'yL�v�.��C�p+(R��h<�~PLͥ�<6��b�"
Z	r�y�-�9���"Ǔ4V�c����.%�	�ޔ<7~� ʆ��J�$��!�-$+G���0l��Ê2��� �p���M$�r[ K9g���-0�,�z)���<�Cs��w.ұ��"�"6�77w��@�3ڏo�tK���X�Nq��D���s_|��/oE=��
M4wk,���lK��$��}��7�mY��)9.6G�D�j	�7�\<$����+tG»#RG���U��iM#���.�,�Ɲ��\�b�/Ԛ��HT�@8�����=A��KRo�B���(��,2�V�t$�����.SX��xm��e��T@�V5����T���
Bmi���G{��u+6��*?��R�'���s%|������!�>J�63�t[���04�X`�u�����Fx�1�!`�-'���r�P@mr���W��,���6������d}o�+љ���X���J���$�ҋ���<iy����z:�H��QfM��hsͶM�,��G�UA#���F�L�ו��܏?��ӼU�*���
����y�7�0��R]9�@_6�J���R��r�G�$���ғ��+��W\n雷U���s��Z�%�6��K���7�NP�e�"���s7m\)3��J����ٯBΟD*K��{ϭi4�J����#lJc-L&Χ,g1�.�[�qf�s4J��>Xۥ�c���Qy ����.�IY
m=�(��n���Vl���%���D�-n���z�S��Z�͚/1[ذy��c���Y���[���(g3��tm�v�+%f�Fd�!-l���A��c�`O>#����h���2&�W
����6�ңN���/��縼��
;��N�l
�d�j��� !�U4�|����r��J2":�b�$4�\��`$�%+��)���` �U��@4�C.���Q��:����1��п�bxӢ�|K���\�rN��cU���������̂��=.-ٔ�S��4-ؕd�wj��?�`���?�ӽ����ѿ�w���`�b�\��%
�(�֚���3|�<B~�g��NGx�ў�0�-,vK6����fxp%W@1��=]����V{T�~غ��'ҿp�/��Α\�P��P���	B�����$\����d*<+�X��$�72�ecH�O�,�M�^��!�f��ɫ�-B�[Uއ�̿5���]ͨ�[���,M!�OA��Ymi����*�N�����k�4�����W��6]!*ٓ2�d�-U3�p߅Ψ-����K�)#��d2R�恡�N��ja"�n�Z�8lzq�^�������(�f8�Zy.��q�H�d\d��M($|HJ�2{UDEL�B߲�6grB������W$��{���3����8�[P��P�c���(7�R�Q�`�ߝ 025�i�%����]k'���Spϋ���|D}@!�@"@��mY��p7J�F�@�}M���ר����{���q��I��?E��C>�F4�GķC.����$�Qb2���%��Z��E���8O�!�I�[/-���,���>޾�@�;����k4�G8D�\@�IϷ�����2/����j�����p�pp�r� ��oV��� ��7A粅��#��͢�it̒(#wPG�Ґ�m�n���_^ݡφ+����Ƙa��b �N ��/j��O+G����*�������c����վc����p�>_!��\p{~pױ��MG�h��q1��a�IF�biJX.��7�̍$�Ù.Dd��7cf2a��z2�]��!���q�0�J*}~D1C6{�O(I'�'�툶P|�ݥ��^�Cp�F�*��Y�|:C�%TT�
A� n]	�aU9	g�6.4���	ݞ���K��T8G�I���ŅG����jꙙ�OU��7�<ꅖ�)J�ڲjw]5Ƞ��ᖶ١
���o�[U~JȮ,g��Q/�5N{o.�Tj�A�n�����c:K:Cu�P>G��:FUn;��1x�3�/�!Z��EQ�.	��pS��0&[Sl`��Q���vy��&R��ɽ�(DqIbc. �QW�)���H�v��+�zS�:#�b��Kq�`p+��C�&Y#	Fr,B~�C>d�t�وj��6�9�%]�	@BLH�"����69r�=u�cI�_������(���|4�r.���:"!:o�����3Ͱ�`$�H,�L6��fϞ�`� �b����ί0����l&�p�Oq�X#5Qi��(�E�O��f���pK�(��?i"[� B��0�O0��c�ؿ�[s�p���
G{(7+s>�|l⛋Y&̃Q��"�x�&��?�d�D�h�J�q���>�p�G_��G��?<.ƿ�sL��.����wf�!�e����)^��(�F���nǀ��
��J8F�r&w�m�T>��PF���:� �
��Ӆ�����K>�RL))����;�c76_n��EP�Ƒc] ��ҭ�a����l9�G���[�����[Hr��}�e���b:�,��ʍ38�Ex�'V4���bH�1�D�����&��Ǜ�i� ��Е�hD�W�W�XL�B&�H��O�O�����I�|����z)���ŋ���oV[�#a0U�cA�`!�����[�	p�Z�����*�*���L�V�ԾO�+8��IȖ=��7��LX�v03a�9�� ǒ��lQ	����҅�gy5҄v~��E�����by�s��kdV~$�6=�;Fpb �\���%�S,�%vk�E�G|/X%�(��Ƣ2�'A�ձiѝ�Z\�='�%�	6��"�l�V�0O$�v	���l�|�2�3�F�Q�V�:3���h�EB4F6�ko�$�����8���KF!oi�e�p�R�F�2[� Lk)�l��0gS1�t
�������5z0����0팰/�����`�b%�ړ}��J�i�:C|sy�o���i�
%��q��R��"�)�����r\�������g������њ��hi�ON�+�%)�oJ��ӏ����κ��[��,&�6p�X��r�S��
���\$����Xr��
�%R �����I�B������	LLM�P�d
�XR����2)<���3e����Km"PpH�PZ�x"�R�(�CVp�VחW*$��U8����T*=�Z�o���/��Tt�5����Z%��^(3o�]z��L,�|9�Y%qF�J��wޯ̬��I��j֤��χ��)T	Ъ�'�;,�Jl���U}�����+ T35����U�xo�;RnB�.���5n�U%��PX��^����ن�@�Z*��$sXA���h�]e��N%"5����`@^�q�Q��(5����u↗��VU�a��1k���Ap0�0�n8C�^#���G�#���|_u�^���3�����W�B�
�|�88��^?n�i�J5ys\X��HJ��,X��J���\��w�'��4`v/j�'#���a��/��;H�I�UՖr�asܵ��`����u��#!�կTjb?��d%��;r/��0���YZ�C���(9==5����B�}i?���tv6���T=��&B�,�n[#|}y���N&�X�<Ņ1ǔ��8g�!�R	������pp�[���A��?|�/NZ�ُ���9\�Ƅ��p�������>ƧG���Cb�ܟО�в��.�a���JDhA�6t��ʛ�L���r ��g2�'��o�p��7J�Cd�4�����F����ȇ�e��EbUē%�L��5��Ż��&sg)՛�&b{�J��-��8�Ʊ�ͥ��F��׃ojIil)��hLȾ���eՕ�V ����rԼIW0�M����(��C��dn�yM�1ռ�0[�o�di��/�u!�͵��&N�BD~`\����pQx�����?|�q������"�z2Cs<T	Y��Qd '�*��M.U���~�g (j�M8�u8 ;��e$�Xg�21�ѐ�~(�ߐ�A`#ǎ6��M�^lE�RV(|��0jr��y[����
�p��p*�#7�;�k�.��R����������W��cZ�(Bz�$�)|�CQ �	Z;�K���=#�*��w��Œ�g��NrL��p1��/@��` �-�O$�W*�89x���}�3pG��q"�>�L��U�T����Y�$:���v���@��HD#8*W���JE��	�'*��DxrQ��mq�@�V���>�NŰ�l�����Z�d�g��e��i<���3���A�dz��)����{����_�+�n?��_���?��O~�kσ&)bK��l���~��_z�1��w��,�7p�w?��a���d��c��oŶ�W�VXa1�T|�BQq998T2�t󵃇��\_�3c�4�"�o��v��[p����"� j�^�Enœ�-O�v�����[��Ծk^(p ��pͽ=%�Z�A�VʞXz�2V�"�@<�L{����WF$�����H��#�G�ǜޒ����kʉn���y�*:N�_�Pe9�<n����4J->�;F���zn������7)�@^?.�m���xK��%�D�:��|}e���zt�;/]+���!PJJ�t,բ�@�y"S�W?lZ�B@*
_:)��n.7R[Q���2Z���2��{/e�'"��t
�jyA�z���'���!v^KJk{n�y&ň�7��)i�d�C��9b�*A�VM�ֽ�m)����b�ʙ�!r&�z�u��o8�X;��!׿�ʬ��K����[à����U?[�P���C>�@�P�d7����%���Rnv����b�ʛz��Z��L6���Do������c#&//)�������rFc��������X|��2���P��$u~�\�WW8���&����T�(��b�m	g��'R�f6��������?��_m8p3�?����e��DW
���ǈ>.>=x�g�}�e
�����ږ�Y6�qF��-��v2K�+��C�B=_D����͞l_���g��н�{���9�M`!c ,�I0�%��U*aP1`��H�|�*�hI���ߐ�\�*v� !0h B���S�k�����<��u�(�ݪV�ӽz�Z���>�3|���r�V���+�ҳ'�g_�+�l�e>���YM59�_�-3���%��j�h+�1�E#n�Ή�Dvފ�GR���0S'Ǒh��d�Q��{=;���ݞ�	Ȯ�ce����l�.���Hp�T�2x`�$�}�Q����>�JSZ��Ƕ^�4A����Ȗ`bH�~�A�^J=�)�;�LDx��������:R�BY�k,$'�������#X��^?u�0|_�$qz�pu�	��'�49�}����&p�f�F�
��ՂmZ�V�4��9�?g�,���[er���l4��GiϤ�r�����m����kv~m��=e�� r&ȓ㯠�6Ityp󬖬�6���7A�!����r�g��!�甩*�I%e,�ט�d�y"d���տD�gy��$�=?�lN%,j�U�u3�`�	�kKVY*H~��R`wOϤ�v|r�~��'����G���H��]����F��v�_AoͲ��]�\�M�+_U(]�Ȯ�sa���|���������_|�^���M�`��/����.s��kz��ig�V߾�����ݯ���|�\Q�����A����������_��|�[�^a��0�gx�t�],�Ó����qz_'G�T���Yϣ�g��������:�؛m;�5��n�Ȧ�pf�vi�=b_y�Ծ��M�g���
��6��p��<]�FfHՀ(�6�8vXm(E�?��)IeY�+�`}m�x�%�� ��SJ���6���\���s��t�X1-n��߼/`L0�4�;�gQL�M7��MY�~�L};Xt+�t�b��':�g1�L�3�=��2hq��X�:{����E�U�@���e�K����᳐�2�7=%(�-�aQ�PP�����it����1�h�4g�O�|�rG�e�6aW�GX�%�J�v�H�׫��`"d��!}��z9��3���@@�˂�)�������C�,���ϖ�R��P�-4u�"s �y��"�NALmZ-@u��]�!��ָ�ޮp�B�WJY�h���&P)){p�Yl�sm���
��%�Np#z�*�0�X�ժ���#�nP"��W���2#�E��������w�ٽ���˯��J����z�W6��Z,؝���?9��/�W��4����������
��|f�J�<�g���e��=������ˏ��hj�R�����m���6�� ���rR������������~����w6U;��?�?~�ӯ<��>���������~v���
�[9���恝"X�:�Y"��ە�լlSdƻ�
n�r�p@���;w�}h�"�%g[��lh��7��o�n�n��Y�ڶ�zŬ�g�:��:%2
p3[�F�9�Xu��rȝ:��s_�,jz>0"p�Eo� ��)����4�ِ��B�da�G-D|���.�T��h�z�X|4w���m��	�׬Tv�/�O}�}����q��`¿�.A< ?��˥Ґ��υP@��.1WL�����1
	)#�v&~���T7=� ׁ��&�y��PV{9���Z��[�m2z�AḘWE0�n�@X��mV��9��x�Z�U,[���[6kѫ6�@�f���2O�Pɲ׸�1�%0�����`f���*������4�=	4D֚����%�1� ����ue��I��ћ��A������"��d�ku�\p[��f0M"��^ؼ�TW��p��r53�i�'��H�KԀ�++���ʻ���=)��g��+���1�iU�vv|h/�kwv��՞���-�x2�
Jۨ^+{������4l4���K�wo����Vz�[;Ϛ�1��
2�W+��y����W�'��o�}������}��g��'�z��t:�_�ɭФZkCs2�y�+�hY�T��jU��a�f���՛V�m�Y��td(��)K��V�jj�n���jf��~����2t���s��糩d���(���	*�7��|Q�zSXI"�e��[sx�+�������L. Y��֨kAv�mH�vL/�e
MƲ��5�o    IDAT���b+��w\@2iĕ�M���Pa�L����i�+1�S�#L�@PT	u���2��<<S�ů9��U��V����E8�ň(U���<�o�c���z��jKQՂ0�?UU�Hv��q1S{�5��S���$��Y1#�A��a�vݲ���u���`���w�>�|��������@�UP"�.-?���U�� 1@οp�֜o���Z}�Q@pÉ+�ge?IYJ��kf���s�2��)'�&2�WR�O�zMd��)^�8��H���gU�5Vz���]JR��I�N�7���e�����&1l@Y�R��tf�G�eZ�Ygg/�a�#ț�߲'o=�0v�f9��f�;F�#�YԛnOkh9��ِ�iW�$ ���}{rym_||n�����ݷ~�j���9�۬��A�ʹ�Wkv���O��u?����k/$��� ��~s���g�aa�]KrF�g�*/�
֮�dCj�o��Ұ�����:
re�,gK�Rqn��`����A�F��avcϧ�^��|ԓ��t��"[�����N?Y�f4a>n�˞-nzV]g�
/�X���$�]�-�˞���$�=�!'e�6��� �K��u�i.=�p�w3E��N��E �$Pe��0#�Cm�����&�2iJf0�����&D��T>�k���x��x.��E�
�-L�SpSB����<�Q�iJ*W��D"yn,��K�	$�7e��F���5b��IN �7�����%����e4�rP����f����3���$�� ������H��qzNXH*H������s_d���h�:� �O�<�[c��e�t-�\��h��6AS���[��;�,���b�I)ׄ�AvD��-�-��J�x>��AV�0�� #���R�z))KD)�d�P6�D{��r�3?(@���N\o�,0��e=�X�V��߳�s�^_ʲ��z�Q��Î��tdN`���r��l�L� �4� ���hF}{|umO��ʶ=�X��ݔ+v�ڰg3��
YgVfP����}/��S?�-���/$�}����w<���l�O��G�Qfesj}j~p?�2Yq��M���,6
6�l��ם�l����!4	̠jk�	+���a_x��6�쭕l]/� ��c=x90r�#�]������s2��pj6��<%�1h(-6�"�.P>Y$�lg����'���M���J����	zIz�7��7��SI7;_�'���F�@�X�2��P����4��pŒO�.O&�&�:�M�/��|�@6A*I�4�}qɄW)�^�B��!GP��e�aŘkK�J�<��28�W��\��?��eI$��B ��ÌI�{<��mS+�K�OV)YV�T/�"�3�xvy�F������$^��6Ye7�m��M��P=p[�j��� �<3v�6*}V>��P	(���1��^!`�W���"�9������
n��@ځ�5��UlP�!���~�y��bM%�J��$݄�f� ׬��O��MX<����&Q�֠)�>!�Z-+࿱1��phJ̈�b�ע�1�=;9N��O{�aCkѪV󙛤���咵��>l�$�}��z�����Nl�nY�Z���/f6�.e3P�V��K��'������B���?�;�<��?�x2�^27���/0��B���G���T�{��W;)7�~�Hd�{�����ɽ�tR~����ϟ�Oۣ��6˛M�����,e�<��-Qf���*�L�Bf[��N��l�٦7�,����^O��X����CS�Pp�1㜪lBmr2�B��Zj�j���9��A�þ�+	K�g�p�,Nr;L��d�`�=�SyYp�����d��$ˁY��E�OS�r���{RGj��|rr�m��!!��M��&d�*ˋ�C�D�������)�.�-SY��$C��CK/�78%K���u��٨)�����ЊY�8�d�䁌�N�s�C�ߓ8%���/JS6������tO��4�4���[��S�Y�` 4a2���N�
|�iɜ	)��	���]NP�bH��������C���|%�$Y6��ua�]"��]�m�T;��a,��+�"���{KK�Âl,�*�nj@����U�L+)'�q��	n��|�?�^ P񾩐����:|׎TP(�i�PF�,�}���j��Ȥ�r��J��~��P�����زղa�*�����F[��ՊN�|����{O�}�>��|!���{/?�~�Ѩ���&�"g�]�TY�Y˅J��Z˚ټ���)V�^�H�V����q�>停�\�������wcO�.�rط��u7s�첦rx�h���
��XiAn's3��pj��H_W�&s��vX�[�\�M�Df��Jn����)t}s��7���FL@��V�l�F\�}�L��$���'vy~!�$�J4���X��i>���Q����>�/�́e\�Sq�9����	V�5L���21��E�㭷�;���W���b|'��M=�0�!$h���qdeLH'��������{ٖ	�MI�~�Zh�1�#�9=�
�=��5[�A�m�Q�>(z_<�x2��CV<g��g���J���A��\F�>�l
ZGL��m�곥��Q�f��1�A��P��pߒ�J*�S0�C��f�.���`�qJ����p)��a{�����f|j��puQx� S�7���@�R,p�W:�k��u�.��iLkc���9���l��B��X�&�KK)-A���Vз�/�u�
�\�{��f6���m��H�vrl�Vӆ�]��.��39<`BK��A�����O������'_z�����<ߔz*K]b�a�S�lF��޴�ZK"�w��vvرv�nEAW6�L�j���FDsіJ���tm��®�=�+��ci�A���:�l�b�T�?8x:]ֶ���a�J�$3�Y��58���Jی5�)C�g��`���0ǒR�I�``W8>q3 ��\4�ZՍG��L^WO�����FZX|%�#`@ ��Ni¡ �'��U���W����j���BI����*~���2"8���	�b
n��QI��@�qEl��� *�O�8z�<���m>���`�W��=7�Q�%w��me�ʢ_�d9UIFVN�Z�R<F!�˴�a�ʧ���P�`ks蹑Š���n����6�:%Y�e����^��W�b���֔��.lֽ�,�n���,���WK���\��䥩:�׌���Fr��I*.n_��`��g0�?�C��l��U��P#֍k8L%e����"б_�D�c�r0�ˮ�LRB��n��|�V���z��5�E[�8o�fS�U�ADh�-;�9���Ōk�c�<��n2��h��l���'w,-�Q�a�b׶�K�xPJy��������w���������S�N������7G��!��8塰� �R88�W��޶W�Ni�kP�e����ƞ��)�ܾ�t��hl�r۵��g�ך��ٿ����z��f7�f�����싌aD|5'sێf¾�ӄd?�m=�)�1�x�TVj�T���9�Aq��.�������|��g�S�������c C�1~�=3,�"@�' 1���e���J�x	E���$�DO�� Ϥ��lH�է�$$iS�>,^��ꇬ��3�_�l��X�4߄l(Q�Ȕ���{Ų���te��[��Rω,ǃ�U��]��l\7��evc��J�pC	dp�]��dU24ze`�d�ykɇ�Q)�y.{��{����P9݇@@�P�r���W}��{��Ҧ�.�֎�)�v[z_ҡK�\8"���8���Q�W��2���L�M4M��+e%��,�q5�h�$(�2�X�d���2f��y���c�� �T�6�H0$-eT��U<@������6���J���V�{0���r�k����'�:��y���Q}�O;V<A���fժ�K���\CC%=��Œ=h��{�|�_~����B�����y��b��ǣ�?}2����������X���/�{�bg��Y=[���p5�6���ƞ]^�h�P$�W������iw� d&o�LQ��{����o�/�h����(�'�.W�����o:�[~��p��g��e���� �`dN0E$3�ò����R�{wO��载������
��"�ʗ,���gV��H����MJӔ���~\K�wa���譄!��C@����0M0��.�A %��P o���l��q��v}z64~i)�a
Jl�Tn�@?u�i�"���@R�k�ۀ(�*�½M�,@eqN���V��-s~H�r[���V=hI3���7rV(x����4HWtf�rS���l�\.v%;kS�2&��rFIO�P��6k���V��6{ra��r(�T���.kY}���Mp�������pA�ԇ�G���Fpc-��@�a�a�:
(��yt�H
Y�[kI A����m��!l�38�D@,L���)�	�7��Te��R&gU�	h&�l �'��\J�0�P��B�HW-m:[xϊC��|FIڱl�c�r����u3[�Y�m�Y(h��v\*3-��o<���?�����i��?��ﻘ�?�l2�o����f�lHN~�XVv�l�?z��^}�ݫb�\d8o���.7�����<��,�u/C�BA�߳vG��{���V��mh3{�����7�ϟؓQ�VHҨc8�DzY�D�����[��b<Sp��%����r�]�1�����N����d|~q.<������,d�l�A�Pr���EmA���Ⲅ��t*��h8���ظ$I	�����q<��y"�9dÃY��l2^r���n�&�Y��o���u�=7��"XVk.��Є�:xy�c�������.�E�"ey*y58qXF��jX�I[���g���ռ�U��R�I�(�ls�`�,${4��K�?'V���o�b1�H��A�S�Ԓ?w`ǐ3��lyze˧����[a4�,jд8� �yo����^����L��,�{��;N�B
��4��=�t=(��Y:�n� ���(�&�TL��>�L�a�h�(�y��*.y�]��5/%�k��p �e��{d��TEFp�@������,��Q@E��-�����:0��!��}�S�.���r�Jg'V�sh�֡�E��s�͚����f3kWJ)�}��9��n��O~��v�����w>��y�L۸f4�;��}ӻ��}�;�mM�FΔ� �2����4�(/2��K�D��N�)g�oul�����%IJ��}�/��>�0����n B�ܸ������ʲӹTK�,��J���`l���֓��A� .n+���]{��6�г�=�̞>w�NN(��SH�n�U�X��#�H�E�\�jՊ<-�3-9�\���A��IC=�OF}.̆ͩ�$��]C9h\5�E���5}ϛ�^��HY� ق���Bا������	�n_p6��x�	����JQ2���ĢP��r��@����v9Uq@5+�oW�ЬY�Q�|������щ�{����^���-�E!RpUba�"���A�&���q^)�"���e�2[Y�7�����ז뢼�@j"?a���bV�{�3Q��$,`��L��ny��|������J`o#����n�����D�<;�w�֠���V��5�ibˁ��.S�B��P�r�pX�>Sp��9�/�BٮW:��֯3��e��q��oj���(�����4�V��ϡ�I��'�tڱ���mZ�]pf36ڬl*6�)�ݩT���/�9=��_~Q��'>��o�X���t��4�G��G�I7�a�y�{��n�A�j���y�U�H�����}�F
�h>�Ѳ��NG~�Yٓޕ�ś�ٗ�>�E)������4o���㚅e��3;�� �|�K��Ж ��c�/7ҒC��.���|Y(�a_e�6�\������$���P��LMN�%�@��y�C<�d˙���)?rqN�?���E3<Q��8�y	&(,����D.�E�^�R�`�����O'=�o���Z��eA&����I���dQ��>�`1�KS:J//���-�����V
��AJ�W�C^LO������u�<��+��R����K@�&8ty��o�p�����hSS�51]Z�?���\�z`���r��-�#]0���ڑ�Bqe�e�.�	�ה,��[����+�6^m2#���Y��C���(~�!��Ǘ�=�� �������U�6�}x�䔃3�x$�B�\��5��=�a��=@`9XU��L�� �P�F7)�2�է�YkTv�<����3�6���t(�b ��;GV8=��Aݺ����E�r��b&x���T*�?}������^������y�����F�o{:�~�:���H�hm�B��uT�er����t\�Dx�i,��L��邫��ɩٟ]����(W��)Sn��7����.��1)�4%��t�����@��#��ʿB��/49ː���*_��3�+�ֳ;�5U�Z(!Q%L=�68,b<�Ԛ�4�n�Vʬy:�E)��xU��vvr��f���'�)������#�PVӛ�L�T�6�C3��=�p�����A���� 
�JBʎi��}�ﲧ2��A��o
�)�iқܹ�sF��� �8i�p��u��?��^�b�f�zE^ ]��b�)hL�j�VC��jط�f�̏a�6eЉ�?j��P���i���Ƨ����le4�z�L8���e��p�'3ѝ2L	a�T�jCp��S"��4Y%h%7�s�S�+z�\�_sW )��5O�7�D�?�Y�OV���ٜzW�C|_�����L�5�at��]�������{�	.$]0^�>j�$P�Q�U"S��9����RTk�����]/�z~� �0r��X<�\��þ��`>Є��ݸ{�2'��v�5��ۗ��t�R/�肃-����'��һ_\p�,}<���[��w�φ�-!����9ɀ���2ApFo�:���۵��>9�++�=���d���*����n�C.��S��,p��A���s`JGC�)�76"SUz|���[enL��rZG�8Nz�D�� V'/�E��,"o0{&�ʹ����0���t���S$YDI��U<��d�2
΃�P��j'H�Պ�dH��qu}m��P�v6�8��W@4ܘg?���'H�i���G���ep�b:���.��Ѿ�+��(Nx2 �٭�[�T��oT�C��-�GPQ֕ \�":t�IK��$��yɯg]f�=I3r�'�# �U+p_��	ԚS��q������պ�]���o,;[�l?�g�� T���ز�L�C#�1�&��L(	9d
V����'��A�J��J��F=+�[�V��&RG���U��i�3� �C��Be)Mz
L�ju��YC�#丨,�N�%�5��ʶ�|UkZ��i�o���kѴ �ǔ�kG�e��foO甤܃�NBޑM;n[�������+Q��r,Z�wmsضa�d�٭��)�
�n��V+;��n������;�AA��g��]ϧݏ=���r1�������� �Ni��k�)�qSeT葐��)�n@�	h��`b�x%��.h�j϶<yixUpw��VCRr6p�a���Z��JTEd|1�	�� O&��z�����od��5`�j�:7�[����E��%,t�¿� ��t8[�X'-N� _z�u{��F��tI��;ׅS�������K�e�'��[���ɮk=��ؔ����iAv�̔�N����O6ǁ �c��x��I�ۨٲT���'�v	nd<�ʠ�a�G� (�V�J��L|^��d�"h8�"� uM��oC�	�L��x�S+��VǶo���U��ֵ�pd�4&�o7^�俇C)z��Q~R=�.�;|��s�R5䡦������W.��r�.�n:��m��	��0��0zy�R_!���Q�G�T?1P�&d�����ϙP��IA.\�����*�>�u?�����.��� �}>pc�@
L����TQ�RKpȫ��>j��Uu�V�ϖ�u�y�A�+�m%8�c-���    IDAT9�P�EU��Z��o}�{~�����/���}��UA>��?��lx�k�'��X�K��h�	�HtG���Z�!U�fʫ��p�'q���'�FΔ	��+L9�;nFK��`�$*��L�0K,��KSS�A`�'zv<n-���G�̠��Q��x��[��|��#�4D� Qd��r��a�'��	�v�}���>��CKʾ���I�s�xd���0h:Nm�ç��!��][�����rf�a���������8� ���t�}(��L����M� �(��:�����2U�v�6�e���N�ș�9eppG���XC�lf3Wu�v�,e��N�8��逅�E~���df��\���Y�?5{vm�'W����u����j���9	2v{}�ªA���^�ׁ�J��ɘ�C�����^Sp�EBy�5�	>[t(˘jb��b�hU��d|mq�&`� ��7���24�iQ|$��^�5|_�4���`��ɔ\���5�no Uq��t1uc�|F�����I�j����7��F��o�֪[����gwmV�X���.��bAgL�%�/�۽z�����?��o���>[���Ǔ���t>���K�L`SZ+xDޚͺ�	FZԑ�q��u�#=ήoq:�ݩ�W��D�������F�D(���se����f������
I`[m,�i�a�B���F�S7_�@^<T�~CYf��@�{�P`蚂?���" 9��O��֞�tlfe�X#��)�� sS�@s>pdpOS��sC�J��,�tm�X�)��i�% �3< �'J�ǧ��/�If��Pe}dRaD�����e��QR����8�J�l[a%7`�J��Fp�^�,W�!�	.F�*�(�45��W����﹬�B��Nd.\zo|��5�؁嬹4���m���J����f�L���2 �T�cz���]���DL�ᏂZx(HΝVC�i�!=ו%��с�5�,0�,+uMN�{AK6*��&;��L�KL�$�͠����Rs���r@y���M&6�u%ѕ/�fCY��qZ��;��`�;���6�d�O_g�b�d�j�7�?���j�f�㎕O�m\/�M1g�b��ł�;����y딪v�V��oy���>��/�[Jp��v�׷��{<�֮Q�o';x)�����"���N�����{��*������:0Vo*��p�4k
 ��f�VP�@�6��8x.�$���J�A�,Sl��8�����c��$���`� ��[dqh�!r	*�	,C�B���I=<�߱Forʴ�m%t�l�h]����5HT�B9�f�5�IX�[;Q�wI�:�d?ѣ4	���~�����70�`*��)`�,Q}���%)S\��fw����|���T�ʁ�$�s2;��(O�ذ��a������&��Ԑ���k���݈XO��,_���A�Z�U��RC��te�u�ʨH_�l��S[=���x)�VQ� �ȡ����Ź��xn�v�B:wP"Ѥ<gUDYMeodzW�מ����aM@��Y�}����P������rق�!(��X)#��	"	��`!��D=�f5�O��F9�Y�O�����Y(،���B*6Iu91'��TW���7A
7/�>�-z�Z���!���� �[��\{�@,&�׵6�ۑ��ۨ��n)g�]��|���u���T�{���K��������_��k.K��g�����_?����W�%�~�6�R)ѿ֨���.w�NS]4˫��7E7��b�7�M)��A�$� ��t��f6M�4��� ��!�(�sna�y,*&���b��Rٛ2�$z	�e��D�{��d�r�2�r�5e8=&�_}�`K��$((r�-iwR:����}��l$�s:���nXA��T�c��X~|��u�y��d�R2�� �f�[dF);������arB͊�xd�)�&�R�Cz:|�/|�eq`s�I!2IO��d^di�)X�h��W��dn�BI�N�9���$�eL�$X���������G)J�C�۪K�	�x�WSW)VA�t8���k�=~n��UfK�Ŕ���q�$Eӳ�l��!Ȇ�c��?G�Yo���b����K����=�kUeas��9�,�2�`M�ʲ��A��<T�p:v�(������|>�����5�����Y{�y�ӳ�v�����|��-7�����򔭣��o�w��a��I��Вj`>Ѿe�vƍ)p�c����VL���8n���sh�j�nJ9�*K�$/T6+a�h�j��~���g����w��T�}�{�������t�?<�����f�s �� C@��͚�o�`&�n�f�@qSPV�,�Ͱ�����USY8IEU�i.$pVϊԗI����LLN�NR���!��:�2<��&3����K�J����MI�z���L3����Dť��VP�W�oT�ϒVZ:b��sc_ߜ|����;ft��#�I���}�*���C���ی�;�؃*٢����)[4nxDSi�T�mr���ӽFX�b�b�ZEޣ��Yރ�a�Y'�+�ِ��
;Z�.�#�5�l�ԡ�ir��@)͡��%h&��k��-2+�t5]�,�Mm����o>�����f�������Δa����p�ۥ�9��&�zV�v[���hj�;���>USf��2�����<j4-M���3�XY�ٖ���b�0%3��41����d���H����\#A^�rY��U���'�\�+h e�Q-���H{+����nH4ׁCvO�]k耤t���+0��[�c�V�n
[�5�f��MV�D/#��=,��n��_wp�?�����}��ל�!yt5��[��?uK7�O��#��f�9emU�O��B��>���#J1*)h4y��6`@ܒ�n��:���R��Ŵ.�N)�� ��B���[�-�c�i�HNZMYJ�%)�R��i����Ց�1�`��WXo�U/�,Mk`"�� #'�2��O7%9ǧ�K�¥�@BpK=�0�I�C��������m�����~�JI��H�5�8]�]	�3=�Z�'� �`�	K٪lm��(��y��A��I(�5JR���d��(�������.�9ǆ��؉��qMt3�w�6d�� k�UKwp+�������.�]���������l%[<�@��K\m���3�b6J�nr;�֤L�	���ŵ]Fpc�9����6 �������ߗ�'t7�V�U�y�ɍL��P�b���f<s3���i�Q���م�rDɱ-Q�T��C�nq:��)��޷ZP� ��2^Al?��Q�?M�E6��Bpk�Y�����]f6vU�غU�\�m����|WJvP,��J���ux�G�;~�/$��
r�������������\��n�u��4y+��~WF�A|�-���ƣ��m�x����%ewn�+D��$����dn��=�	9�k����(>������Ta��H���PŰË2R�0?�DpI�$z�7��@�{� �ZM�����=�=8���U�F�P�^�.��S�()�Fp��J�y���|h�S���q8�饪��y��	'���E���,����W��}6��,��"���u�S�H٭>0`E]kMz�2�S����̆	��U�����ěۜ���`l��6ytn����[��*���M (��!�>�HP��E���f�)r�����vuu#@-A��m��D}�l����U���6�����u�����yX�$Z ������"6��]�����OBy��K��Bw*$���oHzp�����k��1L�^0��=3n�^P
�:���=,h�}��R�3� ��>u 	�:G2���l;�t��<��s��J��f�h����+_x�������#�B���?�;�\M��x6��Q��*�.�<���Fߍ@G�W��~\�` ��~�/Ђ��c��k��=�T�i���Y)(��E��y���"68ϊX��CXY9c�[��$;����)S� ��8h[ҏ#R�*�jLy)�AP ��7���2H���(�r��~�+%w:_���~�,Ӯ�}{�&:P��{x<��Y���h2�9��2/��"�>"��
�������ZYPG�&D>�:���y g�A�N4�4\P�z_쀘.'��^oTP�¢�Ǒ�q��PÉ�6I�o���_�z��噦�FEr�Zp\X�X�&�D:|���ͬ!� �Yn���� �&9�>���Ö7=Ӄ�՟��7�TO�̍5Jo	{T%�]���6k�ֳ�69]O�a�MC>���zJG*pa��ԗ2����&�^���"I�'����V�CZty)~L��dʋ�Ng��TI��2H
��|Ҝ=GVe�f�J��ЋeO����Z�[��V����O��?��?|!��7�蓯^.G��d6�гI�0خ���1Spc��(4j~������)��/�uR7����}D#[ӹ(SS��O��JRY���f�����TH��Y��2��ŘP� #s!B�ps�2Maԇ�N)���|MY	�@L&3?ф*G�	���C�[6`�g�YJ*��=��a�ז�a��R�K�O�^����bA�Tq��d��:F&����~L=�]g�1��!A�FŌ ��2�33����;A�� ��E�À���,�������#�9��T�ZVF_4Q����0=�t�9�D��3�9�l�{4�oBߊ@(tW][^�X�7�RY���f+M� YR�d�R�1L0@��� !dY��0��/Gֆ\��NE�q�V�st`g�
��2�~rue_��7ڌ��6c�͖�v���r
��tYM����/���)��`B~ QN
��{�P�5AAX c��$��$Tv����dj�� �Ei�B�J)\��\��N�*0���F�!����2�Z�i�c+�nE��d3�I9oVo؆uDPg|#%ރB���/|�������O�������y>��������M���v��v׈��sS�F���F��E,�.�O�TE�7YƢ%�J����#{��$����GV���ۂX*E��f;�c9!�h��@"�[=26�W�T(a�h@R��+)(]���#�#���[r2��~�6"'(=�oߥ
u�[�샒(�����ݺ�K	e����(?T�ǄU}��ߧ�dpd���̢Dܿ����Æ����Wv���S�^�����0�PY�/�*�H�M�3!�P5���(�e���c*�.������RI��f�/�h�re�����[,���]��&�\�M�Ǡ�i��I%�d��M�f�oԶ�b�����{����F��=A6��=�;�rv�Z���Y��?�/}�5ѯ�N����X���0���D�~����v���0�Iz�
n���<~�s��.9��aZ�ĳ��W�K+���mO���Tʼ(��ѭh�|�f˕�'�>#L��5�T(9 �a��S��9�r�m�B�η+{4�·��$.6�r���m���������������/(���;/��xk2�go�n
}[�3*������`b�'[և	�H�Mj�
�$`�������FѰVɦ�/������G�,J٢�|�<%�ƴ��.d\xR���$����b��f�E��t'&�����2��]��2�l�|��F�#�K��)�_%Ys2���I�.�I��{�/ é���wz�[�����c��11r��FL���馂�������DD�W6Ϥd�W�x�&ʰ5.ML��0���/�$"�ANIr��o�L��{Pp(i�����Y���n���#HH2Z�aȚ�/xWe&nV��!`ʤ��/�[�[A�3�* z��= R����֜��k�{G�Z�9�w�q(l����?@��A�f�����ݽu�̾��2��p�ҷP��f�:-��ւzV)�2������n�)\Q�k?�8"��(cCz�����B�[��j�%�,��%�(\��g�;d8���(S\O����봿B�l��C;�{�N�ݷ�ѱ�k%{�Y�듮=�Om �)e�TypnY��ڟ���/��/~�#�y!��7?��W/'�_s���G��
B���F��i��m���-��-PO���
�HpK����M��ϣ!@��e��UG���2'�ӗS?��D��F��5���A5MR#�dv�M��/JMACd|���J�W�@��썬M=92�(i	r S#��� DR�5ٜ	���Xh��-�T���� �kHs��0dW^����]������,����CD���|r ) �9]��	�ͼ20��GqJ� Á#�϶���இV�ы��J�!ƗT�Bz�CA�E�x����Y�K��;�E�R�"������y<&���w<e6����g�K[�a]�,?^h�����c�F����Ȼ17%Y.��M��D����H1ꓬ2*���K��T���JI�~���|��Y��ʲ��K���[�Α���+������Y�À�f �%-Wk�n�}��NFI�J�ddx,ā���5��^4�j���ߥ߆����6{9[ =���X4TK�.�	6�����<x`�<��ɱ�j{���k���5Xo��1�&�=���f�Ŋ�|x����=������(������\}��Q�p�����X�h��ܜc��d��$��P �:�}
^��C�;5�=�Q�e<�J7�@2�T�@�D�6B�2EY�r4�r��ϸ��&�p��x��@����9�K�J�CG�%�a�"
X0#8����)K���^�$�c ��-���o^	��I�S~-SIO���cD�, �0�`0 +z���@G�p���C��J#�� ��i
�d|��N �0Pa3���7ǐ!��hU�V�����+dw�H�)m�H�u<!'�8����3��1�j?��N�M��ӂ6ٙ>qE�O,�ۦ?ѿ������𪨖���g���'�� �2�q�J(Uܣ#��0[*�lΎ�-	MP>wC��zn�L3IR������=;99RFz~~n������BrLR�az�l��񉵡P!Ǿ\��͍]���@y�~@`�]!�����tj���2'g�`&c$��&S�<	s��Ғ���|C2�m�>�8�SD���������U�[?����=���|1�������̟��y~/����;:�y�×~�>���b2��|���r�ko�	nE��P�-�_�빵�Z�l�p��Cq� �9���j����0^���}�C��
/�Iu�#�/�X����k�e�����k
~����T:���Q��Bdd�Ѳ�n+N���uRG�z��/ԁ;�o2�ݮ�`HMk�?���x�,/�g�l�����P捃"��z��������h��,:�t=3cahV``ӳ�чK��ޏ��� a�R0�O�*&�L�f�$w/[��M��9AL$���-xB �֭3�I��>>�7���&���P9���Α~��Mwd���2��m���W�0���0��d��A��^�R���k�rCf	E��&���֮Vի&�R�[�m��"u�/K���7Z= e��<��T�5CFȄ�Ѵ��S;>�h�cC�׵>�}�� 3 [V~�AQ���:P�08�S�� ��K����0����@'NԲ�.X]V[-�޵��^����ttd�r�ΗS{6ؓi���S�Y�/1�JinknG�W��c(��]�g�Jp{<(�!)�@}p;���:������� ���OY�hF[/+�@b����Y���W;<��z/�T�$��())v�M�(�vt-ֆ�A�P�e��C${ �zn!���i�
J�C[�O�@��aL��EI.��ن��������a ���P2�=0=��x�~=,���tbs�Ѣ̕�2�8��=s�Sߚ��kk=�F����WG��~M�\�ط�c���'�4f��I���R�4Q�F�d#�\�x��D����$��'������u����dJ��c	dӅ���zL��F    IDAT`��X��Gp��H���v�"��#��%����3L��}TE☂��|%g�� �U�T�y�-�awF֚5�mȈU2^\\�u���[�	�Ea�igwN�谣�u}��i�1�WK���eEY�+x%z�PV�������Ԟ��O&�Tk���	bȃ�/�wP�P���V@Y�ӱ�{vrv��Z��%y�����'#�'������"��l�Ke{�� (@׿���ҏ������ЯnϦ�_{4���'�a�i�~p�H�hO�/N_�K�� ���9�4ߔ�ikR�*�p�����V�~�H�
P,8�)�fz&�)�����ɣ��[ʺ$%_Bc�&���4��t,`($pU#�C�D^F�[ew/�\��7g��Sf��	�ɵՎt[�r�P���	��58y���i4ޓJ��25��4��+�����W�ha>��y�r�{D� 4zdcSV�̇{	�S�̃�Rbh�)�y����F5���xj�\32���P���{��g�er8�������~��0&3[�V��l����g���򓥰oL�ד�O���` �����y��=JxϤ��32I�S�� h8Ƚ��a�}��AL���\�~�s4� ���vm4xƕͨ����֮���c�F[H�n�,�119 Yg��]���v�R��ܸL9$��z�r(�)���$6��g�ϭ{�����֦�-��(X1q%�-��}ܱ��3;<�gͣ��Z-[Vkvc+��4��q��g#�o�(f�����T����?����?������ŉ�U�|�����ӯ<���ڛ��|:킛����M�enj߉,�[�#p<ʔ����"8!<e"��&�66=����rP�A�C��0��0�����XNդ�F CxP;)�(��։���8 ��큉�@�bDPk{�RpS��$}�G�$<�18��y�TVx�IŃ�ۙ�Y^M����;�Ԫ�s+=�2c^b�qL��*=�iR�+r�pLa�Wi#C����۾nb���)� X�w'�ZSɤ ��
�Y$�܄#�End(�ЬN���O�-�Q�B����M��h��F�� Kì{Fp�زӅe�#�3��?��'(K'��ď�1:����g�$>��A��
�a	e������4�`X@EvG��|>SV'�Q8��|:�
$`���P3�ʑ9�j>Z.hJ�bϊ�5���:=�ć��\Q�!�&��Õ��J�����xBD��z�S�V�c���
n��#�.�?ۥ������.�c2tTb��&�����o���=ǧ?��/

����W��|��l����R?�������#�E�����M�N�36`��>�[��4T�*�_n"��䖠���CT·2&��g	t��}�?n�
dQ��yY�Z`^��SH��E�zr��v�+b����Q�zv%��r�0�^�M�ސ,߹�{�)�M}�o/K�/M;I뺹��~�*	*��	����0��*Ch3�⑲��#?��ߋ����E)K�A�2D`$�E�q?��	����9�ESW�M*R)�=6��|#���$o)
7&�5��l"��E��k7�]Y��,��Ta|��������K�L"�M�-I]�m��7��]��E�'s$z�L{�
I�h�,�g�M ΋��&CM@9�aE�_����-�ܰ�9"�x�B��:��Rÿ^��#en2��d4,�����L��4%��;/��[��x:��S��^V*I��,y5����ٰz�m͓;��@�-�h��reW˙=���gOg#�ZOm�y��V�d��
� _x���g~��|�S��R�*���������W�^�����DY:W:�t��6Cß7��m��ir���n���WHMYN�q;��\
!a����L}2��ঞI�����������5�T�:K�\������xRe)p3�M0���4�&*UC$9�{m�BQ�(c��~���(f��>Ѓ[� �i�l�BK.���UC<`2�c!��/��1�K'bg6���e�⇫�Ͱa["%�G !�}�64v��� �ei��S�[�Ȓn
,]N��mTv)�>֔7��^�7Я�À�H�m�d�SJB&��bX(
���l��ۺ7�md+&��KaS%�G�]&����;��rt;5#�
�p��bރ��2ޔ ,��T���w;_JVH~FVG��S�)O��5�{���J��mIc �P�0� ��늲�x�~[��SI�k�)�A�pv��2i-��������JJ�b�=��I�ri�RQ�4�[�^��ё�[��c�:W��Od��|6�g+(�2k)*ӗ<���\Cf�/�:�������-���?���G�ޯ�9���n�Trߡ��Z��o��s��T���dr�ҍM��۔q����$�T��x�!������O�F*�U#�$�K)�s�"�ȧi*Mէ�X�LAP��!k$��7\�nI_>�]*y�9F�*�H0p>Jl��I��5����_wR�H�k7,��,��$e:�R>�{Ġ 靥�F	��~�82��� �F I�V��A[�r���m4_��qܙ��1Ō�Ab�(���E�JYI�� �8�H�>��.�n^�*�	�6�r��	^��r�M粞]�܂���=�(N�#1��^�M? !#���P��ɻ��[�"��3<
���$,a�o������g�s����'h����\��	�����q���U2n��EP���t�@����|I�O@�</��ڰ׷^��&dn�dvx2@�*x'0Ը��Ppc��\ �s{�7�d�Z��p�sh���Vm���|=]��rf�2����n0��.l�Y��>�V��Pp{���ً��O��������Ëi�W���i�$���.��-����~��d#���E�F�%zE���x
B��+c��I�׳�T��hJ���>�,Nv%/��JM��T~
��7 $i��gQj
C}9���kK,4Up]즭~���0z��JT,�8S
V��{������2��}�� ��$LT��s6a6��C�U�[�T�z�l㛞��S�G��.W���n�l�v���34�.][��㣦�NHx7�^�X<�yL��<�����D"�@�wԳ��y^pt�� 4�߻\+�����%]_5�j��f2���M�{ܠb�`�8S9+!UI�ϝ[��5�������:��A;��{��`bZ�ս�>�����]扽 X�C�V�9)�9�A� ��^���+�1!B���K�Ddٸn�6��1Vv�z_G�ݖ/A.ABFӱ]����C98q[uk7�R!�$St��U�:ֹ���R��|i��=�m���8����j9��z�!��A�b��m��l���j�������*	��G_sY������'�����#OF��(�QpK
	�CYJ=��m�~�pQdr\Ь ��2�
:���ښ{����B�!M�H���*NW?eCH
���Tj� ����� R�Ie[Z�*-�L".�^�
�������~�{``�y<��4L�,�׬׸���=&�v���-25zx�tB��a%!D���	�nO���֮�*�1Ӧ�vm�S9�?�Xg�R�}�_g�æ��|ص�vc��̃[���ߢWSM���~�a�B@3�����PB�Hel�x*�^��d�B�J��Lsyk���;�����۔�|�������f݁�)K	�;�3�ZH$q�90�͞�{2�Z�{��i(� K�j��%a��͢��o����	'���1 \'��q��]�>��IՖ�C�*h	A�>���l��.���J�[m�z��Q��m6��{ջ�Nk�>�2�Z�ڈ#(AS�g�j�'�89�e6cד����v9�,���������d�V�u05�%;���A���W����o���-%�=�����COǽ��p�,�* ᝋ&�<AL����t���I=��փ[��i2�_~�[
h�i}Z��d75��n�zg�kx��㱪]#�2��6�oʦR�K�\|��2�·a��!)�iZ�T5d�yF�5t�����օ���	�*{/c��!��qz��j쥶^g�X
��{���+O��f}j��D�Ѳ:ÄMƮ��ۼ��އR�!:Wf־�N^y`�;
n��º˩M9gd�R�^kL	`�oJ}Np�5�K�䧑�"�r�ا�! D�t�_��y��x&�ۚ5e�p�ؘ)�Mz}[Ƕ��6����3M%��Wy�������:��;0v��NÜ���=Ā��$q �2ة�h �t5N(�F_U�И��R�gq���MS�f�a��*����/	v�2%�@���4�n���Y����[?�P�O��Ԇە�Xd���U�Vi5�ztl�F�F�݌�v3�Xo>��0���va��ږ��!J�J�sk4>�j��'~����EAA~畧��y<����7���
� A�W�R�IF�%���5Q&Ɖ��%��d��H2i�:\B*/��8%L�܉9N,�K����dS�nR�
�"��E�}7p�Ϣ,�d �-�P��`3 �+��s���+�������G�9{�/e\)�'K�JV<��*�e���҈甅�� "��;�}�M额v��o��g�?���94�[*y ���[u{����W^�gî]���[�T�
�/�M ���A[&&�׀�DpSi��};h`-�̞ W
^��J6�f���Fl�029�xpb�Pɸ�q���?c-�j8� �@���i%n$܀
Iՙ���w��4tJ�-	$4@�2�uJ��V�ϱs���������[j�x���&��9!�L#r�=��z�L�*>� Cb�t�]0$�>
�({��hZ� �r�9
�2-��P�m�R����B)�@��eq-+l���K&o���&�� ��m��H�����A��5kf���f?�r��c?�-��b���],��x���g�~�G�b�����E��[Men,<���wҼw����7��>��UHنP�܈��5G0�}����[E�ԫ�j�%
h�^�R�,������/9ky�J%�"
<
���hW>�Po�	2r8E�I�
�L��TS0ڕ�އ�r*���)�y�+�y�%���;������[���7ްg1��sx�)�l0����+��N-�DJ=��`JCY �bƬZ�w~���޻�aO7j_��6��������x�fn�Ep�7e�E5���6�26̰Ke�
�NBG��B�^5�+.{76��-�'��\
J�e9��4��RwA�rz�W��>`��'��%]E�)����^�G! *�	��W���.kۓ�O�i��A�U4�ZG/O�<����C�8Ӵ<��1��@M7���$�b��j��X�_��&[Ԥ  �V�\���
ʋ�Mfc�OFn.����R��f�"�u���l7-S-)����[�ٲ�vm��º��)y�Qi���ɱ�ZVYe,?��n��?�?�bd��s��M������^��F�6�IB?�b�l���m�u<T�D(��L=͗$P�{�H/� f�����'=��
H=*Np�jᵰ���V]�2=1I�$��$.=N��H�|����`,8�b3����1L^�M��Ty������{�l�[#CM���x���Lտ�y�pPye"�'/���M��˯��[�
@�t%���2���㛾A������|:����F���fD�������RM�[�Ӝ��}Dm�(�)�����r	rx���@�G
n���U��	n$4������uW��Փ1-�v�j+`�~��6���2���uS�T�����u� �ϝ��&g3t���o|�F��t�%�cQ6�1H
x�Jo�n�w��t�%P<�������:�L��VRx�
���G��,G�^�[�y���v�pk��E8ܔ*^�f�,[�Y��A�օ�]ͦv��ëR�����bbS���l�٪��ɩ���M>�R��џ��|12���O��b���Ǔ��=��sdnhrQ�y	��P������_n�
N�(�^��(m��)��B��WIF���?�Ʉ��Ʀ� #Y��)hi��4e'���̉�WC�O;&t+7�������	iiJ?��r&�Nl1�)�'l^*w�4MִyR�&6�A��,�^[�:z�hP��ƓPg�����*�,�N�@�ψ�GOlxy))ut�(3��	۫X������y徕Z��'v���w2�nm�����)�ݲn^:9)^m9׉s}0�j*{A�U��k੟9�{P(�X��G��l�H̡F/�=���#??=:RpcZz���M.���2	���t.��t�PYN�A �RP���^�hX!��H��g
X�.���!֩�����!�W!G'��[���q�	C�8�7���c	mϯ�'���7�2��jN�"�����}�̍���nWU��2�f�d%�0����u��W��T?2���Zm�u:�b��ZhŴ}�3���Rk>n�,͢4�\��+G�~���C�����k�����|��t��'��w?���fQJ���Ά�	�̋�
��tv<������x܅�<�qs勉�J(�J�(���֌O735g�i��#�����N��\V��)=�N]� ބs��>̇(G�4���ޔ��v�-��{z�{��
h{f2B;)�F����6̓�t�-��u�:F���ʦ�GP�4N��\kT% �V29�?�����+�zͥ{Tq*�[�����mTm�^؟�����k�2��,m�����
�n��B��� �!�����$t�j`k� �1��0�~L�)M��&In�݀����-@���{��g�#��Ս=���/�%)�:!�-�S]��~F�^��Ñ�сA�W�R%;�r��?HJ���#�r1�N�BE��iT&�jd5	иX�>�a�=��&�̮�ۋV�����/��$��d�!�~�%���x�ڣy24�����T�f�-/��YP�`����ʝ+�,�l����F��e��C�������*U,7_Y�P����?�/�����B
�������?����'�^��Ȱ��&3~���hօ��p7J�@n#G��{�FE5����J#�D�ִt��������H.g�$�)~귥SQ��]��L�x��H�(���$���,e]���T@��̌~�9��o���B4�JB�I�b�����X}�R@S�>a�$}[(m��t�o3֩7��PFӣT�m>�$ �����N_�ow��P��'7�v1�[�PpKe邀_D�l���J٢��/�*��-|+e���u�t����pu~)��K=*�5\-1��erOƕ�
'���	e�SE�
[>��{��*C��]�~zn�~���� ��kB�c�xC�.�ے	w�Qq�b�>�#c��k���g���4ݩ�DT���^����N#5?�<$�K=�[N��7�zB�Zv�*����)�K��$1.Ր��H�s��%��ALv��Nk��h(�"?_��"��Hнb��m�%�2@e` �&r�y7eF֪�/��F��yt���m�/m��ci���=7�X�ҭ\չ'��,���Z��D�暆m�-3ˤl@0d�h�$�)���_�P�,j��@n��ӱr�7�l<�9���ޡ��htw�[�}�s~�������dnn���6�
n%U#;N��kn7�c��n�:��4a�i�I�YeF�Rѯ�����Og��1���]���ݛ��؟sS��i�-��|����ćQ>Ǫ��� 7��~7�aXN��#��5��nJrn�z���� ��B��Z���������є=X½;�%�i�rfTB�[^+K�d4�l$.?i���,������TI�N<�`]h��B����nW��߷׃x<�,,��/��47�Es�G�]3`������A� ��4�q>�܄�9�l��J�F��.��ں/�6'3*d��T0";�f��z��~�0��<Up����1�s�'����4*�A�kXf�\{��w�e+���g"sr�t����@õm����S    IDATu����V����m�m����e���T�N7תpC�=!�2��Zo���;@5�����j#�n5J�� �1�Zi{�mX)Nb�bVghc&8Fբ`&��i�%��1Ml��-��o~��?��W�uZ�w�(�գF�[��?b�8�V��UARt2���HQ#���� Es�ce��T�����a��θ��Z���<	����љ�z�ne��Ȍ�43�k�������I^��6����9�@�fN�W�hvp�b��.ke�.���쳘7�g>C�, f���j���zMLxJ�JZ�g85���Ws8B&�Р��E1R^7{[d&�nդYI��	9]�9$8����+�I���s3���E.�����L����vg(��z�]���G��Ե���Ԕ&���A�g� ��
Z����z6�&xk��i�
l=�L<��t�xi���p��2���r53
����a����ʬ7�Z��px�P0f��c�o�7Nފ�E��0��i�8�G��p�q�Ѥs,el��O5}��'�5�zy� cpS/Ӫ�8��37�bq�=4��Ng*��H���2�)C��@�<31�\��L��H }�Ӏ9�C/�Rae���$��N4�Qoݔ�DD��1��-��������)K�����I������_;��(����nx��r�ǒQIR3�	E�udt��Nd�qb���B�s����LG�pm#u2s���M73P0��27��?8��vJ�R?n�/��it�<��1�uC��Qj�@�m�K�H�#n4-`��X�������}�U�}��1nO�S^I����y�⣸e91f�i���JT�!���"X�_���"V�E�>�8�	[Ĺ�<(��
pa޿s�������#琐�����!��Y���JHf�T�}�����c.ԣsRo�9�f����0�*�:�*2v�qpq�멒��aƐj�Ny��E��Y�yҒjG��nO�/�39B=d����j���j#�#l�g�V�ku�ԑ��u�b �
N�uuk\� ��֕m�;��R��nܣu����pT&Ƚ��q������8��֟1���ﱛ�OVNZ�V�NL:�.!�N�_�C;�N�#ax�a���+��C>c!�cAD���|�:)r܇H����xj����/�~��'_�|����d`����
���76N[��W�����W!ZR�"�,��h�V�	K��`D����6�S��5��tL�f.�y=�)�ص;*���ocf�9�\p��vp�Y~i
g�����8��ր����;�6�T��I7jbq��3a"H96�t���eb��v�W�ݬ�8'Γ��J�1y�5��4M�� !S�hW,������7n����������#<�|�ݣ�h�W�7�b5����G��_� ������ZkkkX[[��Ң|+y�1��
���q���{x���`G�Nꖦ�:����Y-~^�(HVq�H�R���������ݦ��b��&��NmVYvG�g�"|�֧��{H�xI��$�떂�֑J�M�Z���)�*�YN o����Q�����LVu���\TAXe� �]�v�I58J�Ś��������u�;�3)��_�e��DB��b���rf��t�v@b~��z�{n��x�Ԍ�I�J�����6��D0�ԋ#F1I�>]0�^)9�7?��
��|<ux{>�������Y����ܨ
r9l��;�˟>�\�ʜ�t�w�~�=�x2� ���x'0���<Ỷa��Lps���ƛ��fu�;���(�ܿ��މ����dCU�-	��o��Z��0!��\�����++͂�\AG��=,7%����SX��D�fhܮ���4�k��Y�!FE�<>�^���ept�2]1,,o�#�����)�b}qo߽�w�z���x��9��|�
I�T1��f6��O���2=�R��ǏQ<����{ｇ����x�ݞ�I��B-~�/�0z���Ϸ_`�`_�^���;X��G&�4�4�?%U�>\H�����x�_<�a���g���:� <"K��h��B�5"��z�J��l�A_|Kfx� H�cp�|��X�8��D��ϑ~7ܴ�&��F��7�gs�����.��+
�D����}��X.���3њ�u"s�#lt�j�3��n�3�-�M]��  ��c� �>s����G��Ǩ.�#��epQXa$TE*�4��^������� �������_�5��|���
~���_>���E��;;�˟�/_F����o��l�n�-K��$�܈OkS�M�܌|x���N������J?ʞ�����{��b�����p<�p@Z��+�6�p<��)�p@��P3��/nqO0+�I�bv��	����Y�B���B�u(�j��&(aԩJ��a������}���xR�����8�)�Ǐ�`#n-��ޭ;x��q|z�gۛx��)l�[�={c���_�q,��y��dST��/��|�3���;�S�(��M#�8��f�AK�"������M�pgm�x
�~O���ZU��G�p�S9#g���o���Ml_��U����mb�M�9����N�ҩ6�`�VwL����E�R�0�P*���3�9�ǤP�[:h�����!
6j\�\�7�P�����!��E{x�{y�[�;tݞp��5c��mš6�N.C�ai�������1���M�h�5$��K�p�h�X�x����a<PU��<�W��hL��oBw$��d`��߯ඐJܚ[����Ƃ�e���+W��[�'0��q�@�K2����8�u9����L�z���R�����5ї�p��)8ܜ��d �|�I��}����zeN`���ǲ�*����	B�9&�O�|,9���.��6v
.����{������dO���F=�Qʴ����dx��3S��qoeC����}'g*K?|�
.�A_pn�?��쬂���eB���߿���e���c��j��$m���cX�XW3�(��/�X7W���g���>�W�jT%��EE��������#�ℾ��K��X.L��8��F`ꖙXSR�-ܜ�%���rU�p���s�-���\�䂝*@w�'@'\)�Ke��*]9)�)u]W���i�:�I��+�'׹�Z�0��L?�|����a�j�H����j�wz�U�Z�3�DB��	*�I����<���n�}z���y�~PIJN��x�H��ȧ�{w�W~�s���җ�����dp�wY�/{�Y������ՊQfn�J��&���z��2	Er����6����d�7#k��=%ո1>Z�3� >�˵o���JVW�1����LНTZ�Nr��K;��`��q�zǎFi�D�5&�4�@�^�Q��7*n�����!̯7�48����pM��ND�WV��e��:L���1D�}����<L��d�#�<D�v7�����?��;�e�ɋgx��ʭ���Bͯ\"�Ͼ���!Ev�n
=���C~q�^GW���Gb��D��$�-@�w~~���4�J�8���n��k�����|��JU�?�ហc��̴6�����x���sM�4���@�3$l�sY�]�ڑ֌c��?�vk�<C@D��"�t=�QN}&������̙m��(Z�e�Xf�d�!��0�#l�Sp�0�q�c2s3��P�Ȋ{c̠�Ƹ)Ks�U�^&HP��"�5CA�� ���h������"�1�1s�&"
l�0͂�s��54��ό� ahR��&�45�����[�����7"V��<����v���+�?w\/��s�[ĸ��e)�8375�%Zi
�,epsP��{g�e�Q�M(��Mq�9��uٞ+��z�=���O�j*Wl�T�`�\L����YR1����S�Yj
]㒤	Ԅ�_�-L�פ�Ƅ��Ny�����{t}�!{��F��@��@��)-�S:�X�H��a��$���t�������{�n�F�\��-<|������2)ٯM'����|w����;O6EUʤ2��R��x��<�{�3�MM��#�Z���Q�N��W�9�YY�[�uty��}��Q��|�сc_L� :3�}�]^]��N�?k�֏�Zݚ�Y%NK�l��M��^��?�5�nX��8�˪M�z�NHV2���Zq��n蠃O��3 ��>\W�Z���� ���a��C֖�nR�CB�њ�[����5��6	$v|m~�Nr� jl|�԰�{�k���j��g�F�n8�Q�`� |Q���(�N~)��o��m$���L�R��I�L�<�9��w����ʷ?%Q��O}ߙ�����g����S��/��x��6�}��e�#3-MF��2s�Ӽh�~���Czl4����O�1���� ��>����ZX�g'�rڴ�e]���(��tSI-..���t6��IMv}>=*S(��_%�I��b �	븟*-��ev�_� �G��I����Mt�Z��	UWȩ�O{,n�����:ˀ�ЋHX�����zoݾ/������}��/���p�/~�sX�]B|��������8Vnn�6���1���w�[�T�bC�(��&)�;=��ǝ�e��~wo���;���7>����#�	?ⴇ84��aƾ���`=Nݺ���el�JC�;)�0��6087+H�������E���PMb]#�>�3���m�L?�\�;�Q��2�٫>��3���긥"$���yMŠ�N3#�L���pu�[n� �@�Vq�-{r߫�V����|�:�|񈙐��R�Q���3ȱ
�СO���	?�+>�I� ��1��������_����?�����N��V/��Q��,%މ=-e7C�C�s#z��.����cIS�p��q��eT�ҁ`πs|��0�ܒa6hjey4��0���k��+'�=A�湮�n�[<����i�;�ܩ�Ǝo�j��,l�.�~��N��&&���A�n��b�*(
�F�c�Ĺr�~��?a��<˭>Dh��)����w��ݷ5���%���!*��zf��yF�Ke����n�-#?ζ�,���omH���������~�,Q�a����Az<v�Hz|�5��;�k��qC��R·�>R`<��P��u7談�Jr����ٍ���!'+B���8\pp[��_��8�1�1�&�sS��k �n�mH�G]4�/\�Ck��cu����f�)��*��ǵh�����Dn�3[B�C���FL6iA�6�������>��jv]����g[B��ʘ�@J�y�(d��(Ti��%X�5Ì-H/}���cCp��xM1L�z�#����?��T����7�o|�F�3��F���
��i���	�fn��)h�[4Z�72��$H�G&�qK�gA��_��iw��X,݄^1^�*�O/J��;Ь߀'Ǵ�	�N>"�]&����0=6'�uN�������zꝍ{w��'7'5d� �|��k�o{z�KlW�ڛ��WNm��;9(�W{B;�~9n$�z"�j/ ����@o��W��ͻx��=e���{���C\U+z�N� �7|�s?�;�� ��n��J073�b���ǻ��'��@�?��nN��@��Al�E����n-���;�tOO�W��㏰[��9}-��e�ݽ���}Yǻ��t�_N�N"�}��Ϝx��������/co룠[{?��a����S�0���={���������Wz�t-�k�P�l��w���;�,�ϭ;D�D�'���d�$ߏ�^(�.�
��&-6�9H�+���p��q�3�G�xI���U���ƞ���"NI)�"O"O@т�Ef���^7J�����������}�������?��oF����e�z�_���17)��N5.Fϻ�m2��M�Ր5�Dp�<�\��iN��ȕe)Og�+�?)/�J��ӑ׉h�)���nd.�R鯙r��Mu����9-;W�^8����ZD���M��M9|M�r�	P�bǋq2X
�b6���i��f63��m'xƳ���f�݁����Kx��=�w�-����5�4�& 75�Յ%����iqA�_�
�C'����Z��է���E'�R%$K�>�@�> :!�	`cfN���zWW|rq��~�-��QAM9k��F���\����tDs�?bݐiVc�ܺbc�G�+Q����n�,�(ee��I�e�u-Mam6g��Tu=S�'U~�qA9�@����3��{ߥȤ���p7��q�T����w%��UI��E4���K��\�z�r@F_p���'��F�V�26VK��sC.v��[�hP � �(�W��CU>3��H33s���a���P)��j(���ͦ���P�@�1�n�W����?�fzn���/�j���W+��n칑8Ͻ�2$7-�g�J�Eo�S�&)h�(Hȿ�3��-}}cN=wB�Ū�5�D�*@����-���;�{�������^�u"'p2Ⱦ�3���il낙�&���g{fщ����TA��&����X�3nnwO�\	��(�X3�����GA&�nN��7L�F����9?{���s�'c1�^����Ul��!��[o�x{_ާ�H��s8.�xo��c��E���xk��Ã�:o��@g��lwV7�#ｏ�׏��s|����A�M��1��6�0�Q�ϡ2,qp�$�"�<�0�O��cX��F�x���>'s$���)�v9\��t�MY����$C�*9���4�7NE�I������,kf����(�U�qkV�P�Sv�����=c��p�M0��$�F�@�a�f�d��>F4Ͷ�ٔ��Ma������5��-C4���i�J����� ��h$�����ssy���#9;�B����S\������{nӱ8fB1���On�-��nG���:bp�4b���X]����~�lJ�+�N`��Gi����B��I��r��mrń	�x�e����fr3�a+�ZP�d�t]��z{�AcYb����<���r�ؼ���(�s�����^�k&[m57g�<A���k�5�)w��O-�;$oc�����1�q��c�
���`7<�|�ffpoq�Wo �)�<99���)
�W2 �X]��ħs
�J[O^h���`~q�Z[G���qٮ��1{.�����;��~���I�Z^�۷�J���p��~�8�:G�7�K�x(�I�����'�KaܸI5�&��cZ&�Ym8����v0�p������$O5�	iy��60볒G�I��~�>2ofp���`Ь1r�L��&��,��|�`0��J�O�F��+�0�k���4W<7F��df(�bK����������!��BQj�L�K�U�A��DA˨��\�d�ك%v��Š�xT��*�J!'�����4��s�B��Vq|q�B�
д�o�+D'�z}��&��F"�7f�~�����f���ou�[���V��&sk3h8bf_x��2����j�I1�1	we��V��
�.۲�W�W67w�|��pCgv��;W�!�+=u�-��5v��F�M~m���I�c���^��iw�6��x���WH�&�2�M:I`�(M�&"��2�f���7r�g2>�@T���{���븯�:��!8Ԓ�	<�G������i������:n�.	)>�uP8�@�P� �K#5=�z����c�)s#u���t�}�����+E�;M�������7ـϏ�����lV��T4���=�/��qY���ƐŰ���X.o2��{ؿ:;���A��iA�su=-��fC�� �0�i�kYe��l�'�G��2v<�t��v��>�%����L:��כ
�Z[�X��7�
�Lp4��y�T�&�D�q<��~IIџD��jU�a�FPu$�^�fx����B�P�4������A
���N6�v�:�鷒�����	�(��2Li/�����}�)�cQ$�2
n�a�|>1�4\�EQ�Pl�Q�Ք�y���5i}	��F�>Y�������_�� ���C    IDAT3���k�}ܬ��a���<h�M^�q�����L�4�9�R:x"�D�77�O&-�QnE��Z��Q���c]��Ԕ@�\6�-vG:Z��G�s  �^'2�n{\��)�z�񹀬A����`�=&���A� V*���� _��:��o|����O��׽C3�5����Y��*Q5淧����I�A���V0{�����|XHM���*�-�b}*��/$��V�(���\U '@ؿ�8)������+��yun�oݑ����gg*Cj��2�H(�T6��D>���w��j�$Ú����4�M����˃]�.�
�#qu�����xxt��'���>9�jt��!
Z`��n��*��&���Y�ç�2t� y�m�4I��+�d-�@RJVR���aP�:O��@�Z3��}��A��I��} ط"^���v�/�v��C��Х��5{k�i�-U?���#iOg6͝w)3~C{4��0�(�XLXS��&�v���<
v�m!�M�Y�@eXNWa0+eB�
����Wl��s�lZ����
�^K�{����@b��� �pȠ+x�x<R��Ɠ𴚈�<H�}O6rs���A�o���{����I�����V-VBb�.���xB�'�	c�F��G�^.s���ƾ�QV}%�	"d�a�`e�,m����]{z��E��˻�45�дb�R�$1Ϳ�.��^W����'�g��8�n=x���5�:F�S},�aޏ	B��.ss�����=Yc_.(@��E�J�r,�h� ���{]� m�u�j�"v��@`��̣7@��G�F>����<n�,cij�@X�pNL�^��:v��u�����ܴ$��,� �g�h�u�{�Ⱦ�w$EkЕ�Ь��>��~��YI*�L}Q��E��5%�X���QA�<�C��ώ��2����{�b�0#a�Mz�e(H��i��sV�k2�1X(����LY�͹�q�YZ�����VHb"u���t=���A�f<|}^'36�@$S)��9��t�����ۢ�5秒�`��tW�����V�4m	�>2׍���S�x&� �l�Qi6����۩���v`B��I�v�G�P�Ϩ~�5j���xM�$�6V��Fi�c���~?*�=j/K`<�I:~�W)#��#<�3��K�?>���<��}c�S��G��Ϟ���p�(��B�nD�3��$\��
e_�,��%Vi<�����[��5�dMnx:ܸ�Ͷ��Q�7�S�|Be��d�#k��}��LL�'��5P�	21z�`�����P�9�O^�	`��.G�c����*�p�Df6���D�q-'�ᦹcr���n�eO�qiQ��~��T����	��1Ka=����e,M�"�K �e���1��p\:G�Q�k:���S�|fV�hʌ+� `�����q^����)��x�M��oci����M+8R]���'f7�h�͢T@�mb��@��LJ�}L(��}�����<̴8�� x���s6s\Tez�K̒�b�Ɣ)��1�0p���5`��o�PTY��I�o�|�x@�rYL�rʠZ�"���,��=-��8����w�g��h ���0y��@*&ʐ���~��$ܧSD�It=�j5�DqX�5�QN��+����b�I93��=e���^�.Հ^̮-#���N�+�=�l�����k���j�A��?�� ��D��]^�ۍ���o���O���9nU~�Y���r���D�O�M�H
���(3�Lc�a���讧|�%�&�� ���ds��WP��&�6~Iz0�2���=��0H�|���izn��cl�-�^n�S��^~�ei
�f�`�f� 	�k��8+t��l��ۡk���W%�a!/NY�&�\Vfb{���Y�z��\f(����X��{#�KH����X+�y���S�yG�::��y���װ����`��46��6�����bi���(1l Z�uZ�=>T��r$N/3���y�^]W�cp�]���0�tL"�~�h�v�}v��fU�4��pj�gJL�k+���H�?35�H`�ӤT"�VA���;}5�ō��V��IƳlで��(k�P-��G��
��K��m�'�5(�MT>�������B^���h��F���y�� 1�9�AUr��F��	��V�I�� |>�Mz�R���X񩴔��
�J��LV�@�e��ϒ�!�J(���J��K����Џ3�e��� ���ߺ�A<����YG#@�=F�#����փl��A���?D��'��V�7~짾�i�����W4e>�V��q��S��Z�:����fn,K��'
��2���[��prv00�`1C��u�*p�D��2��@X��)_��Υ�B�����>N���	�e|��Th�NK_�a:��0������a�(���+G�Ӗ	�n��3�V.�)Of��9i%~#�6�9+86��taqV��&��q�jy�*���������Y8`x�93R�Ng�W���q�
�g'��z�q�ډE�7�L<����SY�'s���$w�����E��m�~\���m�Z��Pm���:6�KRP�4Z��F��?
�����Lj:�x��������>hcD�&��R���R�WC�H��T�r>��-:��V�q]�P3�` � �V[4ŋK��>D�Ĵ{�6!�^�/-bvauz|Vk�wZ
h,I;���=Y��<�x�)64��02D��+Z�>��Y~)9���p��)�8a.T�(7�h���Þ���tp+�Ʉ�������R�A��K��}�u�W���XC?D���UG��\��l;��>JN�)9E��H�8��w�V��o|�o|�����76�;�t�*�M���+9翬�F�?sp���ۈ�h�U������K�I�K=W.NH���Aӓ��±n��*s�b�H����Š��=x˱�i�p:pn2'a�rL��D+-r\�'�3������i��	"��ǌ�I�Og3=M�$XіX6�Pvh�o��\p��kN����G�?��4
���(+���S��5NT� ��K�!fN<��a꣎>G��6oo(Hɔ?�\ ��hFx�T$&:A�R�N�FU~
ln�o(|�Ǉ��9,�,�Ԍ��d@�}��E���RW�
��"I;ԠK�5�IN�{���_�-)s�ka�C��EU2����s�be�l��J�C����̏��Zs�:(]�scP7 b��L�Tk��>�Von 3=#ɦ�rI=���;�:0T9�#�zG���Ϙ�){a!b�:}�Z]�9��A�á�Y��( :��G<�A�U�e��,�i!4<T��)k� ��T��-�`ʁI�QW ���Q�vK�Vև6DC�Z_Blao�n�~J�E�F����2�öu�t�u�<^�ƒ�'��]Z�������o�C���a��;'���7�!܈��jZj�R�]ύ��&A�?%A�R 5����6��i�+KUJ���8�B�{X�N'���oM�ݤ�/����<88�Y�/r�J>ı��U9e*��d�b'�����U�5�j�#�����L�L60	j���H\���D��L����ף���K*��S�P��h�hP�I5{"t#��s��4��t��<��P� ՙ��|D�K

Z`�|�f�z��R���z�"8A��G��o�M�@�;D��7��`��@��f��/`�)*J�!!�e0��3��̬�Uo������EG�����̨
͍䋅%�Ĭ�O̕���zo<HXQ��̭�U�ff�
E�Kbv�~+�;M\'3zM ۝18؁z���C�%i0�����>Z�:zVb���N�������C���p��]$�S�FϊW�4��Y��Mã �\+��3� �üʊ��"<����ǵ"ж�аX��ZM,��`qm�T��8��Є�I
�1�q�� �u���I�"���+e��Ѹ�(����:���S��ـ/��Q���zU���(�	�۸��l4�iQ�r�Q�����8qn�����K��O��������W�ڍ�9�~�U����&dc� �><�!�Ѱ� !�v�����f�Lp3���y&?�����5ev�E6]'���]�Po�N
���A��U���J�Iܗ뵩e'C�\�~�����J=*f��p�%����73^+���^	��Zed꙰�jpM�T:MbߔLy�CN#� b}���2�
��bO����sc��n�^��r^�R��_�v�'���2��ZW�a���U�ZS�D���0V~}*?�Bh��RXDC:h�1��d�d|a�=��tkm]�7b��վ`�k���R�h���){Un�����d�����ƴ&�S��Fft���&`���ҟ���� 3�vW��dV��� ��0�/>SN7[�A��J�9
W�D����#N��IJ[!:'o�ה�/���kwqvx��I����/bznV��F��b��R�X��M���g��053�Z��Ó#�]�K�D#
�<X�!���hf60+���A��}na���F8S\n6Qn�������;92��O)�`$�h��r��z` g��k4�3����LJא]Y@�lNqV����`!D�y/[&��Z��ø�n!��[>�x�����n�MMK��?_=i���^��3g�z�:���Li:5�H�"�hZ��7�(�3>c@��Q�����k7'�勨gd!#*�/�Y�P�v��pN��������L���j����U�	�4�<�qg5�xmA>~/��!���2���yiKE� `��Bׁ�c���'@�m��yu"���{�aL����h�Hf5-�'�
n,f	.�1K`i:9q�5��a��f�YIQm��q�D�{��C�%����W�,�LH`�h�FHIw�xߧnTkaPmb��Y�pP<d6�U.���P�F�/2`�U��t	a���PD�TB�A�ߑP���0��oev�6��+SE837ra	?h��֚*�U���uד�de~����Q�XN������|�c@�^Ҕ�_��1أ"d���vWA[��� �W�����K%�)A�Q���N��$
�`��v��y�El�l	[�v��y�8(��6@���Ť�)R4��/�aiy�pDX�v���n�J��$i��Y��D��y��F�H�:~��M�����-1=�A�U���Z�^[����
�����v�fM���
*L���'_����_짿�Fpn����6/���Z��:�Pmx�����7���@�,5���z�T��(I��%K0v��J

F�I�=
6|������bIe%�i^A�}7[ۻߩ��"��ԝ��f��~�F�ሰV�f5<�I�G�o�!OpL�=�ٟ�)�t<�B��R�d�=��ya:!���d�N	�d_I�`N+�#Ľ�;t�5m��A,D�Ȅcڄ�v[�D�\��%�E�9&f��Rce��P'݅j��'����_qe*���8�d:A���F\��^-��>�g��ƕ��"A�� ���*u�
5��@��>�Ʉ�/3���2�10g�i@(�w���L��I��;�����e)�f8�6yI�Jf�H�R���O���Pe���E���ʥm�{��i��\{��gX,<0�BR�����V/���N���҉�🎷I,b~v�xR���4�9��-�!��Vp�=:ĳ��qrr����w>�{���R����prvf�`�Rq&��RvF���U�BQ;/�H"��!cf6�p4j�����Z$���wt���S��_��k�+��G�{҃t:�u���^#�-�fM?�Q�}>\v�8kTQv� ���^�W����{��QoՕ����x����^�����ҟ�����7�j��W+��g�F�7C�7����37����c3k���&	c<A�,���R��K{��q�:�2]��'�%qR��=�O&EK$v�n|]7�f����;����d�L�}���B���f0B6�d��r���bъt%�̓KR/v�TK�cc9J��7��/ ��eճK��Ć>�gg�������8�1�`[��G�V��	�S=q/�'��$����}$��ɅH-NzF���2@.�����L%�-���*k�V�]�.T�Z���a�8<8x 4��|�|V��s%��fy���tg߈�-ɾ��/FJ���FA� !Dɧ�i������Jin��Y��V*�f�pB߻��֒�#t�/~�����P���iTV0�gnl8�e�זW�x�T^ǳi,n�"H�m6�j�����8�;T%q�������k%���'�Q,����'1��­�5Ap�g8;>�����f��v:-���J�r�MO.��C4"����	����,���}���i#�8�r"���jn�]U;>?*��k��m1H�k�:�	��?Kx�p���"�E�fܦ"q,�[�.l��\|�O�Hp���uk�U�'{��O�w��On,K�\P�����KQ�ޘ��� ��˙�L�_�u��,m��}�zYc �E��48�	1.�4�fe�d�%9c�W��I�x�,Y/�`oKg$֢�8'f]1�PX���cl54]�|h�me��K����<Hx���$0�F�Ї�;(��[������l*c�cv`P-WT���[]^A�RA��J��e�0hz���R<~Y�����,�777ǁ���$	�͎2��D�w0���g�XE3q5�#��f�3�R��Z����R��f
;e>7�t!��jקdp`a�\������	�q� ��c�/�)�a��fIJ��
yM<9�`�Ȁ&�N�FK�s�2Y��l�R.��f�Y-��,��
a�a��sv٤�v7�b�zt�~�o666��BQ�X*)!���4�#O�������H;���Օ%H�51���a�:0�sy�^^Í�e�����C�_Z�R��Npxx�B�d�뤊��"��fg��qtq���:z��|�3���D�N��1�)��=�A�խA_�m�(�@�?��Z�3�\�շ$sH�h�^`$��Xb����/ߝ���7�~��|��I��O���������E�ABD�W37�o���h졠E'�RfOײޮ\ �rK5��p
'}<9���Z�.q85�5n�� }+nl���!#nk�f�t�X��DvʨbaX���b�6���5H����'�����et0Ppc�D�Q�^�,��2y��Lx���$��૶�����_h�8Oc&��;y��~� .N�T�R�a>���,�A���I� ��A��M������)���=B�X��Xi"�9Qe	�Ǵ��"a�A-k�'3)��?�� R��]�������.RA�0Γ�'�ZV�ө��=�9D�D��2�T���xR�t�x�%��D�#�ӄ!Х��<!ӫcvʉ"/�X�. Ą���2:��BH&
�̪*����Ѱ%�����Ѐ��1��@���}S�n��*��°�ѠL���d��i#�������
dL���{�垠1wn����wx�s2,���6��t�7��qsqE��U�GG���	jR<���O����Z�� Cy)f����	�g�ܶpp~�J�n�0 �0��Td#g�I�g���Lb�#���a#�A���(t�����[m�����m!���`q�oN���7�~�����߫��A��Kg�&j$�����5-�,K�0]p�_��f(@���.��B��B����enn����� x�@������{D,	5�4��q��2c���z�
^���	��FΓRN�d��g�H-4ꍯk�Lɟcpk��-Q���Y� >�^gf���x�/��)ֱ��Mc#r�$B�l��=���
ES����707�k�3�)������Q}��m�.-#��ŋ�e0i7Zf�Kd;3%�l����nJ-ҀWA2�M���\f�h7�c_:6��T�p���bp\�tBA��p���2�5_W�'~ U�����1f�����tA��5Qf�&������RY*a)l�YI��j۩��>,7Y)DX��U:��4鶞�ϫg@� ��,��e1.xk�
 �I �ˍe���L6+��栋J�#8�?]\    IDAT�uv�=�..�΍���#��n&r����'�:?�j~��n���MԊeGVO�KHOO��|w{{;q/��@<���*nݺ��TN�Z���+�Ѽ�j1� �����]��	h���BaN�M����1��-π�eND�*|�_��a�-��t����_�l>�'?y�'������f(��G_��[���Z���:�
2	Ѵ���!��\�,=�s�tmH�.Q���ˆ��4:k�>�zhV�����j|\�m:*�S���?�(�1kb���.�f�٩��������/b�T=3�����G�����0�d����&(N����G�㗱1_���S��L.���]�51����&p�~����{��j��#� 6�#����l����w�A�ZF�X�I(.��'��i9Ƞ������%������X����!./��
���Japc|�dH^������Trl�"�NW����������:
�XN���r%D���jt��P�x�*��;�5P��'ׇ�T�=Q�S���S��3� �k�Bg�~O��v#�h����*W������}���g*i*�y/n��zuNA(�t0sҘa��v&�d�G /A���[����Ю�%����ܨ�"�:�!D^�x�g/_`��Kd�)ܻuW�[-��wx �"����l��ᶆ"U�n��ծӿ��]Le�qzu���[����RSܠ���o+�6���0ݬ�(
jKSfol]�j��)`��x���IP�fߕk�U���Q�����7~����~#��w?��=��~�Y���VU�.�Zk4��[���5�B�ېY�27�����h�A�4�x�иx�&������a��^U0���LZr����)�pL�M�$r.�'����4��3"��Cm�������Y�))��d�Y}-�
���wTF���$I:����m������[}������)W�v��T�eq$�\��9��T^����+�p�r��d�>�G>D�4U1�9-��e42��'��he��+%a��Y8QA���q�rC��E�n��L	�P�,�}��`E���1Cb�Y��%��L��Ϧ�2`b�L�,tz�d����)�k[=82&B:d���癹0��a�|F�����w��ra�F���:z6��Ig]�O�X�4�031"�	˰*4V�03r^ܸ^3@�`���{�@˴.�5r\{}ӷ0����<\f��ԻF��LO!�N*�eB�a�;�o���[zН��k#�L
��R������,/�w�A�P��с��ydg��d���ob�`� 3�A�]�f��t�J/v��h�J��_�e�T��(�`�e3��5dd̹��U�h�~AtH�d2������f�{dY�![8�fp��XI���ϯ��ʭ�?�o־���gn��џ��A��������^��ϫ�-�x<"�!}K��&ʒ1R�F��\���4�(l�au�"����E�cw�i��e��/���s�X�D�DF��ܰ'BH�m֫���h���/�ꝳc\6�c�_%S�!�b1�CQ��꠵nU�$y�*ݫ��E��$�0��F&y�3���i�MZM�\��	U��*��з�L���������bs��SD�]��>d=A��^�Dc�G�0���2�ഋ����墲n&�f��'�8?Q�Li�R]�2r#Ca�':�W�UA6rӳ
����Nt~psI�KɎA�+���F;�Q������E�O�"�l��V��%!�<I�CR�l0D��l�N��o <�,y-��`[N��C�f� ��(��2vV��,ǉY8{���d]k22��))>JP�(k�i����9�1 XZ"j��WwtbQ���"�I����4��p��
y��[/^j��ֽ������s4�U��y5�yؼ|�\A�Y�;wpuYTpc�9��n��{xy�-X��#�=ݽq�������p�϶7�`�.�9Z�����p�B!M#P���z�^�1/a�B�����a���%�!&�@H�2�}�=�;I�bp[Me���/��{w��՗�>o��?Ȳ��}�?8jU��A���I��7���9�?`6Q�3�*��n2��BU��u�[R;$i� �ĵ�<Vg������[�{�j�vcʘ��Y�/,am:�$��������g��en�wl�2-.��8,_J�����NS��,f���ĕ�q�P(���T�e��r�t���,6V�8���3{�̍���P���e����#���A��B�7B7���A�$�~]��@���U�;�(��:��),�s���t�V�kq�czfƸE���SR���4��h��p��p�M���OrN�պ�)3�S��}x|�����ɥ){��-AJم���Od�[e��t���T6� �L�V�j�Dc1�P��3KJ�38*�S����K��Z��9�ｴ�8�����Gz�̇x-~�YjuX�SX,Uǔ�7��G�p4n%�M��J�b~�S`�����3���r�ԣ��[(�I.K�t:#��x:�x:�tn
Ssfj�������������T|gg�'�t3kO%����}��E���cgO�yy��O�_����Er��|xw6n�ޝ;X�/���O67�p�9*�����,Mc��p���ZC���}g�36����o��:�|����,�^�ʐ���!I��`+���[󫿱����?���G#o��o���v�4�o1��H�����A�1e�GT���(Q9����9�̴����T��1�t8.���Y�Es�Z�(W��U^����6�Z4=,�,cei��<�l��\����յ�0vb��9)�5KFh�hW��.%}Vf�qgy	OXM�z�1r*E���JQ��p���U�Z���DoH�[7N��qj���G���|OvwT7<��}��'H7K�� �.TP><Ai���2RC?ֲ�X�ɣ[k�Z,�m=��2��Nÿ9L`�"�RK4����/��h��!�?2��F�`�Z=ee-j����"H�jt�8�8S_�A�7ș�ƽ�X*'�Ò��6Í4���:Ii��l���1K�7��6��Ph��`����:���+7��.�9G�#6+���X�� R�9�yܓdi�>�������3�k�Ϥ"�@	�Gf������ngw�����W^S�K�p#�+	��$AL�L+��#QcP�W������2�S����������n�n��=��g�����uMI�����v������f����e���}��G�O�|kSW}OЇ֣����oɥ�8�Gϟk��F��X�G���z'��>�2b�x���9�`� ���>��eMP�=b �PL��j�V�n�@��V�S[��-�Z&��o�8��|�+��3��:l����f�6�[� O��#�G�fl���@����n.�9��w$�I�->0*�X�Ss�9���X	_��)������Ԭ��ܽ8�q�R&��b	��u.���T�`�~W��J�.�)�e�%S�8Qd��Q���閥�!e�j]��u8���q�Gg'r[b3xmi��n!Ok��F?a,�|A�l��@rzH<>f�����W8�A�
�aK^�0�Uou0h�Ы6�*��<�BXXN尔�	�OC2��Uh��?��a��4L 05F6��T6��}4ZM�_�Y4��p嫒���N_�'77��TV=�b��G
j�n6���߲�� b��X���mw%'j��\���W������,6n�aeuUϋ�\�^����Qk�li��1�87�7ql�F˔�v�"�˨0[%F�V�4��[:N�:V�ˍF%���JP/%ٌ��h<n��DH]�(�&\�X���+�Zt�Ji.)���]�*��P�n,�%	��/��`���N���X1���[
p�jC�ܣGt}�9h�wO��4F���CGJ�K��/b��?�g��um�Ff���w���ￏ��<O����<��B�;D�<r����k训�g��e��R�a��bY�zx�Y��� J%'h�3�ZE-
��p�F8�r*��~n�W>�c�~��kj�_R�~_��?���/�|Ԯ��a��~ܨ�J��tB��ƍ�q*�׸��ۮ{n��$ �uz(C��У(}{f7f�o����������Pel����ÀW��a����1	NѬf4o��ڈ��^\v�����<��ae~��y���Y��3Ǟ%a�je����\d���*޹s�pZ��˳s���{���� ,`s
�y"�P�5�u|��<y��l"�+��>��A�͎�*��
��%�����G�D�\R�ׯ�T�R��6��`$j�N�l;n����1����:�G�%9O]N�Zm�V�h+@0���_XY���N���K|��_���!�..M�F�l ��̆���ш-�������,O�Y�|�V�� r�)т�gsȲA�l��r�d��|�Ͷz���)�����
,�����5^�����~�~��T�S�5h�B���cpY<���,��Leǥ=��H$��C��`5�%�ym#)�*c�s׽�*�e��`�L�	���*�Vn���{�[Z�����x��}�.n޼�v���O���ÏT���r��m,/-
��u����L�RrD�K���������|�g[/��ʨ�<��m���{��̊~���3<|��nN��#�O%��$��t���*�� ��U���?��\4}O�j�X���j�,@�o8gn���˷g��G>���xp���oF��ÿuܮ�O��ʲn]&���A(�ϣ��3�$>�4�%�h
.�����Eէ!�Ӂ0nM/��5,Ħ��N��+;%�(U�&�P�CU/��t/O4�Z��Cgp|k�&��zh�FU����#��%��TLX��ǭ�%�L�a:�@MK'g�U�f����^D��i�g'(7*����훷�'P�V������mԚ5t�u6�#73�U;b���h:8/��k}_� �~��$B�?[�1I��*蝗���E�ᶊ]/�
$V*�����3�,��L3~�A�}"҆�a "��5�t�bE ����y�I����C`���c��&NO�����i��F��x�l�������bN!�M3� iN~dRi7�g�D�3@��)ezD�
�zidKK5\��&�)@��$����sxD;d`�r�U�aW\a���?<�s���(�A�ו�eMp����fP��'�L-;ԨU�KEN�k(�*:|ܴ���σ�33?����P��cR�jY�Xtcko[;;�f7n���Ҳ��'O����b[�0[]Y�ﾧ
D��
WEj*��T~��p�Ock[�:��81���o����*ҹi�����K<�z�b��QdП�h	7*gK*��#�^��/nZ�`�?�Z�z7���>�̠���Aª��� ���{3�_�b?��?p��>y?��S�{��r���e)��x�3@Nfn(0{}�nD�k����n 9�0��.0��3�7q?���7o�/����CI��(#����TN�x.�j����>�~�`��vDg!�<��ݛw���DQhV��s��;2�e���3'��VpoyK�",G���.qzp$n����Y��%:�^�Y�
�����rab$�������e�4?;���2�ݺ��?&������#|{�)J���I�A[�����x���"�CfBqD^�k-1 �8��8��t�(g���s���(-8�Ō%{<�7D�M��)gݳ̎��~���N!��Q��?�����ى~6����C�[ q��e2
;[�ꅱw&hIؔ��d2�H�\�@ȉ�2F�
T�Z�}Q��mԚ��	&��0�8n&����ycX6�5y]�/)��az�V@��U���Y�q�E-�ʸ���,�\���Mg�L��A�I�A��NO�p||*m3B}\pS�]�PP@ޙ��֘��"�-'��ܔ�1�0�q�Tg0�w?�}�����2�4޽���X�/�*K�YU�5,,-j�P�qtz�ÓCe�*��]���&��^O��6_����D��B�6Uf覿fX<���
ǙE���=s=!V�u���lw��]���:I�P(��Hb��t�W�����?p��n7u����a��뇭��9�S���4�z	��N7�ٝn��S�^y̩n��}M9�B�@�-m�ś��E�V�����
��NO!�������a�">���^�\j�T�`p��E����5m��c�hT����I��˛Ͼ�o/o`!����������)JW� |0,KhEG��;D�]���|�<ɂ!���"���Q�3 ��|O�X�Y�o�������񭧏���gh�<�|��B�k<?)���ux�-�O/�s�zCȅ�h����*�6Nn�����s��
n"\��^��X6��r��=��A��Y��ݞ2�Ľ#&X=8;���啚��dZ%ԣ�ի��
�"N��!n��Rpѫ�J)C:�?����	jT�E՛��I8�,Nس�@��8LS
�ev,f�;Q�W��p~q���=���#��F]��U�`0Ѝ�2�O�I4����E Ȯ�o6;b�Dc���>��Rc�p���9H(���"����卥����eHd��F6��$�EӼ��.���Ln
�d\��dz����@���u����|��x����~PIemi��,���q�4-�����0�P(DRw
��ܦ���J�g���K�<����).���J!p��ב�5�2X��T$6j}����g791���S����pY.j���"�b1��wy���3��>-�=�P���V�W���[�Mb[����l@JQ�ˌ���>J�����N{
nܰ9O��8�]����u����3#�X��s�jd�S^�W2��">�}���J��hv�zB��{X�- ��QŃ�x���0��u���[�e��_��]��=���7		P�B�<yr�����N[{� �!?F����B���c�	��rg6��j.�l0�n�+��l>�Ã-���!�M��]MLG�6��6ZG�vF��V�*	
�F9�1MhQd)A��w&�[��6��N���f�$�v�K&����H��9!M�����'O���l���$��o�pq�ʠ���R�(;N��L�dg���7�F>)�&�9����E�;??+ƄhS$�ǣ��*��x)Wj�����F>�d��\&�2�Ns�@�k�x�A��Qϵ��L,��3��"?р���H�6�@��ܜNr՘g�t��bo� /�w����j@�lL�:EB���M �	>�Á*�x���W1����&`������<�9��SU=3������FC����(�&���9� x��o�\���Ac�(4��X�t��}]�wC����U�H���Mw�9�|{�{���5:L����=L�x��}&W�T�VXGp _��>���n�K���4Z�&�1Ǚ�p�X�<�:����&��A}R
��C��㑠ũ&Gm�kF�34�D$\��M!MN�'�E�L�C���$�P�R�B%3M����G6������:����Q�����7��P�Q�5�� f�_k��n���ɞ���Ȉ�/B�0��CT�-Z�.�SF����12X�Vj�e$6����P��Ϥ�����Ѯ�Iv�al/������?���L���\�M��y��ݷ�;��r@}��Y��2LO���5�Y�����z���@b��d5�ӧ=��Q��*��F}�h�n�������9��7��/���z��i��ͣ}�Y�w�����ՈI�<uNƌ�>+�*=��F��g(�D���+Ȃ��D�L�����nP��t��#�>��i��\+E|��+4^�b>��sP3�"Ræ}h���}����:��t� n&qp`P>��&��t�;���3��v���0��H����)B8�+%���#���2�2YN+!	׵ڻw?�Q� �~�"Ŏ��\2	�Xs����}�BVD���*5[    IDATkc>4���Y�W%@<_���ؤ��Q*8b�q2#�kU5i��ôs�n�羟1�k� ߇��57+j52Ӗh����n���j�\�0s�Wʤ��p\:43C��E�3��H>���O�� �禦9*�����0U L�X���)VFA�j�ʨ'B*j�٠3L�ut�z�> �5:N9����,��r*Kâ�n1�=_an��(�.0yd褦,VO^�u��4	�) �M�6�JM�2��M )@ֿk��{����w,��&�����������1Mp�Ps�3w�
n�\�:�K��6�e��|�NZC�C�h`�\��]4�9_g�,1�����"ݹk;�\����#�q?��b2�T��~��޻wQbR��u�A�<���WG(-��+Y�m�Z�����ٱ$J(���5��/�����i�n��\s�-ކ�=�ؓi@�R�shog����=ph?�U��e4�Pü]@����6��m�ퟦ�/Ӡ�ap��4�0&�z	6�����ۜ��>s�xHY �ͥ��0�Շ�h�'��`�#0(�����q
���!����t�R��cWq]
����8
�-1���I����Ɔ,f5�gԩ���PL]�0�2�WE�N7"�c��H�J�	��ap�օ��㱈#�����O�^�1�x|���[�L ,��_N�k��
HK���S����]���29:FyMI,�#Ti��?�x�h��V�T�����o��яi���Ȩ\)�~�fh!/nX� #�<j&�T]�SA׭0T�|�ȥ�v��t�G��N7D���e��O����V���P-���/������:D=��'���#9��f�P�|��!5|W�Q���!:��p��$��	Pdx��QB<�>�!��x�*��Y�� e+%���m�=3E]��@��r	⛩�����j�X�;G�n�uoeε�v������R��R̍rMF��Y=S&�3Y�7ϯ�{����6��YO�����Ct��8�e*�}�v:B�f<-NFѨ���KDS��k�vڽ0AK^�4�K�!k�=}��<L�l�{=��N�g�.�tD��6^���Q�o�=l��,W��Њ�x�@&�&'��yڽk�4kRR)�Ӈh��]dKb�'Y�JӺ�=o�3h@�Q۵iOk��ط�~�/�[K	xJr/�Mb�1X�-vȝ���H��jq��iw��jP��A�87/�A�H�oL���W2�DӬ��MG+�#���S��i do��i��s�驙Yz�����[BS����yUoƔ�r�	��(����gDIHYy���uEg��ivKרR,R}h�Ny�S��ςP�U!�	'��� ޛo���m�4�����q����
��\H ;�#��n�|��ypp�����%"�LF��b^��{ĳ�j��N�Ӟ�4��!}F�fY��I�R43��͛n�6�޷��	���H��
+����g5�V�D�\��|9�Qi�FC�$�Mv�:�l���ѸBe`�
đ�0�Q=1�����*˂/��Pkz�Z3�\ !�`}��Y:����)����N�ڡ+�*��]���(q_�8�N�l�jV������~�O���u�E(d�K��T];J�e���8�rZ�{��Rɴ�p���u�o>�5��o���;�_{��T���GfKpCA��H ��.z\sc�]���� 7:����%1stR�N���P�DQ����8����Q�����U��A���ݳ{;텠��f�ktZ@ACam�Fiͤ�N��߷��ڽ��@���0�
n���T��@����ؿ�CpIx(���ӵ#�4`e)��h��;H3,v.��;s��!z���B��F��Neh]e����T�r������H���N��}��jH%$W�@�����wIk;$/t�����d�Iv�<7��� ��H�*R�,��ӣ�7:��ST*8�e��Y{���) �jHǸv�`xtlڹk}��ߠ��I�s�\E�/7��EWL̓2�L���@p&�H�Y!����G�����
�Wj46:B�|�3���1%D�h޸�#c>m�A���۸�����0�B���{!����g���I��R��#c�����V�sdT�� �%H��Q����=�y<É��<�#M��M�v����=����`\6������z 7p !�M�'Dި�q���-Y�<��_C�j�����D4e�0*��h]p,���cV�x$����Esk��in���x~�]Ԡ��V��G�L��u�J���4ow9���_�NA;OL`� �a�BtA�I�J��c����NߦV����le��7�%�V���Si���$�
 735�yl��6���uU��=|���o�k�i�w���%�� pK�A_P`i�����WƬk��<n�wbv̲C2�t�� �J��CZg&hǞ�l9��58�Gj�t̚�T��C2�Z����t�|%m���v`��m�`���N����Mw�~��|KD�Y5R�q�N��l��|�Z��A\�C��K Eְ��{��:�G�w�û�f�2�ُ����<��G���]�T�i]m��~�S�l��T:�o���Ow�}��j �M���e�g:]2I!��x�ҽ�F�,Y=���#ݕ�熨u��-7QP]6�2A���ߠ�F�e�T-��7F/z��\.������Iب
����������o'#��6�I�߉.`&�f0M��$�yx��Ħ� }���)"PU�4Ժt�֏���7m�Ӟ�L���[�>j�A>ꑚɼ���	��7���57��#U��a"�I�0 �r3]��z]�IR%�;�H���Cj��<������kuKS%Őhh�F/zыh�T����7(����	��3�s�o��Iߺ��,
[>怩B��P,r��v���,��Y��e5-gRm|���A
,������") ���K�!�I
D���b�z�}��!Z�s�h�	C��
��T����>ni�M�-���<"E��{����1��&oZT/V(�,�.�I�}�J
e$MW��N�Qiw&M����Hq��M5��󜒕�����<����J�ƣ��od���;�^}���L9]����8�- ���b����<B���聡9��>a���PUO�q�c�ax��i�K���fh��},��s!+��Fc�q��y�	ԋ��C�Y�ܴ��7��-�3�=�F�2o��v�>���޳�Z��ĉ5`���Ik7R-?@�%~ϟ�|��؁J�����`�D'mD��F�@����9z`v?��qH�kr?M7�˅�4T�њ�(���x*XY��:К��w�O��y��jDM8Juݞ�:����9�̻�Y�`�7�$�ѥ�v�{�G�-��fJQX�r\�A���
��u�b��4G����追��L? �3wB؍�.�؈^��w�K?����w��9 7�s�����?��:>�)`eL0$�������)Hq8_A�8�>���锓7���<J�sD����������R����_o�7NQ=_lT�J�o���i`@����,,pD�>&��z!$H�b:�i�5��SȂ�&pR*���������k�l���C��t�u*���顇w�?�����?�Nj�"ҵ2��@m����	�6�s!��5�@5Z��406B�a�\���d�� �a����	��ޏ85̪�\2��]��{���ER�K,DZ��9{���j�����Z�f�.-�g8�{�D�j�P���ʔ�B��d�����*�b����u�=n��c�f�Z��K34�Z�i �� �)[��G�ߺy�~�K�"�_����h���;<�7�^}����v�Ԋ�A	�;��WQD&��t�O:p�8\&ʲ_ �A}3dpK�e쫜b:��uT6KLd� ���ãN������ ��&_�z�Tc�v����Yjy=
Qc����n��t�U��M�K?;�������������	c���Lj��3}�~��!�1�h]Ȍ��Cr��z�(ȴ4=˭t�Đb��ʩ$���Ȇ8*�P&S4j�!��? �'������������#ؚlJ�Tߣ�Tre&&��L���A̍���̶�+�'FX#&K���1w��n�hE&*f�E����q�C�9���^��#��WU��l��Oo�����λ�D�TL ����B��@���]9VU�U:t��\Pw�b�NN�DO}�����=���g0W� z�-X��)\�@��ٽ����tם����p�����(����R�>L�n�f&��F�0aehQ.a���H�L��-&/�$���n����@��� n��n +���V����I��m���=�)��x���e3)2S+��Y��u�{�t����^���v���-��mp�8��<�]\�%ϣ�g�d=�Y���
J��E��
�U��K�I�OS��S��"����hb?!څ�������'�5T�iH����¤�4�p�	D�%&Mc�蠕%��y�&�[��/Q�H��%�����y���֝x�jeN��7�i��@��.7Srf���Ɓ�O�����R�����9���;�_�K����ۣf(�5(H� ����0H�0��c��sG�AF��B_f��X�c��Q�,��v�3��P�n9���ô�>N�#�^���K�ԁx�&S�0h<[�gs����V�ҽ��{�!_GA�����6L)�d�~���LН;���H� n9ՠcFƹX�֜���&�`��C�P� eB60iqd0@���w��ٿ�v�N�X�g�ԗn���PwbpT*8�s�L��Y��}VQEj
�&�#��hc��0n�,d��&"
Q� ��.�@�Hk֌�0���-�Mt�c�T_@�%�v�����~��[��;�l"��a���AǴ\�{B-#�f>�� ǆ!�Rׇ5b� �q��|������>����g�1��!��0���$�tm��ޟ��������g1�%CZHc�\y���[b��m�b
B�E4	R%�o�^c�f��8�ei̗��tڰae>�#�yC5�tڷ�0}�71����Q,t�uCf�#�P��i��"f��?�¹Q�ӦSN"���9�G�v�";���"��v���h`�g%��:f������Q��*RnD��_��{�B��m>�R1��@	��	�ʞ"d�?N���@�%�h��$��;d؞0Ǵ��A�A��&{�n~��8RtL�vL����Ys^浨�3����02�������
n߼��ڤ�|�a�u�Ag)3���HG����LE�;��*�(b�D�
�,�����F�CO��bк�0mĠ{�� �@Dvp?�:�����5.z�����o�ɥY�3u�&�s�ň�*��"�36��D��
K���� ���^�2�P5�۱cki���d��%j�H��Lc�)ep���n�����BjH�t�#4��!_^F��ڃG��Y�����~�C|x�Jȵ�XP� F��d�\*b�lAvΑF�B�Bԓ �6u���v�!%��	 �(�1�����{%E��.��6��b����gK6PpB�;F��*�f�����n��N���i��K�Cw��Wcb+����\C*�n�br�����f3���&���g���O=�T7�b�`��� z�^���{�cp��{������@y�i�ДCʎ������H�
D�A]a�� nL��5f�i�������t��J���_���	N$��ݮK{��Y���O�o�x>�n0ꄹ�f�M���<2�6�ll��FZ.M�����=�ɴ;�&hڵ����i)H���%�@�T��hDm�܌H���,�g�muY̆�QJ�PoX��)�<�x����+��}C�>4�b{ ��K���M��Z�T�;�r�Oa�C��P�@�#�hfa����y�O;��|���=xx?���n ��Y2��Ɓڇ7��� �V����?�N{��L:�8K�Y�OM����%�Y��e�[�t���Wn�������!��]��� �T���.���+�η� �m@A�V(р��Ej�m�\r;�k](Yae�5�4R��)T0#�on�xM!�D-`|`��=�Z�]�p�ˑH���!5>ۚ���Y�D�#�YH� n�� ���@��j Ԩ@M����}3�t�n��"[��.�
Ea$���Pk躔꺔u%*y2O]��BP
i�Yj���nw)t�Q5А�k�@�7ņ�u���!�]�g����I'�D�}*F�p��D"7(	7�:t��ӏo�	Gn�M�um�l�<���7b_t����"�c�����ՁE�7ӯY;��; 8P-pp ��B����y������~��A��2��2��,EL� أ���B���6����&���,�k��<0����7m�@�/fs�b���&�2d�����l�i��}��3��owP��e�u��&���Y�	\ZX��!|��Ad�(�Mц㏥��7Qa�B�'�}{vQ[����6��-�
��ұt=�-��(l��=3K��%&��K�G�	%�z=�SHͧ��t`q��:K���":�T���� &8��2P�.&4}�.�[���K�&}L5����B�G{g'��C��\��
^�� �l��.;�>��s�y�э��s[���Mx��K)NK���c�|��U�^ظ �ƪ�Ѝ����O ���A}
�R�Ų��L\�p�Q��h)���<����ɨ�<�w�����`~��?����u��(��q��S���Q��44�p�`X���xXd��l� ��3R��� �w�����f92D٣��@��4�!��R/�VG>��o��Sץ�R9P�iT�2�u�<V�8;CKaV��h�a(����
���֩>:B'�p�� 7 >Z��3"#�[�ѥ���n��/`pxu8L	�,8Ʀ/���BVp�X���Y��a��I�)Fd�J<L뻧?�����e��N�ǯ!�B���1����{��{�B:��5��ryD�B\���Gl�8��.�#T��|36���#bܐ)ܞ��r��2�bBDQ)_(q�%�v�K{�`*��X�k�Rv ��5�g(ɸ}1I�g&Y ��f��CU����˾�ir4��h"�>5�_	� � t�U
c�z8�nh4`f�iIo&F�Rb�*��:5}�&�t�9Oסn�������!s��V��F��`��7ZTʄ
)���#;4�PN���LA=�N��b_ Bl���n��Y��1����}��㞹pT#7�[#t�����-�@Y��,��!jtZ��� ܠ��mj�M�x%ܭ�
N�t}��eN��a�C! �p8p��z����s(��˱�87�h��x-��F��!��A��XX߳�� BS��� `�4s���f_F����E8u�^ȡCw�Ue9byā<� �h�X%� �����P[�M��{ ֐��t�f�N��8-�J:�%C [ߧ��#J���\�g�Bv�
�C�cp::���0��z]�P��T�;r
j����'m>�N;�4�j�: ����P[�;.A���l��<H;w���N�ↀ.����Y�ud BZ
��蒁�x����Q
����kC}5�Ye�ŧ=�T^4�M%�5�t�5ZB\����O{�d
�y+"]E=�K���2��q〹��P�eB2Go�� lEZ�(�t�f�Titd�6n\O���,>��B��w&���"@�>45ó��?�SCn�(�Ӝ-究�N�B�3���4�S=�H@�@�mϡ\���v�QTΜ� Q@Mf3��&aj�ό��� .�TF�%<�>e���R��uN�Ģ��:�B�MS�%��uy�J���Q�������l�"|1r�)v�*i�k/��$�=��L�Yy.�5i�Ӥ�~�&K��k3h�z��*�T瘁�-    IDAT�e��F��죝�~g׽�))x���>_gΚ�Cf<$�B��q�\sCH�]�`�ŏݯX�g�<�-�4� ���h7���c�j.��1/a(L��>>���=�k'�#�Pv�4AKM>�q��P#�XH3�Q�`�YN+�0� �� j�A�{,s�$'Jr<X���Z.��gH���bP�3¹I�������,*���gL��eU]�
�i{�a �!�6`S��Е����;�,�<����C��Ӟ�57�Ȱh �HT$����M��A{��c�H�Dj[3�n(}�&- lvtK��	�a�=.�Ǿ��h�N �=D�+��bq�Ӟ���i DF�B�/PIX3m�I���f��� �	0�ẒauD%��@/���x���),_
S_���O8�Hs�Y��iú�t챛��ͧp=���B� ��z @��&�]l��C,��id�̘T�Qi�ʶy>�)��P��cW+~�Yǆ���@V8m�x�Q��2���x�N`aJ����!�����j���T��S�J 8�?�4��Б�d�� ��t湳�K��CO/�Q6�P@����HU�4�!f����8�1	�ua�2e��d ǡ
pC��bY�c+Տ��n�g�^{��Q�� n�r��)�s��ά5��'���l��LN��p�C�/Ո�5�� ��T��a��1��/u���k8�-4X9��Ɩz\�)#Ȫ�N r�9��Kȅ��*�D�xf�G�s�8̻	����`|��"�� 7x� <�w�QI��zL�#�l`'��;��[�a�8eqB��G�,y��"2]�'��e<�Զ�nXn��t`o����d�V���p��gITf�}�`�s�Π��u�x��\תժ|=7�7����YM�	h��]t��$G���P�:HM@��f3񸓈� ��QKֈk��`;�J9�A�:�"Q������È� 955��0@�czs^c��ӄR-T/pLVEtp�C4ߏ:��H!Rg�7��q}�|���{�T4"ʤ,ڸa-m>���o�ʵ։�I���en�;�el҅f�f����G�HGQo+��4�v�R�"ua5��9�Taڃq3�fPD=tna���ɺ��*�v�{u�x�-��/Uϭ��l�	�C#�7s@��g�� 6<����0�l��L�:p��ؘ߯\�c��������Q���ԡ,�E�{qG[��@�m4��q�� C�f���Tkל4��?����G�nڱc��u�7e�/�ߚMO�۴�h��-���]���"���/C'��s��G6#>ҩ�����8��nӭDK�0�1x䏅Y?
`�� �NT���9�GB��hN�d
��X5��x|"
z�ٱl2GDp$��tx@E��JL��8r�k�2����Ʀ���k*2w� ���⺂��m��'�-��̎C���1��v��R\�B�
\�xnpyo�l:`���BF;�^<����#dhP�W��@���Ƙ~>�G��V�e_̙����T[Ã�X���<�L䅒")p��� ۅ<� �lڢ�r���s<��a����p:&_�s�(BL�7Hs;�ЕkC��H_���Q�%��J��f�N���<���N�r�(���O}������uk�M��ӟ�4nv`�B�3�s493�ׁ� ��^���SP@�EG��~��7m��H�f;�j�35dp�*x�06��Q�Ğ��TLgp]�;n�v���^���o��Ĵ��U��r�%@��A �2�5�O��E\�+�xE�G�[x��Y����"1�Ƣ��"%<:���t���g_=x^�W(cV)�0�/����������;X�򜵧�?����={����i����s���65d�l�"(2�����B��P��OP��c�DQT�oN qj(BMB�����ح:�$ 7N�b�%���a\����Er;x8��b<^?���}�[��:YP3V9��Dظ���Y!A��8>{ "V�����Ih�' �(d�yZ����=Y���"=��IЏ��s�%�Pk�1�V�L/�10���e��bg�\&��`��$�?x�7<:���8�'Q�\�n�0EFW ��� �����D��"��{�-.1�e�Vc�P��D!]8�c������9��k]�[3N�t ��<��rA�R��m5439A�SS<Q�v�{`��� �<�Gj�2�o�c��%�q�_� �q���p����#:[�^�U�'Ky�W�&B�nn~�S[�'ܱPD���"^��S��� mZ��N9�dN�!8��C���71=�T�{>-.5hjn�"��ajdp|�;�F1G��y��4X�;҅�'���"��]��?p0�
���$�'b�@�7Vs��Lf&D�/�~Q����މf��T���4���i."5�����m��`�9@���,�؜A?w��`�/*�CȺ��QW��m��c��p���q�J5�8�_���j�C����=G�n;tȚ�[���[�:�]��;Ԕ"�+#� ;"���Bk_�s�ƹ?O) �("B$1T
q� ��4�� �H��Ŕ����Nd���
I$_�C�w��ش���1�N4�+$�|bAv���	7`��� �DnlylN�Ҹ`��p<����\��&���X'B�L-CD,(��DB,����]�Ĝ$��p�r2�A��A��*e(�
�=���/�3����p���-ƉPA}�3<<�\-� "`lN��Y�������`*m;�㇛�;�����=,��TjB�(6F]
�w��gY��Mi��ť����&��ժ�f|����B��\\`J���
�pԤ �v@n�>i��3��2>KJ��ƀ� ��}���u~x=���`�44=$���T$*�s\�<����(ds�̪��MNqF��#m��M��D��u*�۠&�.eY_p��DM���#�D$S��E�tT���A?c��gq
q�sS�k�EqQ����k�?F���9h��W�|��k����y�x��������/D�#|"D��S�Ĉg'ؿ
��(��I&<�m��c�-�
��fH��ttl��O�W��}�1�~���[E���<pڢ�~|�m�2k�L��	P`�)�p]�ܵ�eX��wS:Ǯ� 7�)2�����!��A@c���9z,e�������f��ՎS���>��n$�k���w�Vx]���R�Iׇk`<c	�A1^U��ч���P��E�"�mL�E�'),ݠgj"��7�"���/{r����p�nذ��[h�(VN39jC�����l�ݣ
�\|���''�^��Z���L�a�����P�ذaG2��D�'�=t_�@���&�;��<�.jX�~�M�C�Nw����k#�2,4�,�� �X�N1�M ������:^��������yK�6���q�8�N���Kܵ�D��� �i�uUj5�>D�f�Z��8<��<��6����nx�K�<�`Zf�*�,���N"��.�_D��<�9pQ�74�[�4�����J�0`q16kj\�b[H�P���G�q�'���5��V�=�Zs����b�`@o�C#x��=��uR�8N�q���+�&��>�. �1�c�X�O,���dn(+ r�h1Z��C�q)oXT�Dn�i`�{������=���
nx��>������/����7ޖ���<+���I	�c7�.�z�C�|	�I�F2��O��`�'7"�~�N�4�BI�{p���8��	�~�4�8Q�@��������"P��4�'\_�
�j�8%����D���}�7�W�%��1���
`r$�C���k��ro��遀��HOḍ	�"�p	�b���p��IA�4��b���/�l6�/6�T�/"|�|Z�
���� ��@ �$����:��?���Iw�^E��ވ��K8t�B� ���NO��lb�*��Bm�J��!�� �8��\"��p�y1��{�iG��ڊ�D���dCV)(�
�v������닚`�(㢾7<�C�9iצb>+D֭��o���pQ��Z�
�t�uP
L�%��ݥ�ӧE��B��h�z�k ����GN�NA������p�J,p��l�g�|�1�QT\�fH����q�O
 ܒ��-�z9����T�5"�ľ��_�}�_�����P���܄����/p ��[�E�Yi�T��h���[_}�s�;������w�m�n[
^�J�M�s�p_��@J�MFq�n�_�8g-v�!^'>��kq1��3Q�K�;�����Pb�:���V��Ϩ�ŴN'�v�x"����e.p"c�t4�]�A�H���& I�T 4���'#���|o,\cb*�a?�d��P���S��	����<$�	�h�A��La9���1�,�Q�	��e����"���Lg��9����j��ֈr<P�$:� 7�����;@�'"�N���� ����b�x�  �DP1��'\���e�T6\��	�t)�A�#�� �"Jvuo6(0�������+<Hq��}�T�/�j��X�d�c�Ls�!8lF�쐢�]���+:�I���xx�x׌��� ��L�9}�$6��3��#��I�:9~@��?|����*�l�4��p���'�~�!�/�p��t�J��<�b6"R�^�:O\*���s�T1I�EY(���T��e���q�F<�&�f�^jl���%�0,c�� =n,h��� �"��
	�df��X�eM���sO��_,��E���'C������F�ɉ�J���L)�M�49p���(
dO�d�k���\���:3�������'�"�Ʃ��/DDH��ua��	�g�C�x�;F�T���:
��h����",Ce D�
��1�V"��8����p�Psc���Դ��r���"��S1�#���$B����Q:-��ŏ��n�LF�6�=�����q2�x
�1�w	�)���:A�(HW�fÐ�cכ�Cˬ@��
φ�}=�8�u��?:sX�TZ��I����8�C�  $n�Ğ�\���_��T�">�$�~=��B���UT��,�YN*P��dP�t	l��������rBl���m�ݎ#MD�
���L.���-�����O����)��9u�;1��J��̢����)��ध-R�ƣ&�)���9@(G ��@I6�(�hi���X\�{B�;x#!�Fq�Q�ǒ)�ԅ^߿�6�g�`��
תqء��&xo�떨Y�,2"���T$O4�pL��a��)'����B�
���AH��f�"�������"�=�B"2"����˖�?Z̼��N{h��/|�����`9���Z?
(�0�}?/�a.p�|$�i/
�F{A ��$EA�Da$G�/KR$K�SR�(R� g���9�� �P�$	߇?s�U�|A��i�dhj�HRER�G6��ˋ9��T,䇠�O	D@��x3��;�`�sp���"%����h�3O��8G�$�`����T�ൄ$�@u&�2eEaQE�'?��c�ҡ!���kp��#�? ��
u�H�E$�c�x#���P,��"3���i0�� �UЁG(</�]��u
v����czL�K	�H*��4;8��PK�'?���8���w y�C=B7���yʁ��4�d������������>`L�Ad��XByW8I�>��/�$҄2p�<�.��������?l1'��������8D
��p�2�x]��5E���+���t2�2PC�$<�tX��9!��������`,��2��gB��H�~$eD=�)�l�@8JԘm r�#�MAWRU5����n�^�L�Z>2H��� ,�=��LF��oH�qo���,��>��mV�q�q���P33_����y�3�-+�=�ŷn�*�^�b��hh��$��"��L���&���E�H��a�	R� �DA�+
ô$�iI�@�Rjbb'ᓪ � ��Z��l�J�˪�i�,Ɂ�ㆶcG��I�(]�W�0L���k��*2��X�v�ʒ�a�^��پ�9�"��/T�TUU4MSE#��"�{��E��ya�ы$EQYR�>�5���Q\;�Dx��Q<	 1@��*�H$�
8 �e��� P�#��-��'�Ma�#���K�*+V� �]��1�;���Fj��d|J��g'D`�+%�-[�!�°���aů/Zύ�qQ�����ʍS�ޜv#�øX\�\��"D|��������K�g�Ѥ>�"Ɇ\7�g  ���iq�5�����n� =ˣ�1�e�H��AR��""A�@�U��N���+<d��D��f=\�7t2�I<� X �b�����جQ<�A�ф� 7$�� ���E�ɑ����&uj�a�s�1�@�Ah� Fm�zqGTdC<��*&�']ͤ.�1c\��,�%ymű�� i�!����&�$*��D*�Ϟ<����B:�����s��_q�gK)����k륗��Y(��qT��M���1M)e�R�Pt$�5�g�Ty�43���K�2�.�a^�I��yn��8�5�0���V���iYiE�R$QJ�|h��8c ��繮���۲=�`.�KYSCWU�#�D�P�$Y5�P��-*E�燡�wG."+J�2�,�rR$E~�y��@�I��6� ����BY�d�)�*I�UՔd�B���6�} ��|)�TI2�0�d$I�R�1�*��RT��d��0���	�0�Y�x�t ;�)*\��0�S�	��x,�@�;�{NS�(�"�M>�،�����@EUU�PQ��
��%�8�BE����l
��`�p�8PTt�А $�\.�Ʀ��%5YE1��i:#��+���ZR��DH�ٸ�'�A|^�Bt�Q.�J	�I��pim�@��@@
	k�D(<�PB� �YP��\�/E�$#:�����S�eهXJ���<
��/�M�5Ufw�XNJ4�b~�#X&�c<����v�̃�	�\LĄk�WR�͇��?������x���Q<���X&��Ч��S���bN* ����*���:�/i�#�JG�hB��[3��5��s�-�����)�<���[A���i�J$o���������Tk���l6�u�����`�֭���޺U޾}�477�k�޴IZ����[,Fٝ;�J���+��<�N�Y]��\Z����Ț��2��'|�^��# �V��[o��:�NG��j���JYӔ�fS���׺����c۲$���)a *��@1$U�K�T�iHU�Y�j���5Y�I�d�ZQ�-]�j����x� G���B�)���>�?h���_Q��(�p�D�,)��*����v׵HK��AЉ°��j�Ȫ&ˑ�(z��]�=;��U����EM��"���u]��1b��b���I3H���	���呩��T�4ͮe�|YUd�U"��+��מBX˃&I�w4SVQ�G܈1,�A�z1WY�T5�d9�%92YSU�ʦSפИbQN���0���בj� �Џ�i����p:�?�%]�eK�e]��n�4DUJ��(�C)d=H�PLMC-F�A�*r�y�|X��(�.�(wSE��"�6b�d= `��J��ʎ&���+%�BsV�#�eI 0�._�0��y~WY�BY�U��� 9N�%�_\׉� 䄵�T$>P�w$I�Y��J�iJ;��yYR)��S��]�����O8A��>�ד�ka~���\`lQ`�)ЍP1�B+R��D�`6c=�2�?*��O��)���ԥ�<n���*��n���q�g;$�W	�92�@CU�%3#�u}!*�ё�H������iQ��$�<�?\�>�È�mSN�{���ZF��Q�a8���SӖyF�2��tMIa��16��%sƒ4���N�!G������z��<�w=�\�,�Bѳ�hZ)��HuM�U��5UAN�    IDAT�E�zv�v"
]D�<�'��H�A"�Җ��M�:�R.?U��N1��1�A�J0�����'K�Lϵ����7�m��%��@�����W�(G�=!��_ �����<���z$Ij�Ry,�&�n�_�X��)!��E�I�K(.D�P:�ˆ�R5v�&9� p#�q]_6�H�(A�E�7�@�+E��*��+��7�:���6~WY�4C�̔��iEU-E�o�a �{�"��<�(J����f����<וy�+]��~]PK�l�~�P��</x-z�_S��7�!� �t��SR�SJj
�0FwHI	�����1�1J���}������s���u��G,j���,��0�s*�xu|gS�ת�V���;nM�^,s�5�m�b�����|�,�c]��hD8R-�8����Y���n��Nd�f闽ve( �v�HU���.[ �[S�Sa��[o>��;��x�}�G\��a8p4iʀǾx�s�"�q��$�s���h�y�\R�O��AI1h�њp�n�_2p���Av��[Wb�f��~�o��M?��V|�ʅ��>�j�Y�hӽp�1�Ǥ�11��f���C^�Y��@��s�\K徼G/�F�o9A��۱� jT܌�TpkDxlĠ<����V4i�if�`�ns|=�J��A~�x�ߦy���p�S8SM�qշ�Zxr�յ˖QFƜb�@g�;S�E���̬���&0p���[���x��Ϥ��z2�����m���Ŕ���LL��`�~����������m��{��|p��ЅZ޽��
Z������0�T�X!���~f%g���p/����,K��ܒ�s��uW�Y����$@D�����M�\���xeOV�Ȏ��~xX��;6r7��C J1-�j\�����h�G��l!�O�����uF�^�����_�������a��5*��.�H�LOW�����3=Ehx{�EL���M���(n��8sIQx��p���W۫pm2m��-��H�Σ�K�L�WbD�A���J��r��t�O� 0�~X��p������j�� ���ŏ�,�L���y!�vw�oH[)��_���~B��J��&bgͫ]�uMzQ��5�t�[�(��|K�jY��"�\v�Ԉ��:�N�:�Ԫ&!#���}5��K�E�v�ư܈o*���9�1p�o����7�J��ppm:i�;�%�-M��l�荹6�/if*�{�F�P��	jqZ@y#�η���p��_1���oNo���8�}��Օa$}}�I�d�e�����㶟����6��a�Bݝ���e*�my��m�.�hf�<�G]���c�l�Mݨ�K��M��x�a�.�������N�|��L���]	L�1�t55���p5�r�A^��/�F(}�~����9�� �zp��=��G,��T��cy�}~�}��0�پIz=�&�)CI ̸�Ύ�ZhBG]�@D6�KPҨ`@��$nx(t���C}��E~����;t�2�u�Q+���#O�ё�l�ێ��؁�ۛ��|Ӄ��n�d��E��Ǳ�k��
u}��V���_bK)��~�Ch/6�U;��{���]�j:���a�p��1�!^	[��`������M䑾��FS�Q�Z��R��G���j���+��`i������`z*�̥���>/��rd�����J���k�4:�S��^�����C<ih=���U��S�;�X�o��-�����~Բ�������әM��r�&T����b��=ot�����[�3��˥:]Qhݨ�W���IMMM�d*�
.��n��3*%���!,�K[�疇��������T>�Y]��^�З���=���/Bs8�fE�NR�a�'��-�J��L(�^�D�J?ޝ�;d����A	����oS7}������Q��u��?v��7p�'�7�HN������BE��k :DMZo?�������O�oDз�T��"�+�!ӃN瘫������:�=�H{g����������a5���$�-@�7�^K�� �Q�G��n�:��R��`E��N#L��B�İ/%൐2�t}=��fn�6?���{}�"{�N���k��"����ֺ�Ia�[�U��NU6��&K����2�Hy��AS���}U��
�"9��Ma
��rKo^�]O�����m���i�e��%�m &����A<À��o�N�D�n��-����6�
�&����£F&�)	����O�A�
�Pn��w|/=�N���ϑ�E���{��{ա������'���3����2��sgђ�=B�ϛ�ϽQ�����S��~���}��I�B*�I?>�a��Z��a�Y����'�U`��)]*�J&���V�J�(	�E�]bbnn����gV�ˊ@�U�M�1�U0W�O	�V��/���~C<Wҽ���.��J���^�����Ó�.'1gR�q�U��%K����.��߀˿��Kϕvg6N���T׹��Sja���D�fs6�\�e]`�����
M�h���k��#i��^����}��vv�R4Q�$ҟbz���f��,��~��)���K�*��Zn���m�>+ra�]ȯ�K,���s�hYB�Ȉ%L��WbB^�-�j�GN���駦�����/���7���F\�+�P�p���j.����[�1�����{~e��Hأm���Aa43��ك��^F^.�.z %�[u�)���5UJa�W`t:}ʹ�E���[0Y�OCK�A��G�&���R��\�Q�<�=���Kxș����'��Tm�X��؄ �F����Шa4,p�,8�{YF�^/u��T�����tmQc�&lF�8�������b>ʪ���^�ҺQz���n��s���!�{]�UE�e�1�^�9f�Y��R�Ix��6.@��56t_K>��Z��jX<Y*�ϩ�5)E�*����ϐ�w�9<#�e�푇�����x����:�s��N���Ҩ�蟷:�x%Ug�>��Gǔ�ߣ��Y�?���"i]p0=�ј�erM�L��tyD�V,p�4�pP_�y�K�$8Z����7���-�� �pT�P��t�?7{�,]��(�`��(���F�Z����ڀU ҈�"#��i#""��isl��<G�+��^���l�8T]�,^���=ޡuh�pE�90�[I�Y�:�]9M�/7�m+�!�s��=N�<�~��j��v����Y����iYM���D4ӿ��7�C�*|�}8FM�}�ڒ�8ٶz���R�S59d(#5�9T0�ye|j�p�����r�$	(]��>���}c��$M2�� �xR�r!c����-�����}@����;|x��}�s	�lŏ{	l`�w�ͼj�C��s.�*M!����`<�K�W%�o��6/W�MPe��>�LN2>�6���e#6�N޽v�����@.�gc��A
�3AdMU?E�k�-���jXB�rXK�\Z�U��S�n�dt�>ޮ79��I���Y�EN����Uڅ��5��7n�r-�W��B뗡�N�'1�R�NR���/�(V�/�;PO��=��^*�tT\�)�4�׽��V�������$��uz�^E��遽e��u��N���;^ۤ�]�^��w�>\h�ԉ� �D���ʰi�`�-�fx���š�h�����_/ÿ2�UT��*��pClXW�(�4����γ��i[u���AN>�WR���������oi��|I�mR�^�F�}4ǣ)FP�[?4�&�zOm=B���������̆O�rH���T��ж����:��?/�뇻�G	�0��(��y�VA,d�/]��IW��5�Vm�t�ͤ�r#%2�r�٣|~�l^�˘�J'Â'y�6��� wh�D�͛@�ϟ���=��US���6Ԩ��GC�[�����ڼf|C"8���}f���ޠيװ���Ӡs鎣9�ޓ�}'g5�SJ��e��6S�QR\�����$=���L�j�]�K��Bij��å������ګ�!�6���B�������fɹeKt7��:���Z�
MN�b�͓|$\��҈i���|�2��h<?ڰ�����o+4W��-C��Դ�#�1�滉�͹�C�D4�.�����T��~��_c ���>��nl$ x>ؠ�8@8�(q��s=�GӾ�����5si����|$��lYn;��3]���}ގ-�<·H��t�Rq� ��"�Ns�;	7;�'6e9ˇ��`5{�Js�VQ�n�:�c3OU���p�z�Rjr*��;�)
��J*�r�?�� ZQQč,s���v��6`݂�Q��9���.���_����r���;>d��t����*瑺V)(���>!�<w
��k]������|��)O��<���:���O��wL�.��f*�DE����^2U�'1TP�Pxa�[�����ɧ鸈�^|4�n�9��5��?�^=D�8.��j���Jem�5�n���dA��އˍ�����? �{9@�x��	/�oj���ϖ0Y��>5�^y���<u��p��Z�sU��0��U����冃}es>�jx	/6�������/��=�I�Q�V�<]��:
���!~���m�\�����fj�b�\��ي�s�����|^(����!�"���K�k����K8�5{����z�1
��!�ɠ`��3� �;�q>�̉S�8�d���L`��i������k֟�&��m/x�<�¥���i:����44��b��n�fK2�4��c�7NbM� �S���	�h�ʍ;t�Ē���B+����n�W
����h�S�r�kXf��a蟀h(�kN7�U�y�^���'ߒ&�m�]d�O�0P��������gu~��uP�zfH�O���{��`>�Ɏc�`���=��if�u_��*�	$�d�7t�Σ�9-���h-�h',�N�QZ*yc/�3�lqO�x�	bTX$%��s@V���j7��Ƥ��1*��6D���:KO��ϫH��HX���d>�i���J�r:���T����Zlƚ�M<[%�瘾�t�Ӎt�S�j��!fI��wY����d:4���رi�E�A���T9�L>����9�f	6y��W� ��2z�I<�Z�3E��ɢ�0�<����Q;�PClTNoL�5j�l�o˕9̣�5�j=�~�� .���4� �c>��<h���b���乄<H�Iw#��������|��MD�ݵ�Q9���7���?YذB��P�{D��6=Z�8�a�C��Ѕ�ӧͤ�r�y��
�)q�� &B�ܫ�7�+�tX ��j�3�j*����/������'��u(|AT�g��n�)��Uz�<�|m7��f�v6��~�1�nnQ
<� #���M[���C�����D �:�.'��k�c~ƛ?��==p����i[��A�RF�7�v���j$�fO�NR!%À�e�_��[�DD�����4�R�u܄5N��ځ=)���̔�&3��b��|6��#�y���{w&ȶ7'���s: ����M�V#��������u��âV�Ť��:8���YԚЄ�����!��"��o��qTS7�@��?ة���B\�	Y�c�,�Uyقk��ZV5�S���gm��=��i�bY���n�ng�C��T.fsߝ�������	�>�n���>��\��b��)�"h�q�{�w�ׁ4#�,d��%�
�	L���������B�6��b����
e��JYÖ�%��k�7T/�����(����*.@6z�@Gk��#v�U4�����n"r��%j���u���״���tP�pxu �KE2�[����z�'�j+��Du
a�j��??��q���oxz��e�u���H6��Q�wk3��Q�$ySVR!�����*�&x���:JEQ�~co��x �
zA7*L�\�x]RX��t-�լ�yGF�������5O�𓣡#	�ƾ�S<*D�tp�Q�	��|�;�91��b��ixBx�]VGڝ7d<�9�J�J����D��T���k��ۡ�n��%��I*z��#h"�R�SV]z�E�xu5�m|�@�2YL���	�,�7Iv#kĩ�ޭ ݔ�9�`K2�"��'X��'	�$ �����leV)R��J~	 ��_q��_\�9�F�)���7�
�xd�r,��&&n�ɫ�+d�U�Ѧ"k�eғ��x��<���;�����5��
�UN�Wc:D���g�#����I�R�Y����ɑVMZ��Ú����)L��}�&;4|{���|r��f�YW��������g������k��\����LLI�����¬����,�U��I~����+c"06��XF��,���ǹ�r�}�
"9���^��ۈP���V2&�P�y9;�R��ة�̚�9?ȳW'���g/���_��P�<���� i�1@��U�T��ONq�7��_%a�z�ϳE)RF�j�:B�lE`��j+�jځ}k�3�����,��ł�9�$N�q�|4j�Mۄj�c��\q=�.1f>�p6��Z��_�} U�b��
+���uMv�Z�4��w0daM^0W�}@J�1 @�lw[�-]�[��k������_ب�K�a��m9�[������56����*-�bFw4v���@5x��O�7+���jl�'����7Ȣt]���c��kQa:5�4 ��xE��P:����������N\�̚B� ����{^
�x�+�&
 p��b��-T��+�i|K
�&Si�԰
bsL����1�pmw/]��1y��u#�����IN{�*�R����H�%]V���8�0�^�Д��Ua�c�1����&Ŷ�>ϗ8�E�|��2��d��:�� ���Uf��J����=�4��k�� ���Y}�E��tMk^�C�uL����x|���
��Z�>zS����mI$F�@~�`MQn�?AS�2�vؕ%���IZ�e����R)^&�?l5"E[$۾�v����ɿ�J�]B�2�z5�hl��aԕ� �	�l���	/�	y�(p��@�޼a9ҿ9D^��M��$�z��
V{w�Ϛ�2�����	M!�En��,x!���H����`�=��1�������M#��bŅ�Q���b���/yY^�!diA�2c_jQ�'�6��R:������RA6�T�/#�9�:�a^���B�RO[u��>6�SP����T\����l\>�@ w��\�������p���?��yFoZJd�"W���25�؞M>���8����546�Ae�����%Q'k�}�]�+��n&%����2�W�Տ�XO����j�-Я���i}"E���H�J��U<�֣���<�m�g�D�R�����W��j�Kȃhu��~��������u54�w.���/nhHY�, 3���Kڂ��bGX(ňH�D�E��%�9y�5'-[����a���xw���T�	��|]ڊЙ�dE�;U\[��(�.�]��?���Uf3�{����a˨�W�Z��ja�ɊJ$o�\�C3�D�I_��'>��!���o�zA\#���?cN�Õ�����u�,.�%�X��l��r�r+)�V�JT��ґ��<#�<��b�������b��߷i��ӯd�I��M�����~��-xAP�����mK�@�h1b���W��L}@����v3����̵ږ��&�?���鑶ӂDEO,)�+�V�ßQ����sx��7�W��ْ~��T�N�~��v��;݋ޫf�+xAyg�:�+���C�H_����\ˍ,��!���ka��V�į'����O�b0�Q*��V�%|y��]K�R>��=���۽E~���6Z�w���0__���&z8C?yC�o�v*����x��������U�N�L�U���+���&2&'�����|�&�<av	��_{��Ƌ��PNN����@*�j︭D�j*␪L�-�`��&�8{{{���W����������R��4���\H&\�(�D>�Uu/O��Ė+DM�������pDX�!
����M=��!�I=�jA'^ճ�>:.~�9^��{�1�-4�^.K�m�'��cb���0Q9w�Q|o�X�76]G(K�L��e~d�10�B����f�9�b�!:Jv[pq� F��!��B7<�d�����X(�b��'��b�(�rF)�
4��)��㣉�7j%2�J�S�\�߿yH�B^�L��kM�RsY����o�gUW�ҫ�2���߸#�,d˼)3���(c�@\���F�!^��˴�=N"�}��`� ͗��T�����0L}Օ������៾�ޚ�_��3����e56i��A�=�Ns���v�mo�f��{��<����ĉQ9�i������@2cޚ�)�@�ZU����\5 h�t�sݬ�6�cӻ_�T���d�+]��F�R��<E���[^4Ӄ�8aڮ�Q�;;���,cbU)���@+�EҼ�x�9��>��ۿ9��g��ZW�N�ռ���!���O����$�!�3:�M��:lT(�Pw�F�>�~��ο���ݫTъ���`��+d<�ĵ5���w����l˸AQ|z����^il�ջ>t���I�]:^+f�/��)΄D�Wi+����wj=��(W7�,ͻ[Ӓ8Ʃ	kfW~�y]�/�Us�o��{�%���>�Ԥ�L�]RjШ⊢����6"�@ �
�<���2t�c;��s�˻VlP$�RS����=���NP.���J'wfm��oAԋ��0޷��?6f�Eϵ���@�i[��{ݲ���ɭSNI���N����\1��q]��(����}�
1�|k�'0�d���&�X	��}7��,kٮ~�2w�L/����f��?�cߘ������`�c��9���2�N�ϊ/X��^�I��l�)G�����%��`��f��׍��1�u�S% D}4���қ}�Bq�E��9�<*�PB���v������>����-4�1Z���p��-rQt���Q, ����O�O����ؿ�͑�/pO��$Q|3ߚOi �+Pݡ����s�*���?W{��\�ț%����ǊO��RF�rF7�z���n۪We��YY�խ�\)��������}��cva u��bOSo�Uoo3�H�=�V�x	E��$������&�jf���13����{����,��VO���L��T,�LWk��r���*wy!JW��YF�b��;�ؚ�������+ז�Y���ɏs����~ŭe�s��OU��z�w�����֯-a]�*t�M����˺HA;'��Π���̃�M��/6K=c�}��;c�5�|||89�cX-vnUU4x�������S�ڤ&�ٌ��Uƙ�W��&\�b�:�£4��V���I�Q#�o}N,�%��jA�ߐД�'���,b7�N�h*+2V	��쐵TN:�֬ˈ��"LH����]�|��eNig)3��}�S,۠�����P,.n�J�!�b5%��XB�a]����*�'ņM�jAZY�����3��_A�j,ろ������1�1����MG�"�C�ȷ��B��c��!a��x��ٌi�_n�U�O544�CYG���9+o���U�;��]�^(��K�@���t�1�u�3��~�4F�X\l�5un����׮ȼ��+"<]j"�gf29wц�H�t	���Mu�"���,���\5<��H��݃!�+Md �0<�{N�l�4��m�t���[,]@���uE�C����Hu_��Q���Ï*w�F��R9����W��ƞ������wKS�?�^t4Yչ>��.��5��9�.��z�
����K�p�"� S����4����2��1��Xt�"y$O]����#�c�K�>}�e0@{Z�-��gJ������Nfu�Qʅ�����]/��\9<��m�ǉCc�*T֬'��i���2O!&�?q�)&��z�f��8)`Э�9t�b�_wF�:d���d�<�!�6�� �=p�j,�e!R��v�&�l���l���1�w��3Wo��k	+\�U��(�	p���s*�7?~�;7����`�� D��������@��n��Pb�{�<����f�3����5�/�u��7�ty'�U���G��-ł�D�<��<�QC�B>dU��E:`2�%ޠ2=;���yȞn} �=;�P�Z�>��@x�Q�[w��t��,�J
���@�=_|�׺����kl����7Ղ9�D�֧WT(��UTYa�ŜM8�R�����]�����G��57�'�n�M�V��򨉪*-j2(� BNM$8'I�C��hK6�(G�BǤ;�lޘ�"��t"��ւ��T�aUL�D峈��;�~Ef�<��}:�+L#9��������%��2�G��hЎf�Gw1s;}�i�p��2�/+��z�(����]g|�� U'_�"�v� '����������B���1�����ƃiz�	0\����,k���w�&�;҅�e����n��(iA�~ʫLM��E�pw�
uJJ����a��y�</�)���E�6� ������ۦ�$䪁��ȟY�򍭎;��l���	�Fw���M���e��3￥*��}(�L/�������1��������O\�k&&��c�QPoѶ	�4V�W{�Z�8W�{N����̎���CH&� �|_O���v{�L�����c��:�w���	�D;��Ֆ�36Ζ��Q�N��l.���%�7������ۈ��3��8�����-m�çO�r�j�bl"A&�%��J�M��<IK�'�7P��D�KCp���@��t	�$)Q3'ׁs��e��͕��*��:(M�l&�7�"Ν�06u�խj�_�A:,-*"�����6����/���Τ��w���������%��+�
�\�Y�$nc�����ޗ~~tB�P2)�R��TY�����N��Ĝ�3�Ɋ"j�K��d�v83��u����b�F����dzc��M~���7U�\�'s}��]��4,�3&tA^"Ť�=E�_Fo�����d��>�r%�wS��p�l�.ʷ�T�h����!;go3_��Pnǲ�D�X'Y]�Ş�'26Z-<�FD��{�x@������)�<m���Q�V4�9)]3r�wŪNw?n���w�ǊhÙMh�jg����/��Ou��B�������E[[i#���E���^�q`=~����-�;��rbiI��[�K�Wy�a\��CZ�BZj��k����y�����'����U�j�0����#L���=��E�eD� ��r���4���݈�d��`�B]�E��s����M��������!�d"N==�Bm�4g��Բi� �Q�]wc�����a;���U�9g��6A�s�R?|o��q'��g*6t����� ���x�^p�ҿts-�����n���q�b�B����~5	j�{;A�3�^q\�R�������ҏ��e����;�z7��m"���
��Uwu1�M�m�����??5ܽ�s	����� �^���%"{\T�k������K:N��kN����^ɿ;}7�g�t�
��NWlh����
����]�}��2��N���}��n$�[���z�����{jd��F�e���O�ӟo����l��� ��SO�^� <_�$�e�W����)���&���h�ɹ�oN*]s��,�e�uMθ-UG��@k[JZ�!��r�a�K���?���%� ;o�\�@�0-M?77��^���I��CDoƄ?�}d��|�x:F1�����sPf�m�v�L�W�ȓ��D#J�>����8���D���q*�ʂ���p*+��c�J�r|���1��>���W9�8L?�H�؞����^�St��M�~��
�u&9s�I$�y�G��X�	n%W�� ��N��Ɔ�?m��̌$ =��&]Z}:����o���4�@	^u�����+H�WG�ظ,e����!KB��FR��㑑Fb����0��U+� S���{ޭ��$�>9��t��G����|����63�s�$`��	Q8e���ػF}�k��aw(��F�YB�����ҿ�|��[������&�/T�vg%�S��
\�Lv?���^��:0��t�q�7.�Jf #];���-6¯(��ǯ���V}-�|^8��!���cP�E[�!l"��0�3��MLDp~N:&:�q���+\ ��r����c���텅��C4��
kZ]^��k�>�����Դ�V{�u!�aR��q�E����!��=!j�M���ے��Z����<�W;��b(�
33�I<�i�m�݅O�n�d����.�C��+�BV7*��/����F;y]ԊVR]�A]�d/?�_/8{ѝ����~W���(B%��~D{A��6@C���dN}��!���C�f�m*��Q�k�C���o	ݯE�A��r�\��}�VC�@�<�D����]E"hI�(	pR�kh�C6E<�2#?���ܐ�x0�_���
ڻ��jf<�	��ڊ��N�u�P$�l+JQN�Js�c4��� ��0�ǶzBH����x99��}���i	��#_��w_Rb<?�+���_���i�pr�:;�D?��:C �5/o�:�%΃���<�H!��x͆O���as���C�9�O�N���^JÖ5���vN �3|ꀜQ���l�p���:qr�w�BO�b���kf�Z��Z ���(�: ��X�.��ZIHw���y���"#W|�e�B^w@ɓ�yk�t��DK�T�Ik#6��z����s�W���OL�*��)I�z^7�>�~p_f����t=���LV���A?W~�gV#堎��Vkw(����mq����Io�8>��_nx�r�3�Eh��.
�ښ[m&l�}F��r���^���u/�������ƛ���GM6$GBJ,Cc,ώ�Bg�tţQ��FuZ`{N�-��unKQ)���M��+�������|Ce�����J9�)Z�Ş��L	���vc#���m��ɥ�LO�]|O�b�2У���D�ʒ���%#B5"b�+���Nݛ������Ҫ��+�$]l��5[�¡�Tٖ��,rxm�������3j�/�/	F�b�b*1�@�J�]F]��D��]N��doT���@��T(��ǔt��{�O���m���)��U����ݒ e���N����$��9I��`vh#�b7��0�QU����ڽ�A]<Iw%]�0f�; ��(h�W�~
�PK   >�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   Ŧ�X�i�R�I �I /   images/5472dc22-a170-4182-a291-403007edeea8.png 5@ʿ�PNG

   IHDR  �  ^   sQ�   sRGB ���    IDATx^��]�u%��?Wկ�P�D"�3$J�ܒ,�d�e�n��vK�����Kv�r[NK����%y[�$�J�2sI�ȁ�(T�U?������`�g��v�����"?������ܳ��'\��^���k3���6���k3��~�?�'�y�$I � nb I����D)�����{m^��3�$TI*���[���p5���8���S�*�3����g�����\}��zJ)�����/��ٽ9Qr�$I̫���\�YPM �Y���ɞ�?�^��y^Y��o`���?�����Z�W-�'Ib=�����Kkm#W�"�DYFdY
!�a%�z^�C�Q0�C��1cS�A)�"�A,�$I'*H��]�+���.-����ڢ�f�+��r�l�4{C)���K� v�
�"k��]�);�'�et;}K��
� 1��5�(_��U� ��7b�M��U���<��+ާT.�����k�P�W���qv���v���;�O �i���T���Jlۆ�����[�ִ�$�-�x�Q�w3I�H����G)#�f�ϘV�Dqdr�q"3�u�P)��9bK���u��c�ʵ��PP����}+nV !�{~.I��q�K��Jg���2\�l7v�-31�wVjK�a�*���Q��M$����{�̕m��e�R�}ˈle�Fd���ŃcF�%c�Z�s�����99�H�����$񽁲3�(h���a(U)�=e�q�j�T���O�Q�b�2���������\�� �`&HL�N�84ݜ�m����r��xx��C� Il�zs<�g�Ʀ�$ʵ�0�c�qel,q�$�} �:����ǆ��R>�>+�� ^$*6c�1#Ӷ�$
�~���Pŉ��0c7��9f^#�|V�|E���]ʴ�����r��ʱ�/@dF��Ï��a�~W�7o�2/�e'ʌbγe9��{�l�08�IĹ��xs_�s�P�C���F��>���5�9�@��4��6,ʹ��ʽ�߷��g���q�$g��f� �l��+���<�C �s}�E�A�I�8.��*xQ�Dv���<�R*ŽA߰m3)�*�l��R����`����D�3�(��2�$N�$6��B���x��`�F��5��3I��gq����be*+v�2e�MeĥJ)�9�P!{�A��$ʰl$�L�4�DI#��A�3B����p�$�8�|&I#��B�^�e�b�4��9lK�V�6���Z�b���wz�\9�3e��T�q=��r�ML�D^`�*V��K"?��f�H��B�2)ӊ�
��%H">'Ts�q�M�(V��\�T&��¢��zA�q��J9,��,�e��k:��(H~�q���\T(���nmi<7t��ؾ����W%�S������G�����sB�#*�� �Tg�*6,q�z�kY��V�^�s̤�lƑ׍L�Xr�R�鈃~F���4��4�p�-ǽn�,��{N�g�g�v��֖jP�;��T+hk8��Z���f�lvz�aRQGV�����X�hԓ��P�T$�a;I��)ߏ�Pu�7Le�Ib�\�
�)e�|>G�z�N#1�8%��ȗ�Fo��T*���n��P�j���T0�C�"_�l�J���PɄ���(�m)�F����/l�H"��W�J�Ȁ�$	�ǆ	SEql�q$� 
�$g�	7����m�����2`h\3ް�?�T��n�o$�Q�T�y^���h������v۲m+	�Q%��(�1�<W�q�(���#��0l�U�c$��q�QS���KhB�1��X��5��v�8��{Q>_�<�C����B�hz�Qä7�(�`�P�����B���m�r�R������M��X��e3���)Ħiҽ3�8E��4D����0*_([�8"$$Q�R����
����˪8�	��LLZV4
�Ģ�(
)(\�$�υ��@U��S���� �冖e
��h�A�5Olۡ�&�B�۶��a#�$��qNT$����wΪ�/�0�4�{~�\�8D�EN�DGA%�J��P"Eȉ���B\/B�xi���n�+j �M�˖UF�����$�^��Ee��Q���J�����ȵ�(�7��k��f��A?H�=�vs.(L��C�RyQ�KŸ�j�q]b����Te��N���I���c�d��b�ʥ$�T����'!�+>'S��Ib��Ǹ?�4��\A%���	uRG����0ʊ�gN6��$��DV�q��0��(4�D���������7���8�L�4��v[ٮ���`���q3�W�</���r����m�=&''U�\�;ݮ��u�n�k��Eʕ2���$��8r,��Ca�}��}_Y�ͧ0FGG~���"��Sl�0�a�f���P��D ]+?���/Z@F���AE��$�m'�^'1L3�L�;D�<	��B���&��Z���H!TTUq��Dsn��܏��;��{65���\v�����}�o������?v��һ�~8��x�v��yt���Pt��N��2z�:r���k��t�R�{mLO��"�R.Ppم~2P�&��ǡŭ��aF��t����(�"
B�nvL
f�P�mێ)�	b�zӥ��91>�9w�v�9h�
/� �T�:w:#�X!7Jj,Ϗ�-Vnm���
�����(Qp��۬��#��;��(0B���2�t��HLz1�laj�4�.����'�ҳ�7,77,��A�c��Ub�U�
���þJ4�m�� 3Fd D^�T��0��'q���*��������$�/��&  1U�aXP�������)�K��a9vL��v��Y��LӔ�E��A��[P�0��f%J�ĴĲ89;1�*Ra�1�^�y/�8�����X@3�'�2o�� *�b�(*���)�2�Ģ'nt[���Y����08^�4m�`Gyi�Z�����h8�\1��*�|6E0OJ��!�#s�L����P1א/ޣ���u�8�cE����1e�k�g�.�f0��-#�I#�n�m�du?��l�b�p���ٶ���|4L��U.���ͦ1R��U��4]�I���:M����	�� �0y-�8��x��X��tU�;H�8�M�]U9SY|�9I[�;��A�H>�g��S�@޴�A��6��Bz�9'�C�ވ��B�-���@��:�*�[7���9����Q(T�f�e
���i��J1�U/��&���sM��v��\�b���@��6]7OyQ��^��]��pn)�_�H�Y��L�a�9������wYLˆ��"o�&e��4��T63�̬ꎑr9�E�^�Q�)�R�����*	����<1���Β���^��m�QKKK��b�~������!��L�x���u�L�e^h{sׯ_/c[^��3r����?�������ʪ��$��|ޥxƦI�!L��.~:�F�R	-S��j�|.j��vy�����e��2�LXF�u�C�I�������{����5p�U臓�y���|�B��r���v�pLy� ����u�p� �k�N�����-\�5�c�u�n�;+0������T#`[����5X\\§>��e}zT�7)=~V6L��9
���D���7b��Xi�!B�ޠ��c�2$^@���pu�·{��	KC0M�nA��i.���\.S�#LBq?N�
0~���Dh	�T��D��`���(���?K���@M� q샌�eF�n��Y�"`RA\$�"�� �c��;L0�/ g�t���Q[�k���ăֈ) � �qe�x��+�P*V0�z��H�c��䳥�=�OUJ~',���u�2>*ΓI&��g"�]HVd
O�0	a8HyT��]��J������#��4T��Ғ<���T2��9�\���h`ݺu�t�J��\S��(��c ^U��afыKr���I�+���h51;;�f�����t�%��V���@&$_��@Qp �����7��g�t���/�����q��1v�YyI�5�s���@�K��s]�=%l��y��^��x�y�H��O����*e[2�NyXu�5��'iؓ���9��؋�B����g�yv+�K�t�WJ����rn�,���z�c��jX�v-����a||ǎC�Z��z�9���G0#�qD��E���ز�E��H0p�=�@4��p���\aJ,1�d���6��D�x�!��|9[�(�C�c�T*��z��1����4�(�����.�}�ޓ����:��df,Ӕq���Q$�U��@�Pޗz��(���H=o z�P�c>�Ȣf'������enŰ� J �C���
Z'Ҩ�m4�1V�5G���̗�+��!$Q%'J�h��]7o����Ի?�G)���S�^u��r#��G��'V�G~x�i�&:+����ț
q�IC^֒�mІ�oa����܉���r�x8"t�NW�M�� �SSS��g?�5k�`rrJ����5���!$��
7�"��S6���f֭=����T$a�ju�v�M���z0�f֬�Ï|_�֓p��0��<l'�7�(�X&��l,w���3,�Vo�^�� ��]4mG �6Q4eQ��I��0 -R�!8+�xmro(�
����F��(3>�j�h�<�{"���(�����X7>	R�Ξ��P�.bl��n��������B,�������`ڴ��䨸,� >n|�,���熊�J��v�Q���%Q0�\�"��=�n�+ �mА��A�/G��L=��9�Tf\�^�#F���(kn�N���Q��5��U66�Pm7?K��|R��P��+W)`*N�'�)�2g᪲��y]�(ށ��-W���MNN��b���C{~�2�*C�@�r�U�34@�{T�a���|Q�|.�|/��Q���ƴ��j�3e�����\�3�[�6	bR���c]�d�;4�Oꁃ�J1\ȴ�i��2�N��Z�ky�z���=a�\Y4��y<p�\<ss�c�]���&���y'�"�}F���&�ͺ�7י�������=�F����w
��������r�;�+�IB���|&ej4�ǫl��^��v����yO�,�.�(��62ഇ�3�m���́�S�ȴ5�l\g�Y�c>_\5Zā���|����)����ؠNku�L���ع���İ�M��"4&�S2ݐL�9�e��ԛ�����s��H�^'�	F��]���8������z�a!T
�<,�cr��|ҩ��7������߾��-J�M�O�z������g}�O7�Zjy�ё���8w�0Z����[��ڍ����i�1=��%^�n��2&Ǉp��1w�<�A�D�P[���L�R���X ���`p��(�N��k��F0P ]���EI��TJ6��y��-TF���
y���Ba��Ǥ������3<��ؼ�f4=�7l؀��)ahM�
�`r��;����E�Ac���r���O�F��:�>s�?��S}��M�{]%Da;���%f�p�έؽm#�N����I�^��B����S������a���SSh�,��'�@%o�6	�6nB���>O扔�� J@%Aϖ�ึ�9 �.�����r�
��{B��J�ʘ������D���J@���U@�:� �Ա�� u�M+"qT|T���rΞ=+��,�� -���*:**o�w>W���xm���Ξ='�@OwaaA��{Q�SΨ(y]��b��zn��O-c�x]*l&�6�-����X���{Fd���[�Q�S�N�(���1�p�8f˲�@ �Ԗ��/��Q�T(��,ǻ��ё1*4�8^�=c\������ɮKy!`� �jP�zj�K�.A�U�z�ɸ�hh�V��,���8��!���1�{0#�4�ȫ o�w+��?A��X����z���X�705=�f�	�g�1`���2�y(�*�3�O�c��賹�#����'3����F�X4�.����a �ɜ��6���^Ȼ�:�@��+C��{��p=��vl�L&�Z&��C�X�CC���y	����<��.
���/��flT�G133#{/��3�teeE��Gc����"?t����8u���3q8Rv��A֧T*���O�8�7�]~V؄4���gr%a�Y5��kfF&��t��i8n�R�	7�OM�z��C���1�|,7�����P`F��L�M�U��S��|�Co|��O�LL��Sy�:@�_Kf�ϯ}総���0ܲ�s�g�����_�nۉ\t�mnݾ������+��=�ܱ��"��+�H���@D��Mμ/ҢJӁ��Kڨ�a�g ����q���:��M��mM�������V>��" �a|b
�KLL��G~����/>��^���)�:y=��P�_��p������sX\\Ď�������7����Yl�ua��<�|�E/���J�0���C(x���
�j�����eL�U��:@�Z-�޻ož�oÚ�2J6��!��D�@I&��(tB����x�E8r��@�Bl�f�/�#W�<ZD� Ցx� �@�Ey�VC�n��طo�=*	7-�xiiy�[��2Kc�(K�5�C�Q���k�}�6?~��(�v�)k�y¼�� �M��|Q�b�u���+���m���l�Ļ�΂md�e��	O�9w�(�;w�8����3�񊗬=t��z����܇�[;�FL^#�%�@�5�G��0�wQĮ���	�4�<��)�����M�B�� xX���3��y/Xd�8�4P����'�ŋѬ7`�#��>׉ʚ�q��)	�8��@�g�����82>h4����w���	h\2%���CehF�Z����ή� Fl��sS�F��Hwz}1��|�����1�=t��p�ޝ8q�i�9�"Ɔ�0��sb�ƣ�7��e�n��?��={d�(G�e��4
	��Iݕih�-ejD��33k��Oh��|O�H�b�* ̂�iP����U�ݰ����[����|������$����8�|1��@��#�aff�>�8�c#:�g�أ<1�������K"�H��M�"�Ө�gVJ��=�9HW��2V�c�䄟#��z|q.*����H�_���Y�;~�����1�I2�����gN��2��2�A&��<�B�E��ը��Y(򝽷�x��9���{���y�QD�c�W��&�|���~��R�m��p.B\>yEx��>�7ݵ���`a�����Cl6B����XZ�������Ҹ��_J�R@��N����+�)eI+��(� R֤�$��83��x
���>IDP�b�ݒ�>R��_#�O�џb�ف��clj
##��w�=�z=l\?�r���?�u;y
c��hu�����������c�(�Q�T�/��H@'�F���ۘ����,3![ׯ�;��Fl�<��3�($��L����ʲ�F����g_<�ǟ|Z<��R��<�ߏJ���n�w�m5e.�0@�����X�����'Fq���q��>C��@���f��Y���d������b��׉Q ��m�4[uy��S(w��5�2�N�A�_�~=v�ލ'N��BE�<��b+��K!<}v�#@D�ea�2֭[�]�v�ĉS2f~�ʃT#�ޛ
Ŷɳ�ʅBN���ebrg7��B�v:4t��>�W�N�c�F{��F=��!9;�[�máC�@���~���A�y��s	�ĉ0��,�j�u��ĥ�s릧�%&������>@�$S�d�(��K�/��ޏ�N4��wm�sy��`B_B�A4�FǪ2_�fC�a�;-�<׃ J���1[�uyxD����Ÿe����(��c�4��b��陵X$�d�Z+�Ӄ�DX3Z����p���8q�y��Fb�Ҽ�B:a~���Dp���T4�p��7�39rD�����J@'�+�wz��gM���P'ݼ�a��y���v8,-_��ҫN9%�E��˺
P&�0~�7o�`jfVVj���%n~�K�������    IDAT��$%,����v����5x��'P���&�7����"����3hS�,��{��l��֬ŉS'eOQ6���iA�Ua�����/!�(<������Oabr.ΡX�a~��֪^H��t���rM����ܗ\�8R"#�VO��H�,��&jK��l��U�����KsX�q�FG�f�L~�ֽ��������QJ[���׫���������W���	�<F�8q�������x����[7��Fހ�	*�<ry�<��..\8+�7i�+�n"
�}H��N� θe� '�u�d
�d�	��IQ�C<�4�a��N�*�{�I��Wo`^+��Ή���'���֬_���*|�MZ1RQG1����T��������8w�"n��n�t�Xn��W_�^�˽X�o*xteI���(K,
<�~�8&FKPa���T���/߉�ދ�|Z�-���Pt�<���a1ʂDl��	��<�/}�a��u�X'�D)��7��jb�� 
O6h�n:e�IqJbXPFǫ���}8r�P�d9z��x#�|T�Y\=ۼ��,�ZYnڴ7޸[ ,��.�� ��w����\���H�͖-[p��7��CW���nW�T����H��x�!����I��X����
�=�=t��@�Q�����4%�2���(��[6bv�,��Q=z��4뢈)�un(�"'80����7�q��s���x��$.\�$�9b
c�\g��`�刲�<�n'��t-^:�_�[���T����I^�N�(u>3���߶m�$�E����=-��������d�t���$IK1�6mڀ��*�W���9&�Q�4I���%����b��߸e&�f���C��`�֭��h�6��+5���p�m�A<X���/`��Y0�c��|��ljΡ0{�`�0{�� y����� �_+&M,%bB?/��B���( ����`�/���D�₀, ��ߌi�e-6n�(2M������9Yw�C(R
'N�ևYH�L�$��v�7o��=�\���� ˋ+b_��+m���g�I<^ظy�lڌ�/[��/2`�Isl�}%ɥ�6��z �u�����أO�::�N�'@��+/���P�]W������e>$I3��=R�OO��ɓ'Q�۸q�N��P[�ƥ��a�wa�7�s_y��p��ض�\z�����_�����b��/��/���ݣ�d��~�r���@:���!�����������o�F����-͋'Ie595*� �w�:���%���
IQeJ�ԭ��K2� _���LL.A�B�Y����D���J+��Z���P��9�u����n_gs
{�?`���(<��o�@��}����ַ�5�n�p����&����훸���{�#ܵ�xϏ��u�ۏ���=�mĥq�XkE�4+0���С Z�����J��/�h�x��>���w��.���bv;�8ƒ�Q'`]j�zT�$��A�J�Ծ�n�ǳ�=����8s�x�:�&:��;�,-J�����t�ĵ�r^�axt��s/�9�~�y	�e� �=�U@�D��ɽ�(��n�	��S9�����Щ0d#��S�wk��
p�Νؿ���$1*�̻�R��ێJɐd.=Om�q�رC�3�;�s�G����c���Z� �K�iʳУ!3��"yʟd�&�ȵ1����NMO��FƂ���Q�Ϝ9���O�F}Qܦ��t�=F��7� ��O=�533��z� K��JNA$����G(�|^��w_��7๧��1z�Y�6�/͡�1W@'=e��H�!R��}}y�����x��ؼ��ʾ#�1}MkK2����R�r��0[�n�cS3x��02:��5���B��b*L���43��;7���
����`��˗.#fވ�d���! ���µf>��}Lϒ θr�#��uX1|%�F�럅]�dA^~�e�����ZmE�[t�l�CĽO����5�w������SO�:6���y�.�K1*�`�X���/�v��~�Nlݺ�?��j&:u
C-�C�H|*�(�:�t���^��^zi5�ι��=��դY)m��2�]����Lcѳ'{F�W+x��Uc2M��[���$��wWw�qy�4�4�P�(r��P)�K'�4bT�9	v�	{t=w�� ��A|��Ϣ�`��-شe#�.]<�{������_�c�^u��R=Y��?���½^�`j�>�������� ^�(�J����cya��fӄ�gϼ����jy�v6�z���g(�,��ă3-�|]�aIl�+V�M&qIbkGi�2A�Yĺ��J�XS�h��=M1R)�$�D�?Ų~�#����a\��1H���Y#Id^����r+Ν9�/�̮߄���/��?������3�7p���K"�n}Ø�4Z�,7��������~Ղ�T��o}��f����]J��E�#�4(I>v~��
��X�DA��h�s�y|�k_��Y^\�J���"��֪ř�)d�lʡ
q��pw�u�=,^_a*�v��
�w3�D���ꘔ��o��FQ���No���s4v��>��c��$0�z��؎C���.�l��P�<J]�s1
i�"��c��W��T�����]˞������K��%�.��������3h���4p$VK@j]9�۬� B�v�V�/� 6����	2\W~�Ư�������`���خ��z�{�	lX7+�<=y��W�jrO��+=�8VR��[�\���n��>&`+U��K.��cY!�،�1[�NQlH{��0�c8��)]3�l 
B�z}1 ���%�r�N[���&4Nn�ša|�����b�$\�� rJ��^3����ؾik��x扇�oՠ��X��6Z�a-}d��Z�^$����1q�w�\�HBc����Pu��~q����`�r-��Cn���Й�@�)�8'KT��;ti����x�f����7��'�Â����	�=Ӻ���кT�RP��o�.��qH�i�39O��Ԡ����}f�=9Fz��]w����"��x��T]M��c]|�%��y2�����RF�/������?���98���Q���]����O�1r��#F#�f��pm���ߕ�[2G̛���n�}�>|��_Eb������q�f\�x�U)��}?��߻w�V�6�A�W�\l�����&���@�TD�oc�ch�.�G��6�a�Mp� ^{΀�R���$�D����KB1�;�J��rUk�ԛ͔���c��E�M*Y�a�A�vb��%��Ip��&�ō)�/�M\�u�R�Y�N�0�%#��9���>&�)zA��7܄`�G!W��.�èז�ҁè-7�凿�V?�{~�������b]8hIf��&���N��J2TI����7|Xa?����}?�/�kv0Q*�ҽ���I=n�,\,%!��S6��t� �� B~��~��Fd	�G��C���^��=<LJ�(A��fI/��i���ܬ%���0Pb��`��������i��TF�J_ZvH ������Q���q�?&ʎ���c��;X����S�g�i���Q��Y�;�;��s�gs�º"wO^�	gT`dx�,@���;�e`�3�
ntt�n�w݀mۯų�<�N`2�9��
�k9XƤs
4D%B��*e1��W��l�(��Y�v<k��d���֕��j���X aӦM���9P��8^�S��_�!�4fhԑ&�x��ge>�g�pᢀv&�N�8�p��JJ�������`�r8t�f֮Em��3�0�n3�b@��c��6�N�ǿ��o"fހJ�4���5��C��2,ybn����w�]���f0403���*׏���ꉎ�RN^��׉�O��d6<_�qiRe�DX��f/�/K#S�n�z0� e����5�!���9�������%�`�1fu�4
$4#�L,��0_�jg��1?Cy&�S��L���ٷ�!����ϐ��kPv9���ۇ�������$A�Av�L�u��!���C1ԋ�SSر};9"��kX�ư���,*y��~�F��,��0]R�1�l����7�+_{Ny�����ci�bob����'�W߸g�ߍ�����O4���_���=�@�5@�5�aO���S����i�m��u�<u\�pQ��$*Q��y�ݒ�����d�+���<�������4�ݜ��%���t�J��(��(,c���`��n� V"��2>o��Y��'��P*��+g�~T( 
���ff� ��a�M���&'�s�.\�8��J�新c�^O���>��u�\�mU;�g�w)y������ӈb�
0T �p������CH��s�4?R�|I���8`��4�a�	6�!=C[��.^���â�9���d^`�ʆg"a���4����ʔz��р���|g^	�Q�R��0!)�d4*0ifPQ�e`��.�<K�mm��)�gFF������ܹG�*�G K4Z-*�\bZ�Ҁ8MF�czB��8zY�.�F���9�$��,��̌�M[6���# �"�g͎�V��R����G'��i�flܸD��%?���JC�$�W�Xi#"%�`�'-*4ҭtR�R�D�>N�X[�&M�4�r	2��z�6\�s���w���Ռ~~��"5��V+K��~�S�S��@p�8�fF+@i�	k��<:P`��t^��{�B��?��;�åK�q�Ai=�y��r�I�
;�m@�v�v�NQ�c�Ҽ��U�ِ&�i�\;������=@DB6���q�yܜ3� p��\�\��o�m���#ݸ��#{,d,h�E�2����]�D��߿_�sΗd�Ǳ\�L�6�4sI�j@�1F���g��+2�
�ϟ%R_�Z�묌��L#������Ҭ~��)��W��o�8�����޳�&|�+_#�L$s-��+:�����8K%�aL�ܶu+>�ߥ���4.�Ma��-��98v�ȼ��ȳM����f���Y��*f���jya�*>�����~��]�/�#����Џԓ���K��ӎ1����$U,�gN`��Q����߱㴽6��/����&�NlD�[�`ia.k-�j�@"}������ߐ�	�������&�l���9�ӋLN����B�c��8%����+]�lvLC�:m�lT0N�����_�����@ J��)����f-n��N��Ma�م��`���/>�%,�t�O�晈TN(w]�IK�
��8qHL��p��a������_� ��&�������pB�|6�禲M�=]J��M�I�-���ӧ��#��(,fms�,/�$KY����G,ㆤmݰD�ɋE�u��R擁w��P�LX��5�Z�/�f5��	��SW�Y<���m�)�o5��1d��}lF�	P�Y�Vbuc�2�dv�*�*?�veM3@'U�m�U��j@'�S�2/DӷJ䉠�9�P	S�>��s���aʜ��c�R��i��͍ziG,�\2Ɋr�y�&�R��k����z(&�?%H�����;zUd�z��h�k0�H#JwK;������y�ק�"��a�Y��\���a�?��%u��3ڗ�#0$��b���N[��AMS���� )�{��*q��f���%�<{I���Jd��/a�Z���[Q[8�'b|�5�=�]�KkřDH������G`&�P^3��.�,�j@��bP1���LKw�q���/�R޹�8gY2eff47���gF"!vb;v��#cX\���h��{���a���l�I<�$����a� �{����r�?Y�~��s^��GE>����؇A*9鹬լ�+�R�Q*av�:)��|d�Ю7E�	�s?1%��hh�P�)��5�g�,j椏by�N�"��$�P����8����-n�iu:����>�M���>�i�F'��؄��8�T�$���O���;�Ig?�^�:@?�Kf��Ï�B���R��iD}���p��q�����u�:��t�0�����P�MF
@��M�vb��C��D�5�t)	�i�c
�O��c�UY�`��&0�s��S�Kf�͛��R��X��BM����EX,�X����f�Z��5�׋� �ϔ���0S�x~��{�c�NH�Y�q���w�G>z��)�������k��Ad��ݗ�`~���� u����/5Vx�iw��x�&�9^so�~�C?�
����Kc���aU���f t�1�}�Q�����/1C�}PA//-�;�vh��ɼS�� -ԠJ���o��q�� +uQ�4̉���jR��z�a���7o��1�`����w�<d�t0�r��1�G�fz͌��	`T*����N�mi�7�yD�*&`�RE�$B�ONL������H�QQ��J�gߗD�1c�rBeŲR��n��R7��y�N��H�Q\*/6��2�	x!��5�شq��)��Y�_��=���f2�N��h|���1����$2cժ����2�y_	Q������G��
�^L�"0s]�,�w�ќd���rV��{g�]�J	o}�[�0�!��K^G!���ںDf$e��1SƦ�yֆ�9�w_x�\�F���������@���=w݉#���,~	�4ure���媄A����-Xy/�1��Ac�c��,��zs����D�P�7�f��0����B?l��,u��e+���96�1_4l�$Z��� ��G��� �Q������v��h������/-c��B?s�,%���~	�p�+�u�YӞ�9+�2c�����
SA��P���FْpS�ѐ��OͲE���]�961����k+5��a�<s
8���~X���0HHM3�Rj�F3���Я�^C!�Ò��������� �N�U3���8|��Zmں7�ً�ni�]D��a�A{��>����=��X._y����d���g�y�ǃT~s���y�ks�-[6�ÎM;��+'1_�G���h����ų���������m�l#��+J{g�m0�8F�Ѱ��׎Vќ��/�����c��m��_���d�\� ۰�k<{�斖0�e3�7m0_jv�cDʔR!fr�ޤA��8�h�|�w~F9��fL�(�+���x�|��k��\��c�N�,A9؅
F��b��C��~^�� އ��x]T�6:�sx����/��{P2x֔�q���)��6��X��.�w
�e�ιI2���?����7�-���|����u���|����,W6���Ȱ�\T�Tr���P���VBY�f�W��-�rY,nz�'NO3�W�J��,7>�q*�@�d���#[�V�B��Y��7�Ki{C�=��X���#�kd5�ҡ�J!������W�$.z�W�)e�q�D&ޤNjJ���&�oT"uf�3�R7���Y2�^"��Y%@�)����̮Y+^��#GV�� ��ԭHӞ�i�3cȆ��a(��TF��V��m�IBhʼPZ8V�7�@��a>���]1A��Ȍ$>_YH��D����paH&3 x���F���%3���|(f�s�ȼ�ϝ� l?���o�/����ݖ��?��}�c��dޚ+u#�n�~�ӑ�67�,�~JyK�X�랻%$#�u�֗9	d���+��]I��66�*��K�x��}?�N��b�,s\o���roJ�g[d����$L ,�0,�s�7������NΑZs�J�I�:$���y�M����?��5�y�OmiE���E&���2ԹV�RI�L9�4�i���F.�%k���Ȍ<����̌[�kB\?�S�Wv���x�,5���փ�%�l�ҰdN �Gؔ&c�h(�<c1�	�̐�+ł��/-��!�l�7�O>�|(M�E��9��0������o���k�����F�'�����(ɡ�B���Rf<@}�\#�Pn�Nv�4pK���;����f�����G1^�H�W�}g�M�$������6��GŐ�����S1�?���ai���2; 3@̿B4�Ę���
��:��    IDAT���$���w�������PU6��������g����~/8
��H�b��a���W�$��.�4�v�Vx�CcӰJC0�xA�5����d��0q��I�Q�ͅ���x��ϼy����G��Z�<�S(/������I��>m>!�t!ݗ~�.���RQ��% Iu�C]_[[B�IM2ș��^zaT
C��'�r�n��W�zL�LEA����r�����z3�]�=�#��-L���q��6b��f�-�|�1e�����g�5���8� �c9�ز�Z���r\�!.��DI,�4��e�.s�I�zbjR��4u?CC�m:3��f�l[g�gYɬ����J��Ⳉ�v��r�3�*�B��f7Y��@J0暌UG�y��2���5ݒ7K�˼Dޛ�ͨ�,S��Y�,����V��CBY"��ga[Z݆�t���xV	�$��u=��W���Q�ie���nX]��ŋs�<��O@;r������K/\e��<%a��?�dkJ���^'� ��$��a���x�f�E$����R�ɜ��R�;��}��<�RE{�4Ĺ�Yr@ M"�3���X���yo����*&�..�D�);�	�I�aeFOXIR�7�t�Ŀ?���霟D���@�,��$?&�)1uۖ{҈`
N��o�>��R�L���R����de|��:Y�:�+L����u��UB�uhq��2�E�av�Z��{�PY*)s��:�W�\�K�����:�߼/<
+_Fuf=jd�r�g;�������� �*s��F����>u��Sk�L�G�Y\�����c(�
e���R�9LOOp�?}����o�ȃ�<��uɂ�FnY��W�\`jbG@AEx����[YB���-��

��M�\Y��$�I�]�.,7��g�Ŧ�q�}�ǩ�94>O��ĄX����@���d��o��������\3��ɩO��\J��
3;���O��#�`�P�N��#�9]��&�]�̼?q�$�D���[��7߿����D��{�:[C7���P9	�*@ϒh�t9��ItД�?���h�F?,e#]��3#U��SV�|	��G��0�arj7ߴW���1�,\n���R�dY�VTv����]��aǶ��?��s�֓
�ʙ�&�.?�Lw6ߡ��i���!���ӧOiO!�{�)N+t��J&�%��&�Y�?������_��#��M����l��(jB���}w�u��'��K�K��$��K������`����J�/}��-�6�gE�c�<��Y� ;�I���`��v�����C��LkvJLGa�8v #C�-��s%�w�4l����W��r�r	/�? ��DŐ�tE�3"IT�f\��M�ds̸'���t�c�Ҭ��Be��4������6�3J�6i/��|��@�铟�$>�ψ!B@������$\��@c$K���ה;�=N�\e�#���~p�Y?�Ò��Ga������NqL���=B���M���M��:���}.Y��s��?Ęݺc�<?�"�&24�wR��XE� _��r�$�^w�-���c�yT�{]�ac�Ҽܟ�{iP�Y\���9.�'���)ϬN�����J�@;IYÙ�0�<s�{4,XSO��w���$U; �w���LQ�fa� ���o[�J�d���z�D��a�"������19�C#�xq�AT�'����p��'8��+��������U�~��l���y�?\�����!�o`˚x��G ���q���I*��J���n�7���w�¹S8u���-g9W�C��e�HPjS�in-��n�_6\<y�<�*E����%���m,_�����	�
�-��W_~������kw����u�G�ulGw�S�蹱%���o��
���ش��R� ���dV����a�TC�g��%�<�u�XK�X��W<�D��2{Y��+g��V�xPõ�F������4�Czȱ�.=���'������
��]@|�r�ֶT*�l�O|⏰0��˗�P_i�Z~�ՙ���i�L�b�nY)M%�X6<7)7$�6��5��y�F��J�	c�c�qi�9��P��|�I�����+�ݮ *�J憧\�0���:++5Z����<��.=n����oX�^���8���F��_ ��&=
�ns=d	�T��I0==)-M��e9`%���Y��>Z��' �H �ʑ�睴2�8��Ǒ���y��Y��Y��~��e5��P����N?�;Q�<Y�XJ�$�/�K�{R���W �¹��.��X���Go�c�<���� �� ��s�]�9J|&���1u�#��*�kp�y�!�����0[)	���c��>s3��HX��{�B�ݖ�������k��x8w<+��GØIT�NG �?gc�����&�>E� ;24,)���С)]�%�I"\���r.�'A�G�f%�4B���2�TI�A�2bP[����?i	�K8P��uk�<���<I�c/	ʢ�C�Kr��O7L��i�DF�$Z4X�9��1�(�˦0b���0���y-�#�C��?S�d^:׋7Y��A"͔U�d�-��˟�i_�gV>ǰ�ypt��.}#s�}��rf��y�n*#��v���i��g���+cv�u8�� ����~����_xﭻ�\i�������?��l��_}�W��}�* bkӕ&�zcy�������G����H9גX1����Q�8��E���2��6�E�w�����^���סv�fG�M��2ʅ�4���$ **iP���l'/\���;�o}�����t�e��8s�<f֮����e<�9���Wpi~�]B�4
ǥ��{gg�ryH�k9�V��������`+��pO`���pu8�R��q�v;O���W�nՑwx:R�������}���� �v���{0��T.^O�WOO�"��֡�s�8�v�_��W���R�Vw�b)���0�R�,l��6f&'d�Kr���K��4��S�4�J+����l���
�%9|���M&�^3#L �ᱝ�ã�+!���-̾�M�,[֣���L,���V�XXX��PYփ/*���Y*}�D[�+����⭉��	��"�D%�z��	��C3�iZh���1�Vb��Y̚m`ƾ�+�`���P�3��
���$ ��I*w>{֠E{�,U�DL.b2e�Aw���1��W+4L�#��ug#����Y�7��������5��ݱ܊��\��E18�3��	����^��Y	��[���{��9��!���?3p�5��4'=��	<��7�[dm��s��ܜ;wF�l����Z�������)zu�����L��,E֓_��:�nd��|�z���tV�BY'��3������w�`� :BJ�v�,&&�$�e�̑`�2������B��i�'����ц�>@��LYɚ]�m ��^�L��x�i�)Ku����`\5k���[��`�љl����\#���8����J�����bVӈl�t�"��e�Z9?!y��ٹ��F��a\d) �b�N��.�dB9t��R	������y3�/�,�����z�Ov`%�`�q�3�6I�Ӆ�PN#��0�hB��P���W~��?��� ����r��/|�|�-]2��BgiU׆4���7ྻ�c�Hy��g{X�>�	^ǏB��:R©G`�ޔ�|�~'�#n��|��!����ќ����F�.���>�g��C�ﶣ�=?D�݆�0�<��<��C_�"~�~��C���t�E��H���4��~�Ku(�E�8"��
q�h��x�[߁w����'���?�	�n#� n����5�(V��h$c�%^�󡓘^�Nl�p�4*a���_�����bv��<�d���=���m��\��ݥn>"t��- �z�|�+_������J1KΨ(���y}�}�W.V�����j41Qeh[��NZ֕y��q��eYa����铞�咀���P�+���L�bk5�bq��
�I+x���:���j:�T���$��������_/�y��I���Ln*pR��s�1�6z~|6Z�R��Ö�� L�t�e��Ԁ☲#��� Tx��e�ٳH�Q��gh����(U�x�f�&����N��:Q~��:�;��ڽ.�~�˖�����sҹ���J{Sf�K*gZ�ϳ�,CV:'DDC��s|���hu8M�S�I��s�ߥ�f��kĥs�3xf(so���b��jc��5���/��;J��j��yr�4� r6�&l��`��F���&�$�069�A� (�������:���~�[��ޟ�b��i4}���瞽w��U�����͚ж%N�]��jy<GFj��;_Cԡ��W�r��5ȇ�cPɴ WV�=�=Jt<>>�&��ȌԦ���Q�/�c���'�b�%i�0}w�WB%�N�	"4B����z%�D�����11�!~ҭ��W���(i$����J2,/¢/�t&��4G���r��<8�P�`�]wAG�X��i6�$G
�� r��5JG2�
�p]�W��B��1mc�����1��]O�_��6I��.B}c�V�D����nɈ����i�p�D%�L7M.h�G�A�l��%	y|F����w��;}�p8��1	�3���l��tD5�La*�5������^W>v?�%���[���T�����u��j��ٗ�����	k����� ��
Y��1?�[LoB.�G�D
��V�UX[E�D[� ��q�i.]Ҕ�)�JfD�ٺ�%��I�2{zV�����\�̌�@e* f|�\Mqmd"Q5̅$-Y}<�ƛ�<{[l��.�f�:x�!d
y�(/u�����q���� ��a�X����>9�Wq�o/�n{l#G�cv��֚�ǣ?Ҭ�[�	O[UX����9�j�f>�_�M�q�D[SW]~��95^�/p3��V�sȹ�WN?*9�ŀ^v�/\��>���q�\�K}�ƺzi��z���ȌF�j�W���;�� �G`�Q��(�%����MV��s�D:��f�(�\G�	x?�ԃ#�� XJ
7
:iq�:���/��� �x�q�1>�i�2f���8��N&uNDr�aE���x"!$RҒlܢ�2P�٤���^g��;�/V\���?W`����Xd�
҅!�YqV�d��#A�Ӛi����M���ȳ��:�eU����>�M�l�afg����mɉv\��iY�&8�
�H=j�lh�;��B����x��z���vu�(�m
�b�ܼ���b7
�ݽ��6ySZV��~����U:��<'��);n�ͬ�ypƆ���Y���ꔒ�|�TPx ����;��|"V�_��ۨ?VK,l
����WǙ8`��Z��A$R�6(a�ϋ$�dj~��RB{�R��`\�\s���"�_�v�8I��z�w&A��I��{�Ă|A���\�:oGS��k�Fl�>'����n�j����.��A�,q�j�5������Ug����č$X�I&@j�V�"�9��g��p��l���
��ID�Ї����Ux�ߝ;ﻀ>*C����v��oܵ1[>8����*���Ơ�l?��c��k[p���~]Hql����|� M�d��f�
)?���I#�Lal�e�����w�����0��C]�*d��f`wk�3�
���|Mt3}x�_��7>�r8�+V�;�Ǳ���]�ʤ��fe%/v͛�J���j,�j���j���ԆL�"���G�3�:D�o��I<M�`�H=RL���c�"�U�p;�E�uV��3v�%X��ӉukW��!�H��������T\z�9�jR�lS����z�Y٪���O�KЃ��} kA�������X�b��.z�w�߈�Z��ͤP�XH��j���:�3Uu*�M���K�egcw�n�
lN��d
^���E�w�;�yA���Y�S~�7�IS'�g�̟�swo�H�($�q�y������S���?<�`����[o��u�QGc������@�@�U��:�]ׯY�p("�԰����a�����+��[������͜Ƿ����5nPDc�9HX���
����ʲ�	3��7�-8�fT�&����M�a��r._D'�����j�H���z��������߱��s5	n���W�b!'fMX�m�ؠ��Ii��Z��V��ɒc�b��c4ю׎A`��U҆��4��y�#f���Q��a���eH3p��l����'�S�$���`��`Y��""@�2V��.�n� �k�����4XAɰ��%�\'��F|fI<����&���hD�6?�QϏ3ݢ���㘱��uת����w܁�T� 9�V���e)��X�Z��/ϋ���g�v"�� ���h���]OB�F�}�=�{��	B�T�p��,��?U�\;T�db&�,"�����u��/��'JK��B�x�1�L�g�����z����+.>뻀>�b/�W'���W��ɹ��$c]���>���>������;mM��l�TV}�@���|��3466�TΡs�ZUhdbV	�J�Il{K>}�]l;uZk��ő昙�#_d��-��`�l�.&B="��H�3(���ە,Up��?��x%�c�)m#W({�b�_q�^�\���k��R�͇D:�1�:��λ�Y����#R�,ȽP�i����15-v�!%q��lY��L:�x<�"j"^��7\�m���3O�fu:;|r���iVC:aU�D�TD*_@���+���n���X�z�4	�n�ڳ/��مtrH��A� ��UH�3�:BЦ"s��y=�T�V�D�����y8M"ez ��s��m `E� Ξ�*�G�O|�^t��C�M؎J�Xd�3H��ƫ
��\�r������ YJI�ޛ~��H8���'���/�xB�-���KV�ֳ��O���& ̌�b���\*%BY��hؼ4bK�a6si�ԩ�>Dbc��d��	y�2���y#�_�]��1a���qF�
F˚���@�<���I�!ӓ��v&����U�2��`�Q�x���zu�>`�Φ��ĕVs�W����鏣��h؊�V�����SX�)�e7kr�!?昼o4M�H��*O�?�3*e��?|_�CS�+���MgS�9cK��Ձ?�C>[�oH�rGBg�M�0�����S���Dq]m�H���$~��BQߝ����6!?�����U2�~1�`ߚ��V#�N�թ8��a}�\|�Ŏ51���"��P�JQ��lo���Uy(����������[`�4����-bUGZ�\�L�G�\CZ�{n��?�
��}�*�m�`[�@ȯn�Ȫ�~����(�x�e{�֪:��lS@�����r}�?�N�練�({�Ε<�f��X��w�����o�����.�Y���%F��7�~��	&41�%	�В�&R��wKc���Cl=��Ѡ���{{t��S�+��/�q�H���d�f1��!��bњ��˗��aG�3�>1)��Y&n.�2.��J,]��P[P����<��Igs���X��9so������Y(�HM\��1��L�������^��&��F4�G�D��;�m���~|��z�5Iu�����j�T��՝�>v�,g����E�d�7��=����V,!�#9Ї�`<ܰK9�a`��:Mp�:�T�b��i�i*�w>�{���٘�o�w?�>B�%tVcƬ��`�����ѣ|�]w2�����A�o�����ˤ�3�|����/���� �gܙN9������ ��K�=3vu���'�T��AX���A��IA6�FCm�>+|n�V��"��'�Pr��䁉	+�#?R�u<67�X4�$����#��>����
��A��B-�o�����|,Ú�	h/���}�y��l�ȶ��0)�w
~ؠ��h�0��3�B���b���|�#&��s�	W�g���6���p���$6`�n���}4 �’l�\�+�VG    IDAT���֥�`@ <]�b�=��a�jd���C������������z��B>�i�5�!O���'�n>�LA��K���r�?�G6��{��g�}^�C�{�XSR6�C�!�l���z�u�)������e��g f��k��a�r� Q����M��^c���L���K(r3�s���;A�3���gm�mfo�� ��K��33N����_�F@U� �ʶ����4��H3۪����܎�s�	��y�17��5":��ٲMˑ_�-�i��B�{6�b{��0տ��p!�!$'A/R�pc���(�P]/\}��~2g����<����u=��r�|��+�=Y�n6i*�{���Y�p���c��D!���!� H9-8[ۚ��[C�-��$����
n�_}� ��0��	Y�.�S�r�2TP��0#�a������i�sEd=,Y�k��ã�E�?��i��TW���Q������
,Z�5|���t(��üP�CT�2����M��@2WF��A��5�ml�
�V5j�[�*���l�lc�1�)0�ߋtfH��UBJ9�6Ű�6�������Sڴ����朸��U�
$R���E�j�Jt����A"�CooJL[����������K��4���΁������CB�2��7UM��@�/�QY�;��M���"!�v�S>��p��S[o\�XI�vc�f�aC����;$�z2��'�<9"_z�g�4�l�[o�]Jv�6���1 0��� �pȑ�����TnG�RiB���O�Qm��	mr�r�^�B,�t���-��"Z[��g��\ �?7!Ul��DBA���ly-�;�v�K�D�ؒ�6��F^O,&I� �J��D(��5����c���&������dՓ�ϭ�����|}]C���7�#�_n��m�O���lT�7*���g-D?���dB������:2�;�����fT�wL?^{	׹��I��p�6�a[�S����'�A�5��n]�L�j�Y��hZ�a�z�6I��`K���ʦ�deg}J�����n%�\�dċt��k�h�s�
�1U��
��c$���|�|�룎<�r>[��W_{Ӧ�Ę�"�1c������8\/V��V���i��+0Cԃ�юn�5������7_o�m<��]g�,�C���F���+Z��ir�e4Y��>�,0��6�G����U�.75WQ����"A�p�����dδ���X>ސ�~�so�9���Ud��+�)A9Gvx#~��6�w��($�����ۥ��J)�����0~�8V�Z�P�T�d�����26���˿A ��N[�D׺��sd*OU��9ʅ8K�+�fD�d�d�^��Y��n���>�yo���0P�\��>�|��Lb��~���sl���U0a�4�L��|�>�A�|A�(�ɹZxPr��
� \�_�V�m�b��|�o� �M�?;�biӹq���C{}UDbn��l@��Ŗ�'cڔ�h���������C*�A���39t�'�He��x5(W��T������&��N ��P7\��4��]L@�jv<��d�P�&l��moL��G	����\�h�bzg���0׭ݠ~8�eYI�#��`,A�G�@��(�����6�on��>�,ZZ��|��*�y�R�I��}G�K��)x_�\�/�9�<�1��P���0֠v��p+8V���6���
`���W�G.��^�c1dhAj��N��=Y̸��hp���-$���v�LoX��W������#�,�U�hvKJ��YiV��t{$��m���#�����Gv����r��
8|�qlP1S]�f�k�V��)�6ꏎO������G�k���`oߙ�߄�p�7P���zcbö[JTV���^'�l�X�4Lb�u�Zf��@�s�ƹM2�r��,i��?9-<�J6��{�ѹ���#��i�CĀ�ɱ/��[��޿�}�O�P��BQ!����ͬ���3�|�L6���z
�]qJe�JZ���uA{&����<�Z%N!�`m�r�X���?g�z�ʜEUl@���v���L�f�-{���:����kI!;{:��r���h��s>Z���8���!�)F�S-�B���ͯ}��ӿc�ۀ�Aon�ߞx����)�C��h�H�� �C]��޳q�>["� �d�K���1�N�U.a��-�ª�%#� UT����/��� �}�!��cW�3)�	+��Q�L#��QeR��QΉn��ٯ�4�W����/a�.{`��["M7�0���u�s��ƥ�]�ϿX�hi�ں&.���n��1`x�c�^x�Qj����j�>$�}ʌ�z	En7U6�(��p�Ňe�*5$?����2u<\�R�^��D|��+�{Ɇ�"��`(��'E \K���)d�U�#�Jd�i���VD�,�]jh�� �Uq��I�ˡT,�^�R�kl�����l�2�a�1�q�_䩚�:1�����_.Z����+���� 8��/�=�P�{�Z�RŁ�)�C�2��πN�>V�d���:�����\s������4���2�����T҆j��E0sLI�����u����6�2P1�sl��U�2�O��ц�m�v��I���e�1�=P�q��2_)�TE���0I��+n�1^w*�Q	������)�6�'i���*�Y�A� p���O�VF�^�gl7qڄ�jF!���l�����|��	��P�Q��,��q���sr�����T���*�k�$(�&��y]y}��Go�v��&�����;�,g����xXb�%X���k�,�Ό�G�sM%8��7����QI i�;G%��1��e�k����w&�b�(Pm1��D
��`��7�4&�\��M����z��.��=^{�M$��#1�g#�����;>`,`�@mu�-��̈́�׍�)t��A�6��q?�|<�D�J}�9����e���o�w�v����f����w�">#K�8�q���<�Ī�ʡ^\$��h���A1��x�o���w��� ��Nz���p��+V�(�JV��sQ�f�X��d�(�R�Puh�lV�$am=k&2��6�G���D(�I���5~/�|�.��i���V䆇�*{B�M���d}�W2������L��������,� �1�"���^vz8n�T���ҕW�˾])��/F ���'���B\cS�t+�Q����ԩ:f0�]�F��|����x�KZqڸ4{����EM�2
�xJ�D�(璈��h� �@&�����^ZVP�x�!,]ۂ|�T���C:_��i��^.7�D| �La?�:�:�8�ݩk_4�F�@X�H����2�|^b,R��jMY����2����e��D�y���1e�4445ᕗ_ø���kہ_�������ۅƦt"Bg_���TY��?7w�\m������{O_?��hhn��=��:�8�`�z�(��zc;�8�0nX��͂��hR7���q]�!TIV>�s��e�꫒�hF�(f��-��w�+�ꉚX�6�^�'+'
�2#����\;�y,~�Þ��^��
qN �wI�j���+sC�d�C���
��~���n�#n@���M���X���WB3�nZ��n�kzx>�l�0`A)"Z��9��QX"eS��wU7jKQe3��aB[�
�n��m��?#J�s���klP���#e6�Sit�D�q£ Q-Nި��t��+7CL ���]B"Fd�sƔ#j�Q[K�y���9P��7:� �p�qz��|��JHe�/���i���J�,bb�x��k�uk֔�0������� oӜ?�S�kh��LP�>Hh\�Xs<!=L8�@��ߙ �J^DBGSj���웒͇�2��n�Z�ᚚ������aWu�}ϼt�@%07�
"7�r�6̧U��-t{�TQ�$�b�l��,�a���H��йa��լ�sٔnt����q��W*���.�Vӧ���^[�^kM0$/vn�.G���l̓:������o �|� {�� 4����]}h7^z�P02�P�W��]����X��.�Ʉi=L
ՐG��Z$/K)j�{|[�G���R�c�7�"�.F8䃻B� �z���h��,Ԋ5!T�L�,xC��9�}U���PJ`���(��Ӛ3�C�nN�FFB��d��/��Z̚5�ب��cՊo�n��mmB:E��<*�#���GE���2�b|�Wn��(�bfY�V������A����k��<a�$s�	"'=��c�4q�!�}�O���
ֻ�<����ڰ�FC��x\s��䌚XZ?N���sDv#bC#��R2cP��Mb�S}�RtDaL�¯"�kG$����o�w7�lL:L�'�l�T���7a%@ܨ��/d�:���� i
p�EL���$��r�:o�,�7��ܜP��0�л}f��u�X�:U�ZKNϖ0n���`ʏJ��&��r;Om�Ò�F�[L6�&���e>���Aǎӹ��>z�NLr��>��y�θ?%x�}�`GX�&e�k���p�R�;�f9��ꙥ�N�P􇗆��DR	;c�O�5�}qĲ�~�/�v�@T��0V^�gd�[	�S��Ϧ�❫�h,fP4Ώ��Z(�-h�Kn5I��n"=Ӝ�%��p@x��=�� �ᵆ6���kIϺ�v&f�����O�!-�p��i��eǍ�S\����G%���ً�d1�s�b��8�� ��� &D�S)�՗����s���G=Mve'>��w�WBs3U?�E �L�C��|F�� a"WY�0�#�u�_�͖�p�qG��gr�!�B@��1f�dT�rfZ�L3V������j�d ���TF��'oz�ЊU����J�TF��GwrO��*v�e7��>��3 I�Xc�3Y��E��$n��H������R,�f�Z��4��A��x�-U��[�8x�HgJ��4�ɍ}�X}k������4�Ķz�|����˒|U+��G�����NeKX��+V첯����S&�ú��b���.@��[z�����&��r���T=H�����Sa��g�=�Z�\�?�q8D(��2yU�����6�L++�P0��5+V�{'�9��{�L&�/M���7D�yœ�����΅��+������)��#8蠃��s��믾�I?��f�/��%�ѡjj���h�<U��mm6C��ѯ��+��=�Ｍ�m1cKL�6�>�<��C"{�jee��kZ���0�+UrA��;��ԲpH8�xa�hbSj�s�$)J!-Hh�#_�ha����Ȟ�<R$����#��L�ژisƁ,���Մ�����F(2g:	o��<ܰM�l���|h�/W{�n���޻.���g��ʙ�;U����37oa�͗	��7Di8�XS��D(����`* n�j)d�:�
&��H�"ڌ�@�\q��A0�*r���f*@^OB��E�{����X��W.���:�~~&o�y3CI�67 ��"�븙l
�u�� �59.c%��Z�=Gcj3��Qb��kI1�2+b�v%�4�ŖmB�F��򴆨VA(lf��E�#~��Y���z���TrK����"w���E��
[���X�:�1I��M�O!���GI��m�~p��� 9B��8�3�:jf��(��8�3���	���|�x�� �.�������MR�`��e '�J7�5����є�X�j������8�;a�Q}��섻�y�ξrd�l��=d��np���R�*2��K��B�J5Q2���6�i�L�t""��DH���0��2~^{�d���sP��k�
�54!�H:paU08�0Hv�n���N|�pf��{�3}�a�����ߞ���R�]�,��d�ӄ��K/�K/Ek�d�e�Ň0a�d�C����P>��ĵ��}��@�PUPoj�@ C��twnD]Ћ�-Q\rީh��RΠ��\*��A���eu��W�8v<������U�~�ͧNE6����?���&�l\����M'���7��n/�u�
$�PT�Π��ЀH(��˗Jk���E=nhʸe�\�b�@6=�H��-s#��*�2gǶ�K[[��!jOW%���47% ���\�ZkǸ	Hf��s�}��koi��0+V���)������п���m��3�k���
{�|�m�ɍ�Ǖ L��Q�����ѿ?,V2�{\��v���'��c�z'*���V=V�jT�6�t*�����9�1Š�HE*�?�1QԆ	M��I�bl!yŵ S�"6Lv(
"'@�5��A�U��*8c�U����m����[7��Q#T%"W�踰�q�ot"Y�x���ճ/��$W*5�9�l�ッ#������)�t����P؆V�2��ufp��e@03�&�6D5�n$�{����PR3*@()p�+m����Tb�=�m�Ur:�낏�����Ֆ��\��� *r��}�34dl�h�C�d�&��A��U�-5A���(��I/(u����ؙo�s�t���ֳ �@�����)%GGJ8�J8�M#xc�mF&98�XS��~��u��s�Tv#i��1{��HF�*�vv�~�?=0����u?��R�_��v��cZ˜R`��U�̈́�$SL�xx�ę�9�i;0xrP.0���pWb HU���X�rUd1�	�ף�v!�*`����xمg�������N��o��[ퟫ���#N��U����څJ.#R\9��[Tm1tu��>����Z�)jk��l6iE;չ��
��X��l=kW��:�oi��� �L¯ L�"�y*�������D��:6��;�@�Y��t���ǸͰ�5LW�/�M�ˮ���_!�A$Z�b��3>.V�Qy,�!W(+x����E�5����P�׬G[CB�$�:�8Lۈ��fg�ks#ap��E��@�H�7�u���ٍ�K�bζ���O>@����I�Nı�C,,��X��%P,�>��I5��v��M�����M�Ɩ3675����Ԉ+�t&��jgsbE�J%�W@�̑.
�p��}$��o��6x}��]�8��5#m"����;c���˅�E���s��_����$�>s뭴2xs���P�jK�.�?R�E�7ɵ��Y�2���{�_饗b���rb�����?���x�T��t��(�s�om	�r�Y0�if�
O�ܳ\k~�H��H���0�*�5Lb�6$�*�"E����T���*rڸ�F���;��wn^�l Rm��(�&���;mp����x$"b��g�#RR1�kU��紆_	R��B�&�1H0uG29�^1�3Ʌ:�h�mQ�ݨ�5�S����B�T�ؒplo�T�V�T�R�Z����M[����GɘZ�_�Œ�~	�3�!�K=�Io�[$Q��M'3hӊޞ�w4;�eϑ�CD��	Q���:i��Ւ�r��,"�I+ôrz9FJ$ŧ�9�%soxlJ9�BZ�Nl2�3���Q�ڪ��&>L��HsDN�Gި�1�`E#y��[[�u��y>�|�y|Fm����mmB9��S���M��������I�CChjm���N4��4�&)T����kZE&����<9Ob�P��E%a�.�]d�LK����~���Udp��mGu�ӅS�ps�ເ>*���_	�������&�Z)Pf��u#��ZF�M�w�tN��b>�B6�R!�#~t fL��T�^�#	 �IGD�������ӵ,B]0���X�t)ܬ"�Y�h�!���r��Hf3hnmAǔI�|�������%сb�8�<a�h�X�>��au��^e�_~%��f%B�Dcu7��=�(2��{�Jg��
>��B��'��+�"x�!4��A6S�ؖ�)�vީ�bj���k�r�r��Λ
$�b
F��2v��ZI���鏏��=�@�q����������Ť��������H�<��a�["RS���^m�+��¸�c�L�2Y��|�|�_��ޗ3GÔ�k\�>�du{��78�Ǿ�[�;��Cp��)X�"    IDAT
� M@��_�f��6,_��(�Q�R��;Oi���ݍ����L��E�kj��8��� �����oV,���{0��@GF;=�Ǐ��wݣM�ni��Ѓ�0�-]��N<Q6�W_}��
�3_O8�Wg��Xm-��{�طl��q�a�sC�+&7����747֒4F��4�\I:
D4)AF6Mn�����_��l�dF�X�RŁ�9W˪D��N��@�f�RU*v�)Om���T��J.8w-�;��"��~�"�J�� *܅�&@:	{����咪B��: �h5�'a�7�y�-��*8���c�	����$��$)��?{�����{m���3�%�?��9������Emȅ��\�v�ZU�s]-W���B�ҷ��=98���F�Le��I�ܧ����2g��VK��r��¢��U}���!l��>y<�<�M�� !w��Yl�fb�H�*1d��k��3ْ��c5�Q�V�4�i���DM����ƶ�;�۹.m����;��c#�=�?��1�|GҺu���Rm��p8$L⍜���B�
n\�U^?J�d¢��ϼ&��R���`���|9Rޖs�uHЎ� �i%����0	 $����G��U@G5Wl�^��B����qwv�=Ͽ5?^���9�r>�(�\�b��=s:22CC�|��E�R
�PΧ��R���.��9|������J����	3�b��\�T]��W�\-���hlmAS{3b55p���ú�]���!��L��RU�a�kA���ͩ��{�.GOw?|� �.���ނ��'�ù� 	lƺ���]=�����!��Z�ח�G�}	�?�hЇ�7�?��<�k㛯a�ڕ�d��>�PV�H��'�x��7�Œo�6f�t�/��y��?Œ�_���y�`����٧�`��5x��bٷ+�٤]�*;�q��˵�	
!w���6�l~s��H	~{�����o
��&@!tU�nZ��VX���_}�5hh��5����p���%	��(KJ��dN�w0�PU_u��qc�~��'M#5�B]mN��i��]z/V���'�����G�o�^~�6�h��8n��h����>���W������FÒ�_�K�k���U��?c�L�Њ%YG)�����|+L2��~����KhmoC&�����ʥ�Î(G4�2Uu��rf8�`�1j!/@�b1t�~�CV����f��#�C��cFa�A�T�E�̨���&tuv"H����2P	��X�Ѐ��.�,������\*U��-`�ƥ�:���͠	�<o��)GXѣ�	+0�� aN���0���qc�M+ϑ�z�̝18+�c��,���Љ.��1c���e˾�$v��LvlDƎ��H���{L_���oa�so`�wi����������J��!o�x�Lb�{�T�î/r�)gb�E/��o���|������r��usC������
-�M��V}#L����s8M��M��T�.C|8�L�b���*��]�֡}�x�Gk������ئڰ�SI��uk�4�ɑ��w��vx������'� '?�9���>:��7�S�q	�e�S�[- ������Q�]�Ǖ���=3�5HSY0����` �DKG��E�j����Þ����ٿ>r��4i�����O)��:�_��D�RH�.D�d��0��/���l�}6��E�_�,ii�AA���N�	~'JS.u2m
	2s��Wh��pЌxQƕ�-i����QC�^��8օ�QA:��&;Lӄh_@pt"�B��y���Ud���4�ι�?��3��@1G��c�v�A�iם��ڈ�dB�}���hikC0X������ c�MA"��-��C��iȦ�����0��ݝ�@�&Foƍ��Ȩ�r��w>�����{q�����%���Q�$q�Eb�mfc��/��k����Gwo�a���UҚZD*���7�<��,�Z�q��c��w���&�y�'�z�H=r��騳R�bρ�*S7h��ꪫ$���������7v���AJT���۟L���j�� ���Ki�󼆆S�a���78���܋/h�>}*�O�/��`�}��v�yW���S�F1v�xͤSz�r�ܔv�e'\|�E�͈+Be����!��λ�ۃ��1����$lD��4��Fe�� ɂ����'2n�D��$����yn��l��E����_1�����Y���+�m��àJ�a�ZA'a���ղ�	�g�+n����u�Z�.jjb�Z�͍2��3g��+^W��u��A����D���b�;I5�/�c�E�}&O�e�H%�q�J�N���b}�m?�Θ�P���K���a̟;��~{������[�l�2�5��I�*5+=� 
���tV�|��iӦᣏ>�믿�Q.���y�d���n�1x�L��o�EE���ˍ��n��>]�{܄�X��k�pT����A�����V��j��p��n��<�hXE U��^�Ԑ
y�jkGFC��#�NB��&�p˹��'o6��sN9��X��r�4�a8G�1�w�
!���5
��X]�]Y��?/[g��8�V���p^�����}��5�������V��R���O<Q�̃>������i��)���5שIR�J]��K�@�Vq�I,��4����i�SO=��X�z���x
���?x���
T�Lg%�M^�T�`��*:^��7��]@�˼�S�����Gt.���a\�8�������<�:���#�f��Xk׬p�7�j��8VR)�˰��M�2�z��\n~DCU/�DJ��p	���W��l�"�9_{��(�p|��GWO��m�}��C�c �~��*P�3%�)U��ѥ�p�U����6}�^�h�WH�r��4!i@o_
��m���f��g_Cm�8�h-{��W��ރ\2�H�o��>����L!C}�r��)n��N��E��O=�x��gѵq&t��fӦa|�X��.x�g��Ob�FƊ
4���5�Ɠ��NINt h"B��쮻�/��>5+O'H���z=�K�53+�J��Y�fa�	X�x�����z��U-�:����W� .]qf�/>�<fo��$+fڢN�:;�#�|�imz�hoiiÃ�]=�=��x0~=�|m�mc0y�d�]�]]�:/&MM:���^mT��'bAh�S�@XY�B�x���RQ��D&M��j��iS��a�]w�����x��tބ�1qM�<I�d��K%1c���|�i�֊��zNm	Μ�|�)X�d	>���	~$�יM���$�#"�k!h�/��d�$TI��O$�P߀drX�{��gk��a8N�VUu��t��� �h����$��u�$��#u�e�갤9���a��EN�=��ǵ�k�Ɗ�� ����CԵ��{p/��"�{���k�E$Vk����ᦩ��]o�t]R���Ar�f���k�ꫯ�z���?V�H���֩�cPa��9I#�a���Ԛ�T�붝=�7{��9�%0��M�L���&�H#=g
R���nL�8�'N��）��~�a�g�\��ч�~��?8�+���==;~�,���9�u��}�]1}�4�����t��rk�Tȇ������E#0<�a��-岪v��2#����n{�g��Ɋ�ͷ���5F^�_l�0��q� 2�/_�� N��/�o9���ѷa#���&,�v9��vD�[M;�i%� �Č(*]ݒi�Lh���IZ��J�$�	���J�(���0e
��n<�����X�f�>#�mgo�c�9g��WZ�[l��x2��^��hMC�o��!TC�*�o�^�⢳���O{���~��;�!� ���Cy��N���v����n�o���UA_��nxk[�6��� Z[���G�	���-���g*FE�r���<`����U�K%�J�8���e�0W1��"���Y�r1slL��^*���/Z���t�[�1m��z����_/]���v��B�Mx�ŗ1,BL=�u�#�c��h3	���]1e�AW�;��"/��-�b�T�����`ђ/��'#�9w�|�C�}!l��v
��<�j0�����H'ND�رx㭷�"ŖC2�Ѧ����˅��V���E�nB�x]np4� q�W^��"�0Z�vv���kd�KL��18���I��۽�K�ǌ\�d��J��2�P����>V�.MK≔>ϳ��f^���iӱϾ����^զ��>�h���VҶ�~����s睯�7g��L:���u�0{�Y����M���>{�LT��L�2O=�,n��VL�2=}�#�`J��3�p��8����g�R�:�������G���O��Љ+��C���0B!F���ub�8�z�M�z�Bm�3gn�x ���
���T��^��ͿS�M1���K!�],����~���LH�;SЦOM{~)H8?�����~�>n��I��W��/<���[��g�c�m�!\O%?�E�q7
�x<�~�98��3��_��'��8=�0�p�	���+0c�L�������4���fYI\��v�LK��=��sx衇������a�}�A8餓q��?E��a$�$A�R#��i��ӏ���u�B���><��c�46�����ե���%	�]9ҭ�벷�2v�M����}���3���e����W+랻���̝wމ��+��74!O�1	bU=<4��v�'��x���pؑG*�:�����߯�Ы�t���k�t-�13�k�yw1�����p޹�b�]wÆ���'	�'ʲp�b�e� ~��Q�Ԩ�E5F>�z���C��矏���/X�r%���r|�٧��;��o��W���mY���o��y��XI�\�B �ߏ���约?���8�C������7�3��.��:���/ttLP�͖"�n�$�V�ǟxF{5�Aԡ��A�:�\?>�P��g�~:b5&���᪢������L�'L�˯���>��~��� �A�j��b@�KW\tּ�*�Q�ӡ��{�y��x5���A�]En��8�Gs��GK?�y�r9����s�����|�l��C;�C)�-�*�@�:��25�-�>3ko<7�p�ƌp�WUUEȗ�)����de!e"
J8��A�?!e�ԇ'�;_B&�Ess�=�<A�<�j�������'�|@�l��t��6���=�����Rه�T�`��Y$�e<�سՎC���j������#x��'��X�X8�x| .O._�7`�=�F*�CW!��$^��{ӦLl��J�x����ꚙ;{�C��~�H7T2�yM�X۝��0�5�` �
h�Z�I�\+�U��gDv97�χ,[��6�^CC����@L8�~��7v�)a�����Ѝ���]��aG���&��Xe��֋,�de츉����㮻�[�Ǡ��M����~o����a��Z��8���a�a�m��G��w�� �ׯGsS+r�������E����I���c�³Ͻ��ϛO�$7?��~�i�{�-h�0	���xM�6�ñ����7N8�0D���& ��ч�-�]���_	˵�^��,�>yl	׸��v�	��|%�z�3L�a�ӽ>��-�c�0]~��ذ���ӄ3=P��l�cZq�e���SNRF�:o����w�y��<�l�e<c��V�"�䢋d.��7Z3é�&���z��p�}���/���?��7x�Oi�;��������⨣�Bb0����.�/��R.�u$9�G8��
G����<�9'"F�Q����-w�w�D���B�4��3����8Lnl��/�����Z�u��̥��;�+�;�h�u��hmiju�'Hz���g��:�CD#5�9��/�=�M�}�����]�O��λ ��m����9���n{�c�;V�E�UZm��3��3���e���8唓��/c��/Uٟy�Yj��>���TK��JR�������}�y�4~����?�`P\��wݥ$�"N<�C~���>��%]x����>�#��vst��z�����VqLxND����Q,��#�T��3� ���Z�,��MSs����^~� �L�C��j�'���`�]v����Pk��{�*�ƦF�Srh�\{-jcu�s��e7���N�~�=���D
N�
�47#Tä%�k)������{�����_�z���p?:j���~�al}���b�+E��'��Фj���F�t�~��B2�!qLB�B��\6���0B�g!3��h��v�����){��l]I+))�q1f(�Ax�m�$tq�S��vk���^�����y睯�7��9������I�1cBa?Ǝmǝ������x"�b%�����o�/��>B�F�����[O��/?@��eh��!�R���#W�a�}�@cS���GQ){��&�={�m��/���Đ��e�����o��xb��1:fD&�a�Mn��Q[���d�g�<�L��`@�V�ʈ�q&���7!K��u����.F��)���#|�׺]�5�`���L���l�Ĵ�&�Q#i������B�A��=d�O��|��//A&]@sK�z���׬Y�M���Um�>��=!'�t���'�z�!�N��@Xo6_�z`��FC��w_�΍�q�_��_��dI�Z#�s�ʕ���Gt�W��h�0Q�?����
�{&O��_�}�����{�k�x��d���`�����|���D2-�/�'�g������U��k�k�&`uM�|�,�[�|^P	mx�-�2����}�]x�o�#��,�:�I%�����'���㌳���]�HW�4+��{셓N�.�w>�}�!f�+�r�-��˱b�J�����'W�M���<&����H�ǿ���U��;��c1<��o�[#Wz�u���_���<e���(���M��*�5�Κ`������7��<򈮱��&,��:q�x%��s"��Z,z&����w�q;���#B%��#���;��oH1����Q���nD(L���<�n���`o���8���p�a����$��^�Xm�L�N;�t����˓��3��Hg�"���kwW�F��͘�.���J4�����c�j�*%��;Y�9�sf���{����NS[�_�뮻_}�}�a��a\ӍZk�s4�ј)�2Iw���'����N���ի�tI���'�G��n�	Ͻ��Ө�@M�HX�F|�FԵ�c޼yX�z����5����d�`X�RI�#��?B!���V��o�����v��y!��7��;�:�4�q�Y�;w6�3���7` 1�`4� �6o@=�j5�k��^���_]�]@���My��7o����r�^�+��/�Q;o5��A��*X�b�z�\,��X�p���!^�%q#�D"7UIV*"����?� 
�%�fo�3�F1���4�Ƹ�$�3b��c(���A�QLؘ��´ڣ��U�.���L�l��ǵ��1�CKk"� �o6Y���_���S�c���ۡm��u�#x��Ռ�(�"�ɡ÷Ht�)A1�B|�-mM(yJ�{�\=��V�E_� ~��c���fN�����o�
b�P)��4ȝ��F�ۣ���T�y]��._R�rF{�e��V��v�8!4&2$�I������r���U79�E��v�AE2�9>���
ٰ�Ȥo�9�ဃ�Z�fr��V�Z�9sv�g��o�}��~�;��4b�$rL@X�Ujkk����^\p�<��Nx橧q�����g ���R�y�t�����C.ˤ��~�v�=w�9"��*L�in7^~�̟���혠Ġ���(ƕK�z��p޹��g���%%By=�p}��B��}�=̿�nMp]rΛk���wae��؀��n��V�U�4�	����S�Ҙqz#��uC)�:��4~q���������#�"�aVo7�p#�x�5Js�����Y\UD�A�s���z��Wp�������sq��7Hy����{.�lG����9>�@,�=�ޥj�n��{�Alͺ��?>�|�L�չ [��U8�FIa3�o�B�]&/&��g�U){Ƭ`�|���aA    IDAT�d �)����BV��$�H�>�TG+0�����"�9q تc5��<O��s�x2�1�:4y�� app@I��O�U��_-Z�9��F�����B����8��G��OW��>*V���]'ǆ�T4�-�S#�B��9�����瞣DH�5��� "Q\�]����c�-f��SNAc[�H�@wo
��y�Y!w�9M�-fl1L�n���y�x���%�hR6��A����ǟD#[z�f���FK������A>�Lv5�i�?a�����9"�×�l.�L����fD�x�m���TA�;�����?�p���<us�^�^�-��
��PE�����6F�/^v�i~�G��ܔ_x�AWtn��qe��h�1ܹ����~2�:����kW��B�`�� 	�20*�!�Ǻ	�f�Ae֧�>�"N����]�
!J\V��Ф�*7"V8T_#DC�O�i�Ce��rc1ښ�@�B�<��8N\���ٝĘ��U}�O4��rW���3$���߇/�;N�l,Z�-��X���ga������8���0���̚[B(f�Z���h�D�G�H+V}��fL�b�6�w�/=����	gwܱbt��*%T%�S��V̨��v��qR�g��
(f���drsC��TÜ� �E��(�u�2y4���B'�����mU��,,��J=c*K^V��;���)��� ���y�������y�჏?REqܱ�K$�k���]U���G6SD]}�O���6*�`b�����n;c���R榛o��u�- $��; ,/{B��>hd���,�l��LUkW���a2����z��eK��mhjVbJ�s����℟�����=�|�M��O����X��_=n��v��a��	H9J}⏠�z4DM�� 792�)�Bh�'
���h7N~M�pv�x|��Ֆ8��`�iSu})OJ=r.��j���G��$���}vY���h�����'�]V�o��.�|�v�����Y��[��0F���f�l�q1�S%�՚+l��|o/6�a�&0>���$5�����
�M���*q#H�%=�i�$��DG�Z^K"T\ol�����Z�Ye*�9+���E0��� &ut`�Y[+ rP'�g����:������D�Bʧr��z\r&;9�9��B����I�p�����>���S����՚�sӘq��'�<��&Z��8ɬ��qF��`´����#ͥR�gQ����	��:e�$�����Ŕ�[E>�x�O<��kX��ψ�(��&��#~���yCS�Ú��H�q^w>�|o�oYْ��D�R4�ud�rB��h�T���Q�،B�����I�k��&�ճ=H�h'S�4������-J�%mc�����H�r�+������ƈ����?��C��C��?��M��ŷn�F�W����x?��G�ذ�L���v�	�AB^,��c,Y�í����A{LΌRel��?�.T�D��<�(W��a�F�cg�lh�҇Q1�C��U��������Gg dχsߔ*�֘L�^���B�(����6�b �����p晧c�}vG6��"��� A��nMmV���|��x{}�@�˼���}��s`�у,�ׯ@���Z�y�w#	�eb+��5o��&�������}b��B��Y��*�{��C�����5r2n¬G'ALN�ڊ�& V��w���������ـΤ��Xo_��v����DD��3���0U+#n$k7tb����eW\��\�����><���[������;8� �������(�:8�w����T�1&f_-]�]w�7�|J�V~�u���]bR���ށw����t�\����$o��I4��q���T)0��܎���|�J���X�}l��dE����B<�VM�"Ι g�!V�LNm���FJ�r��C1Z�B}D*~1Y3��P�ؑO����.�3:�^�>��E���$��v�y��!)�5�6��B }Љb��N�1Ne�\D|���ԉ�G#����ᚘd��:�G<oLPf�3F:B@��Rl��(�y��׵���#�i��ӛW�TZ���u^A��G�5:����b���|� �2iͽS�_L8ҩ$~/B>/J�RH����=�� �<m���54�">d�I�9 �z�*����o����ͭm��J���d6����Q�3�"�w�t�i[U�%4�4��X&�6a���33�r>׍��d�\���L؆b��I��\{��sm)&#|ny���~M��g@�*���.)`˘Y�H���"BK�wmmz����$�F2L&��`��$�	��e.�����k���O�L�@
�0�c�ԢB)�*Gv����R���'��p��^6��W�ƅ�燾)��ۗ����߾y�����fox �ލh�	��b��5X��B�����a�|�T���c@���,�T�{�;{�4�}*�:3Rnb|(w�iw	�|��ڸ(���NK� Af��]���D8�s�n��ׯWe��n��K�yl􊩿�Uu�M�f�����QR�Y�𮜫�s��(EeL�F_ǜF1+PǬAE�`(buDAAAɠ�:wu�\��>Ͻ���������緦�N��s��g��3F�\^t�r&>3	��o��鑙gf����2���֖Vds�v��`(���6�����S�ByU���[�X=�p��T��΍kP�s;j
}�d��[Mh���Y�@YU�����M[PU\-�W�˂���ʬ��W^)��۷KbLs�$?D8d�Gs��b$\(
z��YY���uKP�M���,�Q!V i5�S��P�ҳgv���v����C�(�\+y�(���sC�n���>|��;P����L¾�ѭGw���ly�}�����{�AyM5�l�!!�""7�����ڂ�Ε8���ok�3NO0�'Ӗ���fl߱����Y��y|b
��Ĭ&�M�ga�f�9��u���!o��$���hW�J��HD"��T����	LH�^%�A�U&Gj���+�<X��R��.U�^]*+)���&<+�xRY��e0�8ؠZVr�RIq�(��� ��f�ʍ�'�����T-��N��RѩZz�<W���ě�>�Nx�� �����O��b�Z�E�j^���u��ZR�;߀C�Td��Z��8���)"
��<���l�H�!��qj�k�O~h�5+���[����n����:�x�*6*z=�y\�����Q �:�����seI	��؎Qw�.�w��7d�F8}�H���F�r�Nf�$�6Vk�&a�0�Ո��YZ-�0���;TTu�����6n�Od�r-qܖ\��%@�2U�P�}6���B�ع��`5#�PJw�	&���.<1��}"Y�Z>[R'���8��U�p�TB/4�I��8���I4�
9���	+r��)�."&CM��Br�(�w�}'�������ZɄU*sJq�dD�*��x&+d�	��w����N'��o�H�b6X@�Nzu0Yr�
�6����M.)v�y�Q_>���?���:a�%M��o}������̦X8�	��c7D�Ӂ�=���Ѝn]:�������>��
�o�A��0�k�; Ai͚ղ�8o�@��_*�(���5k���E(.)��"��(߸\�0y1q!�p�CvN�}�r�
V���V����ʜ�M��	��9t���_���u�֭�T����:U��*mTD�ѣ����._��m���Mm1X�>�.������!":�Vt�R���.�����+��r@��}p8�EN��R���^1�ڽ3>R���}�b�[A�k��O+�^YkY5���	P�D�F����7����ڦ��km3��oq�b%t*�4�mf����=���x*���G�>0��A&�9Q(Ŷ��� ����3N��͸������&�1�v����*� 8�O�D�����+䆲��Dc��<�駟��ƍ_�w�|�w.F�~��~|��gX�z-≌<��y�<�9n�YA%R���E
���u�	o�U0O$�&#�3����%�j^'>&[����r��+4j0�],�-I$��	(��LPc� N<�xL��4֬Z�@��p^��X
6�L�����!cC���:kjnD.�B׮���3�D(�GYq	\.nh&��j��ǅ?aۮ݈PX�S�w7۔~6{���+,+��b��-���D5�x��1"��qR��f�� r%�*h�X�e��.��M&	x�09f��%1�M&��Z��Җ���5�����1?]���Ɉt4&�H�r�_�Ty̅J��W��r��P3�҈�`���B��d�@*�ù�~�g&MƢ�K$���*���@%/��o�^�)8iDb�v��o�ŗ^�7�,{��I����V���F�[Z[b��ٓ�/|&'��ױ�b�
�,3|@��R�Z �M3��]+�9���ЭY��vl޼_�� ��j9�:�AT�栃�%�������y�R�I|x����;�1�S��It#$B�i)�h2f��;��qa��%�6}�W%���q��s����1��7�[j��?�!|�ŏ���3�w`��M�."�4bcv{d��B[i�
�Fc<R��W�G����Gu��?����4�/|��s�����Ę%K�0��@��F��t��B$D�NŢd�bE��Qy�� /������He+kQ��k��C��'��߈�bq�JĔ4'�M�#'���(2�xԢ�&�T��D �xnM-���c�j#tB~.�k����-d����E.���!r1@�18v:������ohjBUM�;�OqB��B��u�^+��>�G�/@�=�VR��ߏ.�:!�#�p���bB.m��-�ѹSg����O���Ǳ��M���T�=�
T�&��\�L�϶�G�����d@'�@f�5�+�	+�Q;ɮi�C�
�z�|��r�����!J�����BV\�LJ��b�>�b�<,	C�`�u�4���̄�((*���,)g��4۱u�L�4�T�{��ʁf$�2p� L��(�͙�pF\���g��H����>��~߈��'=0h����ˡ����*�����Q68�:�[f�|�6nES+�fKE�����v����3
���@��v�(��K@w�1c�`�Ͽ����Y�2Gx���F:ǝ�SHV��t#lV�f$"1�z�����-,*x�1����τ���1��X��6D����#��K��x���X��g�HFc 4Y�p��Mv�¢R�);-&a��s���շ���z���@-r�$�����V��a0P׌Ra$dO�Ya�Ո��h��¥��Ȏ��/o'Đc�>�ۛ�<���4�E{ޢ�~�1��� {�d)0a`¯�ݳ� ��ϝM����}�}�q���z�������
�χd� ��a{"����>���H��C��Z�r�1�閛����,���+���� %�̉��r�+a�"�ucB�c�*P��$�����G8�Z�����0�IgP��`*��#Zߜ�sIf�.�'t�M�	�ص��n�D��!.�D��җ��m/%}˖�=�P�2��c��WЧWOiW�@�~��w�h�W�iuM�>zG��b��M�E��\6�/�Pr?|�@ȔL
R����3$ձ�6}��X,�YL(�q�]�j������{�е#��9���yK��3�3q�����@�}*���a�ɱ��
M'���qK�T3]:w�{�o���H��[�n���ND�޽1u���R�G� ���ǐ!��7�Pu�	����K�%��0�͛�3�|:,&��̀��k��Dq�U�l�{���T:�����L�M�s��'�()*GkK�E�ƍ��Q4~!D��[ҒYd$H��Ml�"���A��̇�1��o��ݱ���G��;2� �LR�2��҈��q��a:�4����s��~���]Ke)���p���qy�ǫV
��33�Q*����-��Z�<�L\�y� ���N��\Nzp܄	���X9�������I��u��U��u|�T��6mQ:�F#�+	E�E�иUP =5	�m�w��^�|�c�C�r{� H��X,�ݛ7���n���'|���by_���C��G�տ��L~^�g�ر�XǠΊ[6T��`)�1y�d��{n"TA$�(��\��LN�[��3���N��H6���c������c��K�V�<��HL��*�[2��UR���/��o۴�Ņ����4,r��s�[���27T��r�|a��x��G�o����}�ek��^f��q��Ew{�5�b�u�Qx���q��c維(����X�R�AÈT�U>:�AT�i#���m����[��_�fB����渚�u�s�D���]7pQ2���~��^U�@�6[��Լ�)|����#u�?�x����0e�(��|4e���O(~�{q��:�� |:�M<��d,��GQn�uN��1�;r(ď^}�����*m0�4��QR��xy�����;4���a�b��q�W�3f�PZ�ڋ��B����kimy/����:�<�|�M�Z-t�����`�k/�ȁ]�f�&��� ��gϮX��
<���r<���b� #"�`NM�q�<��8Q�:�����0v�}���o0~�3���'�ƛGa�+�b��=�:<���@�$�8j�/o��`�%C��֯��;��K������_P�s�-{!���dBJ2G6-�5]��HrK"	�=!��T��dX�[�b��M0��0K5������� ,�$zv�"�?��A���C�=2�D�a����[	��}�T)�=2�Y�V�O���ի�JOH�۲j��	Ӹ5؆��r�	��?k�`k(���%No��óR �Dn�b��*��;F�d���eBʨ�銆�Z���ߍ���^]ˀdV�Y�X,GZK�dD���g�v��(
<.�t�	"ky��cdѬ�m:w���P��*=mr�QTUt�@��H%�+*�7yA|Vk�DN����EƱf��9Uޗ���ܢ>r(�V$R1e�B��*�q���J�	�0h�4��q�fAC�5�R��+&�-F�`v�ٯL/������i(�>jV�^�W_�)A��PDqx�9�؁��+���b�J�)�h�g�s�۳GTʸ��~��$��t�SH^�Py��� �r��W���A}}���yK�ə��g�M�l]�$u��-++�&�g��T|���7�h�*��d%���U���h\+O!�Zfv3��Ze�/	��
��&<�G
ʪ6Z+G�q��i�2�d0�^��TV��x�4&9�x�l.�J�#2Jp�3,ʳ�?p@�RV�F�G�@��u�P�9Hu��#��G��oxLt3&��Y��y �yN���ӂ:É��߫c!�����_O1���@>3���D`4��*�V4����ǈG��M��-*��N�r�6���lZ�S��ғ�#F:B$n�9@/2��=�e���)����T�@`�,å~ͨ��{@��;�׫'�M{\pY��n<�4�޻=/��u�lG?��S>o{�����%!Sȳ��������Ϣ�Uxc�L)*�|r4^���hH��",[��>�h��2-�%���
���sѹƂ��>'���O�[o|�M����'���Ȁ�x�_ ����HE:�^n%I\e@��c̽�=��
=o�?���ɂ��Yߙ���D��
a�Tz@'�����)	쪪��W*Au�D^�)�`eA#�H�!��W�ߖ/qy��h u����9ڣܡ��ӆ��ry,�	���mKNs�3a2�i�1�X�I�0���"D����*������q�kG�����uz@�}��s�dQչ�V+��B,]�3L�(
�Y�x~�*B"@9���B�Vd�Iࡁ̕W���m�D����N��%KЭ�])���+ǉI�҄��`K��엟����G��3�M�Ϡ볣��^��{�b��"ժ>�����LS�^`>-��:�NFaȶ�� h+���6l޴UHB�jh��\|�3�����-ҝ3    IDAT����莞}z�y�ĢE?a���6�!Ɏ$V��������S���[o�!�"� .@ѿU�r�}�9"{��/����wa�����DMu¡B~+)�R�=s�����X��
X�c2�$� Q��K���m�YhFyY�ҧeD>V�4�#\�ϴ�(��+.�"�pZ��=^��~�= ���)�u��x�Е��=��K�?���L�l�Br�H~"]�hW����
���f5e=��1p� ���[2�E�����Ѕ�G9������(�+Bc�!������m�=.�H~�z��W�vܱC/V}���^}�Yw͘Vz�PΦ���.�]��[o�Y���7I����H	k��?����IJ��⦼���1J��n�^d2��������ڗ{5����q}("�v�����gIN$�Q��*���9��&M�q�Y��
��i5�'�~{&�1^����ש�����W�܀�N]{��NR3�c�Ptk�3�i�Z�y�a�И2eF\+V�^%�"H]w�H� `+D�Y�E�|���$p��#1n�X�Lf�۳5U5"�L�I�nx�w0��Ũoj��������-Z`wR��%�,�}��ݷ=~�1=������������%���~�`���PҤ ��Ҋ=���@2s2%|"2��d�q�a�s�fV	8,�/5IROD��˓�I��p�$H� ��e3��0#l�!���`�ݻtF�.]E��b�Jy�I'"`���Pb��RU�^�N�%΀fѩ�
���^��4�p�fv���FS��Q8�?K!E�UxB�x=��$�-{6p����dî�}��ňN%N7��Ք瀣.-M�BZ�5�l�!	J���o~F6c��a�q��}{�J��&\�|2W�#
v(��A	���Q2Г��*��w΁��&�9��	 gV�}��%nP���Եyv{J�2`��j�	��}�w�`�Fn"&��8X�-;D��6Ie${�ǝ,��GA�V���u���.�u�����G�8^GD乡�3җ��>��>J�V��T��b��o��/��0�	Z�-��{�"����M�]��qg���q��n2�P��z��f7!Iy��QR^��H\�wY�q�Kgg+��V]����:K�9#;���	��2��'EN�6?����r�>5y_C�\��)��x�G�����u�b�Vw�~v]c�Rc��z0W�9���b��p�@�b� �^����)Qn�+��>��RB��AB����+�����+�\���\���u|=�됰���Z�$¥b�z]ٻ���w\+�QMĈ|i���F���)�v�|rM�\��9�V��au��6��f�%���l�B�Bg��`�oAe*�	2��9O�g>$�R�
�y�����&0xK��8���d�x��wa�"��D���Ηc���˃�k�GG ׯ=�s�qRH�Ҙ-Lx�2n6pP_��nR�6\t饘>�Q\|��v�+��jE#��BW�W��P�J����O���=�@K�$�N����|��s�EH���1�I�N����&98�`�"���m��	�W�w�B�.X�b �=%�����3���� �;��i$RQ؜!�p�����M����s�8�6V9��1��B-�~$��+$4�ۄ-	�!���SE1�uH'0n�K�a��D�`�O����~X�^b�a ��*/X2n��sL�}j��^=��B���b��&,Y�;,����i�;�7/>��&�ƤU\�f#�����6lZ��:W����ڴQL�8L�������Ń0X2����4�}�,��{1hБ"t� Lm�SO=U�^�?�x�צ�g�eC�f�IL��j$=d�����C�Ś5k��Ҭ����3�38����+aei�b�iO�%�"����ޗs�22����}&m@��������P��I���b����pD�>BZ����������1�c��-"
Dd2AŮ�9Oa��m���M6R�꘠:D8;vlÂ���A2+�t� ��)�3߷���l��hj��M�?G�����1F�F��;%m��3��5�VO4�qDjyٯf> �-d*S��� R1���|�Ck��x4����o���.!j^D87L�Srg�Q�GV����x�͌��0a⳨����r��`�{'Df�~�B�$�i�-2��k�h��\Y_Zw��_�r�G������WM揾������v��	)�~�������R�§�ȈV�3���>3I}Y�Hh?KI�L�xD:�MD�2E��v5EC�@Z3��%��2��1��&��kR�}
���W����l���b�F�S|�<H�=l_�tg�X�*�����i��v��`�I��p0$��:/�jQ
�C�ȕ��={�
���]��p��]
V���$�>ZZ�p�%�����}�>��֭W��Y3M��cP~�D�y�O�I��p��v���6�Ww������/>���Df�s�]�"ŵEn�g&/�o�1�'�U���'���o��~���C(89�V�����d��̉4i%2�,�/,��4b3`�đK�PRH�vV���.��}C�[�k��H�q,f�(�"��'b��,��ҋ��';��4���1��#���eK�a��[��19^@C�3�n(�j�{�#P[׊�M)|�p)���EK�dq�N��`\���3�YN���	=z�����l��ȍL̏P�.lߴNS��V2�ɚqZ��)x}�@Vmv�C�t��Xq�u��jie�d��Ѯ��
o�⢪���}0�f�ق`�N3��$(PC�����/��5{�ܰ)�I��[t�S)q}�ݻ��M�	a�gR��	�j�A	�d2��1�>�46�a���b���KQ1Z��B8��
Y�g�}6�=&�5]:c��/��N,��l��F�����*�(+QJEr���ǲ��l�:nqT���+��M��N���>YQ1��iim(>N_u�'���h6`�s�yV�Jz�&�6��(����|�uK5�m�z�T�&���Si+�\M���J1�@ ���[�%����YTuRc6���!���e�3DYq��n����	Q�4��C`m�R4�����"c�&ɯ�U&�����^������x�#�=��6}���?���5�#Y~���FoW����3��,=t�B�����g�eu��?�wF5Ä�;!r�yS�G,G.y,��*��pPo�#��bpf� 2�lOqM;�"�+�m�O�&����'�����ׯ�N��9��w��qˊ��\�����F��
Y����;�� �{b��{&�B��jl�X�>���2,�w/�x���(�����}Z�NA�d��� ���짓pM�����M#oļo����Γd�k3C�����Ԯ�`$!�:V��$CUE�ϟ��?�����#��[�R�'G��v���4v�L�L�dpr�$k��hȢ�"H�j��n�`���h�߇P[Z������U'��PRZ���߷#�#�B}c���]V���pYӸ�Α�ݥ
V�<�q�54I0j�b����n}}�������N4��.��@��M�6a���8��s����~�z�߼�di���v�n���huA�-C�fd@�~}eV;��c:�ӌ?;{U��v'�
�pYmpظиȹ��Dכ���?��PF?8[͌��[o%��r����1�%�Gf@��COr�D�b�@!m�ۜjs��v������F;K�+�s�w�2��8.z�Zd쭰P����)��S2}���O�@� /l{q�S�De��v���`��5(,)��rfѬtH2"٨���kkQRR�ʚj�r�ip� y�}�9V._%�"��J
K��uS��.@�bH�jm��b����d�t��gI'��}"Ra�}b� JկX��5�-��XْpE�Z#�Qe,��q�e��f7QA�}s�X���:�4-�g;��U����x��w��g��Ků(Eo�Ra�!��.-�!e`ʨ)7�t2�N��p�T�s�(I���#u8n��:�4r���r"���m��ǽ��e�I��*v��4�`{�նT=B�ˋ!z6�oA�h.ljF1u���H�������.�=h�o'r���v�@%i5�yt��LJb-�;=D����'�����Ev�P�f�RY�Y%-���oN��IU>
�p �cj�`�B��st���~����TA!N3�u۫y�ӳBm3�e�D�W�3Q�Cnz?^]�ڟ� }An�O��7�y��%I�c�b�A� �H�B��� a��чsd�"I\C��J�%9`��ҳvt�*�0%��2�D�n�L���1dfi�2��زڔ�+v��-ɅՖVZ>��[��).��r��ݯ/EP0,��("��(����Y؜�0����m���Vc
U�����O�QU^�݌�}��BIq�doNwj��ď?��W���x�&��?��Ѓh�NK
��y#���ːC��v�D!G��Y���R��7�ܰi@"�\�?�/2~����.CUU'\y���v��c�*l� �昏��A�탌P�*C�B�Zga���̥���#�G��V���H�|�~��F�-��B�Z7�b�0�.���jt:=���1����pDϮ�ׯ�lDtTc �Bf����_|Y��)P����iMK�
�0�2�s���B	SV��a�M}q. V��8���X�1��>|,��������i��V���˗K��ǋ0F&+��Mͭ8��3��Œe+P^Q���u�� ��mO�b�N�W�Ed:C���3���b���{�1�RUΈ6�_F��*�����8�F��H�gz�NDCmȤ���(�y�������L6��;w�kcS3.��JaǞHQ
7kB$�E(�F$�E��T�5r���B&1]R��B�~X�0��#<b�$�x���u�dCW��#i�퍑��g�=\P!�n�UA�q&^�I׉���K�}ܨ�����+زe��2U*n�<�zUO6�{�R��!;�UR(oq����LojEfbU��8��C���8�?���mD�a���y�_˃șH�u�9H�R���ɏϯ��" ����q&ˋ�`eg����ᶀ�;"=MA���0��y�Y�g��h���<	�T4۩�PcWV�<[/."���RY��V5����'&F����X�(�3h�8��>��(�Bu�q?"jĄ��u0�ywJ��4�����]$F%d�ݫ�AW���o�X5�����d�Җ��6#6���r���Q\Q�V &���bi_��������t����4��jCy�OPU�����a4�)ށ��뫖��<8=`��6�	6{&XYh���;o������mo����W��<�1�b$4%�e*!��)2l)@`�!&�͌h,�3N;�6�Fs�.T���e4��/=o�݆��V����G��.]�ɨ����f×_-��D'�-����X�z׭ע[� ��bƞm;�+X4���/��'r��Z`ߕ�U\��$��:K�۱c~��Y�ɧ���G�G�|�e�!�a���"�ؽ�Qrl���DF��*�nK���;���6�_��}{пGWd�!Lx�!T���7�E.���B,D/�r�$"� �;wF:�Ä	Ӱ|�j��2�B����ˬ�L�����(��~?�����3�s�ј����b'�̟��<���K�q0�_�Ą.7u2������XI��DV�엋���{�H�|y+5�{�������d��h_cs���*+����W\$�$���F��d:J�24-�U�7�2�3s���6�g�z��'p�E�#j��_~B�N�8f@o�a�P���yP}C�L&�����h�ư|�Z����e��S���ⷍۑ�R�Ć!��C��e�C�D���F��!��T�}k��$o�P�Q	q��<�h1V�!c��9Iz��o��e?�k�F8���1�r�"Ĺݼ�
��ꔛf�$՟�h����T� ���_Y���^5�=��`�����u� �� %^ڼ�7�uT ��J�H�V��k'�h�T\�X4#낆'|n�������)Т9)^uu�>:w��zcC���R�H!�E%�1�P˵�.�TR?���)�J�]�Z-��gUo����9N�Y)�"ֻV)�X�3�2[.�Q�ۻ�6طï�Z��K�_I�Q���)Xjxp_�0�n5�6��ɬ��q�@O1&�/&|&-�ƚ�d��ŉ�c��IBy&�N��|]�r�x�S��)T���D.Hf���*�l�/�&�<�t���hGa�8a���}������'�-M�.��0�mͨ��_� tLll	�ls#���c1�
|Bl�~���j� ����ӟ?qߨ�T��~���^�|�|r0m�LN���6��-�it�!�O	��a�
dRZZ�ݪ�j�"x=�؁������x�س}7��_��z��'�DG�]{��D�Z�x���W�,"�X՝�q�Eg��؅���8���h����y߉��?żￓ�]1%!��b��Ƌ�n�H�bu���uX�����S�Y��f�w�Mx|�$4���A�t�ȥ�h	$QX����L.��ݻ��a�.t)/Db�18�>��9̹R�8�VE$�̄�1�q���HήZ�U|��G7����F�P.H�c�ͺ�)��:��N������ggo<W|^p�_��	�=-o�ai]Ջ^�o�e�18ݾ� ��+M���4m���H��Ѳ�k�
'Y2g2��L��%�߉c��'�NT��(���
�g_�Lwyfd����H&�x�������b��eؾq-�z�nR!��k������D��m�0���I8��x�2�3�c�E�x��������K���͡�A*k��۵�s1jH1a�gkQR����K�G�h����-�K�V����{�j��7eK��{ꩳM���3��U����+^'_iP�x;$�j�� �X��5r�����v^��^+o4J�k����VsJ�_gb�s�;v�y�3HХGgt��� �{yO�L6�5�G�~Ҿ!���y#M-͂qm���?,X��z'8�s�&�<�ʋ�K&�ۦM���o�O�xh�
J�*���<G�Wt�&~%J�"�W�xL�v�����tNg�u������8��6���4ௗ_�G�w�������hll�k�[�.�l��1�&g�nv�dH�M���G��G	�lυ"ʭ�B[L�v��e��l6	�}�V�q~�����c�b�j�WT
�ɀ,�Q-��B�i
5e>���X�r�Ywn߉^��D�x�
6遷i5(b!et��У[5�Ly����y_�~y�1�\�/̘�ݍP$	�� �xNz�S���9;�6#�.$�����rT�������h~�����������;t.A���&�
��C�=;�x���+Hm�������j�҇ۢ���l.G<US����e6l�Y ����G��Ո��سk#��>=j�M��w�Х��p��nİ�@u�n�ֵ���b��a1��^�.Ł:��xa���oDYy!
]hl8 ��&����I�ɸ�Qj���PJ\<m�~�>�	�u{���ǟ��S�7�Fλ�z|��|���R��uBYe�o�Ũ*\�S1 2xP>��
�еg�������0�!� ��o���U#�X��[7�h	!�%��@�JPS�s�~�����j�X��x�oeE��>7� ǣ(#�(����	����U�1�TV���g�f5M��]���A�^���t�cp$�M����y�	=��w���NW��M/M���p��x�2x���FԄ`Cc��i�HX�fM��H$�2;��d�Lk�ht�*�},"� �Ŕ��\4
��	FC
/�xs��u�v-G[��"-�ߵ��u0��3�.}`c����w�ĵ�݀ؿ�'O=��5���J�T�Eߌ���jUc!�M3�����:z�P�k�l�K���GΤ�]J���v{G%�GTqv��M/���wi�R����$Dj{�gR�O�$�p�܏z~@��,w�{�׎Ϫ� ��
�    IDAT�Z��O��'�_7�%�^O�3YP=~����{�T�H!�����W^�T��$��)��Ѓ�bۦ=x�ŗн{�����_~�s�=7�4�
���y�F�wX�|)&=7A�1���v�B�{�E��2K��IO2�;�#3�<GD@F��;［}�L����W6����b����rd��'졛i������V�	t�ta֬���e"<w���هT�����^~�e<��XA��xc� n�����j�{�}�V�����J+0~�xIB����q��!x�GE#}݆�Ȥ28r�@�޳K��j���Ti�]y嵒hs��k�Wϕ����4C�ŴI���?�;ｏK�zn��j|��"�0}l&&L񔇀�G$ac[��{,�c8���x��{�{����̬�߆?����E(��BK���.�^�]0��z@x�Ϟ�kē����\.gmii)m����g�	��dʖ3�r�l�(Pu6�1fsY�ɘc�L�R`���`0�
L
L��%��Q�`0H=��l4��Y��`0�T��Y"Ɯ�d��r����Em4d�df�h�-Ƭ1g��2H�L֤��Ig�t�h̆f����_I�.�X��H�UH$9�,$|���P�q�����8
��8P��\e�^dA���v�B�*�Z�4e��D�F+r+*;��S�B,��[جN�a��+��h�^��[��&D@����y�5�y�8"Goa�0o�+��HX�rV%]:�`����~�B�4����
Wa	rV:YQ\�E���B��=0["�J�Y���]Y�����h��g�>8�gR� \��� R�zD��.+�VEeE58���GΔEQi�T���)�Zŗ�������c�b��~��$����䣹Y������r�� �6��3wme]!._z��E�:�G��)457H�A��A�Ǐ�#įk@KH{OM�ǝ�&��ٿ��3��p<���V���D�Ge��dBaI�l,���VW�9�E�p{KDĄ��J�2ԓYe����'�����:��X4 �x������3ѫ[9��C܏�][pp�6��A����x�Pt�= [��bź�H����ñu�~���Ǩ�y$���g�,$�f����T�7���Z���҇���w�E����fG��R�zC'*�뤳�:R�������Q�p<_�:������٨���ecmW*�搵9gn�H�Vh����^�h$@�g}̪�2Q�c�̵&�����mtc��?�-�t&�z-���q��K��k��b�R\}�p�I��D��W�ٳ�ºu[1r�H\t�%x|�}X�z&N|';�<t����<� �z�x����:���Jq�ॗ^�qO�q����Ǒ/©��#F�o�ï�_�_�G��?��X!Ͻ���X��7��+���Ir�������1B!{g`3�p�ȋq�e�`Ĉ�dΙ�>��lܰI^���Qַ�z=�vE�^=���˼y�b��0��'�3O����r!.��4<>�yѝ�:�t�UW]��F]���;va�ț0l�1�D�����8�����O�p�㏧���ǧ�~.��H�J�U��D�d�>�@6�*�W^~65'��f��[oφ��A0B��,$C&���ǠnH#� ����ȋ��|UU��E1m�t����.����C$�0�s2��ᄅ�j�Ǔ���ƍ�����2�\�Kcc�9�\t��f�hmk�F��X͔q�V�$mS�k���TJ��RRb�oH�(:��si��|��\
[9��`��*��j�q ���\&���r9B����ɔS�w&��L���X:i0d�\<�3��fOi0G��}������t*.��<��dNf�M*.9%�2�8�6����C�f[Q�u�����f�6Я� ��7�"�	���o��g����b	�n�{����v��E9d4�f
��`��hWI��
r�����N�xm��v�
��6ذ���o߉ʮ=��&f�c��Z��?M�06lڊ�nR�+�B�Q7=���F�~}�}�6�ڴC��Gs�~\;�|�pto�Z��D=�vñ������� �܃E��h����Ǉ~���\u�5�߷&O�(˦�����hK�[J�s�������+B~n
�P>�ߓ����^���:��MCg�r��<;�q���b�
�&�=��Ѯ񮋚0��F@O�=����N?��/��[`g?����^$kXŚ[�u���"�5c����9 �J�d�r����*i�HK<A2�D���d���	<;�)8l9�Z�3�����иw֯\
c<)�'E|��G?�������^��ႋ.��)/`Î����lK�5�BV�mN�8xS���Z��L�(V���-�� ��I©�i��.����L^��g�E��$	d�^;z�J�71?	��LM|>FGdt�@�l�b��+l���޵�����o�U镾^m�W��1�����T�yd,"-:�P��zE@T2����#�ಋ��#ݎSN:SLI�Uw���>�܏~������_�`�ʕ���1�7D��.^�u�{�TWU`��a���|�+��ާ`v`���ĥ_��S�J�9a��"#��	���z���G(*2`޼����޵g7���#�b1�r�(�i���J�w3�2�S��5��P��:���.#����X�t)}�q!��7�N��ŋQr�u����gr����xp�����[q�gࡇ@��V\��a��������㇟~��w�7� |�xf�$TTc�O��#q�������ba|�YC�ys�T�k֮��sM)λ�*͚;�d$P�e��&P�⤡CpϽ�c۶Zdf��d>��6;ij��鮐.������1�������'0�����\�����K1y�;x���`w� ���s�;^��4�����O��wۓ������G����͉d�M�7T��߿��c�.X���&�!d�[���΋ݦi5˚�c�7k}��_H�}����<)�g�#��� �|��D�*C.�d.��Y\���iM�l2Z�q
�$a �E��g��	�4�6ʖC��1���)�F%Ū0ɪ9ح��$;�&��U5�}�Zح9�z��ػ{�XV�y|�JřP�(�KbHڐ��aC<����lG4��N#�Zd����sϻ\r����L	[��!cs�h�I�NA���
TF�s�:��$�t���qA�f0Ӥ3RM�nؿwZԡ��N���0�^#��vl݀=;w�fs��p`��hh�ǱC�ŀ�G!��c�3S�r����_���V��̅Ւ��iA<BQ����Y�L.���FYT*���Һu��c+B�vd���P��bk�g���r�c����*�(���u�oz���ͪ��W$I5���@�sޅذq+~�e�xD��H.]����$XUUVK����$�sziGkR3�K5�frJ�M�A:�%�0��-�EC͸��K���{�~�,�u!:WÐ�`��-p[,8�O?��7�
���M�0�9�=�x�?��p�t��=�����$�[p�>U�ֵ�%���|�}j��DV1�����x�M�Ȅ�,M���t{�J�j���� �7��o���h���U�H��2vFAB�R0��<���7MGHn��?*��K�h't$.�S�zއMK�I�j`m{"�ӷԧRGQ��JC_c]�0�����ߖ�k/��qw��F}�47�้��=��oǔ)S����?��w���^������vI�g�V{�`�|y*����9�g�0�T|����������~D��/���w.��pD�ATWw�%�\�l*�׃��ǣ��#o�M����Ask�$���\|$�g��[��.�FY�_������L�w�y���xL�:�~��B�z��+/��3��/��w<���b�_�i��G���O��v>���0c��n�u~�m�=�"�~�a����+׊�Î]�eO�ҭ�#V�4����uמ����M��Jj5/�3A�k=�U�w�~�M}�~�N;��xd�=X�|7~l,,�E�3(�<V���7�`a@O��s�p�U��-Є���b�?`�ͣPѩ;f��6,�b��T���AV82&M5>#{�&x=��BGj�S������k���xޝ�֭�:��c4J�:u2��` gC�M�\������l~�>�ߥ3����;]�*�o�'��n�ڕZj�����􊀋Ȝ5Km�о0�D���ds�Q��b�"cȈ�i�>b��˙d�I�h ��C�M���6���A$�X��bdSc"U552��G%�ljhT��i�sr䌣b$�)X�)����!��~��4��B1F ����otq�9!��{�}8n�	��T������'���(��1��瀑#o��Ͽ���z��?u-(�j�a��qWf�MdE�z�xe�ص��E�ݽ��>���W# ���DĆ#S�,bZPXR(��?���}��8���T_2�/眉p�	+W���
hQUQ�-�0I]"&YIb8�F/u
�P��9��9#O(]�r��rI�����8�c��c�A �F�w��=�Y-)�]���(�r�Yg47��/����f��7��4�
YF�t�p��7f���"��Ը�M�v�>V��	�3K�����]*��2�>9G��~�k׬�$��IfV;�h�����VTv邱OO����������&$�l?ЊpΆHʀ� ecbY�kIU���ŀ�M�]1���@�<&"��$��ﮪy�*���,�Z�M���@��Ã�^w@���4	���G�u�\�:Sf�b`D�K�+UoY%��5�\ޟ�H(s�������e,��}QWS��{�9��9Y���m"��`N�]G8Ý=�	 n����ĵW]�;�{���h�_��/<x�m������{�0o�"�!���T\�X��w1
)*-�}�R������xﵩ=�9���k�v�J͚5�7lO�E�-��՝��؄W_~A _�fL��c������;v�r�҄DDO,v�ɳ��SX�X��I��߄�a��f�;�b拏������w?�I'ä��`׮}H%R�Z�ҥ��(�~�ilݼI��t��ڭ���1Q_�jn�y��46��qceͿ����9��}b�'���i31��O�6�����hT��-p�U�q�0��q�h47��B�zb""��).�ME����عe{�t���w��W�ʚ#�BT-����l!W�
���%`7�����G�E�ϊ]�w	Jx�u�1m������a� �2#�c+N�sRЌ�t����͵��>����/�ו#�G7����j��n�~�	'0��hh���Nl_ɇ
SZ�Ω�,����������`�d�Ԣ�F�A��P2�	�C|z�|]}��9�//3�t*	�9+���V��P��$����G����C^'���U3G��v�Y愔�]%h��Mm���(`��`�_�q�&�v�0�Dը�Y3<��
Z�27�d2&��j1�ي��Ѳ?��BaU��E��}��2�>e����}�>���0��4���w�>ralؼ����G}]#Q�M9d����ġ��
�M-H�S�(���5�����n�!����ؼ~�8�Q����Ԉ6��%"�p{AY��T�D ����W��O�.���sX��wh�7��4��)J����R6l�m܀�[7:�j���Dz{۶���m�$ �d8
00#g�D(����>��߰r�*�Ƙ$���v�2����l��&�~}��s׮x���d���DYE5��@��Y/�#V�v�ڔ#���MM~��̲Ͱ{\"�ʀ��{Ǆ�5h����+���	�`�� ���G��)ִ$h�/�e����T����TV���f:zܾ�ܱ�X�����`rc_]�⃞�	�Ey�V��\���4�y[M�L���Y��w{�� Gh6��6�59 �o�җ&s8d��=SdEޗA��HGi*�1/{��).$�l�׸�����d��=J��5q�CF�4��Z�L�<Mruj��)T ��^����r�c�ls���׀!��g����뮺UZQ�&?��4�S�N�ͥK���>��9��7����1��!G�;y��9X��b�1�EL~�E|��������"%�ǎ#&>D��zM��<j)"c�����^�ĩSJ�1���d.�UX
_i%��܇@(&�U���,�s�T>K�ĭO�N��ʃx��Y��/ѽ�ҋ^��rlۺB�ɤ�n;�mC�_|��S�G�^GH���cp�e���984;������z���z���{����8�Գ1���ū�qc]J*����s{\v���ǨQ��;��ŗ܋�`X�O��SRVH�5dHOF�ܓ�aЀ����U"�ZRV�@8��~�	��(��D.�V�Χ�z�e0����٭��o����QL��
~]��i'`�"��)e=�P�k��٦�;�VhO}���7�?�����h�����c��=ztw�Boij�9Y��%�j:d�����@����/��JZϘea����U����ǵg܇�[�p3i�����P�>f#�\U�v��Y��_�0��'�3���y��{��yce9��Y>�r1љ�J� ���q�1����>:�w�f��F�SV�&��V0#%n��=;��t�S&a����۽��i�ՠ�`v�R=��|)+YB�U�bwʪ�g�&�t�	'bǖ��E���e31��Sr�܀�.>&(<޸���L6�|=�5"���ݸ�ҋp�Y��Q_�_6����$N$������X�r�|n��>�@��U�{����-m"�Kz�|�ǳ���J`1ۅ%O�jqVsP!�.� ��#2��B�bB��_n.��2mQRR�E?.���DB��PLn�\��]�h��*L^2Y�8��\F��h *���L���!���V5ϛ��ew�u��B?r��7R�(��D�M�h��G�AZf�9���B��>�Z����>�����-n_	��bHՒ@0�>�W��.o�K�'R �w=���qk�l;����b�ʵ}�;/`J?�0Z\{@�E��J��-? K�A�J-����^���a ��}C>���t$3cz�e�rΥ"?L1N��3ٙ��5گ͓Am0��q��R���=c�W]~�0�O9�̚���_�ѣGc����`�7�����ʬW$�>���رc��f̘.�ٵ�\�!C�¬W�ቧ�⋯�G��.�.>�;˖-�:��];wb��c�ͷHK�a��Gd.��}�=�u���BFG�<
��0���\s�\?�nd��8I�A�
�:�Uh��5x��G����a�s�p�I��I�����˒2����V*�%�!\uť���+�w{n�u$�=�l�u��8x��]v���x�L�2	����w���oaƌix�������'�BH��D�C:B�ۊHK#��f8n����-%2HX�[`02�Vm�ЮSx~����͇�[��r��N�6,������ʂX���b%k�ŀ�L���Xk/^�w��7��0�w@�?�t�	�͇LΎXJC��;1�Dn�f%���~�9����xn���E@߳��X<vv����.$�75��R�ސ������zլK�x~�:�Ԣ����rxeߞ��A�|}3�zk�����3O.P4�(�Grr��(Ly%`�î��RĀ�h�g�'8:�+�y��y�8(�	sW����2�B~f�s����&<�������C G�P>,0�<Fc22DE8��2t��C�-���*���T~Ϫ�/��T:�N�R��a�Ӯq_P ���nij���ď-	U]9�F.����0s�t���A^Fs���t�Ba�/m�&/F4ڌ�b��c�q��/��y�e��z�)RC�9-5�����Y*�
y24��"F7#�Y^�l�H8$3����{q���Q
�;�<�̳X�|��鰹��}6_6�z]f��$�Ӆ�3�ND	�ťEb@��G1-"0C+^�>�.,ԏ&o1�� �Z�(�!H�W:)�?C$�����F�aeJԯ�`�i�bD2�Z��"n��HW�=    IDATm��6���3��SB-kIl�jTƹ�1�MD�+��ܮ����ɇZU�V��A�<��%�I�R��|&�|��~�(����?
 @@������s����K��������:�7p�������՚���䉣h:�szA\u�E��Y���?����p��+ѧOW�u�(-UʆL��~�)����ߋE�~��ٳq�	Cq�`����֛q�=���+���L��n������l:$tP��"M�WA@B 	IH�
��|���"/�HoR �l�}fvz���9��������u���3�����|���p߃���CmU5֬Y#�*v���p���2_�j�$�n�Gu���o�~ӇX�䧢 ��OaWK7�?�d|��cp��7��{@Xl�m�=�F>���jj<x�����Ã?��Pz�x֬~����8�cQqk4)�BcMyp	vo�y��G}~��2����p�7�9�)���s/8K�/�d慗���>�<��#���'��[0��WV��!�����4�\ ĕW\��?���Ft�"�|4;g�.��Tw[r�b�;��&�ݎ%�2R-���h ��'�x��N��}��!6���=��vҙ,�����	�buc��mX��>��a�^�D5�,�FEɴ�ܰYM(��<��+��l��T|j��i�ukk�_���g46YЇ1<8Α�2e�N����(?ز��� ^8;�ׂ�4���V���y�u��e&��	���_�C�����CS	~�d@	���?Y}1s����o�?�����W~��˷A�p��݀$���o_��X�t-v�t�ʟ,Bp<)R���Vl��(JS<Fc ���񣢪�hB�F�&��JM��9�L���양[�z��c$�S�дb�	�VϬ�.���Iǣ@�"� R�(c��م�xE䆓O+�T��i�Hз�����/����7��S|�qJK��M�bZ��r<B��x<�D���!�L��ȬD��"d3g�}��2ǯ��B$Go߀�}xn>��#�r՝������?DYeb�<�"����� ��{�\R����"�N����!+���~�ߥ�������y�y�mN����Q G������s*��DLdq�Q��!+�CFdCXD�*L9O��������%��B�5sV.~j��orO(ĩJS��Ő"��]��9ؼ�����򜸦���.�=u��_G�����L���O�ߩ�>&@�!����kc��7;x��2��s��%`(~����Y�� �>�{8����f��,ʋ�ر�w�Y���1<�QYIP,������o��9眃��:��f�����{ｇ��޷̃����O~�x��8ꨅd�b˖.���+�5.<�dYo￻�����r�J���=12�@e-qD@4�ƕf�i�0����p��������,`�F#�^/�)+kK��?Ɯ�M8��'`���Xqǝ������G����Rx� sodP��lx��c����������w,�3�}�?��;��y��p�%��C�-�\�3~x	����X��A����%0Y��h����ݽ��p>{x�~#��wҬ�M6d9�$��sY��8�̥1��^�]wo��5�#A���Ѡ�w�N��N��&��M�a3�ȣE&�@8Tx��v����W�;�7Iv���d\����䒖{��4�6ǟX�蒕�ͬ$R�?�2�ٳ�x<����F�=G��O��+�)�S�ISr�����������)]f:��w*L�ל|��^@��,蒨�j��::�N5!���O0f�Ȏ���忮�����ֵЩ7/�i�J֮��u�X�d%v��ĕ�ވ����,��.� yc��x\����$A���xJ���0 0��o�C{W��ѳb���7@^/��8�G�aʥ���Di:��ʗ��ҭV#\nb�����j1�߇��(J�|�4���!A�f��n����kǅ� ���W����h۳SE>;�`̛3[�<'o���(���pi�gnd�NDb�����ۄTb��(,��y��Ȭ�i�,��އx�ŗ�n0���O�ŗ^�k�_���zV�G69���e�E
�R�;��I�؆�H� >��%�L���{$)�E�r�>�bX�S �	G�u�Z�b�� ��6Sn�S�V����R"�+�:�J�ē���:�tx�ʗ��I�J��$�/7�V��*��)9ϮT֘h«/�H��e'�����$��NS��{wR��=�0��?v�u��wQ�˓|�����3�����kL�,���BP�唖����<YcT�ȗ~����WA=)\�\6!4�``�E~��gZ�1�`���l]�y�4���{��Ő��{��)|v}�G�%��μ9se}����]��P�d��W2_�]b�h�d�)��r�����)�>ܸ�%�"���k?�����Ȩ�������.{�{�O��WO����382���*	꼏�����`�|��u�m7`fs��>;;�Q[W��sg�ޗ�����?^{��;�����.�V�o�.��S��W]8��g����Uk��G�>���B�@�3��7���*X�,�LY��}������
v(��ؔI[���� ���݆ǆa��3�Q���h.g�'L&���
�\�	d���`���T�#ns��.]��zKKˇ�X�Й�Ͳ����D�� ]�VԘ��H:� ���D�8/K/̴�V~~П�`)����6�$ҝퟩ_�}⏅s:m�>ql:�o��ɜ�yxFk�k�'|Y����"c@Mf;���~�sC��`L�<	����3��@' .B�I�����{~.��ϖ���=�3�P�4{�)�"�OڴѨhw���vQ&gDQi�̂�v��4�X^^*X r�㩄T��tr�D&ØJ<b� An�r+�"�!#��7fNdeɣ'���9��|^���F�(��5<�Y�?gc�R��1��/���|��?|6S.��K.>���T�TɦTRR�g�{����}3Kل��N��xNcCg�v?�@��B�1��Rݏ�p�-K��`s�['���N���nv��5H�ZYN)�-3x%Vc{T��/לB<��Up:]���=j��x�>̙3OLr�{:�[�sU�'{",���8�lS��Rp9,��ME��y��Y�n�a�䧫���,,�Ɍy�P)Tp��k%p3=�|����{�<*���=d�U~@�V!?Y37!�_�ɞ�Zt�����׀���f����}d�x�!8Ӎ�&�]�y��~d�J�����il�?o7U�Vh~F���N"`8�9g�g���4(�e1g
�����$Y5fY#l���Թ��ޤ^:�#�~��PD��D���|&w^�[��o�T�\�Dcaٗd�a�B�N�E��Y$"C��d���+F��"������\'�K��I#��T2�`�˗/�1��3ϸ�hB@�I��"�E��BC�g�|��'q6��؈ te��䥤�N�GFP\R"	i_�0JKke�d69�=��qTW�c��Gr~��b<��_q��{coi���X2#@`%[K��E�lu0qm	x.��,��'���(�w����{'�a���#�sx$ �F�W���.,��ҹ$҆��&��X�Bq[b�/��%k>S@���� ��X/���C����T9�6#�/�3yb��t}��t}�<]�>����ӵ���Ѓ:߇7��-��)_�Y@��x�
k��sfi����)]���F ���5�Wݫ;���739lm�&ss�Пݢ4ƙ,���nTT���W
����n�H(���˹H�R�r�L�ZO$���jsIv�ty�ۛ|j~�|�a0`��~�����4b���@9�e�Y.7 ��D'��L&]��e�8MM�̞ǃA�1x�����>�wFPdw�����X�W_�3^|�Yu�<��i\}��غy=6�_���<ZZ�<�&��âEK�ߛ��tZ�Gav��Ӗ�1ڏow�w�7�}�f�l�@umJ�*0:8�b�[ 07޺&������n|��U�uÁ��\kOn�:Œ����##h�h�������):�D�}>��$ҟIA|Q&;�4f45�ɑI01�8����QRR���4�FG�#@����n7L+eؽ��@H��I]���K��
 (��u�	�ԫN��
gy��Z �gÓz�y�(yɲ̢��gvb�����\���!u�?.T����ǳ:�:z�!�-��OR\ճ�	������oD���?�	������&��'�	ڜ$9�,D�!�Yq��15��n��gBѰ�GV�|.�LΉ1�}����P��L���8�7	.D�TJ��"�qaE̚�,j����yf '����)ɄtoH���lV���G�n?1[�;M�Z~���@���� �ʘ�_r�Yx��-X����b7Kdq3A���U$���U�l��.�:�N�︮D���C
Z�s����	�]����7�aq�*�Ddl�� ��^R:�,�BA��`
�x^��%�J�_bbUR^! X&UL@D�Kc��Hg�ZXݯ�|-��,:쎚�&I��D�Y�����C��n����T%6ɐVn��63J<�a�5���7\���YUCA���������p8����Ad_o7z{':[�
]�"p/x����Rau�W��G���'���M������N�@e��,�K5�5�9;�B���;z��6; 9�r\X:<6�A?��	�i���((紲:�G���ڻPU]�e�WcOg/~|�b�E��d�N�8�fRB��-�e��l&E��H�Ehq�j�p�甦�ǩ�y�� "4�Q.Q��(�I>z� ŒɴBwGc���0
I��lM|����|�́Ɔ�ܶ] u�e�1�����o��|��w��q\t�ipZ2ؾ�c�t�"���N�bǆ142���y���χ��)�f��C=��h*��+/Ķ�`�֭8��+1c�<A��ba���X��?�g�����ۏ+�������j��kw�&:SY`�E�$�"7�;R����S @���nˉ%����>�O�D�c��P�l*�L"�+.� ��!��#�Ҵ���`�PUU�\&��*��f�R�z��!�O>ނ���Ϟ��p���;�e�IC�˯�
�����̽�l����&ɬ _Z���64�.�	H��k��"Ը���w�^�� �0A�¦|�e?��f^�o20�G}��!��J(��~�E�$�g�OJ�O�e&��O��}@�	�-ϣ��+iZ �������J�<x;��
��ː�m�x������I/z���M��yM�oV�l$�B�s�A�߫J,D7�Sd���/-u>��M�Yr��F]u Y�DGh耉�����������\��P삼�H2��S���I$])�a�w��( =�Ș��	 ~J@ ����8�Ig�x IB$ �����j �`t$���: B֠H�i"7�v�x�R�u����"�P�7IwM ������#��vo]���.�cÔDŔZs����߽9�ؑ5�Et�T�
����X@q>Ð�t�O/��3���{v�b��sf5+Q��>eqɶ
YRI�yk��T@獡f��ߪ��t�����Aaz���A�5_gF��������e����_tqD�8���3�3���N�.}��
�Wv�""�CTi�Yx'�h��7Hƺr�j���c��;��݇kn�}�䣇BqD�9��� �H���_^x^���=)����h@P��"ɛeF><2�<����b���:���ܓ����8S�$$r.aK��0^��1���&�J���2y�^Ax�=X�+QY^.����e���;��Q[U�K/� ������_���_;
�?�X����|�4|��@�+�$+%G`|C#1�^�k�۸%�37�OaC��N9�Kx��_b�M���nr&�\���it����۰d�ݒ]��k�q�.���	R9��2�w����,�l1��b@��186$��W,mC��:�KM�Q�/AmU��:���󢹾U�>�{�-�"ؼ�C�wc��hoۃ��J�ҝ;�^��8Y}�.ǹ|IY�Xƾ���p������}C�h�9��	á0��1<�v���em*�I���EU��Ċ�Kȵ@�M�&jГQR�����3y�'�Z�z_�B4y&KiZ��V�A#=�fկGLM�M�;�%��S��ǉrw^�}r�Rf.�Em{jkh6�F��|y�x{u �9�LV�z�N����,8~�XbdĕT����T�.�O��v��P����7���s!��{CY1�\��vI +���{�[t3$�;��dL��L�ŦU�ɘ��%xv��k���؁�6�ԅ�� ��^!�̊�=,�V#R&R��y-ɾ�DX|��G�?�(*)C[;U"�d_`T���}��Z,��#�+�٫�X�r����b;�V�#"�q(�.�{%��kQ�D����9�I%	H&X1��@f�8���"���ێB�h�F���Da3Z '�B1+�_Q	r�`x,��^{Y��Mx�Y�اS�`��6��}�kN>��������?�M}$+�ݑHd��z�m6�wP��<t�l�^�5q�*EҪJU�)��Ғ�K���^�8�h�s�`8��WPW�A�m$�$��F�#�-Ɖ��ip���� ή���
���`��2�d����]�
xx(sY�FSI%�~v��o��%�/G��n\|;Z:{14@��BYYF��BW!��Fo[��#�/q�f2��������~"���7�[��ãҬI���|c�̛�6���O����։Dڄ8�h&�lT3c`�"��u�����EÜ�]�w��DPSU��r2ֽ��y�y�?�g��u��ḯ~��̀хT(��H.�KfV�X��z?��`+��U���p���ߍ�N=g�b���q����~&��2!�%���ų�;���G�s�;�<����>'�=e�u���O;ܑQ�UTHbB�ζ������-���:�w��U�@/����:�d_�� ���@׮ݨk���C���������x��׉@C��-mF"w�0��*dS'��o`H��6R$hwK��|�	�p��wi���#H��m]�$�0Sh)�(����&���(�K\Z�f�(K�%���Y�v�u2�4;	S�L�%s,ԙ������y腵���>��*��;���,{�TYZ{@ъ'Z�:�]��*��l��e��)��y��菂\��%�%u�/9}��Qa�����Bz#�5�^v����p*-����G�6E^�\�),&8cKZ�,����@q�_��QM}M-�����P��)�$�e��Bc��ӂ��N��#�lI�yR�d�2�016��7��%����W$��4%�UIY#�6�����cTnc�Y��F���п������D"F(#�_d#��ɕ\P�����|�j��F�2f�'0�
�:�q�	��΢P|�Ԧ���� �{7�F��3&�K��]���Oy/p�ּt*yZ��>K���?��������uOKg$�c˝j^ݝ���i��$mG��j:5��r�[�����֭+�`_x����S*�O�p'v����.B�C�
��tV��4�F�s�l=hS�����W�\��9�礚,l��^��N���%���q����'�wcx���fg�(0����iT"�y,&�o1jd�C�2˝=�	W_y9����X�a3�}�����R\Z"-w�ϏM3�0�m��غe�T�g�����D�eg'R�����=0:
��)U��XP2pFI��*�eo�b�ǟ��2�jOa��Z\p�����Ʀuo���M8���j�U�]*�����2��$#Q�c<���ՏakK̾Dsid�Q3Aw�����c��MB߉$��j8 /}�cA1�i㒫�g�knX$�<�[�U�cp(��/�-JC�$�2�(.��[�C�P/�QU^-��H�G0@4DyE�����%��%EnT�zq��E8ha�Ԋm��H��Ea��D�_���ؙ    IDAT��<E�`�����6oCS]3^y�M��3�꺛P3�W�x7�۴Y�9���6ߕ�ȃ�b�Ō�͈8�A��dri��F- ,�e��*>���0ata��lA� �g�*\���������2��2����E+^�^4Mv�GMnj������f+�kJ��f�T%`�1J&�if��=1�)m��`���jUf����|�Hh	��10�؅�|7r&,J���_�{��ס�.i���qL��������\�];V�Ľp�a��=��K���q$]�#��!&��Z�do��K,C��O�E4>#Ì�B[��D�� ��I��2�*��L�4ͮR��D����<�Y\�:�@.�v"�cwFy菓j[/R5Ƅg�b�c�t�� ��er�@��HZ�B�adX��oLRx츤圱(����8lF�\(�&^q���L�mOkO4�f�Λ���M����E,т�F}��\�e[����X8/�[��',��I���8��7�{�O�����P��3������_���1�ǪW��f�М����7�.p����&7��i 4��P٩լ@d�%fPX�����X�b-�lۍP4�h� ��L�q�9�/߇t'��\�5�'�ܘA502��s���SO��p�x�e��0	`��e�Vy"�C�(���c����i���ƛhk��E^*���7`s� F� '_�S�X��<��E���ٽ~T�W����[���~	�S��#|�ѻx��ECM1N����ױ�f4�o���#�+A%�1�p�i��(E�`���*ה��Ȉ�<[7��1�/�����Sh#22
y�x�OXu�/��dpâ[���[�׿�
��H���7//r��l��D���B?��lF�����K�PS����Vt���n3�Ŏ�xC#�;\p9���rX��V~�$bAI�I����k��]J��a�*!�� ��{����dKk'>x�#\}�5x�����_���=��{���c��w	,n^�u(�C+P:e���O�@"��d��/�Bs�^���$�u�F9��*Uk^yˍXg��"F��/�����#�<��MEۏ�j�Oe���(3om��m���\��01��n	�&�3�M
�L��8�9�t݊��0�[�tdUM��-۷���	だ|��J	��ڵ���`�It�s��b��=������������EbِH�.!��׃#ʗ��R�v�����>����=R����bP2"�I���/A,�Fc�L��eL�:�d�8��Ǫ���Vu+�0����+!6mt�V�ĉJ������*�MmT3е�/�vβ�'oU��]��Q���*p���hז>_�{8���i3�;�K|ץQ�N���m[��絤@V^@�/�$^z�U���o�?�q����X�bfC� a�ZZ���G����k%���e�.f�SQ�������0hO���u�>�ԓ8�m��K��N7,��Bt�>kS-��V��������Mϖ;�pӓ�V� %S�����s' �-�TZܸ��45������-��h+�܍���D���5�Ջh��6� T��o�Ę�g9Ӓ�7#4��ax=N\v����ظ�-D8���
��/�(�pԀ�k۹瞏��-������g�Ǳ�}������څ�`�#!��qY�v��D�Z��͙>?���//-;���.�~�3�q�����_�6|�&̹�Kq�w��=;���|�f�=�P8,�F��_=�$^~y��fc 1���� ��N�����c@[�v|�����Î@��L8����ض��W�=��Hgr��k�3۱��{��X`��^��v��"��lj����<���;؃��T��av�Ld1�ر	u������Ǜ����b�o����K�KFQ]�Œ[�����O6}�d<���2�cA���S.#(�C=H�C�B����"���Ӌ��|O��+~���0ڰ�/bp<�g�w)F�H���Vi�Q�W\>�s��̥�rc+�3I�$�,5�ZYS��b��	��IȽ�MY��ȳ��93������mb����G���?EJV�vz�Qͻ'�5V�{��UE�7Mmo>�:O����c'>�x&��� s%�I���M���ĩ����=��C���o��{�����H���x�5�u��ߕ}�'���i�O��F�7/^���J�r�ɰ�lx��g���+��d�<���Dv�W�e���?���|��/�k_��M��⋘;o6.��r|���x�G��X��~���z�!	��l�����!46����h�1���7����loϐ|��'m�D2�h2%���t��Y��� R߼xW��V�[S5��뢮a ��D�,��:�wT�稧	 M�*�%X@�N�ܙJ�C�g���Oڜ&g�)�΀�'^G���`�P:XY	s���-��D\Y8-p�^p�����#�o����>C@ok�3���f5�:CǞ���v)�қ2i�QVk[�=��h��W�>�p��d�(� =Q�U��c�g\{m�|y���y�j]_�����ԍK�kz3�󜟴p#d�b������M����v�_�����G4���I���?f���}?���7�t��,]��l�	�ӍP,�`8�����qʿ�kb/�>���v��ȍͥp͏��Ք�G�^GY�_�7�����b�Q�u�r�a2CO%�ظif͚�o�M<���x�����
��P]ۈ��a�TT˼������XP�o���Dc}=��u���.�?��2<�����+/���`_Ο�#?w8�n"���Y�P�������_Q߸ 6'eN��ƀ�s[�������2��7۶��gIe�y7�;�����w	x,��7�$\���<��J���a48�1�ϖ~4���.X��g�i�E�X?�v����s���v��s7؈���6vb��+1:��@�,T�[P[��O���~��Dq���B<3!��!-ٺ�9n�O9��RHer=v��aw{;��4>�ъ�p�;�x�����Đ�R�#�h�s\�0X�1Y�YEiE9�t��qR�vҹ��I&�z"=FN~s~@��HM�G���(���<���8�N&�·�l_u0��
����̪����u��i��z^�����f��{�!�2������nE<B&G.5�1�C���x�Mh�o�s��x�g�����Vg�{��.�&�f��K����.�&�#��7� ����"��_=�{���K��_��[o���'ǃ.�����wq�=���G��f�a��S�²e�p�A����I'��o|�8\{��]}�2����FAu�X�k`��J!�����O=���l���a����0�l0Y�m/*��p`��A\
�-�3<��R�~0�8��@L�L��!��
��5L����\]��MD�	�$%뷶Fwd�J�)����@�k�Z�&��y�D[_:[2��}E~�����鶭��q�7b��n3����ۓ/��{����?,�)5��)��4CZ?��m�ϭ������QZr��I�
�-�T9�Z�2���������������wZ{D�č�_��U�^�7�r}���b���nZ��.��<`���@�D��~��;Ż�'�� ��ۖ�®�.�-���963^��(4�Vg�jNO��W��j88�˥�o|3�j����9��Q .����8q���������;����fs��_�:~���������m I�Uf��GeMbsXZ^+�K�ׯ��Ζ)�T�:��#�������̟��(�]�e@.��n������������͆�nA"�����M?FEe#�F/rE͊�vD�.��F;�u�p�!����Z�w��Ƃ!���߰sW\p��hUS���%��#x���b���`��%f��Ub4Bkk����W�T�ݝ�t�ݨ/���w��Z���*|�m'��$�6���#>EEi��q,��z�"��.Asc�(�uu����Fq�W�.�e�ȥU�r�F�%eU���ǟ^�+�>'���9�O��AIy^z��`G(�F,��Ȳ�J�t�|2Y��'sF,x�^��|y��_��ed�!����Km�z+Y�^����ҕ%����&7*Cf����u#�W�.���}Dp%\&��u\y* L�E]pm_��@Z���';�x>�G<���=.�y�Cc�:8��/��$I���"+۶����/�9�]�o|�زen_�s����ŋ�qӢ[1���x@0 LNibtӢ��%����o���n�M*��{N,�|�5�7����֭{g�y&�q�����o���QG��?�ֵbɒ%8�G�Η��gKnV�-?�U���~#�CR�74�c�����������֯߃[o���+���d�.1Iq�#'@��銽"�>B��LUe-jHr�M�+'[�23$#�L8�k�)��?ђ�<1%�jO�����ڿ�^� �dVM��1O!�?��J{��0��3��&r�f+v��[�W�-�����;��E��Rt�>���cl���QI
�RS�s��5	�*{��M�A��(���t%�}���Q�Ӯ�������ؼ���6ٺ�w*t�(�N�{�΀���$���'ש_:z]��K�	�(Z�:����r��n��wŲ��o����k�?<�ۗ��x,��[v������(�BA=b���qFC�
ߏ�r[tU�fX8>��#���Yi3��lݺJ�F9oN�\���R��8����Nъg�y-]�
�Ī���L( �:�V���Aye�������=�Yf�t9�b���A}C�.�?�K��.��߇��A��p3��&�w"�3Ȕ�T!���f��쎳2�,v���!���bDE)A!��H5�*�Z�Uu�B�۲�c̜9KW.��M���O �� � ϡ��ٜUU����S���DuC-�{:��@֊"���A5��G�������~�lʍ�x����$��~�r�	�;-�����,E"��`/r�Tq�DC�8�ω8�Ə�����3瀅͞�V���Q_:Fdl�cqG��G���3
���hͳ�I%΄���]�H�s�cq��IQ�N�k��D������H	��r�����|��)sJ��X�L� �]����g3���T,�^�M>6�瞧+��_���
#�~m_a�F0V�Ң�K�="��0|n�ԙ@
�dg��8픣� �	f͚�SN9��W(%E��Rd�0 �]^TTUJǏBBd@��c�={Z%ГN���$����;��܌ݻwK��䚂H\��,���;���@�
>���C)���� lٶFC�������EF{E%^|��TT�▛oā4�տ����A�������|�2��a�~H�(����rƔ�(�Z�02R�E���I�l��ڗ�K����?����?& 
�'�t�T9��ϻ_�������zr�{La�� Q��P��)����),c��`w�z{��h$Z:�j^fz:��:��r���K%���:E8����tA�7ߧ���u��^̧{����c�7���m2���B4���˾F\$�s��R��� i'mMF)%!����s�E��y�۔4��ދ�3g��.B Ŋ5w�.puMZ;�Ő���=�}��>�x�=�t����=����˦��-]R�8c#o�����gޑXT ��97��P^R��s��I�>	�>\���~W��:a�^r2���2������Dڐ4-�����͚�,� R刬��w�!����܃�y�q�~�l���Z�D���AOW� qi�
EdN�%��g	Gǅ׫@�،f�x�عy3b���y(.-C�h`g1�l,[~�oX��/�A�,����
�΄!iDU�)�ܹ�O�R�fԣg�_T�i�����2�စ�x�5x�Ý8��Ka��g-�P@�1�ӌ@hT ~t�c+��H����C��~\�OL�����`^o��s�80E�]EU�X�p:��J����fua�����ݭ8���PU]�?\��� ��J�����<�h��(�)5b�@���u�Q��M̘]H��_Mj�3�����������c���{�ڟV�K"A�����ǝ����TY�Y/鎨�i ;���t�R�qX�ߝK����v��i����.�h�w受����k���D{���!N�,��J�l��i����^T�7H��4be�b�׭+�eܒ#=�u���ՀT�����b�)A�F  #82c�6���h�s}��̎_80�,��w,Fq�>�}}](/+ �-�n�1����4n�����J�cg�IJ�z��:�	--�#��cX�k�?�?k����_/����d
%!_ݯl�Of��Z�n�G
mY	��t���Ǘ)��H��qW~�@�z��PNi{��#Q&h,�)�ˀ�wa�ؒ���n����\�G"��9�r�=ݝ����A���( �����{���{~ ��ZP��`6)B3�B�?����tp�X��D[��	SA-���w�_��M'm������b�,���:��c"3�) ���%���<=��p30�->�Bgv����vYz�
`X}��Xp��A8�@8��`�Xv��>1`���T:#�@W�c7��P:��
����e6OSf�l��O�3��'7s��D-���Y����IX�U@��|�P\^!҆��2+���JlٲE,MˋK�M�B.�@�?��K�-����ozC#�����4g���A4��V�LL�6�oFiD�)8=~q`�P��aE:F2D:JT��#A�<��֍3�q�yga��X�����q�I'
m���w��6oo��W..l}��ho��������>�����f����ؼyV��o�q���%�a��v+vc��"��p���
�6%�uv�M����?���/�k�1�x�pF�&���Q�+<6l�Wmm6m����Wpŕ'���`_��| �m��H0�ߏʚj�f#ð���iժ6T�5U�E������7�}rP��F��T�vz��L!HM��u��){�4-�B���C�O��s6��ڊ�"�D�[���n��8�a��(��R�Q\��8��y���/���/�x�W������K�Ĥ�A\��(�w���&����%I3�m.M{V.e��i3�1�k� 	�Q���>���n��LNx��h	�#��U�(FZ�����M6���a���fA2=R��Q�-.�.�Â��12[Mdǩ��'���afc�=�Pl��&�Й�
'R&�V/Bq�O����K��f�XJ���M��V�M�ϧp�՟&AϓE������$_b�O��%櫖��/q�DD$])L�;�R���\JzS��{c��&3b�4l.'2��=��!��]�\v�~�zgG���gϘ!���)Aqz���^��N˂�z~ �Za����.���n�V�X��1��6��
�{	�L���0?�`pQ�2�t=y�[���A�ռ�].�V�3�s>�z͝�oj�m�ݎ���Y��?�K����x,	i~��?c��vx���"�L�)�!3��u���a	���E:�_��RHb4�j����mu�T�J�����w��L�Gt(�Q���q+´9������7K�PUY#���۷K˽����~�-);���q��s.:^�19S�f��~rdH��&�&Y)�p������٨�DB��"4W����<l{���q���A��3�/@�5kV��j10�DY�����ᗏ<wQ*���?0���N9�L,���;8���4�V�l�Ԅ��m"��g����D.�椃UV���p
c��x�s&ID���j�Ɔ�E]e� �,V,���C������}�ňfrŐ����UP���ED6�K�QWW�u��3�2.��+� 7�_��O���g(�Á�g�����(r��R0�-�t]4�.'ia�:�6L]�y� �[P��'V�t]�O��-�k��a_��	O
�c��f��&��>@	�P��,-^��P�)� ��7�a!$��hj,���]����C	    IDATr���pݍ7�QD������U�:'���PU,I��(�lp!â*��I�ب���}�
��B��� ,T�L'��!�4���aDyQ�p��������qI�����G`x5啈�"(� ;@Ŀ��H4�p��36�	آ)�H�-�K����ݽ���Q���L�G�6#��8V-_���=c�����2I)���-#q�N8�Ƈ�6���W6Ѕr�oզ�w@�N�T�;���Y�Q�ۨ0��)�]O���:�ru����lZ���o��uK�=�j�i�葁,�>
]�Q�u��3��r��k>mM��ϝ9Sް��K�	Х]�g��lW��p�h[k�i=P�2a����8诧'�����ga@�[��զK&?}@�B�u:� �^���L���B{w4�G]�@�����bfϛ�E�����V�Ɖ'��=-mBWk��?~���غm\n���7�5IqM�
�����M'��l�ǈ�0�RF��w@:p��-��t����B�<��:Ϲ�d�������f̚��Ʉ�6n@qI�t������J2�-S6�C�n8��&�u�
̘Y�Ì���P�+�t�Ņ��0\���	ꛮsV����F�0:Ё�
?R��-��T���t��Z�r�t'�g-���*|�l�@�3ذy�l�No�j�����!��B�-m�r���QY�C:BO+f7��[�<^6:���>�w��G��)��D*�ёA�w���Fp��9�+8����qZ�{�v$�a1a�;�+*����a�;
��m���_�Ë�9�ɚHd�5�����s�((���(F���q�'c��Yx��W��� �c`((	�����}l<�d&�����j�]���ѓ
�扁�i�� �����9]�0]`���	�^�~C��K@�����	�EU��["�f&S����lFGaȍ#���,ĉ�>�>؆���eؼnd�����pc��Vn��3)]�B�����+�D��"!�Op%�iV~�>��J���͌D,	��#��$�ŕ~	�0To�;)[A&ƶ�_�L�H\�E�S�}. �_-o�F4@<Ĝ�j���p!gReq����vi��·������*���㿂��!�GeU=�yg+�Y$�%��y��KDP]�G,2�-O���"U
���u���D~�s��LOk	���y%x|2��.�����\�,:ZQ[]�`8"V���#px}ԬE2@��<T�<����<������ƢѲ9�3���:ۜҬ�P8O%@������醆"��0��7|~��n�N;�GJ.ǣ���}��ra�0]����&P���p�
[�zR�":y�o��rg@ׅv�q+)Ľ��]����~���;w.���zq�Z�b����}�Nq٪���Ǟ��P��g�:`��%[d+���l���ՌD<�X,*z�ۃ���	��Xn"CYW���w�Q��:_v��ԅw�WT�`p\9���
n���ۃ�۷	r�-���&lܸ�X%�b�C63��y
~x���ϼ�U+V�������&��Y��Y�q�ܵB�K�i���4�I�h+��eN�q���\+��L�����A��p�mK��ւw�~'�t���ݾb��������ꤓZ���в�C��������Sغu3��n�~�f��x���\u�%(�o��w�{F��1<:�d��̓ʪZ�@C�aDB#�2(�8�}�7�d�=�l߹MF]�_�?:���=l۲w�� �a����G��B<kE&m�)g��dAy���0�s���n�shl�D��Ũ���[�9&�Ǥ�PI�4-�f��g�.��4���zkjbC����^�.'��0����|��,4�oT��&Ļ0���H�#�W��n,
�)�/u�z�hmہ��~�HE�u��3H�#�z�v/2t�E$�LdMp�|H�`�FL�\h�dC��G���cQX�v`��%��{"���[�Xʎ(�}��(4�b� ʊ<0��hiEY��e����>w�t �~;F���[�p��p� J�������d"!�q	��.X-NX�6�搵1>>�!���j<��2�>����꾇Q;�`�u��g�� 9�����Z����DuF�=����V�Ч��v�ˀ���<~�.��x2�'`U{�X��a�tvvc۶v�%��`��T�@2D��4\�3<v�kWQ��_;��#�q	�T����?t��.��b�i���
��WY`�b�;�O���2�Me}��<M��	�{�Ч��'�n�?��z� F�{���A}�
�`P*����f��D,�Df�e`e,$�h`=!�`f�R��\�Ɔ����,��e����~��[��ze���'%P��i�9��!���x��~h���83���H�NKQI�܂��<�	�:?�B�:"TyP�����h� ��V\N���00�F���� ��ڊH$���/�����Ѫn�kD`�����8�ԯ��'�ǣ=�Ӎ"��s0��������k�G[�y�$SX=&��U��`u�����Aس!�,Q�x�������#0(��-���������OY�����������QQ]/nv�~��7ϕ꿬�C#A�ٳG���ڦ@�e�hj�����p�����*�!��oŶ���3 _Y���5;������`6d�Y�=	%n+�6����εw�Ï>����Å�1
-�W�|,~��3��N8��;���.������F2���lGh, ��P4(�T2d�L���[��	8�~T�TKEHs�h*�Պ%;i~�5��i-�lʹ��P���v��-�b>̀�0��+�+���<pӔ_�c�^8��7#~��~m����\����9;M�`Jq������p�e���5 �Ջp<%l	v������p�y����cD��O�+�\:%�W��x3��$Ey�G�p#cx��אM��r?d�|4����>AG��X3
�l�B�=N��j�Jq��Gb˶=ؼ��Sh���Q�,I8����`�&1���rZ{;PQ[-1 Kb��[04�If�6d�4��!
�_�F`l�� �^}!������{�P6s!�b�gu�h`L���y�X#uUu�g��diR�i��(� ���'p�̲w@�������1��?��2�b@0�Ï<����D����V�YTzMC�̓w�t��cfy�s�Ԏ�ցH$R>�y�h��vu���>
s��B��˅G�m�;$S6v����1I*5�u�9ӫ\��r��յq��+���A�z��E{�^���S,L��婖|a�N�d=���K��Ø��sQ'�U����t�Й�3��~� ��ε$[��1d�}�2����K�ζܬ�`��;��;(�.f�Kf��̴���;���{���e-L��j��3(z�R�b�(Bt~R�LJ`��.�`�c��"��������1z��L()/sf�;��s��c�$U|ow�8?��L]9~z˥ؾ�cܽ�>X�@�׉��eTU��5,�
�=��lVvnn����r�2��~8KkeF���
k.�*g
Mv\rΩ�AWo��er=����5�?�4�\�6w)��b<���x藏�W^Cw� f��8�؊K+14��O�����H�AyY����Cc8��q�E磨x�����__DGW��o'(�e4#M��ɜ�ِBtt���Z̮�D:�J��BGw�T?��M��8��3qꩧ�����Tg^x9~r�����8�H����0[�nX�6���H��(&����G�>cr�/.Eum��Q���]��Qh��$H4���$�J��c@��xO�dN�'~�����%�}������#��{ײY���&��n���D8�� �)��f�ᚫ/�ko����&�q`0 v6��� ���<�u�A�G�kߋu�섿�V�,l��\��v�2��@,���8	g�u�?p���b�ͨ*+���n��Y^���.���a 	_0�j���Z|Ӊt�P�3��;nGC�o�ۉ[��9��2e��� B��X0.9�8�&���p����(J}N9��>�,^��ۂ��mș�p��"�DÖ���,9�W�����mm�8�B}�XlH���n�=��3v�精Hi���?���l��ּ���׸u}�"��,��O��"	3��|�+G�g�N��d�?��'���F�3�	d�f8\@��%���\w���-��������6����E���93�Eű��C���YL�lZ�̜ܵ:(�����t��km6�5�}ѫ�R�s> n�ٶv����'|U����#��s���~�t���Pt+"��C� 9Уt>�p��[�M��e/H�^�+��]w�#F	��X) �e�W��3����6�X���Pܶ�)4Α��[�j�A��*z�ج�q�N��P1�-~rVu�<7�X"��.��R�kR�2'R�	D�������3[��c��ې���Q��X��C$I|��3QY]��KoGmE	���jսx���a~s�:p6f6�"0ڎ�Z�ƙs�[�������bëo|�Ǟ�<�s�n�h0�����I,l����
�����+P��(��ln����O�����k���W����G���PT\_i��#�J**�Vq׮]p���٪����с�xN�V�	���`��DC�����@Dw���kA1��p[�/}�4W�bݛ����H��������b��{��]�W�^Z��;���-B<gF<c��Y�h(�����[0	�WL|R��D`��`5��M��D\�u�ף��Ҥ) �P״�[֯���=?�O�?ETF_SӭV�r.�h��z��ݾ��{��U�5'�^�ۊT.���*f����c��٧�￉7^-�}�Y����1�
�,86*x��p_s���~(��X�y�R�sfA�+c��������O<fpǊ��/�G�5+!���y=�g�~ių��[Q�Sp8|V9�.��b�Y��m�#̙�b7�[?��'|?���:�ʻ|0�@��O��B�z���5��\+��1l^RE�����)��-��nEY�+�>�W�\�݃A��1�3�O��������{Quf����:�)�=��-wpY�Xu�r�/�؆���=v��A6��f� c7��%;�;��i�}a��K��ѿ����ܝm��H���y�н(n�m-�dKs4������{�GU�_�gz��$�$$!��DT�4ETĵ��Et]i*"� MA�뮍��bY]{Y
�tBBz�dz�;�����M&C@��>���;��$S��{���)�s�I��K)�I�l��-_&8�zo��7`O��i#J/��4�l��]3?� =���*�e���'�!�%w��HrTS�jE��E�G#�n@��H,�u�6p6�n�F4���G���+�Dcc�zW�?+W��?@*m"��|w!Wq��}&�	��^�N	R�H��M�ݒ�<����ԯ�.�����eD���\�Eq�2�o�^��h���¼��1g�=C,˗���W\�I�Fa�Mw@YV�>�O=�4>��SLs&�^o�Q�Q�#�#���@&�	--�h�;�Ƃ˶�+a."�6p��Y58oT?\0q$~�r;f�xr��y�-A�$����ÅO��[���%�Ϻ���O>�W�C	��Wr�Mֲy}
��q��!��,3
��p{�J�:���)]w���>��I��t���f��!qjWt�K�I��ÿ�S=r(NR���~�DB�:�>�5ܽ/�K��iU�4��	P����B0,�Gi��>ۍ�<�;�-Q�6��Ck��(u��o���k�1���{J�R�Yv��ŭ4�{�c���MD.���K$�*��X��ϸ�
Ģ�����C�H�����H*�����F!G�;n����ڽ˞�_�1��H2��&*ZE��;pӕ��."�^~�]lٴM��eK��Yn-�*0���8\oG )g!��;���>��x����G1��{�Y���e������w݊�B%�������=l�k2�p޹S�G��仮�����s�����-�ɀ��'M�,֯�/��������C+W��l0:�~�Yl�B�Z)x3��|I�/���_2���Df>Q��{��\Y�RE��vM�7p��OWM<������Z���t�5�ބN�-��\p��m����_@]V_W�����A��_I)Ψ��� �2=ڜX�6�ўH'�`3��3�@�D�M�� k(syiٴL�$H�2��2�'�䟙�S��VD\���3ĠFԱ��B]֩��q�<�?9�I��b�B<�DZ! \��Q��n��8��+[�j5.��R�`(�¾��܋��29�iY\�"�n��I܅Z �j�m�M�ZL().�^������,�:�>��&P��*���70���f�)C���F[���	0BB{��5�i�J��/�>|������w��˯�j@|���8k�̟�w;�U�b���X��9|���8uH%��y��zL;w��A2
Jp�fgۚ� �n����EF�����>�]�]�|��Dȁ�O�'�5� �`��ulf����U�U�nFX �Yxj�Z���1f3]k2!�H�����u����	��;�,,CzD"�G<* �p ,t�󒜯�!1Q����ѠV�
Y9��b��3�����~����Xݯ4�6|�HL�8G���ٿ�]^1bZ=(Mو�Ԝѩe$�#�p��Rw��$�g� �$�ĘM��M�h6�b�B�ס��f�+2�!�3i��|2Z��e2=mi}u��S�N]�/�
��5�IjMc�Z��	I�������@'M_���$���Mjc2ER��d�i@2�ǀ�|�x�.������+�G�%�A�0�.s���A�@�^���7�<� p�ʭ�z���6DJ�C�t74��Q�QDݍ�s�Ř=k&"q੧_��W����������	������_;1��U�*��H_>QA�I@�oǘ*6��:�n��߻��h.=�2���W��!&�Ć'�g�a8�1d�塽�&�W\:sf�@,L�Y�m�a��'`+�(�I�Q�I����:}K��ˮ_���Л��+��[�.���XJo���tz��t�N�q����ɒ���)"�]��M�D�('<�:e�\�`��)���D�̇ !#ZtrP�T�#�E�/K���2�x��S'~�E�:����*�ׇ��~$�������5�)CgY��Ǖ�H$�j�RD�t0L<H>�$�����t@��v���`��Х�zɮײJ/d��@��4hP@�sI-ХC��"U8T�Þ��e�%A�ޛ2t�5��c0]�v=f^�.�R?��b�x�yT=ƀn0�pɝJj$D�7�����9T+�~�T�-.DQ������{ly9\��x�K�NTR�c�Q&���F6S�>8e�����ݎ�س�rm��tyYg��ۜ�N��z&�����%Ky����_��	��W'{�ڬ��z�#x��W�ƶw0c�d�?�*�cGb�Y,F>�2�F�Bn���@�k�z�[�~W#ƞ3{A�Z��3��'��3�p޴�%e��jTj8�+�hmw�׃�X��)&�,\�?�ڇ���	��Mo�*�����v���(3UM����lKs�2RfgM	�bԫggq��#�۳�f�4:�$�aZM���\R���|x;���@~~��zǏ?c��8��s����Ͽ��������X�#.�")�@� ��$���hqh���缘e�x�J	�Q��7R	��
���Hֵ
�����!@�l���R�go�ԺN���k�M�7 =�ω���@�u�N\j��)���O�~�&��0�ģ����$�A% ��@�4r?�T#�5#B�k4�`Pu�`��[q�%cY
������Ĵpj�XE2ƣ�4NU����m��d@��W���oc�����F�    IDATj�=����Y��������{x�շ�קn7Un̬�v7cL?�ܰ�m�(�,\�Vw :�
g�:w;j���x�ٗ�g�!�9�IY��N4�J�/��?]~�u-X�z=�r-K�&�O����0�Qf\4g��O?�}��,xBIˡ�R\D)X'�L������6C��7���N�k��˔=����)C6n�v�F���e	
�Ķ	UZDyJ��l)���*���68���]��Vm�|��׍�g�_@]VW{�6	�3�+�m�h��M:-~1��a���͞�3��)�5�3{�|�"���8 O���L��N.-�~l��袦ow'���_н�ܽ^79:I&�&C.u)9\*�� ��H���UZ�H���D�%@�,wӦM�E?��J�}l�&\|�Ũ�o�����r6n~5���h�f���#=�2��Ak�r6A)꓏��=#�E��ÿ���Q� N�d�Շa0��5���(��[o�ls��=(�S�n��g�yYV�9���;a�ڸ�M�1���F�u?m�)�ⲙ���/�駟�����x
Kʰ`�=��b4�
7��������p�Ё�~�iPiSF��j"�b�uR��D2Y]�+V����(��1�jjp��(�X�����T���ƃ�񆫡����j��je����mB�?ށ^~�7�9wރ�u����K\q(�[��9�&KJ���^SS�R�b/EE}������ I�KQ�B�@G?�2O!)�Kiܓ���b��m�B+Gñ#�}����(��a��2(�A<�����O8�b]m���/�����C44wb�%u��hsT�lD�*��"�F���/�(k�� ��#��D��m����qۈ�)�A�d�C�6�����a��p�A�cf�����z��uo�������MR�S��uU{�Y�>m:�}w���Ԩn4RI��4
JY4�!̺Ꮨ4n8���?��k��f니@��dU?%��B��Q) h?�f��K��������Z��yl�+��;ۮj���Q�q5�����m7����_�'&M�U���x̏���D�zx����V���V�T6�\�9��7bˆ�V���aν+�F�|� V��g��$�;���A�^�ɤr�1h��G:�z��5{a� �n^�A��yk]��ox�o��f!S��w� t�$�m:l}b����?�c�҇�	u6|�(dL>�l��o�� ���lћ��� =u��%����xO��zk鮐*�]2�	:6v%�B�Ji�ӱ��H��Y��tU�
�h�$K¨�;����cb�=sn|��3��y��� ?��`0XQY^
�R�%�NG;�)[$@��RJ�WtQ�>E�Ie!��h~]��t<�'�� :o@� :l���J�����%���t�n��}���]:�� ����[��w3�8 ��,W�F�7	L,�(��	зn��e���{���M��`��騫k�>yAi%6o}�$�p��PX|������p���CNf]x>Ə;{�@����K>��C�ڲ��D�;��31d�=�2?���x�8r���� r�������C�3�d��@��X�c�3iΙt�s���mo���DXH���}���3�	��Ͽbђ����?�oQ>���<r �Y���q�Ö[$��&����҆o���ǐil0�!$ı��_P�m���}p��3�j=��J1���,A�T���`1YP�Њ5k���_��5Yq�Ms������L�{J��Y��pP��ɀNeg�ٌ�%E�{�hlh`{"��"��5!Vhh�FRU$�2=���F�������f8-;;1c��<v�]��p�d���G2 ����z|�ٗ��m@I�R�޽qhpʈ����o���ԚX��2&Y�n%�PV���"�!;�T	b�^�Vk�J��B���]�:��+=�'��@��/����R����ĥ:tFF}�ƙ���~i6�H�=�r���Ǘ��.`�����q��6�2(h� y"���������fϾn� �܈pB��B�#�lә��@��q+�f��'���+7�˝5H��Y�UA����R�t�	���F�~ݹ�s�Y-�ɧ^���eQO^>�D��	�`�������1o���hr�( ���g0b�#��Q)���1�ehh���8OmY�«�(���u8x�j]6"19\n,��q�T����h8��\<+��������֗�Oh!ȍP�����Ѩ~�W_~.�z.>�������F�cZDH
��-���O�X��RI��@<5����o ���z��6YU��C��&���/��XT`C���j�����6A�{�����3=1m��O�;��w�9d͍MG�^oUyi_i�o`@'~�F��{~:��F��]K��Q�@O��{~�x��G���/-n.����<-��'�\��i���^KJ�1M�g�.V�Ks��X���RP#)�q����h��ޗ�xt��U�U���h[[��>�h7mzS�NE]]���`Ӗg����%w.Qh����\�f��d:���̸p��ݻv��LO,$ CU�>��#6:�2*�.��3���S�?O���fg�׶����
t��Tht���+�Ɔ:hT2�^����@�xw��8��ojGG���y��_���aÆux���0r�i�8�q�m7A)�#ۢ��jCnn6�Z5�T��'_Bc���B����g��*�Vc̨��y��}�P���(ַ����C���^}m;�F<�8n�s'<��x�@��L�l"NB�ρ��`W+t�>/))���BC]=��Ձ4�'�/��O6� }{$��i���PX������F~���c0�b��=�0�T�}*�+6mz��(���x��ٽ�5r�(45{�Ta�-�WH � �P�I���doLǡ��"t<��V�b�Cո��,Vң�>�T�� ��$Lٹ(�S$������+�t����`lMJ�{�+ǡ�z[+m$�7�@?n.S;6����ޒ+Z�:�������~�iyj�S�GF)R�t���J3.>�'����/����r��Is�� ���'d�a@u�������'pϊ'���G!� .(��6G���՜���	�<����i�u�e�
��ϼ��^ygO���� UH���{X�P\�Q�W^��������'C�߉S������S����ݽ�͸��Kqˬ����m�=w��>�> �E�Z�N���<�^d��}(˒a��E�,�Am��Vn��c�)��h�֝V�m��ހ{n�GV㻟B�U�� ��1Ϥ{�(�t�ѭF:[�f^���2t2��q]O x z�wAI��p��#;��Ż+]�C4��pJb8�i$HvW��j�h�	��"ɨ�`y�KW�<����i�-P��6�r���J��i�wvv:�y�Ğ�FQ
�=�|����������	��� ݮN�Q���z�EM�$PtԻ���Hg���@��� ��\�w��G�T�L?G,L�*��S������S�ƍ`-Z� K�N�J�N����#���-hhjE0D�*�E'@'���i&>˨G(��
�3q�W��p��!^�������ݷ9��`447aƌ(�[�2�MMM�8m$>��44��_�a<s�ԙ�ao�Sº��Ъ�W^|��6\�Nl��V�Z��'�/3���a�~X���x���O�C�%����bn�f&��k�b��p"�õ���W?`��_Agȅ�Z �5�H������\0kRU�R�d�J��dCs���؅^|zC�r-�{=�z~�u O>�W�\~���6������Zf���MIY)���c��hL��و���մ�+䐫U�F.���`w�����hzY�O��cD#W��hf�`AA�
������a�)��/�ѿ��-�*S6���G�4d��R�E4D�VtJ$����H<��n���TZ"�Q_���z�{&���ʣC*�}K�XC���I��w��e��n@Lw7K��'��*`�c����{��%)�����U�ʄ���QB�vh��S.C$D:�9����Cr�FY�F�Ȍ ��C����\{�X��������EH��P� L�R��)l�!��|�tܞ"�=��x��w0y�Yx��;�j�p�q�M�pތ�1���8K�U+�?�FvA	܎������^�D{g��]���,]p;��}&tz�������>�L��PRo(�N��R��\�I�A�>܁܁�'�d��������!��BR�[5�0��\9�\̺�bVV\��o����0V�
C��}8�f'�J��Lm��@O 3m�NTz��H��)`�Z6��d��HU�T0�n�����;j!�~O���w	���,��ju�ta���p2��k3�:�O��v͸��'uY[K���5� �X�T>tt�����i*�^�)����������鯣�'��+��zzf.����Yz梕2�t�$��	�	�K�={��$@:*��Sɝ���$?N�<Z����Kb�����D��6l`�Ѕsƾy�t*	?�n܌�ѬE��2P��;�;��F
i	!H��Nv��Sأy�)���7߰������M�\ޥ쁾y#�;�<�nյ57n<�=�\,\�Fc6b1-��f't�l^����r���� �2�-���'�����]��=�M��8x�j�Vk���3n�}n�����>��0�2	��ɀ>�����C�j�񵼾P�(ӷTe��

�ߟʜ��� �Њ���Z��ÆrvNi5�m����:�S/�\|	�}�]|����d�p�J�W^Zv����������a��@�橅��	� �R2����YYL�:ഷ�(ۂ9�_��e��+$����S�hw�B��1�^xѥ��������~��#N�w?��_k�P�y�T��,�J���@w�@řTv.�
P� �jS&��E����`B��N�	�
�e��4��Pٓ�����b��@�C�}K~����a�� =x-g~�����ث���{'=I��-CgƳ��yLE,E���q�%S�G|����&@fb�aʰ�=jzS ��A���x,<��B���k�1#)Ƞ���U�4��iB�[p�u�Y2�g��k����'��#�q!���V�u�<��I�\�(F�*E��=Ҍ{? �1.WN��æ�k�S�`��߱�,�?���������;k�۠4��	B����
ǡ1[ B�:`��q�W��K&s��`����=H�r!ǃv�x~w#f_wf_}��}�m����`�; m.R�;��I�3z��=��>���� ����Y�V��y3�@/Kpqi��q1PY��QI�B %d�� )uz]�$���Yّ�z���A7LfR�	:y�Pi���?^rλ�L�t"P�}���,:	w��a�����i�b'�ԁw��J�]'1UF>��O�[��0�H�͟���{$�~4���:�R��=2�a������;�iK��=��h��	��%@�2t��+��tp�B��d�t�9�H@��r��ЉQ�`�B�-[�Ĕ)S��؈`$��Fa��'9C�I�t����EF2e\ԯ1�T�����߯�mG��=������XL�����e��%e��ɓ�{�U�u��!���[��9��1�M�t���+�N����Ŀd�<2�j����
�N7�Y9�n��X�n�K����e;���Z\w�5x�����_"7ۂ�l��D�~��Vtf+	P"&�����Ʀ6D#q6�!�ɢ�"�6�#)D ��V���`2PTR���b�9p����.�y!���b<�ʧ�n�^44��D��k`��V��q����}��rrPVV��N;���Fɠ1���q�T�J�fH5dG��%y��<⅐��\�L�A�yj��a<�������ŗ�a���<��r�1���嗷�pun�k>�<�?�=��>��������@EJd)�?*���:1�S���MA;�����`9,����
�\�R���)� {:%���R��(�?��>�@Y
����R��2ei-�t@z�p<��\�G9?5b��}M���É�ܵ����GC�� uᜳG�M1>��7x�ב_4��I;;;�'/ ���Z��7�W�����g����|�s5��B���*��Z#�SN[�*���w]7�͚�p�J�oa�ko���j�HF��N7�]��M�0dV�z���O�{�?����������+�Rh�r'0w��_<��b"B�������v"��ADm�;�JCR���2 ��<��tI���;oƵ���퀻�<��~ڋ�1�9�o�e1�T1��m����E�xy�vdT�T@��sɝ`O2CI��.m�b�L�,�8�@� t�B�Y�MH���{tK���_tg��hI��ě����ZꕓV��x���IP���P�~�Q�˸�G�>Z�
��ɫJ�

�
e:U"lQ�(�<5s�ď��:���;e��].�����Uj����l4���Դ�w��)2�Qz�4n{��Otr3���O����[�uc&�w_��%q��J�3����7EL�\}7�J�T�R�K��M?~J &8:���N�!D4� )#4�\ɤ�?1ł��Q�G���7���P	e�/��"����K9C���&�w�y��N'��67=ɮ_�(1�I���SEP&"�B!�A����U2���j(胎��#��u����'I�r�]�@cc�r��	��h�� :m��QA�Z�t[�B�ml��Io��	�q�_�b�x�F�=�ݿ�ǒ��2�\OQ=�tJ��ڱd��첱����o����=S�P�(G�l�ՙ`��g5��C���gRPBY��ӎ���0�P*D�<���O>�a!�������&`�O`���v��	Ag&�=��啕��=��O����ep�;�o�Y��S�]ͳ㴰�J-�����e�Db�S���w�����\b��;�v �DA�����v�Yf#&L:��8��Κ�Ͽ��}ϭy�x��� l�i}���k�-m"�F"\gl��K|t>�8��?=>��i��]�EE(�[�j��$�DYy%
ۜN���DT���^�F��a����"=З~�k�:)���W�V"?nCNӖ��������/��%�FI���MLT�3z|#f0'��h�ryX���X�:����݊���9�ס�B�/��B�F����8�X�1���X~�-8w�p.8ݺh����e���,��� :��m�Yr,p����g�?Mg����/��2�O9�,�3���'oi�b��e��h���uW_�+.�M,�E�.Gm�QY�z�J������Ýw.��Ӆ;f݄���hxx��뫟��)A�/�@"�>�q��qD�HF�(���U�w\{�s)[�'^|���9TfT�,>w�ܦQD�gUcѼ9�'�Xr�*�ߐ)�ڝ~�D'������SfN"g�j���=�Y.A�j"�2%��j��T�H��P"gʻH"&te���/��K���m�R�_�{�{�S���b�L
Yy�erR�"LeeK$>�8�^А!U��F�l�"w�Tf{�֫/��%��j2WY�W��p9� ���	3i~S8&E>��%���i�z�z�t�w%��^/���~ף7�
0���(��S ^������qd�T���uq�����$����a�˵�$������q8�r��щ��P�j���ي+yl���Vr��f(C�q�UCGaӓϡ���Yޑh���3��ˉX�z5��I�6�0L:-{%�tC^8�L�,'����.
��X��]��YL�� �C.�"	�@Q	�ʣ��y<�����$��ƎŨ������m�e��ƺkQз�A���p��'��O����vq��7|�y���\�`$��:���D狎��=�>��'\�"�W�
MM�(�,By�b�+x�p��YLf׎}H��Ƃ,��e�*���@u�&��\iy_t��PW}�'���b>F��=0
��.[�&j�BIrI@E@���y���    IDAT4���r��3GV�O���!�6u���-D�+S�{U,�@ݱfx�~9u,�^Q��ф
�( ����c>�0�m9<�J��emO ��xz!p�H�L`+,DEi9�;G��Ɂd�T)��p"AJ��T�Z)B������^R?>� $@ۿ���u�;�čD��"��u�b]��޳�v�j����'�n��Ԩr�kˇ�@,�^��>�RU�]��|[�0BPٮ�Q�F�3�Ѱ�z�Vu�C?��%�%�a@�m���#��V��@#�r@.пuĔ�#�cΕSq��?�<��g���7^���c��w�����-s�CSP���M(�ec�?�E<�kG5�;���r X[Oe��p9}X4o.�6�+��ݿ��"�� ���N@��!�LB�e���I%�6�6hǒ��b��c+{�}�#T�|�I�*�^'Gg�1̙u��z
r��}���Ͼ�	_X[Q)�^g��d,�"@G�be���I�Mjuvf��q�$��Eh���HZ+�1$"��`Q�]L���O�t���]�ϓK�dQ���Ci��+��
a9�`�NbU"���~��oB|��L	jhQR�R$!���f5�C�XE~���g�����t$}�t��{t1C��
;��:R�������xd�,���'[șs������{���� ����ل���̢�u�.Ni�N�СCy����)3���w�8%���yӐ���T
���[�d�#�T-�������G��ax��֚�%_�
�j��K��?��t����q�V�z�aoŀA�Qٿ5�� DE5
6h�z��a���e ����u6��#�BLYmʑm˅��bB�
��pۆ� :/�˖-�N�ŭ�͆�bf���L��1�H8��c�b֬[X@� =�"`���W�RS�V��M�A���A��2�7B  �|)��Td������ޤ��oo���A���#�P{�	��(��/z��Gj���3e�%hjoB{S+�Id�����h��`� �#M@�1"!W���'�y1+�McaDC>X�jX�J(�Xt2��*�5B؃�?z��%0�/F�>FC6���ر�0L}*`+�B �`/����I�����E#mP����r��tp넀�*�y��Z���ˉ��T�U0�{�$�ByY%z[����g��{�S�ڞe�̪��z��e��K����e��u������ғ�L@W��f����!K���D�m����Gmu�GRk�ʘ��[�h�J��$̪��{����p�ecMw,܈ow�@a*�r7��i�P� �j9<!�v̹l
�r�5�����]�I�f�|�c@c��@{���\1���,�YGz���O�K�SOm�Ũ��6f͹����o�W]>�P/�������f$�Ehs9���LM$^?�z%1?�a�Y��X���%/���v��}�Jy���V�a�Ʊ���,����Q}��e�p��Q貌�"�69���b
�>S��UHC���H�+�ⴄ$�"��������}z4E-R���38���CH~O��
�8�)�/���x�� �,��Ŷ#4�%a�|(Y��F�I�IA���a�6�~2�V�(���3&�y��!G%\$@?�r��ؚF�Ie�\���:G=I#]7v/cc]o�aF"��Ǣ��#OF�c���Yo���X;I{.�c�{�1p0�*�H?O�� ����P��H:m��Sˀ����$���Q���3�$Rm�LY�;������	�	�h�6�Տ<�I�&u��S�ĺ�O�X}�L%W+�^:	�Ļ �z:��B��׈G��`(�3ƌ�i��¿��ovr��M,
�QUU�.<����_}�7�ڎ�%�������D���J���:�.4�43��rr��g�O;QP����c��x`��8p� L�,�N�0:O!yy�1����{��'�REX�R�������Л�ܞ��ж4��@�J�t��*-���@Y?��J��<X��V�`�+�R�摰���քl��M$P֯
�k�r�C�]R^������$�A����.O'�Y��ݝ�uf.���������䘴�9ې�������$���#x��W��ן��Wͭ�u��xƥ�e�>���-�9B�7Ι�۟@\��^o`�{5�'jąA/�9�^8(�\�)����DU������N�aEy���!���3��w�k�����{Coy� ��8��=+l��2J�'Ҕ��u� �~�&%�cߑڀS~���C�Q����f%.�h
n��,����kq��АY�A*@���Ick&Mr�/����g-���7����LZ���.
z�*Ba/,�:k0������K�2�����m�aʔ	xxᝐ'��� ���0�7{Pз����4�}����ic��xOl\����0��'��沪�E��;n�%�wo5�-�
CZ|*r=�wCB�Th*֤�C���UE<�f2 5�aܹt5�u�6�"M@.#��T2Ǝ��B^}u�0 ��B���R�˞ꡋz��� A&r7h?��#�J��˙����oj�M�����2F��w��9
�s�I�������Hz��H�EM��ʉM	3��EVQ�T��+BD�$LoPS!�bitj�=mG�5�y�/x�3Gp�.kmi=�v����,>��C���9�D�R�ɢ��u2@���vj�u��N��dn�ϬpQ&��+�K�I���9�Ө�F�`$�~��$@/p�6��n��%'�|�H�]����3H�_�gM� ��7F���5�Gm]#�1����$0�L0�K%w*�R�O�N�:�@�G��Ղh"���8���?����b��>�VCҠI�2�6_|�-�����7;��[�FY3��"'?N���@���ΎN��١R)0j����=�y�N��������r/�)(R囘JMZr�K��)�ڢ �2v��&~��a�{����T%!�6)�V�A I�8p�K�4�U[[���vTTB��{>�P�F"$�b0è1�y$@��{:���Ir�յ0�T0h���2�hVAc�����5�uZ��-�e��R��dQ�2yVf]{%��J�Yx������<G����w��y�.�'��_����z{�e�=��Ί@��g,�,�=N#"�l�V��)+��
�.����OQ&��3������+˺K�t�++@�R��N;�}!.m���w�)��33�㞗��@�V�i�n�7��,I�q3��T�~��Cڨ����	�]�DX#=��fM���8�?`��hq���*��N�¤(����$��f�9�2\:cr2���^��!,y8X�s��C�Hn��G�ߌ����1����_���>Ą�n�]�͂�n�m!:=4�<�ChU$L�#+`���:]�=��ȳ�⫟��z��p�Ŏ��"<�a,�=�������
C	��<�H�0�۠V$���!ڱ�?�O�Oca����-6>�:��FZ�:�*�'��+����`� �Gl�����8�.���O�&:g��Z�*�KS
]���E��'k{0O��R7���r{ﺮ"�����=�����R�'��'��K$�ۅMRA6*�S�]p���].�Y ,�M��4��5P�E�p,��H�D¢+��޹����6yP���ٟX������p�J�bϨ{δ7POϐ��d�G�������4.m ����ͧ�>����%�
.��&sȜSty��M�1��M�z@QBI�(U�5�{��D�Q�U�G�$S2����'�w�W�����7s�N����`�)�q�N,w���C8�1�7YM�wR�����o�1�#}��}ƙ��_���V�?{�e�95L�z�%cȲq����)����0f�$47�ؕ̒��@$��%�ܜ.@onmጹ���{�>��ofևW���@<'��M(dP&V9�����3� �&bəҵ�s�E�c�e����ft8�,��ϥ����{��Ͷ�׽{ѷ���l�=_ ���? [q1*����EI��HV�w��	�I��b2�����:�;Q`���%�(��2 ��w�ԮAC�;2q5�r���桠 .�N�䱵���9�&�16��:��䖍�>r��Yju8Z}��*�t�-�q�.�����*��}cNL�Ű;��*g1��!�uO�-���<Z(�T�SZ�{�2}�٘��������GeE�������~��3t�K��P����@��+<M�!}}�����=}h�g�c�ǵ�zW�9.CO�ȏKZ����h&��z�B���
S&���ώ�~�2�	�z"q�i"�%��,��{q��2�^q#�J`��-�g���&-S;G��sNj�$��;0q�@<��[��jBs���~�ڏ�FŖ�K������=KW�S0� 1r�tp:�b���1��0(����0�Ԑ�u�[݊����W���ubŊ�8wBg�_~��Y�T�P��$ࣖ���{x��p�ð�/s�o���V���څ8i�'T�^'������:���x���ﯿ�%2U���g@'bz2����	D�Tɽk���L�$P�*	�Y@��.�KIi�q��R=�ަ6�@�!:u�2��!h�~O�$�$�Jrģ')��C�:&ѵ��hI�S "|N�z-sdHjת#.��X^����}��������:�K`����E<�d�Sp�9����!���h;]�%3��(���3��Ř��9Dס�1a3/}S!v8�*O=�Ԕ]�h��-�3[tl7�'}&���1HߏFŨgM~� X&f��6>��'�������j�?�M-���gq��Ir�2�͠��ba�����>*�ʹ�*W%1h�@��LM)]�#��ʫ����Gka4��h~�e?>���逭 V[�{sK������h�I&c�9����;��H�9�wt �l�Ɋ��� IP�B^G��_G�LU�kL�6L(�l�yL�#�o���Q��Z�����F�{��CaA~~�a�,p!ۚ}V6L�\^,u���KB-#���kU%Z;�8r���L��g�����a���TU���B>���7�x�k�q�������$�T1�S$����Ձ�Ç��FT�7j(���R�c���*j�\ڧL�ig���?��n�����a)(BvQ��AD�c���uG[=Ə���xZ����ÇH\O��N%ٳ�sU-\��N�N=�(R�����=FՓ��dk��>I3�Gf�}ҍ!��Le����22����I�4�^K)ٝ��h�[,&t�5���ZnDp������������ǟ�����"�w�F���I+�^��u�QY�"��Ͻ�7���O5V���C��69n�u5.9,�2�������
Z\v�w:֭�Ң!o��k��X���Z�Y������c�㖫q��AMx�"	�و���}��*�TU�ɍ@����������w�Ƽ����A��}s,���?a��R�H]�Տ�,^�V_�K�P�9��qR�Q���P���|�ï((��'�?��L��REr�"�s����	�{��}p���`�UJ��EuQ1G�k�%E�t�'��c�V?�CN��R
q"�t��%Y������!�I&X1N����&��2�#
@g�!(��Ǒ���I�s�z.�G"�=�]��Gd����N����4j5g�T"�"�;}a���.5�3Pv�K{��3K޿U��D.z[��Z�d.��T&e��������a���w�t�4wiF<R�yt���>l�0vA-�ƢK�KX������`1�)?)�F٤�So� ��������Ú5k1~�xVc�c�7x�n،�6V�"�O��G�%;�������̉4
���z=>/2
&Dt��N{'3��(�J�
Y��J�������.d�f!@'�pKN.�������o�R�4x��!Gii9�;4���F3�F.�R�H�
�$SjM��>�4�E �'�M�{Q-ɟE�c2Z����A�fn�����Z�=��/��m�|H��F���m>�tؽ>��٥�*�`6�aЛ8.�_���6���V�a^ ����ʱ�#(̲�E�s����n��8md.�ﯾ<����5����GLH@�v��9�{{3Z�-��8�(��b�F��	!���4�RA�nG��.��F=��
m.t�\Qw��ZeW-��ò�����O�_��t[���^V�+..d@w:���GyY���
��3t�`[;�LJ�+��.��/���@ti=���ho����`Kz�,��������/m�'�O�������ra_�f3Z�b��p��3з��/k��`��J��7d�א����VŵWLōW��)�#������_���`Igkv.��Y���'�̑zc<��쾧�펝p}�q�y�o��e��r���YP�� ���FV�
�P;��8�,_���'��ر�+{u~�s�q��E����Oa�����?�;�?D�dl�jx=.�����Ŕ�C�j�q�;����Ga�h��xZC�UB��_��)�/;¡Í�h���r`wRk��-�h,��"��\tq!�,�������K�.fPi3���,F#��k���')���i�9����%�TI��uQN���������zb� :�e,F��"���
c�g�&ID�7D|�h"��,4G��6�M�<��#���֣���C�g ?Fnk�vd[h$H�ĩT,$���/��*��VbO�߳��Kf�,�Oϒ����XZ����x����2�Y2��S����3��,�ʻ����\Q�S*�M��6����h&��QI]��d�JB2�]֭���~�̙8z��G�D@v7k��V���P��)�����}���L&��!��ea�&��Z���No.t5�r4j9:���\��8�Yrm�h��@Ss3
K�"/�g[{��+**��k����:v��r:N�@�D`Ӫ�io,+��׽n��F�j:V��f�\�m���k֬�޽�Y�n�ʕ���od��k��O?�4��7oތ7�|���v�3�|L�6/m{���{��u���2e3�R����/�:Zp�� T%
rsP^^���j4=���,���k��T��7=��mа�0����?{�T��d̂���〤$E�W5���B0�T�:��9��~�P&H��,%8r��QA��Ag�g3W0��dB@"������ 4k�Hb���q�h���M�!1t�)���4�Ú��R� �ny<d"�n�Icq,�K�:��յfL��6�=_���|��x���M�ܻ���7�4�{��;�>?��G��Ϧ�P
�eI@!6���OHBU���ɭKA�K�<�}�k�j�c+��?�Z5��5��P+b0�#�w�M8gt?�\qdg+���P��e����9�@(H�/��}������c'��5���{��-��f�CXf�B���W�2�L�a��~L<c8V?p#�V|��.,\�&[9:]AX�t���xx�<�U�B7�w-M.ĂA�i �ӂ�>�멲'狯�/�};�Y�H�h���ցR��N���G�ǙC���Q�\���,t:��Zx܌4Hݐ��P��l:3"��W�rMp{��u��eBI�%d��Ҟ�d��UBy�%�e2J��B�����)#���)�-�@��ɒ͊�d]MID$�dɄI��S�*)�W�V�p�5i�DE���!"�+S叜�I�"(D����T������c(�sC"[D��D;%F�5������ ��%@'��*�ICL�l�??	��ONz�.E+�{f��[ =�����t��LU��6[�%@��Q<��<"]0�}��r:�Uӿ����Ϩ<,:�����M�D�������՘6mZ[���0x�(<�v#��.��!hu(Ԥ��2�RG��lb����'Ű$�v:��&N�a�N���/gO�����E�����%�������~�BL���� �m�N.��))>��&��H�8�Q�+���D���8;�\�b!    IDAT��JI]-�6���������ASS���)���Ç����'?��#W=H��6�U�Va�̙|�/^����/��"����cs����o`�M�`ԙc��K��O��JeB��S�H��vACr�%*���p��(�NM:5J��oY_��2��3&��AKMM5���z#��^{��ۣؽ���!Vkya+����b��$�{��HT����դ(�������?�\�BJ�_ 1�js��q�`��iǀ�R<�d.I۶��}�{XwzB�	��� 'Ǌ`8��$�C:A�����A2Ǡ!#��2��Щ�����ꉂm�d��z��g1' �� B�8{���1���i�H� �Ϥ�m��v*�g&� ң,	�R@Q�*�����Ғ~xt�V���0J�d��A��P��ШHF�y�ذ�~L]LC(ĕB���t���Vp;�x���������Чo	�ۛ0f�(<�� {�3��.C��V��(��'���:�kp��+q͕8��ag=�-]��҄�67F�1�~ �|�s�,�2���F&@��� SE0$$a���mO<��m}9�UH�-p�b<JIKN;Mu����1r����/]��>e���P��,x�F��cZ���@�����
|�
caq�*9��"�)j�566C�"��$�dhI���Xj���0He�x���|���ƅ��x=���be�,	D����`��ⶉR�/J�!ݏ�ۧ:�eB�\N��t�H��K
�
y(		����*���>�Z��j����t,;C �Ѓ�OKd5�4J���Ͳ����������d�M�&��*w���"#��gÿ�d��g��dFܙ���z:��/��O	t��CF�M���J=_ Е��s)��*����h�fO%���*�S���'Y���i' t�zޜI)��j�ëx�z�$�rڨ1X�f=���rW��:�dZuP)L��R;�%���=)p @����_�u[�z����{��U�_�gz�����B5@@� �H��X����)!@��"6�"�H	)��ZBzv7ۧ�^>�{���Nv���y�<�ݝ�������[�{�a�g����C�����E�i��p��_�ld�~�mۆ��1gC�G���.s��:��xޛ>�,%w�|�����<��M1�(��ȃz���DA�0���rl��#�y�-8���E_��[n��׾q���3�jw�A!�b͚5�g����>�H&Β;���<�r�,X <��O<�)c=��#�<�(�(�I��&�D34wu�b����5w��,ݎ���uv���|��L��-#&K���B�v8�{�wq����G��1�R�����e�h�1���xM�9��xx�����H$&�i�|�bɂ�H6W�����KY�6�͍��p�3Y�FQ�ف��]���F�t�K����-�����+:ʘ?o�@�r;�$?��^�6w��M������=U01U��%*8W�~�=k�A� �o�7o�<�"L�D'�Jd�Ȍ��9$c#8�k_���(��o�2�ӣp7��AQ[�t�w8�$����Zm:�����7������k��
Dg=쏢g�z	��z�e������l��gx'�f�✟� �l�#{}�d�`� ��A�=��2j��At�Zq�/��^�7/�{������P�٤6C�|�p���P�6�m�q���d^y}^y�M<��*4�vK�X�7��d�|h��0i	�b�}�@o?��p9�e�I�C��X�u[Ŕe�h�l�n�f��� ª�ю��v�a��=ff�k�[+N�V����=��Q�v	+�:=�d�Âl.�\:�#��"��ɏdĮ�.��e����w�#�V</�t	�~n���J1�"oIo��B����̩���/Q�F=Ɉ�]��Ƃ���f�+�Ka����oqY/���l�ԜטZS�,��Y�59�HQ���ŎdLt��Ҏ�}{����Q�4f��R}��}袺S�x�����M!��?-�O��Yjz�S�ϧZ̻d�U���7j	��P+.�:eYR&H��.�K�����Rf�R��RX��?'��3tf���y���%��R���e��c�$�G��>����%�l��Htz)�Kt��H�k�0�9�sM�b"8sđ�a��.<��C��`�����6����	�I���ͽX��'(���-hl�/Ȟ�(��ۤ�˾�Zr'��F���X����n&�PØ$K��m�s���x]��G�u3"�!_���2�FH3��!m]-3Lzu+�^7��	�����%����ߧ3)��vJe�I-�qc��P���!G@�G^�ôysዄ���a6��XW'����ă�X�����}�g^��������������������hl��X,�����%g�\�⣏��m�a��{b����hl�#�ʉ�I�\����)'j�ظq�\�L��	洈�tشm;����;*�kٌ2i�v�?0
_  �s:������~D�
p#�E�̙�`������/3j�S䆀�ҥ�.NY���e����|��\Ѭ�-�O�R[�5>��'k���Y ��Yc{O�W�]��߼�z��'E_h�1�G1�R6m!���	fϚ�+/��d�b	z�[Dcl��C98�n����H��+g0Է�3���� ��L���Â>eJ�]��ւB�(�l�׆P< ������1�C�8���Z�+�0�`��PH&z<:��Ff���'���P2#�����
����ؿ�X�&J��,^�r	�tLuH���v``dN�G̗�����y�����wN>�;���Ӹ��eذq3۠�;E;�΃($𳳾��VF���&q�!A�/!`��@�$*�z��"�ɥaw�K�e�dP��ԎP(�M�{Q(R�GC+n��Wp�5 	a��i���_����կ�['�(�����W\u�ϱa� N=�t,�����qݍ󦺆v���P�F��P�=���Q;m)�"�d^�9]��G���-������?<t�bSSS�e�=k)8K�\J��k>�ؾ�w�}�>�H�)ꧥ��mu0����p{Q�a���Δ����P���E@�K��у����!�̌`�|g+e&���B��V�pwe����T��T����U��OV�S_�vA�F�j�a\w��� �D>U}����	���z�ʦ�8����
�������T�Y@����]}��HW_s-���W�h6b���b��7!��P��ds!�e牪s:-&8�6��1)[7y�t�l*�eRJOM��A���w_��^|{,��t��� \7RY ���h��d�δ�HT�6�[[�ibB@g况�A�K��z=\� ���Υ��$��$��t<��&�*$��e䅝��^���)���Fb0��2�Fu;�g	0�
�ډ���"����$���8jd�!�`5��H������у��?N4uv����n� �Ɋ֖z�)}}��C����k�~=;�q�_ĥ��t<��Q?~p��ڛP�<K>���t`��磭���ٺ�MM�w9e�?𣩱^z����OF���A�F_�v���tZtN�ｿsv_��7��[����hj�.��?��>�~�!�;�6�98�t&#<���8H#�h4.׌��̤��L��NEG{̱�6��Ы����*��`���}���a��K��W�j@Q�LT�?�P��=G=Sr��Ⳣ�� �b�L��l"�� �hmi��O�^{�}�
u͘�L�js@*���eB48
��}9C��b)�\1-��lt�.���ff��d���v��q��D�"c��P�+k$;-t�j���ڗB�i"��f@2V\K%X�&2R��5 ��~�\��T�H�&� ���bD�%���5O��R��|:%��y瞍���^/p�������hC0�R�=Q3>ܶ�Ry�<|�v=F���h�}!���!���(Pԡ�n�9 �M���d�JԪ_��bN��[�	[�q�W��w?ބ_=�G��u�x�w`����2	���;W����h�t���Z��:q���p�������N���Ơh���2�&�.�v��Cho���+��q�@"<��C^��?�^�1�b65�\.k�~au�ko|��֞ѯ���ôﴲ���%�5��f���54þ���_Gx;�� �K��#W{j4^Q���Xu�L�f���W��RG������.Hu�c�I6�����(U6��ҿʂ�� zu�]�}&�D5��TԀ����ڨ﫞��T4�Yr'+��[o��w�U���c�"X(����5�o�H�}5�Ij'�H�E*�FgW;� vkC��ѓ��F� z,�٢�@X��k�hnl�NwWּ��~�M!�x�[K�`�7�l���C8@ojk ����F�}J����&�%�,Eq#4��0��1�^[���C!�F"��2����0HV�d�[�Y]�
f1[��X/eK���Szo�{�:�^Wn>��v+±8�:��ؠ�ZD�-/r�6�L��dY��?� �ɂ��Na'ϙ;�7���T�}+���xm����04:�[oY��h�	'��hFs6m�E�W�+.=�������-Q�r"�����I0��g$
����R_�λظm����Sy�ݭ8��".���E�.[������~;��Z]��
�>��Ci)0��a��M�5�9`0F?�(�� �tF �s�ٳd{g��v}W�����5��5�׷�f'��&zmy^m�=��ڄ�v�7��M ���p��0$/�����X���fs�<�$.��B�g+Q����5ￏ"�x)�ɬ��l���m�ȥ��&9�@�.���T�bZ�/��6o2�Ln�TuJżI��s`�=�-�
4e���y��F)�M�d�B���E�B���e�#d�JKߺ�텗��dJ�'��	�Ztgd��8�u��҈~�4<��SX�n.��Rlظ	ϯz�hV*c���xHo:͸���Á{�M&�_x�M^�%	��;1�};��hj�.�AV��J�K��W^~U�����v��_<�h���W�@z�3)�u�m◰j�3��ފh`���.�2	�~����o�ˮ��]�_=�"���蚳�XR�-��D@kT�$�ԪG�*�Zd��@:���m�=��~�OK�;uJ���P��M�o|���������?xZ�`�[284ܛ�0�bu���=4��������M�R���:e_9�<���H ��)����W���L �O���^��`;�{V;��f�j�^��3���?Ɗ�T�^]�sȴd��9tt�������7��x�V1mپ�V��s<�.�\�l�d���yr�<��r)�9����_��^����ER���"_T�����$�[%�����\G%5�[�fdR1�_/>h��k!��9��f���嫹���n��瞃p<�w�}�5�6���z�V�G }xt��-c��jA��Q�����qC�@����DX0�|Ab���&	��,}��\��U�lMFO$8h�̀�Ş��)��c���:�gÙq:�^�2P�к2��"gJ�r�r��9d3E�;oꚉ�P�KZ��M�����݉@d �`?{�>���G���a�80���9���x�a�д:a�6�������_��M8t@*���􁡝���).x�����46�D��h�k��˯�wg|Ѩ�һ�8�ؓQ�܂�n�^X�>`k@(ĳ����´�2��F`����R����<�����;ޓs��x*�P8n�t���f��U`�jO�]o�V5W������������a{�`a���.�A�c�^�vt�y�,I��Y���{���6+he�nС�\F*6���/�!6lN`�5�b�=ȸ��ϼ �ۃl!!�ڒ.��^��U�f�((����C$J���v�,Hg�(4��R�u�d���1P+r\���L�X�JЛ��s`8���fC�U��B�t:M	V�y��	�V3�$:k�Bi�tˠ�j1��gPʡ���{�7��Ųn� ,�ǋB.O]=�9����A��p�%?Ü��uF����l.�h���Bl�'���"�I8E$E����~�g��ln�B ��W���mN��f._v�f�(��|��c<��ߠ������{�Gkk�?�|\q�5��y�����'�|�uh�n��v��ҷ�}*E��b"\�C[�CSHō��;�n��?<�w���1��s�O���y�������`����ӝ*�a�:�;�c@�����tM�(D�$�S�<)Wܔ�Y��Qq킛ꐪA�?�]6��l{L��
p��z�Z��U���"�JCS����D0��٣�?��C��I_���3JW���C�]�S�]�j.��S�W,�
Z���q� ��W^�����d�>���o��`�$C���%KA�c�8�YFK؃n��u��Y�o��,;��{�����8p���rY�@�8����c���Fl�ޏ}>46�Cg�!M�7�(�-<6t�C$l	�,�s^�׈s�̎�8�TS3
��Ib�n3�B4�C>��k�8��+^mO��J4
�A/o�f
�P�_W$����n�)��Ҋ�DQm�ى�h��b�q�tA)Μ={��3��ƭ���!WТ�{6�Z+,67�������(�������?�O>���_x���{��UO����~t%>\��/>&��l˯���m�����g8,�tN��O7P��n�YD���o��Yx�����������+�_�Y����8Ͽ�O<�:|�2L�6�(���1鴈��@6+<-/��q�W�ף��v�C��i+�^���Гi#���ger�.�W��ϳq����Q��U2g��E+D:������	)t�~{m�=~,
0O����~,P��?�b�Qi���tN1X�yg�j� b_,�S��3(!���k�����"l�1��i����!�����x�׿Fc�2��f��hVN��^�����&%�(Ǡ�6�3y8D̪�@4�l�|W�}�e�:lm�cQ���D4p���Kv44J�i2[dD[W�*-�RFĩ`4�`}	҉�%���E�yoE#!	��}�)زq#�y����p��<��6�v��H�Ël�~�:a}ۨL����A�S�3��UѨ���R�g���4��w����Z��0��ر��H�P���Sxm��hjj������Ï�S��v���w�y���x����/Q����b|��'�ܳ��?=��r��8�3�mn��oDA�����'�F}K��L\?�꟒��P.��'��rvs!���3�}����_��z_^�.|f�Ea�RNg�O�52%�{��/�����P��2g�,�2�vP�uT�**��}�:�Q�r1g3f�b$de��Z��醠���V �!5����#�M�}b�}�ܔ�[�^���a�d-Z$_�o%ZS�['���B�cVK�<ՠ�@��s�="Qz�-�3�ǹ?�9�q�&�B@Y��AX�l��R�"l.�Z�A���%�f��F�T�!9�`8���I��ދŋ�^{/Ċ����ւ��pځ܊m[w�#���-�wb�+�!�����#ėQ@�6n�W����eYO��'����b��x:Gc���G���|��Z�%S�}V�� ��1G+IeΓ�!3t*�1H�(���9 �K.�A<��bV/���Ns�;f�]�����N� x�q�W��ى<�
Ͻ�*Z:f#[��`s��mB]S������ނ���|�q<���8����c�%w��7_��k�b����	������y�:�i��F��؀��V����PP4�y�0P���|a�?���6}744�c��o�u�n�>o_�~���;`�#+��$d�2���3	�3�*^�֎v�%�(���&o��͖R"�|u:=���q��lYMFtˎ�Hk�f�G�J�Qq�R���ul�W?�f�[��5�i=h    IDAT���J#��{�����Ԏ�)��W]W9yE0D���eB��$�ʀyI��J�[Mv�M�\w�"�t�Ϳ����o��+W��Z[���҂��}�i3�8�EkaGo/:��*j[6*n�.> =��ȹ͜�!{Q_�(2�fN�R��Seq2�6�E���G�- @@��f�Y��Ҋp�/-�ǅ���cQ�A���Vc�=���KG{�\�����&����p�i�
/���������Ҏp<%�!ie�Y����ˌy_?�:�Ã�s�ԁxw��ٰǂ�D���0#�Ć�HU����p�LF��-M"K@��;�����Oz�gp�y�u�`�-w���"�ˣ���-�&y��5����O�KZ��<�8�}΅�"8������oO���t&y6��N�U���� �2�Ʋ/6��Ń����g���¾���g��=��K��n�D�lܧ���P�äI������á����n�h��gB�Q�Sa�@vv��>fʢ��A�Ʌ�Ay��[uOk����MO�~�*��(F	8V	Ϩ����@$m��ઁ���c�ߪ�>�LifMj�>vܕ]q�T3N�x�J���.փ�h�m�Ȥs�뎻D�ছoE*��E]��q��4����ދp���đ/�a�;Q���4���7��)34~nd�'	d��\n�a������3k6F���e�6��d	k��0��p8=��Л�rcBa�B��쎊V�c/�77
V2x�qN4���Y�z�M�0ط�X��wB��K��g* ��ףl���+��\���ßЙ�R��%�DT1�QI�"a�,�FfV�L��,G�6c%ys���Z�0�h���#�V-�ӑ. VO��v�����_=�(��v-��h�Sg��?�f��ݝ8�;��o��uk�E2���Λ��]�D&��鐙Ձ�;���n���lf���H'�$bI�(�b~��o��}:Z���ݍ??��&�t�o����:�w.d��Eǟ�Re���d:���&)�4e�� ������A���.؝�
�`0V�tT!hE:y*P��9qh��^�<�[�5k�Sk�ͫ�z��-��G-ɮ��j�]Ԗ���W�Ƙ7D�PE��\��L��a2ka��P*�
q�}�b�=��+/����q�|�]ۏk�Y�.� G��}w?9��Xr�8�Ѕ����K0�|��S12\�t��'_|M������[o����X�x��⡇�[n�����s��b�
t��X��L���K.]zfΜ�����Η\�-m͸�³�~�+�X*�Ng�}6�<&�y���������&N;�$��q�wbG�\�&d�E�r%���P�8���Pv��\m������C{�B|��GhpYP�&��Hۂ=样o��#.w=���A,fDR	��Z�f|��F�d0k��cy4u�į���\�/ԷuB�3 
c��y�sϽa���s�ѿ>���	�^{�M�]vz=�k�E���$��~�V�&�٦��J�KEB��p��ߝ��ɏ���G?�-��O���o�z��w.J�N���ʗ� }`p�H �k"������
VJ\�cr�im�k�#������`U�T�c��$�>ipQ�W��j�^��Y�|n&����ѢZr��R�Ϧ�r���
@Q!�QB�:C'谏y�-�I6D@�%�X�d)��җ���F1g�X��zt�?&+��(�P�d1�onl�,�=T��	���$�R�/gMʏ�
���L2�B�Vι�7oq���Q��"#]2nbs"�
8R�H���	)�3��y���Tx�I*<��*M1���=[7b��u�}�\C
[>	II)CKPeelM[�Ziu:����5�Ye�{2�v�$�2�,,6�R~��l�(�:f�f;�e��ds#������@gr��5�k���e|�i�lj�R����I�%�� ���=`S�B=���ۺc;�0����/8��p�.�pU �����}��T��vJ��b�4v�}��uK�����V��Ex�+�f���ȕLB��8�P���|B#;����2�H~�s����}���<I��^��BB�,��eO��J��˔I�[�^��H���Ts�*`��`�'(�NEt����}:��*�K)TY,+o��2Ţ$d���i�9�
qx�f��m�l������w��ÿ�=��쿯�7dq�����݁�38������n��u������p8�Œ��{�M �v��2���ģ�<��<r<N����ƛV�λo���ؼ9�s�9��U�~���ہ�����8㌯�lɒ��Ձ���ۢ���;Q(h�l�Oŉ�e³�>���n̟� �l?�"�WF�]rr�s�Ti}d)���p�9a5j�O�c7�G���n�K���w�����p O��tr)�&s�De� ������-���ς��F2���GX�} <�t���xJ,�WFFF��>Qf�[���M�nF:	�Ū���(J���.O�oZU+��|�8�`,�,�Ļ�^��k��c�{O�wOl�{襷��擾�����|�0���>�n3��zpt�/*�'d�J�������^��V:��ܚ9R���Y��؉Vz5P������{w�v��{���:��򅜰�.\(��1VYa�r�>&�[I�Q]��	P�[n�E�M7ߎH,�e�o����G<���،Ysq�M�"�@c0���P:�����vf����!;4Ǵ�]�1�/>�C��R�%���������� >�d�/�6m�9�LV�l�$`K�TVH8c ��5���߯(�Uj"xmXN�zWG3���8�;'a����^%D ��7,�q,��. ���C��[,*��"�(�#�S�Rr'����:\��4������wN�[����d�4���9磩�O=�
+n�-m��3;e���W}##hn��ͅ���&��>��R6&ɮ��M�x��w�Ea���-:�6��EA��Ԭ��-vH.��f������)A��xώ���lHg�(괰�dζgЏ`</�#��N2#q��1+/HٝLf�����-���GF�5�e��c���g{��,c�z�B�����V�ke��B��6��p�M�6�UB-�ͦ���X"�y-J�z��P�Om��$+U�<���1ѭQD(*��"�L����g�:\��E�Ll�����+F�C1�0���ւ������;wʄ�½���m=ؼu�ڛ0sv����{�E����?BOO���3��r�B�|�q�/��c�$�_z[�l��y3p�����AEj90���"����w�qb��OH ~�I'�=��Ǟ+ؓN���ܭZ�J�<�X�&f���pB�5�6�Ao���hTLo�ed1$#A9��F��0J�v�6sF��dto�����Fᴛ1<ԏ��F47y�O@�D��z�۾�G��c����:y�:�/��6��F1'�X&�S�\Q�)�`�����O�����]�ޥh�Քg�]�(J�c)�͇�?��=/}����7��T�f���WW~���6-Mk]{�#3Vr
�}>���`��п};|���R�����7c���To^-3Y��Z�Vs����ZRۮ���%]��W�V�F3��L�W}.���{����!c����P[�sx#TOH@P�(*��^k�y���c��(��n��7�_ ��W܌y�/��:�h]�f����/ jLz��Y��F�Չ�0]sy�4x=R¥n���EC���͞����z�m�,��4�bڴ���{�ц�x�w��K@�&�(kl��:/B���`��z��Y�%��cFN�&0���ݝ��نt2�l2
�͈z��|F��h,,@L�;�gf�ʜ���m����{�V���d�����_�/G�� &≘����荍M��a��Lv̜�F�1@k@�����QV;:��K�adp�$�]8n�B[g2�"���,	��l���)׫��l�s$��.l4�I%��L&�����&�[v��dA�<&�'r��,ۺ�~�kl�i�m���F�ǕX��	�Vf�#� ����Q��d6#��\� ����8���F/=	d�}�,w��]u@+��/����-�Okە��DW%a�Ț���+S?c�,c,� W�\�j�ܳ���efM��wA$g����Lы0����wRTC�B������2���y[�JT�8l&dY�����oVT�e�b��0�E�Ĺ���:�?A:�J�M?(ZI���r�"�/�>ϑ =HXc��l��u/�sH��k�9M#�X���
��L*	j�7����f����|6�H�-*+�!�XPO�M:���I�l.��7�2y8�MH��`k�4�l��쮇�B�L���$0%�OX��&Q��5�|����Ud�ſ��jW����u�1�b>��)g?��N�r���Gcj��8�~ѓ/�j�e����t�8�>�H�7:�9�[ }`G/F��QGh1��@T#��z������f۵�. W�"k_m_�'[��njRꯔ�k���d꟥]YE�S�8)��G�a���C��ƴڹ�V��m�n�tr��"3&�F� �=�7ڍ+n�|���Fp�h��F]C����Ԇ'��O�!�S��Eb���5��X� �`�I�����B%1t�hl���b�1��� ��d���Lz�[����a?F�a���C$3YxZ��i$��(�Q��=k�D&��$�\�Ã�?y}=h=K2[[K#�� �6}�N��8.��Ee���#i�O׸<�ו���S�c@�k�kG�^oE��(�
��1
E467#��f���SI���!�H�h�cӖ^��N�BXr��"�V�G� z���D�nr��Q�yy���.����T�K���Zс�X��Dю,"ѐ�֨@+�`�/s��G~��X�s�.A�,�j2Y�7X�3��'�5مG�mj���A�X�?�k���R{.OY]�>cP(k�N{&�H�Gr&:�) ^��,3�	���R:�j?�d�g�2�������]ZxU8�f�Q;�cr@W���*�J�=�`��+��\��tZ����{��o�fhijF`tD�7>��$s~~�.� ��D����Ћ\G7Y���أ�ϫH�2�ł�����SM�RmaՇ�?~mljW"e�HWs�q}q20Q��ȹ�UG�)���Z� !���Tc�Za�3�e�*��"�ʽȤ2B0g`K�&9�,���ݾ	3:[0�s;�]Hƃ"�L`�q��aDS	)�;]n�,V��N�eD��k&�u-�k�HX�2H�K��\:'��l�L����+�<f�f�5d�"�@�I�xDo@�+�q�@>	�EΧ}O��g-���Ń�����|������FR��S�~W!��|#�ё�,t=z�]��+�#*۽r'OU"�>�I�S�J��M�
���'��K  ��]��Tp�<��Yz�@p �����U�]���J�����k���3��sa��0W ����Y��W�$��K/_"fm]]�A]}�Y�bфd�
�hi;X�V�Qe.���E���2��r��� �z�Q�O�э��v|�������n!�����z�O~�P4�WV��C�8
Ͻ���-��H�|Q�[��1g�N�e�������F�u�XW��)S��?>�����eW	��󰡰�k���Jɝ�0�Q��F�������\Y^gY���%2� 9�sf�����8�e��d�'�6�P�l6;�_q�]��/���^X�z��xf�K�/IDDh��S��0�a��ǖ�ۑE �^��	�L�N2����a�ٲ?0"nKV�Q,n9��Q6��==��J��Ή9�kh����x��px����a�?��Q�����5.�'�����F�8I��_[���%�i�[�B�TM��P���*=C��S=d�����tt����w�T������iR�{���i+�d��(�s�$+�H/��!�Yr�(�:: �Y��V
�8�Ť����=4[x�N;�e��/�y��� �uu��@�A�n�}F��Z�:�i����uf	ny1��|�Z,��T?�o8��H5�׊Yz!O�e�d�±`i@6����g�)js�i��ב^G����yڹ�e|�{h,UH��<L��9h�Yh�i4���;��O���k�$�I	�#����X
�x
nO�(i��4u@g����L�BYڔ,�3  ���,?sf�hO�FG�BI-�Q�B�o`�Yz�fť�A)�۪��S����g߹�S��:?����עg��h�h�rT���E	stt862<�=}���>���q�e��,�q�����8�?`����DV�x�{j���w��k2�Z%��M�������_�SmNc���������
�qK�"�ʅ�z���e(,}�(T�rt�=�+�w�{;v�b�u7�v�9瞏�7mD{g7�}~tM��m���2�A�g��9ʫ*�.�4�	�TBX�SbF���~�b̗w���9D��-���މ=}�Lظy���b֜�����q,�݆XL�R��*��SJ�J�j����A@�qjj�Ⓩ?�������Ö���L>�3���Ҋ�Ug<�M(Kֶ� ���IO�I0g���=ߟ �Ϊ3�	�9�ì�$cX�9g/��kcS;6lځRق=.¶�Q�G��-v�tt`$s���!sY1��3q��Qf=P���z1i�0�5��N�L���m����W.�I+՞z��X\f�l�̧�(�!�+Y��BVJ��`Z�M��;=��#U�\�$�,��}.Y��haV�]]c�h�s4)�N���p�og�"~����VFˤ^mN1q���SքE��O����{5���R��5� i|o����~ٓ��d-�.�5-w޷��0n�)����#��0��z$ SD���I��{��#`n�Z�CCH�Zet,�ʎ�c����Лh*�EY���┈�h@2NA'�L�eD1��fwK��6�l ���+�_��CY�
O�砂�v³�
�9�'�Y�rߥ2���f%:��X����B6�1V��1��{�p�$�'�E>�{��Gm�b�����LqI{�w�%x�}j�;0g�<tL��<�,�]�u����mBh���Y�p�7z3��,��8�0p/�G�-(=uUP����l�	�3���lf�E�0
by\�'H�哣����o]r����/oj�ܯxr�������`�yx�l�đ$_���hdtd�%�8��۶#8:���zrY�l��R3K�Zc��!�F���ˉՌ��}J�_�;���	߫6(�C���A������ZZ�����^�s�=���eᩜU�s����J0����x���ח����>w�y7�}���ۤ��d�2���:�\���ՀX")d�S5��2T��(����w�m���ʕE�rv27�ʢ$�P����(e>�����V8���VdI�ZQ�j�'D�}~f��|�fs�����C	�|o�))�<\0�Pd�	x(q�� �����\�� �����0��(Y�hhS�Z/�G�޶m���̟甌H���|D�A��ܘMl��l|�(�ju�q�#I�hi��B�@Wf�x�ZE�'/��%��gF˲(O��"���&Z̼(�S�ge�W��Y�3��3jE~5�����?�L")
�@m�-R����0C�Q�%i�z��b�Z��a��0P��n5.�.���r�v
!����g�pY�"������?W'Q&��t��F%'�55R���Ɗ���E�}dVp�zmO@O�A��%Q)LU9T�ޓ�&�|'�(�c��WS�]��一���O^Q���5��tsIHYJB�4?% �(I��S��GU���9~ɓ(�S������]�-ǖ�QѧU��0�x?��r�R�5r�����f�E���T����V	R�(�HR�P�i�>F� i!Ѓ�Q��mfttu
��u2��v���O8�Lo�C{�sg�c���������]��I�����p��/��7��<�T�()�����47���E+.e�MT    IDAT��Az��+�M(Q)��ެ�왳W^�o ���"Iq� ���\6�� �6�-g�o�E�����/��69^~{�_�xǕ��e������h����B#C���A�m �ˮ6í� �/�����R�U��)����k}��':8�
��X�������)�{�����آ� s!�����U�4������1��.ǵx���bd�'Lv��\v�Ux��50�]"�h0Z��N0��D-���Bf�2���Xj��l�,k�Y�c����(e?F�����4Hfs�1�*k������L��pC `F��>�<���V�`pB %83���`��=�w*���܆�owܺ�p����U� 3�mc�NV+?f��J@%X1���PH�p�L#G���v�R֔�ہ�=;D�u��y�����ǻk�㪫W�s�<�5������"�L!�ʹ4����>	*tZʶza1Y�q�@j���GD7Zg�(�q���eػ,"En_�ؾm�����r̭��a@J�v�CX��P�;��$osK'��0:ź�>�;k?��U���ftL�s�a���!�L��\�:�*�ʶ&�(�'`.xEϡ�cU�
�Kս"̤��	�,�������:�2�%���T �U�#�B3�r���cF�$9/z�y�'���*��B6�'�L�mP�U�`>gˠ�����(���2'�S|⪺oTWA��$�r���BS��?>�T
�{��,�T`�\�1�0�ʘ`�p��|����q�J,4hA�+��8�&^|M!��2b���X��;���~ه�w�"�D�R�s���"O������m^�s̙ք�o��G�����1� ���]�܋��i���_��s�p|��x;����}��� ����>���}�)I�T���MS�i���*I���K�*�X�K0&נT@����D�x~Mlm�o�p���_�o__������'��aL��(��R��P!���F���T@���J���fP�_eUAH2�J4:U\��n-���Q��*���Ы�����߮�?u�[]2��P"J���0���ﯰC�LW�~��h� ]=>5Q�ߒFqYS�S�c���{��v��h�����&�u�H��ЛlrC��B&5}�Y�c��J���Vtʧ2�d�˹d����,*�9�2��L����8͍MBh�짍�q�I��اb��
��H�����b{�,���!�2�`�gE��y�]KqZ���|̗C!�Ć��btx N�M6��]!cѸ����:[�pG혩3���0��C!�"�H%�4,z�����js�[�*���}><��Ӱ:�Ηel��؂�`z���։8�/��0������?�g�܁ �,ND�XMV�מ��َ��!|�/�['}]�F�����N����S9�[d2AW{�䰥�ܬ({m��'�g�͉��Q4����oHX�w��[���1�TR�8�Iy�d�=��Ȧ�`9u,�U�s%�-)Sc��E�ͺJ:ը�&@-Q��t]%���JzE�o�/d���eϑ�a������YrQ6�	��ϛմ�W}}u�=t����M�u��c)[�����(��r����v��󭀶$V�ҕ��X����+R�H�Ch%`�B[f儿!�P.)J��eO|5�'jV ��9yME�N>S-����Ub��TYC(+�GʽB#f���))*�<9*�)�V�ق�ϯ������-�>&�TF�\3����ҡ��Ⅾ��YmH����� �Ϡ���`w��+!��|q5|ᔈA=��%,>�|���P��x�M�� ���S�]^�2υ�q;.���L�׽�W*�g�h�TT*1٣aN&!-������G߼��ӏ������k���\�,�a��I�EE�����5��N��N����Q������(�;̤�P�:?ρ�E95Y2�d�Pg��f���%���m��w��
iG]d*��{��A'�t�Ac=t�"-Z�y���A���׶�j����i��W��X��h���Exi�"�K��#��s�l�۶�2���8��	�̾v�d|$��7Gw3a6EC����\e�S)�8�6���1�Nا�Vau:������tc2���ˤ���C���t̞9�.�[�F�h>H�����+0Կ�B��u�<��v*�u1q�e��a"����3[^�ȡrc�<�����.	#��"�S$/��������@�ބbQ)�m��Ö7S&�6G�(���yQ���{ԋ틫��#�Qa�66�c�3V\�gɠ��7���� f�	_:�h���'��k�B__��#n��|Ի��� �N��`1����o��m�&�cdI���p{��|�m�BQ�^|�#��������������p��y<M�z�	q�br��O���J{�*9�*SS,@Ռ��e^��Q�L�*����U����W�����+hu?�LE��\T���\_�ngiv��rTJj����*)���N]BW^;��-���Gy�j0(��*��-���j��z��-:��f��5�����=�	V%�B��=�l�U�
��5p�i��,g���|����=V��˺b�NR��҂���%8r+��J�F���اf�^���AP�6���	���Ȧs���DX�g��ͯ���ߊE{�ö-c[�z�T ��fw��c���r��-j�7Fs�h�.��I5�sv���z����I���(6��B�K��K Ȍ�Z
��z��PV4�sI8-�|)�hެ�+�����;�R&���|?�ݫw���������,�3t�vћ��>����P��
����:�_E�X�Z�1Y��EVn8��4V��a�O�c�_��0���,pg�W}T�d�;�k�z9O�ѫ�Ku��:˹��Yr'��d,��N�^�U�
�Oþe�5<01�K�N��e׮P ��K������؂x:�ь��f�w���11��@
3s��9�>���@4�9t��%wi$�R>&x�������TN�W:�E��~qU�x�?��ᖹS�:�74��}���HVLF.�����F����s9l�sjm�G�6\u�������F*�����j@W�O�;�A"7�6ϟm�T0��gB@�9��N����::��*{ǥ�0���(Z;:q��~�կ�����лsNO3�f;�9F�zq�:���q����3NC!�ApdW,]�SN�.��r,]��Y��y�>z3�x�=�u�]p{�h�hǒ�/@[�0<8 ��m˨�C6G��s�w���v��MH�3�֍O6m����Co�b����q�1�a�ǽ�y�^� G{�^�>��?����׾���~�ۿ�7��?��9JqJY�b�+ ]��g@U�n��!kAJ���P��Nؚ�(�">S1Y��^'t%�P Nf~+���jB�Osk$pM�=�jm������U&1�����
F5oNI�����`bc���Oʈ��h�WT�,Ou@ѓ�p'��P������ă���+�W��Ӈ��l0TsIX^�Ck0��7�af�PTF+*j�J�p1$V(HK�ewf�ՀN�	q�b��G@�j��|F4:�(���߆&�	u.#�8��x��08�Uȁ�+)����=��?����@�`G&��
���Ī���a���}�~��?�e�q��� _E/���,Ĺ1�i�_q�3hU��b6	�I�r1p�5+�{��?���͟�'���޿�|������9�>���nI�,�P�PM����#�s+Vxcc�@'�(��)zk5}�Zz-�r���՛�d�����V��N��6��9��J�j)\�7���Y�%@�9rQ�</�:Ʀ�guϭ$���S��/+?n�$>�u�=2+L@�d�W^��_{S���P�Z����ɦ��k.V~�\��;$�z�X%��\��U�V�x	��DZ��S� �&�#A��`�ob��}ݑ����|�h$.�Z�,X��Vz�jB@�\@&�R|�\x�8S=�����w�6�Xɝ��%B����T6%�3G{�@AƳ�z��!<?�o��.�'�ل|�V��)��/k��֎#��*�|w^z�-�R%��Ze4����6��t�.��,\���2;n�w�n��W���ׯ@S}~r�YزqZ�[qѥ��[� ׉�_^|6l@*�V��<��oQH�+,q���׋�ӻ��b$�9��x�z����(����ⰣšG������?c4�C��=���up68p�ݗ�� �W<����GWA�� GZ��V��H�
Lq�S ^Y�ՀΟ)�;�3V?_}!Y�U��S�U& &����]�~��L"7������T�`��Ӵ҆���T���s���+O���g[SAP3av����6��
)Nm�HnI�/��!�(d���f��G2vu"�+dH�o���<�n���V��\��\�Wl�YZ�NYq5d�+�e�V��צ�N'�M�	�����نlZ��'ᕤ.��X)����D8m>������1�����6��sf����}oO?�M�����U������{��$r�6wb{�(�e#��X+cv$�)ddV2y�l�1�`U�D;�IH__�\{RJ�I��g�Yrʠ�]�r.�R.]9�E[N�=zm��3�<���<��*��ܰ���+k�}"Y�RZ��d�"����-�8�w�P �mh`pƌi�0�),�}^�SJ�*ީ�Ê��E僭&yN��O���HU�^���k��v�=��\����x5ȏe��Q~'��*��8��D R�?�̬O����V��&�xXA�x�:>�ƅF@/���1�ՀN7�믻ED�^�����d�k�dJB��A��N�f���	�Y&��-�1w�n]�Ļ��Gz�d�+7�2�%S�g�R7N���p��Pz�[߄����LgDv��Q�#>�I�`��5�FzckQG��(�1������}(���mF�ɸ#�w4E`�z5���&r�ҥgo0����
r��;�{f�>����U�^�\��^	����űyS���P�����lκFtϜ-��T"�;o]
��F��� )�O�O?�$R�.�t	�:jo\|��2^H�<�� ���yL�.��a�X�r���G��-H��7{���i�%W�#d�3~�u��K��fn@�sȚN��wH���G�Ǫ�7a�����ۡ�hp��a���(�U/|����*�yF}!a�r�U
���(��$ʃ%V��v����U�I��\�:PM��z�.+{���|������L��ޥ"'�Ԡ�KQ�2�TUN�eW�������$����2��S�Wվ5���+��JC���3�C�H��
�K�U~?v�&^t��Kis	Ϥ����� :8�.�ʊ�� a��'��%�g�.��:��� g5�s��,��]��U��F��L.��xg��;�3�.��о��i�77����㾎�O:�_�\t��5w.����m��N_���!�͘�p�~��E���"Σ>9l��9�8����+*���3�a�%�P���QםĿR&VaiŜVz�R&c��w؍�}��C���3��1�U�V�~e��֭?7�(-����	�����x�Á������t��8����@&����yL�d,�a9�6��l1O�aWK9�ѩ����Yү��Q4%���H�X���}`َ��r<2��h-Ww��F=�U�Z5˝s�
�]}��d�%��WS{�z#E*)%b��w�nA����n��7�B*WQ���V��"���;u�3)��ϒB,�CJ�}�[2c�m�V<��S�g���+��_������c��k��G�x$�X"�����x��g�sy��A���f��+X6'lr-��d���:�����G��H�<�\(�������7W��^[Wf�d�sV���{ls��B�,U�����������%������̞=[�Nc�\.�"����C>?\nl./:�fBo�ch8���yvW#`���m����{�fv�����
���z����C��g����N�6k6n��fL�v��'���W]��i�1���ߺ�w�fYYe�s�=��T�+t�t��D0���qfF�t���Qqt TtPg@E�b@Ā�M�&u����+�[us>������:U4�}����<��<<EUߺ����{���Z���'�(N�oT��[����)���8�d$$��LVx.�<y��c�{�Htcպ��O��S�<�N9��Kxn�֝t�''1>;��%\x�ؽ�E�s6fg<8zx�M`Gl�O�`̄R��J�PչK*Yb]9�g���i�;Q��TS���]e/�G^�HX�|7�us۳���B�t�� �+�}S-G}`S���`��j�r�����PzZ��#�]�k�)�l3AP_��vv/���8��~��&�T��g}���9	�b8#j$�{���:&���řR�QF�^����+H���T��=�L|N�r5��?M�Q-�15>rv��_���B~w�:��_(g�7��Z�s2V/_����.~�ۇ�o���s�|�|���#m���x�"848�_>�8���#S��j���$e�T�p���L`���2q��r�C��#�HA�Q���ȿcqGr"ż�D� <�������}����-�t�X���9'������u��K�zE��ǎw�:�����9�?�W��ڙU_4����	���PoTaLyZ;Za�N��^���-r�G�c&5)$$�I��y85���3�(�Cq*,�T"un�:�r�����o����j���I@wZͰ�I=Z�2�$�8��s����H&�@�1�+`��Y�FV�d63H4!��^�O�m8��Pb2W5�FR\&[��}�F��I|��6!_���B�\��=ΒKa�3�*qS�ҧ����9�b'�[���V\q�eػw76=�$6l<Q�m۶�v��fUͅ��x�%��\#�᰷��U������GGG�r؟��lz�lTd*%kw`��LW�rd�Vay)cZĝw|�1��կ`�� bш�L����W�/G��I���M���I��) >/|��.Z�3�)����c6�����U.��'��w��o��փ�7?����D�]�&�-����ǰ����/|�\�D�\�Wo�駟�w��=������m�}��������?�	b�Z�:����-�X4�+�e'Š"�����5�$���*� ���#�x��O"������b��T��/�A��%V�"J����f �i�8[�?�����5�@;�;� �h������e7)L�_���X�Y�n���Z]m�k&�ΞC=����5�@*	�|輌}.{_��E?�F�;]Ū9w]�	v�PE��X���iJP3�W<��¡�*ET����Ss{����}�z�CH�ck�hQkKޫIr�ʵa�X��lʳE�a�T���	Eɑ�D!3���et�K&[�!N��,���^I��qRk�[���ύ��I�\:'����G�Qr��f��NZ��\x&�`dp?^}�Y�-X0A���]��6�z^��/m���i4���0r�zQ�R����@�]��X�QM����	���"�Lbxl\y�@G!��LS{=���Rl��O�
�E? Z)�ШQ�р]/����p����g�\�v�#'��q�sQ{��sQ%��r��ı��ã��Tn����KR��E���j�
�O��@��r�� �v�@����]cc�z�{���?���	�wd@�v/���<�=�hg���7� /Y��\?�MX�����Ap��f��缛h��vu��5�ݟ�JP^S0�똬8
p��q1�����LG)�������FƇ�Ixs0_�ϙǕ�V�*�A��>��/�n��7�����/~��x���B�&D52�	�����V�^��E�IG���F63�5���|Y��ʷ����DjF�</V�v�~��W���9�\��fvJ�ʕ�'x��G��ϡ�g5�~f�Rh��qt:R��e4��W7$�SO�â���e��A<B�`:Z��������&�D�,�4����f    IDAT%��(�y�� �ߗ���O�V�w��L����r��{���j�r�c�c2�D0<:�cC�H�-�!��^�_�͗Iv�X�c���ǭſ�Y�df�O܌'�<�m۷����7}?�����������0>9�������X�z	�'��:�&#����n�� �I���M�i�ʌ����݊`���N��5��� )@ֿb۞~8<��;c����E��aڰ�Щ
ÿf�1���.�
'"�0պQ�4�ѹyf	(� ��0d3?�㼄�	��]�	b��* ^w��]X��"��'�J=pn���ne�R�e�,��N���1��y��&�N|�]PS�E��5U�oos_����޻dnZ��.�/�;��]Z���{�AM�lL�E����# ���g�$�IzkP�%,�\�T�dq�����0�epD�gE���C�	W�^'#_:��ĠH�F�o 33�F9���(���eq������||�_>(I�?��}��7�B�T�s�oG8Ԃt�F �_�鲁�?���
٭:�]�DØ�P钒�-�҂��rrN>��*oR%��{�J���e&]�׈~�a�U��X̓�����#��1O�Ƽ^;����``��1"�R%Q���*uO�ϊtW��
,��GMP�j>!�z�a(T ��Tf��ȱ��zz�é�a�����̈́OK���d����>f�����z��U�k3p/�f`f��<�dɲ¨R�W9��E!�_"4�ꥸf��=4���cq��I����/��ŭ�����s�V���
�4I6tDf�8uCR��_��]B������S�|O?�Ŋ�L���?�j6
f�*�s����p0(l��Q���N,/�|뛥_�k�	��?�0����-��T���v����A���g���~��^���=!�-��/�Gd%�"�d�;��l\��:�>�[���02<�+.�;�����>��5!�A�T��F��̟�o����e�fB�nH�����$���(d�ր��4��*�5^_P\�hMhXT� ��e�Z;�����lVZo�x���FjzJ��/}�%8�ܳ�^�-��o~[��}����_%�ԇ��ʜs"�a�Q��`��8��S��L�3OC�� ==��}="�ID�HE�\^�{jr��c���8p�(�P1�O���GZq�脨c�AQ�c�EϷJ9�`X�H0"�6׷ �7�V�
2��|�
��ri����2[���׷F2��)�ywBp��Z����O�Z��G��5j�R��D�9�B}��~������+r�NAsg��0ؙ09Sb?�B�?�����L8HJt�#��\IG�w~g;-�y��J�J�]�
U�L�"=�u�v��+R�u��uCa�'a�Yt��uZ��9�4�5�+[�S�7�)&<rq�JT.�=���G���+����.��)k��D�=�$.��bA$���������q�_>�0E�}1F3%TH��?�k�G��#CB�?`IR��8A*(� ���vC�w1ġu��j\���?#	�H�^^+&CD��w21a�_�QE�*�E��.B�R���z�Z+�m�Z��̺߲��c�0�,�l�P|Ax|4ݲ���Â�����SS3[��FN]�Ӌ�ߋ##55.�;U�H`hfNΌ��E�W7Q�L�i�N���H�\�[��ݽA�!ֽgw5��_ۍ��ۜ��<�MLс�3�38�4�����,���'�߀�����EL�J�Fɭ����t����9j�_ӑ�y-�v�]:6��>�)$���[nœ[�G^��!���@��]S1N��%�RU[".��5+%���s����
�}��?��d�<^9W�W-�<�p�=�\,^����'qɫ_����k�~��-I�T��|H�wI�:G�%����L	U�hkMȘd,����j�,��뫤�DaB��r�����j`���c��c�ug�� �9tBg�d82�k��ρ���� 	h4q�}�184$��sλW��,Y��<�����$a��B�!lW())����+�l;��PP6���I���틥d�(Z�tlZ�z-<,�� 了]��a��Aî�Z.  7��d�s�JCZ�C��y�t;���8Nɶ�j&*싚idO#��*U����I�XC�g�҃��5
�p��e�r��Ri�U�8*7�>�U�`��Sg?9^�K+������z�h�ߙ0�2U����ݽ�&z�{�J�F���isV{a�}.�3�/�,n"	�ޜ�qs�3yMj�ñ��Yԏ��;U,D4�i�E���ȕ@�>K��5	�9��'�2�t��|^YwԹ` g��k,�:��*)��+jt��)�OJ$|�H�r��x�)*�6���4��⵸�O߀��Fa��5~p��d�����߇+��3���pR�~��&ء��V��i�6��G�<��mAN+�p��7K5�[[n�N�U���:G��,3��e��dI\�Dפ�l�ay��[d���|)#�B2�}^g\�Vʢ���3����=�N�^�)<Z���=M*�������S��-��~��A�&�d\�S.)�$38~�>�{a/�m��rl�?ֱ>�3Oda��y���ޝ�7����B�c�V���8?7�&��������&��T�n&��OL�c��U2��YJ¡��y�I�`��0s�Z�|����Av�)�n��DL|�k_��c���'nA��7|�l~f�0�Y����Q1n��*cI��Uf$&%��M�)<��S�l�R�^��^z)~�����			q<>��Z�?�8�}�e�I���g>#�6�6=�r�F����	4�5�ʹȱ�%�����3\B�bC���q��g��%��y�B�������7/�YQA.��.���y�Z��0���g�=�'^w&a�'�V���I���i��M�z��y�.^�c�3�?6��̘T�0C�B1AA�tLL��&G�IN0a�g˔@U��Pj�J|�U�)ژzn"�i]&0D1���������Wme�Z̫d���j�d|�0F'��%�����M�QG��!^/=�=�&�s��:�|�^�$�Z*�x�� �{d)�,�^%��|�K�DK�`�95ܪ*L���km��*���ua w�̀������u@?^`}Q�>�MNo���4���P�j�STd�o/�&�id�aQ�pa�S'��MT�΂�Y�5��~��Dp�Oן��Y����s�c�+~���<�8�L�վ�
1"LԹϰ�#��bQV�
n�וֹ��k%4@[�:�q��@�����߇Rf
��yx��'aUO"�:~��O�z	=��E�r���x��G��_�CC����c���ر�_Hq���c-ȑgT�E�.B��-�L�s�(�J���'"RY�!�7�*y���2ҚC��2؎t�F^;��B�V����^i�z2	C-�� ���((�a�l��6��8
��&5d�Xl�'Ǧ��=}ْ%|8�� &�G���MyP�Ǣ��4�������Y�;xK tsP�~4f��,ua5�!)�y��=<�[W@�=1EBqf�>	�N��>g�n�?����as��W�΀����o�%���8 U��U�!� �P���p�P�����٥���A�i�|>���|�8|�(>~�'�w���	����b��ƥze F�n<ph�*c_����хh8�p0"0���*�ǃY'���D�Mu7N*����q�B,�l��'�-²��(V<�D��Rl[���<r�����8���dzj0h���4�F��LZ!>MJ�)���-S<��`���+&<&"*	P��{�{�5��vfY��&�v�g������ �3Y���X�j=JuSY[����+b<�Z^�#�ID���2���`���3���@6���n7�H�(�K�w�dj(���>L���P��k�P'��4�2�{x}��V�6U�*��tH�� kX�^U��\�I[�~�NM{eS͗��D$��(U*"��/^ך�L;d-kҩCs��f��ҡ��]�ׅ���糰v����ɂ�����YQ.H�_�=�v��T`lSS����L��������cq*uUo�H�j�ս7���"�}=s}�DZ�>�U����{0�3E���{;��jU?��:�8ɭ�w�jMqbjJ�I��{"��<86�����&R8d�9&=NW3>��b�Q�9��Gw2���)�W ���Gb�d��atr���wallO<�,�'Ӱ=a���w�`S��0�j���d�mI�;*�#'����h���d*�H�EFT��K��~2�I�@S*�A��2�"g͖��'�*��Y�p���r\��=�(��D�_���g���=-]i�dx�h��7��	�I� ~K
�f�>99�ild��eK��ᐅ��1:ra�1cS���Ct��]S�qZ��Y�;�k�p��ug��ݝ<��D�&�͵J{����@4l���Z�}�@��d�J��"ň�sp�xu �������6d��������_�/|�H��J�`��K�,]�QdbKMZR*U�8����>ě���ǆFqÍ�F0��?|#|���x��٠})����,4���(�E�r�,��F�H�5���G�b%ȬQ�a�U�:υ��5�!6��f||�d��30j!΢�em6���`8$ɉ�S�L�G��&
�4b� 6�_�5+��7����iT���!��7l��d�.�x!��PU����7�2P�H=���y~�>pJ!�'B4���z}�X7�|�u�{m����(���=��h�Y�`�l>_�F�xX���5,�u���N�P���kί�e"=>I�,?Y��ٗ�|HHc�ń�p���[;d3�m��`��![1���ho_��)��w!����TeF���q��̠�y��D�]�,��ׇ��:_��Bs��6M&�y����kR{�+tknbF�1V}�ٺ���~�	�{OY��������:�L�x��E�R����o	t$��u!*�?��w@_��������z��dD}�f߫��ڐuR�*s�|Q�'B�T�^�$�{�jٴ��-7�l��d�P�����Q�M`f'�����c {���$宩x�����y�G3��DHx_[��#��r��?��=���
�
z��^і�۰�s)re+�*�.Zڐ.�Pk��A9_BO{+�:�(fӸ��q�~�������v&�t��~Ë`4&k��U*�Ē6A�|N�h;�ϧE,��9��#�[>_T:ф\�5n�/�!r��P�����6�a�����6��HA:�r�}�s�pf�Ч�R�>���K�Z�� �<$��ה�k�Lȝ�O��HPs��	=�w���������#���2e`V����#���RAde�d��朹�]t���p���h��*P�T�
�P��i���
x�7�݄�	W�EA*&��G����!���1鉰�*{U�K�5K���"	�,6�T�"_ �!����h4�w�!�T7��)��6>𡏋B���r]$)O�/�Йa3�v�J/�Ѓ�6ꬳ����a�q�V�'��$�0A3�w�� �10����[�dƜi�����+��� �53X�t�L~��r�9W>�>�MbgG�{��X�r	n��11:��e
d�^2�b� �g�y�X����A��Dhj�KPr�.�?���Ǯ��X>���7�t���1 ��	�^��֬�}<�g������&���
'��ɥIěIE6����-�ka ��y���.	�]G��㴭�W��{.-�x����t���Vw� Y�>�l>_�A7`{9�@T���� ��r�d�Eq :��I*�dӒ�0��5b��/n����&��FLA�f����[hzIB� �Y���d
vV[�3���-�Y���߻�N���,n?v}�$�M���A����VYR�)�*_/�qsU�*\�	���4�x�S��k���x��o��F�u�����Q����q#�^�D��6��*�
�>�ƽC�υ�OYV�`�M8*A5�=95�a2.��Ӕ�G�	;���x�+TSR�����H�h�8�FM���BG��ߋbf
� ��℥]�J�q���w|��)���l�Xo~˟���6cf���b]H����F�/(Ē�pɢN��Et�%����$P��o�6�FƱw���.#j�J��Z��`z�LL�&yX��\E,_ڃ���:��Ʊu�3���#x��(�?����ʄM�R���1���D�7K������#��D�a�� :�����C��B���蓓��x�����u�W��ۇ����v�7�b:!�G��/6Q��Ke�kJҏ�+%9=&���(��ʡF B�=%�72G��R*	�Ǉ�K	AV[�0D�T�,�o B)��g�����){L�;͞(�"������&4̙qV|�xc���᜞�� ѳ�v�"i{[��Z�:^l.�H�Z�r%��J����NA2т���j���������*e2e5h˃/U�,I���<r�~����ʁ0��_����o�S���ྟ�=�	�|	� ZA�*
�IggEx����]��gO��`OO�����2Յ�f��t,�`�"�u�q3�p��U� e�*�&&`D.�z���Osi9X���]MI�����l���Y��^���c����$;ڌ��ԕ�;7�Zdl31��
Up�:��\�3���q0;�Lx>+$��ΦP�d�H��0����c|j�E���
�a�1x�qT�m�e�$�U��kMW*�q�>�H �ɨ����1OWU�ʉ�?1>*P;�?�bN�ΰ��l=�_��y��
�9%Y_�DW�#N�\�#�ˣ���R��#��D��@0���d��v����Ų>�.(���n�Ꙣƽ6�Ȁ!���X	�$�r�W���	:	t��嬯��Wς*|~%�Ti��mI:�Nf�AĀ�?�Ȝ4y9�TGc^۵�֛T��82�j��(K��L�ز�y�P�MP\�yV麷�����ɏ��_H��܂&��sR.um]| y�T@BH��r=H8�]�V����(r���i2����#�C�<��U�Ұ�e��N��#��hdnF�k���1��1ؓl�x/�R��$�����G!ˇcG�����k/8�q�q���=��_B,D����X7|��{?B0��>�i$[���3�pt,���N�L�,����j�*�Q�%�������w��3��C;��S�1=���;a�8�T�|�0+e�_���yV>��ϠV�#����}�]v>p��p��𮿽��~Z�	lذ�DoټO<����r�v�Rl�9���{�噽864��\�<��Ӹ��C��;w/��m,!�%�?��.��(�J�����;wl{���K�<D��׍z�p��^�
���Rٴ<���{�Zm���k(2�� 2fen���4^�{qԳ���Q��\f�+<�6�0�du�.��p8j��/<�F�|�a�� Ê���X�:��p���:a�O�lzF�~�D���@,E���U1;	ǚ�q��~^���E]$��x8C����
jV׃�	j�t�J�Y�!-n�UI4DO�Ti���x�w����O��*|�_��?�1::z��zlx+NX�TjJ6�j�"��I	ad�CĢ	%�Z�J�KƒjL��㥂|�Nn�k��h$"J�D�V�+X�1d:�c쥩�բ" ��� ��ƙv��(I�âg�Y-�
��A6=�k���G���Ǖ}�6�>!r�^]O a|bTԛ<\�yz����hƶ υ=bD����Ė�RyV���<~8:�"��������9>"D3xP��Q����sK�+�WV]���\�i�K�_��\A�����B$�R!�M���� ��]������S����|^ą�������$[�G�&��R0�fp���M[F-�X8\V��X%	s��(/�v
�S�3����<���(Э���^��suWj��u"�0�� ��[7l/���tK����7k^���Ϝ��"�i(r�b�{�D��E�OuƊ �*����2wol�ĝ������p���^��(��
^�cz���v�ט���Pc! HP��Da2�k|    IDAT�������J��%��cφJ�Ԝ�����1����D�h���ӝ�{��Z��c�D4K���#��f��ܚF��?�	+{���3ؽu�y��(��&fgom�}?�v�܋�=�v�>�ѩ�&��[��r]�5��j�2"� ZA��T�T{ıc��DڹX���M�/<�|.�E��H���A�M?R�Gѻl1V,��֭O��x���7��n�go�ÃCx˛�$$�����U�p��>��O���k߅�����{�/��|�y���O�٭{q���h� r�:>N�����,����/���F�_��3�/���Xv��c#C�P8(��u���te������V �R��ZU0�W:b��\�����0���d����G� <�z��`�f���I�h^�h����!-_�V�4l����X�3�x�zîTju�g�Z�O���D����$�6�}���*e�P�CC<�9J� eY�ʼ�$�#��@1���]np����?��5��G>���F�J�<��E�����]`e�/�ڣ�����\V��d2�����sq��&��~��������=/�}��b�Nx��y��g�u���o�{�g������%��-.X�
��~+��t�>��<7�pxK%�s�3��ș�-��H�I�u�$��8����3�!�̦F:�&�/@��G&=��O>S��D[k�B^�_�h��$i`���&�JdEHd������&�*}��e�vn`���y,T���)�ܩ��#㸊�b&��/ĹՐ�H6?��N������RMi糅��Ǥ����OMNI_���5��U�_(�x\>�}��h<���$-Z$�$ꑳQa����T**A�|���A[G�����i�!�[ԧ6EģVq�euӃ����=�b���*��W�B�7I�L��IF�y
!r�T����;�ꀣ{�����
��Cn���E���ϲ;�X���&��=Vˑ4���	"i�t ���1�K�ˍ���H���N;�u�T�̀=Gvsp��+�~�ﺌ;H��w�]:�M��R�q�WĢ���������<��I��[~0[|\�"��c&=�L텤���ߐ�"^����}�8�C��8Bbj�]%�����I?���	W��
�^E-
J �f&p��'�s���gl���Qڳw}�vԽUQB�Ǣ�>\���كo~�x~�^�2eLd+�[�N���/�eؕ���8���IepE�Q&��l��Ц��Y@B!����pR&tض4l�x���l��0xd���w⪫.�{��g�z�'��;�oA�-[��W]�7������k���d���ނ���*z�:���?��A��(�-�k^V��9*첫��c2�֬��";x�`�mۑ%K:+��	�eE`UO�V��zR��Ql�iF�Uz���eˑZ2�l�Z���
ǡ��h�ʟː"�O�\��m
J���}>_�Ѩ6�Qm�X�4۶�J�f��gؼ��6s�o��F|egN�r�sE
s�����
�K��֫��3���}�?�]���F<B[2)dfc�]�b7*�B�M("@�"��[6#��#������d��d���h�tF<���^ր��>���r�и�}p��Z�!U��O�~5G2�	a��w)�._��Ͽ�����[?'�w:5)7�}-T���:W���:�Cy<LbHȢ��sj�+���WV$=J�L���g�� �VnlDb�0�E�NlS�
�'9��.:�G���H��(Ꙗ�=�xo}˛��ǑC��Ν��V�e��L�%�¾���eqƙ�`���|�n�:y�v�؁�N;k׮�?��T꧞z*��>9���?{�����6�|:�,^�#Gзx1�862��=�$R�<��ؾ �V�O�e��{���hxY�)�=nx�,ɂ�����9�m�[�T����*�\&�EmmH�c���N��#���[23��MD�����$p�ȱ8 �h���$�Ĩ���\�� W`PA�/�rڵz<uA�xߔ}MZiZB��U�z��V�J�N,�c���] m���p˱���]�.������V�;{�2��|��tݽ��W�bd�պjj����ؚ�kb"�M��2y����j���_m$��fW@WCps,y���	�|�qZL�4�H&�B�k	��)Pm��,�/�`�R3��Y(g( qjd��ًfS)x&zzzd�GQ��-H�&��R����ɂH�d�E�t&�ݥ(�gR������-~#I��vMi��$�P�	Ǉ�a�PD4B�21:x�0.<�4��u����h��G��C͠"\�pX��U+��_���<��D�,Z�e�P�����鑪�݈�&�q9�x$.<�d�Sa{�H���9Ba2���jqv�m���H�C�f�p��^��\{5n��ø��_����e�����{�p�9�a��m�R}�?�G����q�ߊ�;v�O>�<�{��]�{�ȕ��c(�l��1�d��*��_�a���߈8�����>��z���(,�NL������>����/��m�pL�1|�ggR0�T
Yy �(��{����ig338봓q�i'c���8�o���uu����yFf��?����enB���{��������
�p��ad3�/��݋C�ajbRT�֭Z!�LL.��=t�.��0XLN���&0��!�hSs��:�n߆}��ɆLș_|�����c�ҥȧ&�+�7(n�D�l3٬^B���3�qB<���T8͵�����XS-��y:�F�XE�,�3��9p ���%�D<�5��avzZ���=�3���?�1֯_����z�y睘�����g<��Sҏ"S55=�o|����p�I'��ۿ*��u�]��|�;طo��nϞ=�����5��~����ÿE._D<�"������U$	�0L�X�FbI���$S(���ȕ��aH�Rf�
vtX�|us�����X������8|�
¦=]����������S"�I���_�jx���=6�#GF1>Q@�PԠg�bE�\@��
��- ��
���/!
#�3�����f�˦���`,Ҥ�sB���0s�̖
2U�r��
�Z�S��~	W�Y��QyQ�������9V8�,�]vؤ�4Kd��i�=����Q�$�B��VK�E��7�Ri	����5�������w����4��h�&�z��\iū�Q]��lQQǀJ�uV�0�D�N�����_�1�����%����NT��"J�g7.�+�ТcD;Ԭ���%������2���1ARZ*]�BA�"��˨҈Y&��ZcA5fgyQ��Q��u��;[U�b3�9��m��Ht��
Ej�x�{%���V"�����hr($�!�a������N��5J�Ve��38��"n���o��������n�?a-����/� �|�?
���?�я𖷼	׾�Z����q�o�-��~��aXQbm(V}�4,�XiFe�I	�'���	&��l����?��o�}$�h���o��ÿ��W�B��=_(�IR�7��m]�]��K��p|��J��^Ɗ%}8���0����El���ضm+ҙɬ"�0*�:V�^��֠sQ���S������Ü�SK[��݄(�ϑhU4!�Z�J�)�ϬP��#��ܬ�(�ך�N�� ��`tl�JUHl|�	�3k���M���̛�0��9N�|>̹tJ~����4����R���#�F5$�V��C�!�����Nx��@�+sj�3P�I��"T,��T�h|~!�����)WLO����X�ՁW_�*�^�
�����~�	��Dp��M7݄/}�Kشin��6�!�����\�٥�t+V��{�D넍��,�Tj�\^�ed��g�¡~>mj��൧�� ���i �*�c�@��c[��\�Q�"��MMUP|<(�-|���E,E><���h�X���G���c"D�Z��9�����x���x�oơ��8ҟ�l�+D׸q�L�
Y��}	�-�#�|N͙{}5�[E��QĈ�˸�r�z�̴#��{Pz���ȩ`rƪ�L��5zu���Jz� ���I��9n�b�!�l�tsiF�iǜ�x��f������A�
RM����yGOCF'�tT���Ɉn���K084�0��!��$�1;�((�������1��jg|��r�ys�L�4�2E���;����Hb+�V(I_�2-	b7iӕ�3���"W�=D�7��r8��k|���<G�*x������/�3��͆$�l�QL��1�|�,j�[��e1�VE~vZ��z�!#�H5d?K�[dޛ�7�h�/�,�;/|���RہS2}RTJI��x�<:�q|�W�:��'�����	4�p䛵J8`�?��y�[Ձ|�^<�⋷ނV�g�lyj���N?�L�̹�o~z�<�l��v9�p>r����ݩ6,��^���h�a���(�"�?d��~&��}z��������v�>�-������M��ǁJ3��]jz3(3��MX��BLD�hK�p�i'������{��Gd�KVmwON8�D�Y{�'g�|��<����VU�@4��%{��Y�0+��Rl�E�7~q���%�`�y�`�XY �t&�{Z���z\+��7��HvJ��8 ��~(g��Ĩ�F�>ǖ����w�h'�_�� ��Y��K�p��B���L$ZT�^�J�;��O�j|�'�=F�G���A_w��yx�_|qN;��a=���X�l���GG�%�)�[~ԔCD���W���E�2�� 2ż��t0A����6���ZjT���!��M��h�3at�}kU�+R�,�%��T�����VqIԲ�x�%g�#��K��u�L���Na����O��D<&�.M�j�\x�؇��^�L>��^}5B�.<���A��#�� �����8�s��_>�ǟ؎F�~��2�e8�Jo�p�0�4S~*f�2���.,_��kز�Go��5�~�����u�za�-�K��E��w�u6���{��e���R�/�w�sx/�%u��Y�+D���XN\�g&��Ab�,N9�\|�y���Vl�;,'$u����Tk$��U �}��؛�r�I��ʜAJW�z��x�f��19]�+��!҂hPYУ�{�u�
�/�lSX!>�^�+�����b���$�dz,�M�N��:q�>�>�U���d]GPk��Xǃj�-H"��Hjf�Т<������~yV��=fZ��>�h��41C��X��
,M+�h[;
6y�l��*7����-S�p(D�|)�Bf&��.��H��a�mQ� �T�	��ԍ' 4�At���Y��\p��(�ӢvI>y@g�u���{v��ʕ�����&'��X]�*��e�򩧷��w���,v�= �9�eS�U/����e�����''�/�sϵ�����S�Ŷl�,P�4$��e5ٯ���+R��E!���$ZcX�l1J�4�>�t?�ggd�S� ���E��[�������h?�	��ég�-�$$\)'/�WH�aS�@j6*�Ѣ�2�.r������g0B�P���|/>d���?O�sj����E�]�Y1ss]�b�T�|��!�Cx����?��"�n�>���/��l6C�W��:�j�_6�G8�?��8q��uFY-rޚɌ��92��w��=�I��d�"�g��x֫�����"J6��_,���;ω�I"ކ�[�K�?��_��ѩ���iҖ��%\E�殾eL�� �h�����(ں!���ăcq4+�J�FC�>���ϑI�P4��e�笠]i������9���t-��~}߽ظv9�.�ÖM��M�gۈ'bbiE"�p��He�x~�N��v��`<U�o�c<��8��3���^�l�N�~�o�4l;�z�(&UT�"|nʊ�M�z9��Q{֮Y-I�~g�$�c�Fg]t�y���b͍Sɳ�V3mB��!�W�	��M�~#�Z<Z��-���:3���E�J���	�˧��"�I��,M&�R�E�~̤F�jy/n���C4�?�b`tFxu���W�O'���;KSח
�sJs�_����Ά�usD>�jV����>��8z�l�Uף�����H'HH�f��GmY{\�k"B%=tuĚ� c��^�bIf;��&zUU
��"V����a���-�}dAd�,���ut��P"Z&4�d�pf;S�Y��ȵ��aR��?�G[;0�ck��	�S�M�B�+Ā���d�s�i�)�_u����}�\+xՅ��-��K��Ϧ�E��>�B>�d4,�C�hD
GV��PD%5-d����WLhZ;�8p��&&��K���,��;���F�m3�,G()�	��o���QA�cc����_��S[���@�A˹JA�#}&5&�/���R�B^���d�r��(�<	qo��R��Űg��8��h4(��l���]z����@2$V���c���bwJFt(u���je^�FPHZ�/))�uW4���Ư��H	��2�ͨ/���E3���i�QL����cy7����]�p������)�Ku�Z���O���"Ѥ�67h��#��8�C�t@�&�p��H�IH $�&I
�ㅁ�2w��P6�$ӷ�c@f89�Q%�q,_�TFԨ˾~�LNL��ƓO4�`)z���%��Ʂ5�9z������..gG��&�ZGE����q`e��K�ur��h�^!A�؇��o�	�*"z#���&9A]I^�0%l\҂���!�r�8 o#��x ��������
�9�ю���ٗ���ڃ��ێ��i�͵�i�q��o ���݆���j���.E�D��g>�+<��>��D_�Z���+��r� d'ga�*8��d�:tp/�y�ո��xz��~�7���� ���D��E��x��(�U�ǍZ���l���ȳ���)5���f��`��S�9�&��;|$���_ŴWϓFQ����1~(Ĭ���������Eh�VB4@8N� :�ίނָy᳷=�Ƕl� � αM��UB�A�Ӣ#��u.ϒK�F?ǹܨ�<��9?A��u�`�ǃ���1�%Ϛ�\x,<^u�� �V����ޚ�Λ)��(���s�S�����sP�*lp��ҳ3�o�D�X�E!=��z�_��+/F��i����g�a���&��b���^!����>�*0�Q����j	�B5/�OA�i�Q%� e_��6��eՀQep��$��d�=��
3d�Hg{��|(�5��;��m������o�(I��%����滻:��ךL8*�$:��$�B�����p�LD8b��!5;�(�qlp-���b _k ѹeÇ��)�#-0	x�!�C��O���=���~8�h��+w���'��T��:��j]�����Ը#�j�. �\��>��@����]���a�sݻQ)����G�x�tI����D+,+ �%�Valb
O?��T/�\�GG�1,���;Qڭ �9}JnG��&��'��	V{NP����	ѱ2���쏐!��TZ*�Ϗ�?�X$.3��!�ϥ�re>����u�������xj�3`���9�`nʼ�l���r�B�����	'm@*�X�
H
�d"��E%�-�9������j�1@s�kI$���SP�ެ^�Ft���Fd�������!���vczr
�d�x�d��rM��<~�
��%)Ef�nO�?�TfB.R�T�8
H6w�X�w�]������12���r,��*B�|?njܸ�����	��*v�8��%��u��!�w�wp��pډ+���¢w2<n4 S�q�ů���,�۶�_���W�v�8��ۂ����ꦅk��Z�|�R��xj�s�L���Q����H�0�����c+gr�����]r�x������ox?��"�;������?���LMga�ыbXs�MXd���Ɨ�RU�*���̙Wޟ�    IDATI���V�^/�;v�:��`���GdԺ�D0wB0'�:?�Z�y�%�΅#��0Dp(Mn�߃@�D0��h����7�Mox^�}߹�7��PNbH��hy�k�<����)��&��mv<?y�79'G�C���I��������Ww@�kI�0��L��f`��c>3O0�!��E�	5�H(�w�0h���ͤQ��dȃu�1��4n���X�Mt�ՃO 1@ο��O<�g�ۃ\��5'LB�d����eA�̔L~?���rL�I���EP�U�g%oz|�>9�\�>_�!hX�j��q����
�"����kv	a���� �/�Ɵ����L�'��{�mE{,�V��Gd���s�Q;�KY �:�K�� ���T�'�}�yz���#����9
����X;�4梔�7 _��2�1��������yos��|�{����;?�/bQ�܀�fK@7}	�"^I"I�@1�A(��]+K�K�\-q��)]��%�� W���ē�!h)H|dd�!��V�?t�}�Q=&A�Vk W� � %Q��!M������I��O/TW@wU鲐�3@`�K���y$ے�PN�̱����i��v�i�Z�#3K�qK>��5#�e��p������ؼ������022�H�=D�+�j�]�Z�	�ƙ-��RJ˶��I�Lg#��s����<��c���jF�BGI��Z�����>tkKB��S���۰a�����#	ه0<� �mg�;kA�R�'B�<hE�
D%+(cDf��*�+�[*yQ-t�NM�ȅ�T)D��ή.i-�0E M�kJ�Aw��޹h(p��Qº�\y٫�����M�`Ws�=:�	[�<"� �|�>t-_��T�w�ǋ��7|
�>�4��v ���hA��(�	�7�"[,�2))�d�U˃6�&l�b�BJ��j�L���i'��b!�����}�d�zJ��_��#�}�h/ҳ���M�@&������dNU�^�r*Tu�й1/��ͱ���pyE��7]��sW�rO����p�Q-B���3��乤3���'Ǖ�5�ֶ��ǐl����\'������%�&��I����ה��U�7G(�9)����	׹�����&L|�lhޔA�[���6#I��S�kֺ{:@��ȍa@%І
�E�AJYu�ꉣ^��5�z'.��\:t��D��}��>�D�N�UP�� s]^>�4��%�f8������,�јU#�#��^Ip��r�Y,�**��`��V_�B�dH_!�������Q|�k�c������H��%�BHea�J�@�;
��'����A�8��՞���L��Դ�A�5��N�����n��{ѳr-�&a��̀�slo�#��Y����{���S�?�/=�B'q25�annjE�\m-!9�(��Ge|����\
��Y�g�q���X�ƢqQ �8����ȋr�wpp�/(A�cټ!2֠�\�@����>?�v�g�����LV5i����g3R͋��L*-�4��9rza��(������)��L��e�nblR���c�d�e&i���`\S�f��y�eRf�I�ы9��/=�p$.����k��/�0Ûe6)�����\#��0RXE*�xK�-	ޱ�QlذQ��d��ߧƩ�Xp�T��6q*"���^���f���Ju���K64B���`zT%�����0̙<4�JDkIq�)8�@F��E�=�<8>5��lZF`$�	;�14i�W4D�)����u��,�����q`�n����� Z��)cljR����Ä�
Ἃ_��v���,7�vJ�k�
��R�J�L���}�S~��&���4�� ��<��%k$���6!���9l8q5�;�L:| /�܋ٙ<F�gQ)Ta�/�h��P4$��6��?�`eN$T��9��c7�.��<�P�w���)�.I�4��������E����ދ�,o�O$5��I����� �B��D<��A���1_ .SLf)H�$O�|���=u�M?���zLO!^���x���"9/�[�eO�mT�t�	\O�f^�TZ�e�T����~˹��\�.e�㛣r�>�ڿt@7��	�2Ӝ6�Q-�Df�S+�3��dK'���m͍��;���T^\}>N(G�HD��ن�d?qHn�A
�}p�B~�r_,�
��uU����S&����⚯TD��h�gg�a�R��?�+��>�#/�Fjb��2Q���:�|&�B��T��c��tK�lb���صc�� Z�*g6���[��w�2�+6���!_3p����s/��hg<�4$��F?�W�����W���q��~�eۧ�eoo�JI�"���TI�����X"(Z̦��q���ى�Z�&ջ�c����x�8Y���v�UrQ�m��-��eQȗ�5�8�W��ȕ��<Ǥ3���e�fq���`�I�R�.p.y6�S�5^�Y�����i��G.3+=��+�"1N�qt�"ҷ�T�V��^�C�7lP�}�:���SA�Z���K���]j���$!N@'dO��V��j�=��K%���^]��T��GG���'�~�أJ�i
c�5���/��z��V��9�[�eM�_z�$J4�k4��*�vz��+��h~̺��̝3�c��͖�Ix�U ��}}D���@z&�$���r��dBP ��2b�:�4�3�����V�$Ԅ�{0��B��92w��<��,3�
f
6��<��oācS0�	8��9����7d��y����Sz��,��j�u�u(~�(RE���6������E��HX���3�g����]��AWDP��2�+�����Н��#��e �I�[��%�8�s�?���!f�y��0�]͐q(��E��yt����d18>"R����Ƒ�hW�Ω��S�B7[9�J9���i��$���m'X�xeO���&T0WI��B<J�mQv���_/ii���
�;}Mej߹n��8}�Φ8��/}��ʅ���x��0G%ޕ�,�v�:�����}v2E��,|�#�p��?�t��I�0E2a;	��(��m�h�d�L�E&�X�/�B"_,����P���x""W)�T(
��p*t����C{��nF[��o��elX��~���?r��=29�}�~d,`ۏו{��
P\���i�[J;r�����)yC9Gd��!f ɎE8pd�@�\��>tE��`k7j>�h�c#�l4�ߺ�?t�O�jfo���{��ɩQ	"��m��$مf$K�@�11z�3X��C~�_�l	�y5?�M>���$�pL qn��r�GhE�����T�čN������s��Rي��^x���HFu�4h����-K�� �1�"� ���'���jE�eh���]X*��\��qA��-�Ϥ�
X�uo�1%!�i���P��ˬ7f�Z����ב<&jS���l!:ϝ��c��v��J�=6>���qtuvKR%�q����a,_�5V�P.u����Z;�05�������M���%��$�\��u�Vw#�/����|YF�m�_���i2�"�B�orrZ�Bx������ڱ^���吷�*�ItƣHZ!�*a$A��F"���=(�3>"&\�ӂ���ImI4�����;N��/����	7)�Kn���z�BbU�M��k4����<ޡ�AĒ�6b���O67+h	7.�6�7������ϙt
�dR�@��3*�mڐjU~'b���:���ϵ7������&�����47�/��_
	S_���H�3����Z�G��O���t���C���>?�+�DK�RA�1�J�^%�T�ˉ�3g�|o�9��T��m�$��n����
�e	�*���,������q�c��s];w����ڪQqFh������A������-eaԲ�\WQ����Վ��Cb&n�FKK��~�mC
"U�5�@zKDQ,�P��aӳC�^qB$�_��׃�~ZW�Ж�\!S,O?��sa�G���nr]��C&J�4L;�O�����w��O��]�f�H&b��Az�ƍ��?,�c��>l߾]� �F�+�9������wxh�Q!`��Ղ:r$.�V�b;������-m&�0S���/E��Q�J#��ۧ�����W���Ѱ�㞷�~��ϔj��:z������S�J���C%[C�h���G\��86|H��HVI#V%���%�z�G6C����EX�yqC��*o��J����1�[�M���*iGw��	q���p��^��SLa&&�eSi�h�M���X(����abdѠ%���(��s�AB�R��kq`R���A��,x��A�%���D��F>aVf��.�##ajTO���[e�����E@�^L!�-%+�k)b5e����q��u�g���^��.ے,7�6%�z�	!��!BM�	�!$�f&!bB7� �c0n�n��w�������Ȳ�03y뽵�e[��{���Ww�6{C]�
�$o�����O��t<�jj��&`�kUު�v�$��uF��jA0�/� C4�If�0���fG*Wc�^�1,&Ȋ��~���''��C����`������.��`�XU)f��sb���� �D��fˌFʓ�����iE����ذ$Xj���D��No#ƣ�M��[�D��$�	���og2I.�	��lJ���v�	����� �ѐ�q�+&x�u4�B(¯Ջ�5���x\.DCqXE�7�E���qJD�-�cX�f�%tu�w�U�V	}�D[M���yXK�=K���]���'M�gz����5`W'�
�١ڛ�h�F�b\pD�1*����"��l����t�@/j��
���N����@5����w��Y���Y,�+|��m���2�����	�����&����bf�n���'���ּQ�_�jq$�fU����5��i�t�E��.]$�qK�J��!	8��Kd�)�lu�鮁�߄tJ��]W�I�	��&���N��N�X*�x��$O{�Βz�G.���5D�N4��@ۜ�`�V�bI��lF��,�=�*(��F:>���,�h���o�o�#��`3��b�<���Dz���^·��m\z�%ذa�`+(z����?5~g��,����ِUD ����._�~��E<�3���^����x4��:�#���sԢdR	��j�΄��]?����)gܕS�	��Ptr�j1�I�7����=�j�a��>&�[/��l���	<���i
�SU>^v$�Oe�.|TQW��`J�Y!�w�LV�<t�xT�T{ ��D�ϫ !A�R�ۥВ� ���Ĥ��B�	�d�b_>�l�q��Xrߟ�c�z�(�&pY-Ĩ	ԋj���!dE̝7�rE�јз8N��^a�D���v���ѐ$B�����a����R9�@J���S�֤h{��I�z����j�d�}��K�����-v%=j��h�s�<)�x/�s���IT�����KY��ě���U���>��7
�O��r9�S	�
4�H�Do0!�L#g�huJ!AQ�h�8���T�>.k�"waf�n7��� 爻i�3���X�`�>�T���attFC]�����:�--�ƭ[�,bf[;�7ry&�)4��Ŏ��{���F����X!�ՎR�;B�l�cxpD�Q�:,hC(8�pd��yl۶;w�cb2�4��u��SU�׏�6������\��Τ� <��;;��L�&0�۫��d�]|*4h�H�b+�	]KBZq;5�-I��R�+�"y�(^��t�G&:pQ���K=�"��������g9�N�q�L�C愄�,�`�Ӡ�����<�JJ4��:"�$5ʜ�����)��t��H�:������<>U%�sz�g�B�'�%���������>�H���u����I�ڸzB�*��&j�D�t��ʏ��d*�t&����"��m���A*�G�@�e����g�On{!�@ht5.�N��q�nG�,�TR��e�P��,O�p�y�V'J&�Pkm��&�T>W  ��x"�Tt�\��=�������:�ɴ�6\x�IB���q�W�<�ڵk�x�}�����n�.'�JP�XJ����ܝz꩒���~w�m��O��7/\x��`�8�h휏-�=�xH�m��)��<��J�J��û���Ɗ7���E�Kr��`K�+�(&ݒ	�H�Z��u+��tiY�l�4`�!O�Q�͙����P��|E��Y�M
�Q�U�7��!MH�/¢��@-�C)�ꞯQ�Wr��Zr��q�]=8bP�����/����D"��'�o|��HF&���\
ۻ6�m֣�jC&�D,�����S��т��Qĳ9,>�3�����;{P2X`"e����DN����\�c�s��?�1�{z�Zݺ�K����s�kCmm���=c��Vh�p0"	�� ����W_-��e˖axpP�y���L@:;;�����)������=�%�M���yW^�2"�T�}NV�Y���vH!��>[
���~�j���ٕW�opKz3fcێ�vٛsZ2>>*�����.r��pD@f� N8�hR)l\��Z$�1C��FیF��˟af����w;��"J�8vnZ��'��}^���u�\��%<��K���g}ɔo�؈��{00�+P�]�X,��"���L��2j��M�`5۰�^s`��c�:\v��q�g����v��x��Q��@�b%,��q3�2��4fI�XQFE��0���E�1y�����{M���$*�:܅��r�V�B�������.m�>]�mW�����`Ю��V�Yv�6|�*~
9��I�	�L&?�R�6�?B�!�"�)���a���	j��M,�t��.4�
�|��A���(�MFB���"����/-�X�.�2l�������{`v��G�������&	�� PqOh������ǰ��a��kO��.@��pJ�	���h�r�yuX��'�`����ņ��1<�SVT�d
���
�x_;��.�.l���+�A���s��Jő��+����\>	��麫����k�.�+/<��͛E�9G݁R�￟ġ'�z>���n�E�x�g��s��3B�;e�)� �r�~��_�������}A�m[�a����˯��g�C��yp0#Q�A��V�mYs}���;<�Un)�\m�xȗa1m^�dhL���*���պ��`#A�����n��N9��J�`U�D��hi^h/�F�b1ZQ��p��RmV���a��Z�$�D�v93Qю_ϛ͛�џ�(��銦v����I���:m˾䎓����F��8.������n�rtoew^���~�y�4�̨��#�/b,�̹���>��(�t��E�A�d����|�p��|��a� ���M�p����G:�U+Wb���dk�iFm�N����ME�YF�4��PO�$��T� 3D���_�!����^D�Ay�۷v��$茒��Z��	'� Ҥ윹���¶���E#q̝;_<�<t�^���ÃK��'u��並�c���ґ�!ݸy�Ο/ԯ��a�6w �,���E�*�͊;_;tj3��A��!I���G9�F���8��c��$�\���fQ.\�p>����S9C����/F:<�������劼O�Ǉ�?��ߵ�֮G,��W��M�
f<��[X���݂�� w�E�q�˳l4�P*r��Z�w�f. ���;~�DBa6lچ����"��9�1W9�z���N_�z��D���%J�*��hIѕL&Il��%�\(}42�q��mO����t���s�>=�(ʴD�������jW�# -���b�
���%���)����*����z�YVl\�qm��Q��=i�f��Y��(Z*���nJ��?Y˴D^�5����������AL�h��)�A$���(���_���ׄ��I�&���t�:��R�T��U�?�h��*Q.�}�G�-(&�B2d�ػ�	�w���w�����02    IDAT��7ȹ��<�\}n֯߄Ɩp��X�y ϼ�%�:j���0���S0:\�)/��c���K1oF ��<�֯�sO>-t�D$*q���E�s�w.�X~&�]��<�tiU|F�2�~���%2y��������_v�E��ٍ���8��sp�a���jP7c&ƣI���k�CW�
���.�����3�xo�o�p�'�Y#�>�PdR:CA'�|�]�=<h��	��w1�k�L�D��n��7�I��ո]��B�}�lNLU(/�.'��f2u�9��Eu⒀MV�N֒� ū�~14(��_�І�^��X"�~�^/��JqL�5�� �;������זaǖupS�xr��:�^�sYd���z��g�9�7lD�d����M�57�+_��5	!ɀXkJ+��V��u���o�+�3^x���G���+�s�E:gϕ}"������{�v�J,�7_:kʮ��b���������'������n��H���7+���`o,Y�~=/^�/����2`�B�b��wW`��nI�g�q�{�4G���6`t�_(�D���b$����M�VV�˗/��>�E��q�����`g��E �+ad�2�̘5S%�� �L����;�B�C���#��ـ˷aɒ�����ŕ���[�6�XIc�� �vlF��`��`�_��,z��~��������q\��kQ�Xq�/�ƫo�G��C,_BKG�"��Q��O�N����-�I٫`FK3z�s8�����N�����CCaĒ��1��T�>�.����x�*yA�<R�!%��_���9�Ó���)�I����P��^0$SNj]�]:U�R�Y-�wO�'�=��t��+�p7^L'a��"���"畆!,��<�F5m�z�y9�L"O˞�S z۳�b1C��ádS��M¥�~�{1y�&��I�D�E����(��͜�q�D�Eu?49�{���y���X�.+�O��f:�M�������z�{��ZR���b�L��.0%��`n�EueQh�%�@&�}�᢯����`nG�(J�@'G>�b	�k�N|�~'���p�w����~XZf��)Q1��6]%�{�:-.�Dl�˞}���m� �>��_�Z8\vwwW�mF1��D�ȹ��#�q���<�m�q�q��\���N�׋��?N�gG�l4���K/�h(�dA�}���4��B��w��8���u�����𙯮����hV�?�@x�xH�4�h���XFCV3`c5���n3KW����	V�N(�!;Z��M=l���5�!<j����"�_����L&��~ٷ���n��P�4� 0�v��qGL�2�0`���?3p�c��ˋ�kE,�����S	��69�O�����7]��^y��8~'�}�u���d5#ϑ�ɆX���9�1�����`"�ı'������w(T������HR�I�#;�L��������D(8�|:��^}EW�z��с��N�&,XD��h���k?��t����h���[n����<p?6oވ��m�45�k�����El\�3���!y����_�o���̝'כ{�D2�W_}#����K��#��x����\(�S�u̞��.�הּ�(FF����
W���>��9���%�7�㵷Wc0C� �L�dM��V��.ǘ�4s2a5arx7���1on-6`�q���_�s�L�p���Nd�a�j*i��<l}��*�AĨ��_����a�Î���ql�ُ�����_:Mm���G�ʛ�l����-�0<1�	��ѩ-L��a(�i�	����k�sO�(aDc)����z5NI����t��R"�IR��A[���VC�H��c6KG�&"�P�1��k&$�TqǮ�Ego��	}*iL%��9OO��%O���4��v#
!��^�kYuy�h�1C��T6�'3�.�u	v1�	���$3��Ci������,��L|�nS���M�qK4M��4QG�W!��k���)k��oχ|IM\��+A�_M��iӓ���=)�mH�j�R�i�����!&V4���ԋB5�N�d��(N9������0���bݚ�2-�8���E����͗�ѹ/V�݆m�A��ڇ�Ӈ<�7����ĥ\���GN��$�C���G�ϊ�����yo���RdK�|�f�[,"�E�&',,�?��_�LT�:�����5���rME�.��흈Dc��3�W�9�,D�T�d<����Ӊr���u�<v��+�ݖ�8;�<�Z�I� ����ND��+fQ+*��ړ��lD]��:9qۡ���	�<v�Sv�D s �L�f�d0'
������s�N䫗�:������5��@&����H���:1-�$�B��A^k�,t)�O�{rb���Ϥ�5�{�p�4��丘	��Q�/����-X�v#y�Y��E{s,^�LvĲ9��D���x�&�p�`���%�x�Wa0ڐH34bd,�@��8*�4�j\��O�E]���X��=DCA���xƌYR�8���N�l���\̯��`wz�����ߵ}~�Q�ܹ/���^�W]y%?�p˱���c��k�n���6l����ǎ�^C1��OH}�w.��9}�#شn=��f�����Z�l�(\Nv�6�Y�^{uV�Z�c�;u-�����a�����k�`��~�j�14���:s��j�Bj�/��TD>����m8��������O"G,:��.�6?�3X��-��AG{3
� �֮�!�:�0S��T��'��X��[��;{�/}���c	����1{���X��S�+8�+����ēK�E�*T��#�=/t��G#m	��� B�k:CJ��^Ą��ұȥ���82W�:��j9�v�b�j����^���U��$p"�iФw�{�R�S 6�O.@PMȤ������N%���	G���� �=!���\>#����5�>H����(���������j�ȸ�bG"�T-�Gz&��G��Q}1��R������2�$r�t4�!����@2I���h�����q���o&�=h�(1W߇6Q�5vP�p���7���"�!;r��8%\������k6i�D�T�vn��B��9��	����A�GI�,V#^z��z�as5�?<��=�2ʵ�(r�Z(
x�D�P�̸
a�u��F�������X��K����BB�夔�<�7@�)�mpG�u)�2ݨd)I�l!b�
y��۠���&͍`�
\�E��ގ9�J�P4۠�٥C�yIU��7K��i��%���b�o���x,�J���"������>��R	�P�P�s�+_>5^;m9�Z�[6����&Ó2f�q/���N%���ǨF��3g��DX�i;���F��K�U���MVZ�M��+��\NF�<��͗�*��/`}E���0��߲Ï'��H���>�\y�Eذ~-vtm��b���?�Es;ᰑڥ��Ct7*�e�|̱�b��yX�r���cpy(�͘�[lS�~'=׷�1P�k�):`r�V���c#���⅋0o�\E'�N:���c�v9�s�t��"б����sG��^Z����W_[�ǅY3g��o_��;n�K�s�Ʉ��V`|tw�u���B�d�:��������d�q�%���߾ �7mG_�N�������ܯ�ԄF.�xL�$�L������<��
:l�:�s���k�*���vK�|8#����$t�g��5��̀��wO�M&��~W]v	<^[��xn�:��o[t�^{�M1����g�����U��߿�W����0
�Y���Y���]zD�P�6m
�w�݅��Q�:��.�2Y�d��^�����<��ƙ�WAm����^�1��)(�p6�Q�ߚ�V�"��.'T��Yf�F<�8x���D���s�	��h���3���J����m_��~�nÇF��q�|�i��u�;l�{�2� Z�A�gT���q�����/�E��Lz��� L��!�4��"
>�v�t�2RW6"�[B���S�_CلB&�l2���z�~���w�^x衇�a�v�RF�L��5A�qs��~a��T��������^���j�bkZB�)�l�	�+K/���I:d�a$�#8꠽�n�ho
� ^�P��
(���Q45�a<Ļ+7`�^b$X���=C]Jz#�Œ�Z���X��(���0!>9G%�cZ�_��j���?㡿-A=Ņ�a���rE���.|;l8���8^��кsyo�����W�t�~�Ͱ b~������@�PB^gB�lF,W���Ҹ�� ͧ����O���������PL�P�gP.�Q1���*�\�����m�!�
��·믿V�r���c�T"-7��d�6��169&;V�����ŋ/;lqp�!P߀��L�bx��G�j�&�N�@�O�BF�G�ɧ$��ޥ�dLμ��S�y���J%u����D��R��ay�L�v;]�x(-��L���_,	k�uh���`_?��[DI,��at,(��s��x��;%��Uk�kB�hG(����E�Aҏ�����|�\���xz�cx�����A��Yhmn����Z7��`P�o�K=��3`w�����cǎp��.�o���@&'Feձ��(�e�|�]?ȱ�+I���>_ .��Lo.G~ց��_��&8lV���)�s�� :fw�}v�$�`(��~�u��{G^��sro?�hl�9��X��o���,#Jq6�u��b�	GCQ���/WP���� j<^���L�P��F]��h��p<��!&B#شy-"��t���<^_�26lZ/*tF���q6�8��شa����|s�ar��hm���(���q+\n3����u;�_���������}��Z_��HN���X�PC���)1�a�Z2*���IXbFĂ�^x=��016.��?:
��j0$kE�`��y��g�KM��_�2'���J`�CW&��� 8�7���U w4�o�׵Ⱦ�@J��<EOH���h����Z�.������,WE�ST�#�c�沲�^�^�vK�ӵЙ�(����w�J>�����|�d4Գ�n��OX�j̶a�Ʋ� �ŀ\�s�=����?}ǭ�jԇ֙k���:�):b��ѷ��v{�=���t�ܔ�f�}r����M@	Yt�&�A�L,S%���Z��߀�D��=�P(�y���%�9��`F�,�^�	�Wm��D}I$�6��(w��C���f1-Z�6�ؑ�.�����S���'��c6}�m,��΢h�Z,�Y0hU~�Sb:Or�J
ig�{.X�8�I�1o�<446cݦ���H��0��H����oAIg6	�[�ʴ�pl��}��y�7Vn��gg<���B iv�q��*[G@_,:�=4����~۶��ͤ�X�$�Lxደو"�dk8�����Ft2$	��/Ip�M�����m�d>>��'�,b� �

�Zf����.7��^�����&���Ƃ�����$�qLg2 �
���Mv���Љ�l��i������ ��BƠm�[dDĠ�qy�3e�/�i�l�C���C26��D�.[��8m��I��T"���f4��_>g�z�oلg�Y�\�\��۪Կ�tx�y��e�h�hᖷ�~G����A:��~�+X�vV,[t��I����|l�fϞ-v�,�Y看+V��w�Pm�X���j�T��^��|�$�G��c�!�"/��ڀ��X uo�9�^��٣�A��yx��wM���c`�����煶�:S�Ո���FqX̂%�x��2h��h4�����Մ���\o/9ͦ
��	��,�7�;�cdl��M0K�M!��JGI�fN�j�Q�4C@Yc�a}�����E_��K���xF�]��啨�f䮐�I�)s�bI'��g��Uep��}��"�kz�=Ȗ��e��3q{��s0��\2P��3K ��g�ə�<V�dom���/G��<��t�S��*Aj#tM����[�S S%̟W,䠓�75蝢!ο+抂�)pM�"��%���+����-ʺ�#xN й������ԮoC�f�.E��ҩEA�=r�,ЗL(3���8��q��G����n�q	�_�݈$s��Й�Y���>�3*�Х ���5�=#��8����?I蒬����U��V�U�yvK�:!RJ�ى�;��_��m��b�#0sF;��G��g����+Q�87����?B��F������8f/������ۆtt3�݈��a�k3�8�X��ؼ���*�x�Q��0f	X�H:�Nb,φL��#eS|�Ͳ�*��(����3]�`�I��:Dֻ��#��z�jj1:��[g�U�6������%��ݹ�w��-_qu�n#h����K�y��ႾP��ͨ��fľ;�+/��O,A.��L:�o��L�"<���>Dbaٕ�k|r�M|u���M��Z�#KaѾ��e˱�Օ�kn��p��\^��?���X|@�1���=^{}9�M�d� �� ��Ռ�V�>�)J!V$�Л]����E܄��F-vlL�W�֑�V���3 ��U��9bd�g ��T� ����Њ���p@�o1f�jE�ߋ���`tdH��\)pr@}{���Zɭnnn�#��I�*(qRT����E
���@��a�&%TA�r��������Y8�k�\O�"��	v�abf��`|d۶mC,����١V	
L�p �;�Dtm�A���uuc�pA1�H144:$���&t/r�2z{�D����&��Y��)x��I%c�;�3m1���p؅IA�v�� ���o^��hE
^h2�Lvl�B�����4!�L��?�X��l1�`Goo/���_�\�35Z��5���Z��''¨�oT�EUqڣҗ��1))�s��P��,yk|�t%�Xpdn�O����HM���il1��`�;Q[G������gd�+�`{8���:��万+���?*���� ���hxS�����{�3 ��B헲RZ��N=�����D�[|���b)��H�(��F��P���1�؀�*�t|�ɷ&(�b��e����s�Y��Z��^}�HvO�񤨠��.���]����R���0���3~��۞I[��4�%�)-��ޕ��Ǉ� ��i/^ۡ��T�~�װ��M�t�$(�d���� ���]�m���i�y��li��Ą4_l|��9���2���V��B(����E�&+����F�� ˩M8AC���A���ފ#�g�y
2�0b���N9�|���L0>��"Q�,dWUA�J�@��7��j3&�'���sKq"Ơ�s��Ֆ�]��<'��{<��G�`��]�Ѧ��6�/ؕw.9�zo��ܝ�D�b��xB�Ռ�� L:J鬸����K�����_;cC;���P��d�)�.���#�I�󒄘0��g�㎑��b���_�!��y����BEg��w�㍷֡e�|ēe���Y��:�����3�O�>���w؝^X�iW�f���c�I|����<�st~cr��E���&�$	���A(GT�����OFK%&B�h��'�H��jR��e
�Z1��,G��f������L"
��}%�\"�x"�@�_I�r�Ja�B�A����6���8�f����$�I	�U�qA����D�3��p���/]��J�, �,��c�8:2���!474��� B&�ư}�qs�5g�pMFâ1O5�d���/Y��; ��W}#��L����0:2��
r��0�?�\��l:%��r)��<Fޣ��Ao(����X�K4�99�DS�b`h@����]��-��bN%NTD��b���Jaw{E`�� ���x�#ﴰ8�㾚'8�\T�h��J���"	��Z�`p�D^S�O:�i��?AmM���b�(���B�Ҟ����u�=�>�cId
Eq��p'BN���(�~�{hҭS��)�\u��q<�=�t�e �L��A���D&mA�Wg��    IDAT*S�^䕳cr�첂�'��a����pF��|�6�mQJ�y�Q��lV4@"��~�{b>���H�z�.����/�L���H��G@�é⊊rˏ�&D�W5�~������ZO����L�5}�D����Um_-�k�4�����������i��3����\N�瞌�W㥧a�%ׂ��<��?��:a��]����	����T:�I%j�a�9$��p�\΢�n������ࢯ~�x~)6� (@׿_��Hqf�A���x�	���<_u��ڦY��Y�$W�!���+",�N�]��c�cR-[�H�D�9-`��:�O(���:���L�9L�t�BF�h>�2�(f���� *r��y�b|�K���4 ��LN�UT�\�x��E���G}$����Յb�:jke\�Gѵm'�� �}o#^z�=�ۑ+�`q��;�q∣��瞃��w�޿< �lR^�����f�T��sy��V%��8�ȡ%��c$��M�e�I�+�5����@܅2��fU4p$<]�v�AU#Jm��1#wE�)���|�>7b��b S�$d�Y��)�AF�C&�E2���b���t&�5�+;x{�.�=�`kX\E����k@�v��<5`"�/d&c�:�.slL%�Y�3h���[#��`�L0�[�Q�Ҁd.���q��8��d
��\0Z]p��spTvY����624�r�  ;j��˝Eܜk���8���Bu�@I����;�� _7A��X�s;E�:����ͥ��o��0��T�Yo��bs�m�\�#�����d��zNm�JJ�òw�)�R���0L67��d9��������=�-��%<��@g=(my��2`���8K%��$��$���$8��
M�`���,��p8��'��+钨�v�*�j�����Z��aMv!,~�%{���p�^��+��(���	�ȸf��b�R�fa���DV;,.|6�Ԡt/qL$\�I� ���^ N��]N�x-��s���yY���!�V�,���mvd��O��-pɬ1QhE���غ*m���D�����1���?)�O�>{v�R~�`��i:{�A�?k�lb�Ǖ��i�-4��!����^@qT&�303�t�}�QHN`ś/��JL�=cb彌����X��`dRL��m�����ZB'��C#l��YavY16:�|$��.8�>^y�qtm� v�Q$��t&��Juu��4=�L��T�T�[����ؽ���)8:�D��sJ!���ONIˤs�M��4 k2a���Z�,>I�<K�΄~��'���w[�y��3	��^��$�o��F���0�&��3���%] })�\&$#z���wA*j�����I�s�l46�
���XI� 1p�yh�t�!t�ƪ5��� �*(.C�6���|?e>��9n�Moh�-qI�Ug(њ�,%9�}ŋ�0�3�U(�A�H2!��/8
��I���`N��諻�]cu�U}��D29�e��ʝ���t�9ᆢ�q�oHP�NI��Ɋ�"~�\N)��h�]�ۺ\����	�H`�q�L��z0��-D��+x��8^�.]�&����^��˼?���Y��f�k	�]���{g }���<�Ѥ 9�ә��zkQ6Y�%�Nj��8e^+%����j5�(��w�(:������,�������b�2�ޏr>#R�"�k2��N���x�n�$v�1����i���;L
�$3Y2]��om�&�����n��v2�������@-L�2ҙ�P'�[10<!�?��<LV��`��L��̥{���3gc�ʄ.v��X'��
�#c��]��+���:;���o����~<����B��G,�Fm���Ϗ�@Q5Ak	]�x�J^{&��	}�.V�l%7e@%�2���Y2Ȳ8Sןg�*�y��9���IĒ(��0�lS4W�{�b1�.��u�C)���M�=�t���Ʊ �� X��:�EX�)�򥲈߰X���1	]K���.׹��������0ӯ���]B
?�uמ	]� ޝk9Ĥ�y���|*�r:�C��Y���X��0t�!��R�b��4F����0<G��N�
z�Lf�V0p�G��N�G4����:p_|#<������ނ��L���S��,��N��c��ٌp������f���vN�aF���*,�NJ�9�Ķ`�*�]�@{;6���h���i���X��L�W��c'����w��sA<�ri��dS��ɉ���I��%�an�`v[���
�^�&v>{t���<)޹s�K'<>:,8���B6��_��ރ��6ʘ�u˙d�^�eؑɑ�:��:="�iw�d ɑ U_ev�)��؉�ʂd� ܫ3@s$���.��#�M/��p.{>%Ԥ�ţr�Ű�f�q,G��"-[E��z������>�Bfұ����3�M��|2`Wc��u8X�b�	d�i���5�U�*yx����Qȴ������ɘ�c)Jn��A'�Kܫ�e�Z~�h0	p�#g��m��J77����*(k����f����-�Ŭ��T6���v���Q[�$�t��f��;k�ĳ�c[� |��(��"Tɕ	E�\&P_���f�`br��pZI�)�F�I������;_:�PQ]~w����8��f�2�X�hm6��)@$�eyd`0��j�֮��C�/Eӌ6Lv�z۝p9����&
�,��kq������f!��cU��\0ځ_������[�@}��FeLL�"C��C���6�'D,̨ ǂ����Mj��]'u���/`N�l�n���⮻����x�x��W���[\��[fBo� ���A%t՝Wy�Ue9R��Ѵ@�9�M���6Eg�
>��y� �JY��h.hF�ϯ�rŢ��f�BM�H�+��;�^D��ϥ���ұsbB���\���􎯔%1��aqM�z>��G.�ݫ�s�O�N�y�t�L�j�>m����tG������CM��	���t�s�w����lL����0q *����X��IP��E�k��$t�Q�Y���Yu��W�s�K92�Z��cx,.x4��9�~ۺGP4�`�yQ&��nS�-ņ��k�B_@,����.][W�����������N��'��{�b`�̰��G.��ZQ�ܰxg�gQ�F���z��-�v�-F���L�`���h_�;FG�5�`q7ݘ	��m����������ާ?���۳E���h
�|�b��L����i���LKT�̊i����uW��7��� �e
a$�Pp�{�ٟá�*^�8�N$�X��;x���W��(U���t��� ��	��6l����q�PHu�3TU�h�����0���"�׭%2�X��"�Ȥ,���$����S0��� 7)���1��+Nj��a7+�Ʈ}��NVt�<Kg���i� ���<��8\NL�n��O�Z0ػ�D�-��|�hX�/>��r�S� D/�;"��S����edk�I@䳌�}-�ǂҗ�%J&D!����)^?�����ɵ�׊5)���˗˲Z�D�3!P� ��@}+�n+�_������� 2�������~(Ah��5�*�&�ʆR� ��#b3v;=p�U�s��G�zf4����Ҥ���VA�o��%����W�Kss#��$���t����Ҍ�_�u��a�6�� \|�0�\�GSbS�e�E}�[�ag�L|��+0wA��1<���y갽g������L��^�` ��#�	%�A��|�{��RW#o�k�E��<mټw�y�(8�q�(���!lܰ&�o���7�?SJ�8g�ڛOS1�5j���ϒ:;x�q>��Ő� C�D&_�.�K�t�'Y%��Eɚ�P@M}������n�V�*�q���r9�f��b��?�4��|i٪q�EE��>�v��<�W4b�"$�`O4Z��u�ڸ}�E�n����4��Y4MO���J���xr2l�U���
��؝���ت�����C%�@G�����5{���0���9�~�n��q�	��������N���N����uJ;�XB*�/~r���V���>��6��q Nɺ���:�T2�R|6�A
1�!9׊L�l���Ȏ�.�<_u��|��KVL�3�a֙ $a�um�Jđ�a�׊��Oe����9j���3%��H4]>�J��ۀ��~�Y�rx�N��j|�3[����p�M?���vXL4bQ
@��	�:�c��1[�7����a�-"<2>!���01����؊��q��~�ֵcl2*".�t��)�YjQ���Œg����FB���*77�������"<�fD�I�$����N���I�AD.�̄�+�$��W��2D��73p��LL�90Hǐ���������+/��o,��@?X��3g��g'���PP���`�48<9�E��u"G޼�"��HH��9�͒е���F��V2��~)�g�r��9�� ����c����Y��*�Ι�QL=��al�ԅ�@lv/�Zg��/���p
7���X��JDbY��[�޶H
���V�b3��օ��I�#zdR:�)�X��f) ��-��#C[������|K��&,F�/�'��o����V�y��r}.��$1ܢ��ՎP8&r�?ش�rF�#��1Œ�IP��f۶n�}�y�����|��ˑ����a��~X}�`r$���]�D:�KO����S� �GdO� %]G�� �Up�O��0ib�"��g/��7n�>��S�Coo7V�\�H")y,Z�(EAZ�j	��Q����q�ũ�#��8>�aN�T�㲙 pʂ8�G1K���L�x~X<2�9�t�S &t���zp*�s�����H�y�+rF;U^'�����_�I�{6B��J&	^7U�VP(Wײ��2a>�h�6�u��d_-	�Ak���?�����v�h����U<��Sœɨ�g�F !^�f}��_?�4��y4�y���Bp:XPD��j��'�z&v���Wׂlɀ��.	�@�ci�,�YPw�Y\s�Ř�Z�M．���6��I�@@�g�y�<�;{����F�x�3���ʟyF���Mܱ�6�����x}�h��*��m;഻�� �.Էw`0CJg��Y�U%�Oe�~����jK��ْcQ4�G>��M�#��t�i��e �\r;�umĬ�������O>��"�]c������@D��-�B1�����q��6̙3Wn*�䂴���+`�R��<�Y��2��i����%`���O�d��4�7���e!XLF�3)y��6���R������;=u�ƒ�U�~��jv�}1��u��UvI���Y�������Z��D@;m��jdB.���#�Q���p�'�s�;����6���O@��*���6�� Mu���"�yEO2��*H	0_%&vYL�t���U{'a����@�쬢K�3�ޛ������秷tE���f,�g�T����ϧJ�`l���zT������w���>�W�kj����:O>�"n��n8�8�Г�n�&���˟�u�	��<��Q���Lcfk*�0"�>�q�MX��-�n]�{n�~�}��xǪ~����蜍��Q<���w�/n����dp��	��I�������de�_��o`��{�A��-@h2�D"���ň�[���\�SO:Bt�׮Z���0�fv^zk%�Z;1!U�&8�g�Tx/� �b��D4&����qNi�JWj�]�I�Q�0'��]?���Aq/dAK���hnaq��zjj�Ū�~�����E>���i{Ҳ>.�����y>�;�z�ʄZ
��xt�?3��������n���,������4��έ��� ���\rD�sɠ-�f�EV>l ��&���SbF���ȃ�]6�;I����"��=���$=�����{��(|��>�,����8y�{��}\B׾�(��J����&a��6S�O��R+dR���Ch����O>t/�6~�"���LD�O(���^g��8%[=(�0X=�[�Э�УL��[�t�`#3j���Ytx��G��cK�͆�uob4�Z�<�p���l_���v<��SrV�l�"TU2:�^Y�ʦ�Hz5~o�ц����ǋ/���_�97o���PA_~�%LDbH�9���t&�����Y~*��y�ȷ���C��XK�dW^�%�uZa0�0<8���DI�_���.�Ϫ�׾�9lٴRn��~i�����0b�8���:���"��!�ݽ�^(�K�,F��N&�1���:�^'hl鄞Jk�pf��3���O��t 	��턎��LB�P4`I�T�|	�p�nL6':�h8�5�闿pG��C44H b�#}B�54!��h�JB�����6H`��TBW�4������ �t����J��8�³K1��_9�<���+���=�O?t�$KypEfJ-q���E��ªY�^���~Iq:��?4�V�Jpe�P�z�QONx�UbW��Լg���ɉ��?K��UvX���Hu����8�ē�o}�.}���g,\x^}�-|���q��
�Tğ��nl�ЇD�X�,|b�!��?�p�f�؄;n��N����7�2�ǂ{K��ēK���{���/Gs�u��ٹ��m�3Ͽ":�:�>�'�v
���yޟ��&x<�@� (�r1������H�S��݁�@�n?|3���r�x�p�4K�nvxP��Ne$q�k���5%�4��LU�#5W32�6��V�	�@�\�/�ƌ(�F^�\��y��6��R�@�0ihv-�H"����3�|��8�?Es$U�ML,t�Ҧ�e�����^���4�'�1��#q8�>|o�ا$<|a�TTB�-+��gjpdX��Y �2I�j�2u�ב�X��8y�	c�\M�suT�;z_=h����}᧧����I	]���v���s�4u����V��o�5��&52Xi�`�\.g��<\6;"�}8�E�u�p�]���ε$-��2���J����䄪�%�0;��FP��j�<���@�\���h�n����އ��|	��.d2!)�Rq��[q��J�ͳ���\~�l�2�y��ַ�%y��F@|M<Cb'�+Kޠ�#	�J�g7� �򚕫q�q'�k_�*�����4e��RE�:�F�kʎ�S�C����{}���c�x"�b�;��p~Y�Q=�^���D��FFz�u[�٣@�E!K�CDE����B��K�Q4w�8�v�}n���)76~�B�4�y�}�Ѝ:?�z��b�f&+�
��N���mF
�!�r(��b�*b�|�e�����W�_M����1w��8~s��ᩩmnr�n��-����N�~�&�tWR��˓ƢF������J�F�g�����������ߌSO=�w�xϝx����s���	�4�A��9=���Ϫ��1_�*(y�yg�n}���-yk��g�8���[g�.��&ׅ��l�UEix�<P��)7%��(�v8�1{I�09��?u�%Qu�I��_lU�wΑ)̦�[p�a�ŵ?�O<�w�q�(L�y�8���)ُh��K����C�L��,ف_�|"c�X��K��o���p]���Ux��ELb��ƲW_GSS�����6�����SO>��{�y:��F,�1'�E]Jz\z��Q.�f���9�q�ϮǓK�.�7\�C��c��xo�:\��hn�^���6�(�P���Z��̈́ĝ(�9vVj��F�*�IQ��n'Ȍ�U,�W&���~se�,�	�#ȫ"#h�81)��pF�hf-�eu�9(���^B/��H�	]NՕ��c�
A�1)m��癣l0�?��9N
� ��t]�,�!�C� ��������T��يͮ�5'F�%���vUEs��d"%
qZ����a\3���%k�0���ch�S��������ߥ-L���IB�_N'H��?��l&�R&�sO:�N�[o�Q_�����å    IDATE�!�:q�cq���FY�\��;t�6t6�V�}�]K�:j�Gq�����T�s݇+�B���h����XT��O:�$��i��d��Y�F�N:�D\u�U�����$��ڑ`@}E���;Q�>�F���}��'Qxޜ����w���M�sd�^��P1�`����R���K�>���Ȕ]��b�Id�8@lhhX:�Y�R�������>����DRr�E�Ո�����a&����k�COO�\Lp;��cg�t���AMm��#��:%_K���]f�,�bF�dneG^��:)DM�*C�DR8����q���6
��]׀��I���W�3Y��2����A_�����!�H�Z@�0��P�\%�� ��	�=ұI�r����Y���%F�Ɖ�\�,}�Q�Y����Cǜ9رa����x�Υt�Ii�j;t	�DnV5���&V�� ��r�S�H�H��IC��N����xj "-�PV��f�(7�x���̙|_��0�� 
;��wl�{;k�,�D�Zq�q'�؟�txl�:�Ưn�߿�N���[�ij�gO<�}$�|�ؾ}۷�����s�+؂[n�)�c�X�拸��kp�g"�̡�{n��6������hl��nrȡ����d��V~��x��������[�\�����眍�}�͸�����.Ǜo-����G�;�y�I�Q���W��3�B��_z~z��ڶ ���hj��\و`���Bd�:T����.�g�tz�YM���2�2I U����7o�LC��g7NWA@�)E0����.�v�����KWY�ڜ���	���J����T��qI�
q�	�3�۳d����� ߙP4)٪��I���+@*?4l�[�9���"��k��)�L������\S&�J���.����9&�u��j7��)-��Zaz�eA]�%�g�矴�>��Ȥ�	�5�f�&d�S���d���&e�(@GfRظ"1�QIGpȢN��Y<p׭h�� S2���U���w���ъ|ńB�,�2:��r�b���gP*��K�J�a����~��31t�^�'�������Q�+
�N����׿�U��"��k�����=��*ϭ�=�7��dI�a:�tL!	�JH����4�1��:SC	���{�Er�eu�����~�Y6��{�����22�F������ܬ��A9?���nXmfQ�;x'�)���L�s�?O�}w/;�p\��+�#��c��h���ndu�B�����ʪ����/|�����`CӬh�6�7��N���[Z��0�$#�r�8lVβ�0h�7��8i8Ty���*��PT�U4xY��l��b�$x�])�ȤR�l^|��bX-2�C$��	ǉ&D!��0����<��iQ-*�A<���i��ĨZޢq���1�f ��z
�?�4|�٧bjKѽ�r�Zx�%rp�M��*��,@#U'[к��G�(��ο�Cw>�A�z�a�\�ol\�3g>��M�E}�#'C��c���ٰ%�E�_��p�2v�sԄ��PI ��a\�;VG�B*�(�1��$;G$z&�S�A��Q�k����>��H
�.g�	�I��T ����|�y�b����#���UOo ��n��>TՍ�U�܌��,^��n3`w�G:���`E:�ِB �3��7�@�͸隫0f�H��t�>����PR\�X<��Fc��8���p�W �˘�a�f����'�X�d9�:�(�����ɐ��<�?:/����s漈{�K�.����;�xS����F���g���PO>�2L�"�c(��F$�����T-o��$S����U�G��T`�Rt�T�8<⸖H(,���UZ��\j�o�XQ�h8�I
����Ĥ����?�3%M)@*��?K��"��|(@1u� �d5Ģ%� �q�7���MƌX'}�r��:�;�������ۥ�'���ӫ�֤�b�K�#�!�N��Wl�D+�7E�Ϸ�I9��|��L��=��B�	O������^Þ��i�zN����)�����.3�,2!?�N9� h����F��(�T��0��|'��bUc�#�?Z`� �C�%t:��I�arXм{���ʝ&t�؂'��Dz^���RQu
x�Z�a'��g�}&+Z^sq�:��riy��P ,l�M�7c@m��L�fN8�L�|��˵غ}'�5H?`6#�!ʽH:���Ȅ���˧,\�sV4��$�K&��G�[�@p�Ʉn�$�� ��r� ,�$&�����I�VXD"#��N��@�Q��0~�D��;vl��'OS�ݭ��x�Rh�&,Y�����"?����iA ��Y��!���I q�^�Xmz�N�������E,ɽ�ټY���R�,VDc	t��ňc��(��D$�$s�G��L.�<_V�)r@h�>z�F�+	=�l<������0a�`�|ݕ����0��)ؾmF��d<��[�e�a�����Ұ�ҕ�P�����pT��v��n�T�'L�](H���S��(�*�[D���2Q�*�tE������8����޳|o���XNA޿��k"�J	�5��b��7n�����[,_�o��)�}�m|��q �}a$���	��Z�_���1�{�q�"4n\�{�vJ�lذ�}� d+*���b̸Iظi�$�믿�"�vm������+�fC ��Q;����+4�4��v z�A�9J$���[q�C���O�Ηs�7jİ(�U"^y�{����P7�[��z�J��r
�@-�
UN	����~�(:����ʪ>FӒ���И����$�c�]9')"\�kC���ɹ(�[?>u���w��g����gO\�:�VJ&�"e�����O�!� �$����Y�}���Ʌ�l�B���F��� �)�, N�С̰`�!=K�C��T��eW̃$���F��F�IYW�]�HS\��"��=�p� �c�ZeU�`�ҡ���ۥ�-����,g$B?Sw�{k��	]���EH�S�г)D:Z�v��C�S�O�{�TX��X2��N���S�`$�`,#�����݋�ь����
�	dS9���,�Qd�1L��F<f(�{�yԯ]���7"�M��t�ue�PE���y}D�`��3��BU�Aq,�|�6�Q�=�J�΀Au��e����o�s�����L�,������p���5͌���$�ɔ��Ѡ���B�N:�ΐF>A"�M���1�0��=��| b�w�X�t��F���
�����.��d�"\z��X�a�p�?��+lݲKoB(�μ����Ѹ�\Æ���.��j�Q���fZ���N4���M�(xCs@k�Ac���I"����BiY�K+�����,:��@���f���X<��ZI�
��G�88x��=x���X���ؼv�P�����gQI����oi@<AuU��*��I�R�
Wv��9S�C�߰+�T��σ���	;��TA>V����A6��>���S�D&��g��>3�Q� ����C+݋���g)�_%�����`�֭xg�;�N��m��`���F���8d�t�	���{�1� �4"A�2�#���a��`3���Ҁ'gߏ��6`�%x扙H'���ӏ�g/Z�cF�CՀAp��������w߽���[�w���*7mڄ!����m���p��w���b�ɧ�S��~���[���X�v�M{��N���?;�p��pv�j�Z%q���+��}����R�)Œ��E
��}.e\�0���a��
���n�H��c��Qr���;�3�@��V@�����Jc}��_W�?a�p���	��)eG��5����γF�Z�2#igј$B�dQp���Z]Gլp�9%�c=��_�{<
O]��o�p�$5Aw
罐5��j<�� <j�¸�|��'��5����fB'�`ߏ�
��I�"��	�  z�;�Wex-�q�'#0�C@��U��̎�^y*��F�p�%1�\2�ēYDi?ju+6Б�/r:�$t���r)�<U(�R ��C}~|�]�-�������r�
dJ,�)c�8^7�d��8�N��
�f�޺Iku)�~2FS�4��%JF�{�"m��B7)�zL��������x�1�7�bB���b<����NLVP9�T~"W:�&	��4����;���rn��fQ�b�ew9q����7�X����f >��C�����S���ckK;&;��v~��+a�zE�4a̸��񆫠פ�f�2�o�"T���f,Z���9�gg@���n?���њUk��+Ge�@I�&x�Q�t�X\�\�*�*#&P���r)LC�c��:j��{��p�o~���<��G6���,476`�����DK�nt�u���L�3���F��
PJ�q_Ȁ�
���v��xJ9ǝ9�4y�#�5�	����,��LJ�ħ�(�6�[��@��5+Jcґp��D:3v�*mF��s2����˦��|��uX�~�HA^q�X�t���q�'aws>���ڰ	Ͽ�6n��ؼ���΢DS�7GE�\��ä�v�c��м}#�-��?|?�7c���X��{0N�p�Labɼ�ԙ4zx�����X�r��v	����/�&1�ǎ��Ukp܉��+����f��&M㪿\�����j&�1�X���VD8=%���c�,��V�����l"	���f���u%����"{t� ��FS���E����>�N� ���d�� G�ڔr�جFʪ�ؾF�}{�����6��بY�=
>��x� ��uJFвS#�[r�)-�:�;�OvT�P��XD�.�K�{�y�y����	'�v	���p�`A8�O-j�J�@OJ~����f�)S_2�=YV�+�:�wM��?ա﷽.�ׄ��ޝ������Q�iM!׵С~��
�B��8��I��ɤ�=m:ԋdO��0g�|��Mx��`�����b�XG�2���Hg�6Bq&w-lE��FU%��D��[\!�8��
�9�6ƜG��Ȧ��ߋ��fp-ǂ�Όja&�e���<?��$�k.�i�����E9��˄��B,ϸ1����Ԋ,U0�:����{�l����ew��>Xv�����������#a��.UZ[K�t����O�r��� ��9lvo_����g��DXA���ګbi:u�T{�qr`8Vf�6s�L�<�$�W��9ϋ]( �ގ�˷��O�d)C"����8q�!0s��% k�zP�裎�W����{�$ �Z&"��I�^F��Hv�%�e��5�l(0�>=gsZt��.h�302�$�CJ�t���8k���	�aw��F)�q�՗��q�q˵W��{n���r4�܆C9+W-���9|b�%�B��M.$ ��dʝ:�us/��ݬ҉3X��4�	L�7��;\�[c0��O�2��@��yc��( ݥWǉ�v� 2F����\�8po[P��V�!�� LF_͟�-[����캤��8����9sp����/�����ӹP\Q-V��|J��<�v�Q����(V/�M�kp�5Wb���Jw�K �jf��n����0d�0�x�����ь���r]�Hc��Ո��8�Wg��S�._7�����ow��/>�G���{�K��.���0Z�r���|A3="�q�sHSc��O(�j�A�UUם�qJ�j��塑��N���*؝N��pz�k�6�<e������uW�n�U�ɠ��E�k��]Y�y!�+I��8$CqN`�"e�&���>��?�EwA�+B.�'jW�T��� �,:e�K�Get�c &C$�S�+#v�\)�c)���>Y�R���g�W��` ���c�^�o�Ix쉸���M0�w:]��K���X��טۅ��Z� �j�V�S�?r���cO�W~�b�oBW���!��y�HB�_@��3N��'t+� �\��C��q����F��m�Y��M�d�D�E����A�����}:��VO)2Z �9JBϤr�(z^�E:�ˠ�.D6���;o�ı#q߽���ݎ�˗���V���~�1����x�T�'Ϻ��ld8����;�\#'��"�[��7E(����N���ɣ7Qx��_��}�G+�_���H�6�R8~q��0���ީ�4D�&��S+;�\�NCc������gp�K�Wv,��}W\�HCغu3Ǝ�%KK��z��(�����T���nx��X�h5�vwCk�����v�S�������x�6�Æp���O>�c�>*�h���!�	����/�]˫ �Bg��j/�&Z*~��(�@P��Q_5�JF���d �X�E��t��A"�A�d�(/=7s:���[X�x�x�A4l݈�&(T�U+���;L|,�b����@ C��$Pq�.t蹬�$� 92�z�����{E��T���#���U�Y��E%�[�׍�E>�χ���n�R�HԸWǯన1ed�uK^}�5����~'@�ꚁ�;������«��ˮB��8PT<@l��s&R⌗M��QZ��]wߊ��[���1}�]p�m������+G�,tv4����߃���7� T'�NQ���U��)AiE�-[.���<�w��|ƌ�0���q͵wbs�N��Λ�ӕw`S�nQ	.��W
�A�NX�[Z�Wv��K�����9��{�u�V%�r�NN�Ɉ!Æ�Ǣ� 8&5-�ד�� ��+���|D�&(�+ᇝ���-��v檊��ű�Q���[�A'�nZ���*�p=5�+>����)����X
�V�+�z��|G8��K9{te�dq�$� (}�LD��R�G4m�iNu�ʎ��	L����y�{��fE���Rjx�a�`6��r�[Z��n�L��J�'Kb�ZE3��&[����J�ƕS�^�{�[Sz"�Ȩ����v��������Z������5I(\u�>�Ϗ	��c6/�2-ҡn�|m8������W��օޮF�m&I�,�ISf����セ�3�|/��."i��5 ���F�]�����VH\�5!x:�mԢa�BL1�|�m(7��_w�MP�j�V�1��������Iy�$?��F�Y ���H&�����iws�<4V�y=Ry-�k!�7@o��ry�|����v=�X�vG��RT�\V',�Z;� �	�AMZ��Tv}�'��\�H7�K��<w������x�U��⋅�T[S���&<��s���SN�v4�BEU�.Z�h0�[��a��uV�T�JB��^S��.��-;PTd����G*Ƕmې�E�j�H������1 ��{�@$r�/�P�)�0�K��f��%`򦯮��/"�we`#����2"ء�)NC^c>�r������w4lZ�;o�Aϸ����ö�-b,"d7ٻ��I�߯$��1�nTzb����8&W�%�l+�����g �3P�-��JB�&���`U�5��:�C��	_7����^N�f�x���[�yoSя�e�5��?�+����ز�^��u��EK��s/a�1'��#�ß�|�hh�V�E��'��Yt�H$ø������O���\��"�8�Q��,d�;&����:j�B� �#v� �A:���_t)�9�(̞='M=Y�ml�ŗ^��/�S�9	��64����(�q�x,S'�U�^1�����_��_���V��:�D^�Y�`�y��1h�`B���2y�Do��Ɉ>��1%E Խ?���фN>�R쥸�`w���N+4�$�fE`��(t���q�׋5.��P�����!�J�ȈdA�
��U<���;6�)p[�Hc��G�<�W#��0��8�F&<u�M&v�{�h���b���X��/
g�=J+��ETQ�ť%�~7�5�׹
b7��O̐� R�"�L��$q�ŒS�=ԉQ(<����c��I{�d��1}�+�QJ�Wy�������.�Jȳ�    IDATC�	�%�ǚw��#&��'���o>ƦˡqG	�F��[h�RD��U���շރ�U
�ŋ��,��jCO JCI�K++��ݝ��)C��VM
<�7�<q,��o�+�Α3����ןqFŒ�Q��P��֙�>V�'���%��9�~�TP��,�h�?�d^� A�;��<,�r�����_�RܴW��t���bi�5�˘�t1��	��}<���X28�ȱ0�c����ePWmm-��r4�O�>�{�1�88㎘ 9@ƿ �X�e�9f,�����Ԃo���77�qW'*�F��v�;;���ø�Cp����a��C��ۃ�O�Bg[+�|����Î7�L����J1��W����Ѵ��)���a0Z�3��F�c�Y��]X�Kb�rX3�jw^h���Y-t�JF<t�-x������W^��'���7��� ����J"TsNI�;IB�*�V���ⷮ&t��9Q�\��E���y�LŮ�� ;t��(EC���-����^��ڹ�`��]ho[Pv�|���lll��| ����o����<z��ٰO>=�����GMŭ�O��<����*�i�:�H�c��h���cqۭ���I���edOk��A5.��rټ����NY[P��m��\��P/ZZ����f3���P_�Æ��%K�h�"l�фÏ<���_���ذ�:��(��]��5Ԭ�b���!-��Ի8�8�HIh[q�Wc��r�X����]�z�����������E��G�w$IU���a��1�%�(Ԭ}��Q�2i)<G���$I)HI_d�"?<��붉v�� �sϠ��a�k���d,O�\����쐙���[R���n�uz���������+��g�Ihy<ϫr��r���<'MfE�FG����	-%�SI��:������1��q=_#�����ԙ�Y��4I��J<�P�>���)j�|��:G,:]���ٵ�Y���O���{��Q�\���w�?����(��Մ��C���0��CO{ݽ��$���k������n��:e%��>k��2���f�VD�@8���^����+L��0�Y��W. �s���N3B�fL9p,����_~�-���`�B���R����U靼�*�F�y
�"'8��(ar}��#9�ģXL4�Ӟ��B{ 
��D0 FW2;�V�ĩ_�9����hm�X�2�7�D:���.�Ig��.�FM�\y-+�,2Q,��/�Ô�I��)'#�}���0�?�<���z,X�@r �Y#F������a���h��Ɉ���-�b��u�Dr0��Ej�⥼�%vF�^&�-��p�����-ͻ��*K$K%P����֮ЃH�!��dA&OW�*+�7�a�����[k2 f'k��\E�2�3P��U_٫�Rst��B���&��Y���gA��W��B��ލSO>�7mBkk\D�s"�K@�t,Žya��(\�4v�J�Pw�LȬne����Y�r��v9���J�(�D0��]�l��yy�7�8�q�nTl��Z����\'�U����-+&�[n���o���A]�4����Y�`��	5�`�q�C���`�z`�;do,�I���� ���ѣ�	��j2����|Vƹ��S�%Jmp�;kPSS#_���� �I9����|��g��_�Đ��p�7��O@}�6lܲ���\v�������nO��ƙ�5�*atV�F�w�ݑ�p6t�p�ᗕ{1��?�ן�˥���s��~Z�Z�����&�Q&t���e1x�pIJ�v톕4MNl�Bu������!����`��� ��߉����qh�����"�V����W�-��� $R�V#ht
��V���dS�iQ3b�$wZ�
��Fm� w�:��$�ΟI���g�g@F�y�Z[e�n1`�k��X���X!�'�5}ԹF���ѢC<�+�1��)���؈\V+�Oy����r�дHQ��@�����H�{v�ʵT������&a��RU��^�!�F�*��@��h�`bm�0y�0<�Ƚ���),���6)X��9��nz��p�`Ԅ�«o`����S0�K�Ә�י$�����:�U�����i3��8�7'��a�H���Y���	�¢Q֋�j��T4�ׄ�}Q�w��is-�ű
z��ڱCO'��h����� ���VT_ ��X�}�/2�O�x�IK�4>�uLO8!	��OL褅1�sƄ��F�q��6�����fH ���Icq����͸h�b�SvȡX�x1"���l& �O��o�eW\�p$w��|�1�._���Vt��P\9�x=��$�J�[�K&����->|;� �3	�\�Ṯy`�I$92���ppLW5�Z	�z��#h��.C"I'&r����jZǛ��21�ݢ؃lyp)��F��	r=5����x��ixm�l4n[�k��=��;z���� ��IX8�"�T�T[%8	��aW�����d��U+�*OS�q����[�p�wv@�=�ɍ�P�R.t����t��z�`�����S��e|�!9Y��Ca�$1�����QYQ�K�x6�߈��P=P�|�q<�(p�\w�m0ۊMdž�����(�(�M��%)'�B��Q�$���bTA�GZ4"�*@'�N��z�]m�HǓp��^�{ 2������b��w�ŗ�������|���'��$�}�V{�b�c�f�Z���
�Y����J-)���].�|x�l��ˉ��!M�/��Sl2[Q7h�L�x�(y��F"�Rd�� 0S���P�?���"P:tz2��N�R	�Y�2vl�p褱��3���-�����TL �.�mmزi�$rJt�5J �ė�uFl���Å�-�{o�:�Hgm�ѶP�
#v���ΤΠNP�ҭ)�B���;/��#�2FlE��P��I8�MM�"D#J�1�d��4d���	��q�ѓ1f�X���[4lۉX<�H,�T<OY�$�X2+�9�V��x!��*���Cײ;���룖h�ʋ��?��߷kW�q�J<���xBO�z����ɓ0r`9��6L9�@d�q�74�{�xd�P"F?,Y��]�h��AG ���aH��4���W^oY�b%O
W_v~��3�I���x&�C�#��P�C�I&��T�����{��s4�H4&��X,���SC�Ho�"�%3Hk",�.� n�dGJg��V�U�{��'/Z�4#�(v�참��й��1�g"()��y�f{v�eI��c&��k@8Ё|.��ÇJ� ���`.��Z�`PeeL�:��4*���V�Ub�w���BF�F��DiѐQ�~ăa؍f������T��:}V��T���+�:���*�	�w��£�$&r��R�;�#|�`��z#��%Ei�:�ac��i
��j�*�2$���׈�6�&t�N�x������~�r\��K����F��n0�Nt0�`�ٿڌ ��n\�hA;[n��F垫8��Ϗ���V�0�"��?�V�j� *^`���U:��@H��7�'�p��ظy^}�uz�d	��wPv����v�YO��3�ĤC'�ڛ���@6���`yZ&uV�����!ЍZ�M�)�2ɨt�}�v;B��x �V�f@���Ɍ>��%�=.��vA����{n�i���?�g�����b\p�ɸ�o/����U�X����ܑW>K��* ���$R� 6oX�K/�4NT��/ۀ?���fy����:�tv�h����R
�H4.�n�9X(�p�����,�롗iGf,B�$��0b];q��!x��G�d�
,\��hD�Y�fąa�喫�~�N,Z��sV�Z%Zt�����W^Ǆ��]�W�|�7�c�ైg�P<���k,�#�.W���Ƚ*t����v���RVA�)0����H@�2h�s�1�q�'����>�4�QҞ �N�[y^�4	�@T{��C7����c������ �TN����42,)p$�{����^���3e�a��?q���2��xR1��a.4
}�z"�]̏#��5e�p����q��cԨRPJ�6�k�.�Z�F*E�X�j-|�8�kG�*+�Ήt8L�^�JK���(C����=c:�����7�����v�TV�*���$�,�x�2^���:�8|n�w%����I>��F#`�/.� ���."ݡ�%��{˱�݇��
���U(��H���<uن]��	��ѩ�2r7j��l���нEN�ضV8�L�-�-#T�^'Lf��s18�z�h�`0*����%�
�G4�}]�s�jk���aX�`=�5t �q��$ձ@C�d�.����F�3�D3�F��Ǟ��`1j�q�Eӽ��]�}��
c􄃑�1����28�eҡk�6��9y��$���cB�q�e�J�UA��bP���5)\�OEp��#�o�?�}W\z>r�*����f�R)�g�׋"�	�iY!S�S�)�r�.Q��y*ձrW$3��P�hU`��Y���n^�~��>����	�!GJ���rVw��#ϑ���%�C��B��$���f���v����A2��ĉ��rz�����Ͽ�_n�Q&0�<�w��eH�(�i���h~&tZ�R��;�%e�U��� |�-HD���{� ��OP�ܣ�Q]3@D��4���G,��nD{Gj��λn���Dö�mt��Q7x�>�O���f���}�I\�)=
,��B	+\vnv��D{�r9`!�7����8�tԄ.>7���RIFT4��Ģ�fA��?�7���^��C4��ФB��]���T���K��d�"|����p���ƬY3q��g��c�ŷ��/7N޺{|���K��y�`[c#�:�<v*���o݉�a���Bc�!�� ��ʵ!b�	���p*H=>;��S��"�9������H�H*��w��q�����-<����������E��~F2a�]8�ȃp�=����zrx��w�y�v�jnG*������ti�8�An}���9s���8{q��w����D���W��~�ǽJ�I�2��CȏX�Nq؁8�7�cݪ�X�l::[���Q^Y.�Y�|5z6�J4���=��[1�n8�M!� �p(*��[V*E*)k���<�jJ����7��?��:���&.y�HL��(�J�'�lo���~�:�Pv*,�����M�"R�酑L�s =�Ju�g5�;�୬E{w �W���2y�E����`ůohz0����G4m:�wB7tBia�N��ݻ6aܨZ\u�YX��h5!�G2��f0�e,GjGj��$p���[@=αpLP��5UrAJ=^��yl[�������	)��Jf��P]Z�ݎ��&�l&0e�[>�^_v#�I�x m6�p( �ଳ�����FiU:z#ذ��6�#���܁��tF��fHp���f��U�fTY�<�a!MɌ<5�ca9̿:i
���,���sq�y�C�ˊD(�C< �G"�"��&5ڕG����U�lJ��V �P�	]��V�r��+^���_W�y���Q�����.�B5jp������]A��g��՝&w�,I�g)L�DK[;>��c�"������}���rL=�d�r�3�Clkl�#3���<������nhw+	K��iZ�j��;�"D��TrX˼�>�6EN�h�s�$˂�tD�8�Wz�x,��و�?&�����Հ`����u�]�&���#؏�'�
���_w>$4�H��I2b�F.6;q�t���5���(ҙ��h�{�e��NC	��%T�`8,��G�=�ф�Æ"�J���遙��D
<j)���5�k'����	lcI�.�"��`���V�t�e�f�a�������ĸ��� o�� �Y��;z4V�Z)�~h���C0;<��'_�+6Ao� �Ѣ;QA��4\���":ä�j�S1���&�Ϟ��2ʮ�n5"���a���f�i��~��Z��λ�h�D<�������钦��4������Qc����s�n�^�Y�t����|,��K�T��Y�a��j����w������:�H�2)*`�C�U)k裿D�EQl3��c�B<ԋl��W	�W���1���)|;;z�ze4zđ���kQ2h��f���u"��xUT^*k9�v6��g�D�ׁ�x/>���ރ��WT	���
�g��ׯ__��Pd��M���lv***p��������N��U+��lش;����ц�:�n������_ �����fن�RZ�0&tv��ݤ5���C@&��"�k߁��Ÿ�oWc�ү���C�bq��=�^�F���r���d�9N��"��d5)\f[��a���j�zS;�:#��STR�!U�D�R�3�&�Q�f���F������Q+f-�`���8��0��#PVY��]��n�R|���0�9Ho�Fo�?���n�l�	(���M!�:��q5�}nss�{Y���@IH���k�A�ⱇ��7݈	�cܰAh߽�U��uX�p�p��ʧ2��_�$L���C����93 ʾ>�X�2!���jU-��Ѩ������~�y�e<ꯓ�T���	��￻ﻹ
�2I($p�ϛC�����¾_� ��O�t�X�l5֬[������G�������7�vn��n$r�y���D��SR.��'
/�h�ՀǏ��܂��.�	�T�`@8�tl
�"�Q6b8=>��C�^�	�m!I:��S������������?>�e�h���Ǟ®�nt�b�q��&@+'k���=�l���GI�"Kj�[���Nc�ŢLDv�M�J����Q��bE��A����c!ɏ��jYap��<���F�?�@��e���s�F���x�6"��p�7�����w��� l*�E�Iѹ��G�C[s�.�^ $W�:d��k�,�����;�{q�}�U����Y�]��Jr�9E�IF� "���R$?������
�=�XH�e��H��f;���8��3e�ܳϣ��]X4�-p�p��g�(&���y�eY���4��G��< x�ifRX���I:�}��}�~��}��������������QK���Pb��;��:�v�H��(��`��`�^�?=~�`.w�j
 ��F�6��p�at�z�a�K�deQTQ*kHz�s)�q�_p���x���ㅧf��؎x4"+#R��9�|���e?��x��'%�ӗ�v���8�U#kde�7x�0�wuJ2i�D�s�����o���~�%˖����&g)\�h�G��J[�E��$�oly(�q�G�'���6��]ԄnГ���ӢGs��{���+�l�g0����ys���c5���Z�f%��/�W
D��vqQ㎌��j>���o��דƺ��(<�ÅN��&�`q����$BQ?LV3�{����a��a#�ECa�����n�$�d:��"	"��z�`A��rZtt�*A,W|�i�J�q{���'�����p�������!�����c��n�ڨ��~ϭ����"�݋M��b�С�<���"���j��J9Ʀ`	�p���e@��-�}�J�7�
6��׬���ʸ^�jq��b�v?�)5�(	^ղK��#t�(��A�H��t>�~�bq�q�ۺe�ص<Tv[7�c��Ex�������=>��X@I�9�]9�*�A"^�p�fuR0d5)x�vX:���Sq��Ѩ�*Î��x����,q�>���]><���0� ̘1���]x長ŵ�q�L�~��7���f��}#���[�t��V����XNW�n/�:x%�z��X�aZ�v��+/B$��e+�sG3�i�(f3z��@�ہt&&R�,��z��ɗg�����G>������{�o��oB��@��ky)va#=4\YŃ�������O�⯿��a��������ł8����so1Ye� ������j\B(Ek{'j���BQ� <���08K`�)�4�3#�W�݂ �y�2��P/S�Q(`N�V%�-�B 0g�    IDAT��a��E{,#��Į8��j��m2n��������V@�v�	c�W�(�3YI�b�Fʝۉ���U1aE���Zj��{n�o��3��}?k��#_W�Ol\��+���L���81P*�E�f>�ڞh
�Py��S��Z�w6���4�� �Vɔ)(�˅[w�lu N�D� ��5����Ә����+@�lF:t��Q-�Ӂg�����ُ�����jV�y�:|(+���g��y���SN���^��?�\:m��O�6M
9����2i6�g�<EE()����]t��J�1z�,\�3����Z�E�5b0�s��И�<���[�%��g�NI�	�~cpzgK��{Մ��mw��c�}7b��O��ѷ�SƎ�	l4���cƌ��G-co�C�edr�\�l��?R�(����a��m����գv�$1�xK���QCjB�V
�H<*���h�D�XT�2`d�@_j��R��z8�^�Ef� �(M:l�A������Vd#�)����ل���=N<�h�X�s?��~I���h����ju�p`�C7㭗_BG�6s�a�noÒ�qȁ�e������X^O�ص{�54h2ʈOF�yH@W�ߪ�u��οM'��"@\�
X ��
rcnV����j#`b����ݺ���(���;��쐝fC�vl�ߊ���7�z�u�z~�9().D)��YX�q#����'L{���l�z�8~�dd��������>���*R�i� Ă��4��3��Ǣ�؍���ûo��^_��$������[\|�W��	����9Ee%���7Ћs/8�_p6:|�8��tte�j�z�	���3Y���9Y	0�gSw}��Z|��<\v�E8��c��c���xa�+�E4H'��50����;lH%Èƣ}	�d�HBW;�K�R�l��L#�=~�TBW
�~#z���5y�aT8L��Sp�I��d��8�7������%�PRQ!v�ޒb�o�*����H���/Z�r%G�^b���y�`踃���o!�7��*��]�Xր\a"$ӞB"���ߩrFpg�:�v��6��P( "ƽ��ې��
�bj�sЋ�rf��I�ȯ��q�Ap¤S��lWU_��t���+���AyA��_�"_��:;�~���T	���g:(rzQP?�QU7P�=+'D��)z���T�4Zй�U��N@,D}�zx���l�)W��
-�<t4�{z����&�f��Ӏ!��d�˼��h��A���=<C�<�3�|���()sJCG0c�ĉe�z��cҤI��`�LߏGyD���<w���?�n�$v��L�p ����^-���SN��9/��YO=����o9��Q�a����ew�{w�K77O��\C�$b��JB��{s�p�M:v�)�L�ikDu��^��oX�l��`'�����
b���*��0G&
������v�:�h�)#`�|��r;vm�ļoV c(��[#c�@0�2��f�I=S�?͑`Lv2�ψ8�&/���#rWHTV�r�����p��EP�v��M���,.-��ȫ�#Ԡ���#�`��f�	���h��_���+��V���'�1�@K��n�+&����rF������u����T��N~n���@K{�$�`8(����|�Z-�6�x�¨����ݶt c��L �����y-\���h�;k��U:��͉u$o�	���,�x�t�:P�uv���ӊ믿k֮Ǭ�ϊ_4���a#p�!�����׋��*���=^���p˞���#����Z��;1��S`�������:�����wBg3⌓O�'}>��V���>�ɨ���+������v�_���� ���JȮ��$��z\wݵ��HeS(-/�1�??��$�uC���$	�H��3^<A�� �v�-8rJ�;҂ԝ������)vc8N��
4�K�[�	���TYE��"����]&Y�@�����z*�H�'����W\p.<�(lY�F��5W_�q�ăBKk;l'���[�,��야���7�[rB2܁�QT�Ł�U��f�X����h������������+R�����~G���؅�fA��������,Ȱx'ؓ�)=�u�P@)x*�z�r)I��3���Y����&�	tB�bҦ1���dM+�3���W�)���?*{�����������������?	`�w�u�P�0����uuf>�3p�ic׮�v�m(r�"��z*��U��3����l�T�V<(���ҡgDT&������>F��%x�����X�EHKd��F�������i�L��ܹs�1o�kE���.r��*vtt��L,
uQb�����F+`r�Y\%z�h��]���t�La�;�Y��%���g�!�XJz�<t�C��Y�P��M�ǎͫ1rp^|�A8��ޱ��6{
��d���X���ܘ<N�$��IZ�TF�|-�{v�z�	`ۖf�q���a�T�[;X:�ʮ�"b� r��k�����C:���p����q�r����XJ
�Ȩ��6
�S ��4�n8I`��c���Bg.��T� B�(�~�Wj�Y�?���i�!'0L�R��P;�v-^x�Q�v��uW^�I�GጓNB,�GÖͲ���;�ѣF���#�-Hyx�����-�z������j��]�iT��f�x�	��u0 �.v2�fr�d�F6��	B�\����M�c����''|o�\��!�h�Q6l8\n7|�a|�`<E�6b��av�,_���3f?-��w݇h2���P��nԌ�Au�X�f�<�H�|rlV����[�a�z)��r�(�Q?\:����΁���=]��/O[C
�ͻ[�ZS\"��N�:��=��"��mTO�֨�p��PY'ԝd:'q�8�x��k$Q������N���o���>���[d�:Ģ3j��푎�-/���0����lÉ�`B��	HBW;��<�����F�lf��]Sy��iB*��Y�N�s��]���^���p����z�E���i�\�K ]Iv��B'E�ta��=(������8j"��d��BA5��������'q� (
�����u�Si�S�ns�?Ϭ�j���3˂�?#��e�R�i(`P���z�ڥ�
�A:x�hPFԒEҘ��IH�.}.��P�)����ρ�~.�N*��@i ��w>�մd��;syTe^;�W��NkA�����1�Y�>�"/*�{�}�/�9ݾB���"��KN'@s_���t�\a �\��R)�LF-��<u�=�tY�����ހ�e)g��:!������=A5w�6���.�%�s�xQD
��� L��B�+S��`���kVoGIu��4�	�a������zk�YK65=�3z��?6�7�ү?��١;��|MR]��o�*���>�r1�����lA*�׫D*���jt���r@�t`4�G�w׈?8w��D�H�Vo�cO��0l0U!g!�ǁQ��(r�**��_n��v"q؜n�"L'�����N��B%�M�G*���b��Ha�,i��i���8��6��[
���.���+��!+ً�#��nH�v����E<�����[�K������g��".���S�>��"F��&�D��7a�����VVY�)S&��^919�9ѥ��|-*��H- rB'�)_��B��/Jo��I�}w�jܡ3��߫�����G ��������_|�~�9�6��]]n��SG���o���V��_��G��z�.���:#���<(l{{+��N�������`�}����|u��2ͥPS�E�U�`O��|�ۚd���	G�m�~���GU� ��.��.4���ls�M�5��h,*�P4$�?��`@e� �F�#s��N|�:�F���0[��;��)��*�qC#���%r��!��B����?(B�^�.�O�.b6�Օ�����[M��2)Q����H�qǵ���3�����1���G��d*�`,"*�=��	�K�Q��OJ�}�x)��pH��ɞ�uZ��Gp�	����^EW$���) %��M�#��C ��ΫQ��--t6�N-��8�r�,�ʫ�w��?���[Di�{g�V
Te�t�ܗ+nr��[!G�2��I�|�^EjYgP��{�S��♾�c���u�?��?�����(�Ay]R���|��/�{�`��G��]�I-��=n�u�w��p��������a�WQ[3;v5#@�w��dY�^���Ly��TPx�Y�B-/	=�ՎN9	7^�������@G�%gTmTX:j�V��
��ج��� _U�����Z�P�rga)V��\.��H|�PH��X��8rא��.Rx�	���j�J�?��7����wݟ7�%�t"�ͮ(�5w��:z>D��	#���i���� �oC�ۂp�\[�tp���ޅ�N_�Iw�Gq�T_4�ol�%#.1Ie�˛�t�:��ѿ�лa+�E�dAŀ�Z[Q�����>��n�����DY�AL8�%���j%)��yɞ�m�N�9��F�+3�8u57�Ѝ��$����B(FgW�輓;o5t�H<,\a�ǋ�Z���EmNg0����-�P��Ø�b@����W������g�n�`Pm�$�"�C|�)J�	�f[�P��12��n�d��F�Z@(g	����C@e4��+�c�G�F~�_�1�8���M$�ͭ�q�:fW�X����gwğ��A��k��܇��u'���6 ����]o��.-^���_�ǯ��&�jiG	��f"	��Z�&�wn�y瞃�n�	������?��V�4�����s~�+L9d<F��w����" H1ra�ʕ�������o��b ��bx��lu�2��S���nx+i.�c�ַ�aEO��"/F���;���k�Fqi5�&'"ty������Bt�#��0	R�
�bb*���1X�s5���T��%	���J��Ց�ޡ�h���8�'
�t9AQ)�u)\�ۓ����O���>x��6;�J�,'!U��(�錦��I�Z,"�G��������p�QS1��7�O��ʃ��ۊ�3ZdW��Q�[DOI�����e"��!Q$�Г��$ Ws��K���V�>������g1ϯn]&�4�\u�^H�L�}Fe��獮��S.�p�%��m�_�,����(����G�t��T�|_Ǯ���%x����kt�N�j�!��*�]��aqke���ނ�;w������f���.�k*�1h��p��%��1�)t�)�*K��$7�݅b-p����&�٧ÿ|%�
�!���d���)1E�R]$��Mx?��R�P��p1v{�����pDi��6r2,,�'a)*E�l��NY�_����o/<{�����xZ�s�AtA""�~���k��f=���ǐ�"<��=hmX��k� �0�7�����,M�jѵs޻v��]�����	A�=�G�� ��^AQ�G%�G��5!�dA�(a����g�s�w����v�z�_����WSU�����}�z֚�����J��Z���`��,���L�:�b�����t*�G�x������U�G&���^l���IOx~�?������[>�/��Mԛ=�US9���ƺw� ;e���oܸ4�pΜ���.�C�.7�ڪ5�nl�tezz�T
�J�jI��j�ҁ@vtԒ�y�O�`k{�`KcAh�Q/o��y��/þq�m�8}�AT
�8z����HM�ZT�Q���T���#=�4tB�w���F��M�B�T<W	�3�##9�f�T�"�}��AT+�K�<ɗ�z=Ӧ�Qv���rc�L~0G�b�-�v����Y���U�v��eM��|�_�G��Gq��o���/��~��pumM��fr#�7;���2�\D��CP���c���̹KB����<��F�~�9O�3�x;��]���_�4��/�7�8&l����+��?|��/�7���x,V�;����G�ތR��f/���Y��x�t�d�Nm�ﰌ	cjnVY���&"�
k%����=RE�Qs �J�5p��O4��`rf�H����x��c1�?p [~lm{[NE%�hd0�Vm6�$�eQ�s��ȮB]�0b��k5�Oph*������]��uXZ��l��H�A�D��o�̷��½Kg.u2��[])�1�"���������V��)l�Z�ҩGM�����ឤ�p*[ľ0��(+Am}�wO|��{.~::m��_�J��3�;�E��۝��g�{D�;&8�_ݢ��]ߎ\��@���
�XR�����N���Ө� 
➮� 
���� `���	}D{Q����p��y,5:elV5Z� o�c��adb�p�P�nU��v�~@��V��@q@���=�c�n�����_����S��v��OިQ�~�_���yp}[ª&qO�^�߀�-m3G�ɤI|����Q۠�|u�ҩ()�M��v^����vU�^8&G3G �P�s]:�W��K?v���W{�#��mWkh�kȤ�����%(.���BX���N����Z�z54��h7$�ǰ�F���ǧe<.^���<9���U�T���_���)��9|����'��QF�B/�@R%�>��?�<��:�ƻ��A����b��D0�TFA�T�B�xPnI���Ҩ)͸��r�c/]��n���p:,��
Eq���gI�A-�.��C��sр4ٳլgH��JhL8� %hG#�^��3?�'�~�J��Ŀ|w}�"��$�K%�̷rbY�(P��c]c74U]����I��洦�{:%��[�c�;D���썂���w�E�	��-W�g�+�N�s܏��^p䇽ޕ�T�u<��Y��9���Ocvn��>����j_�&T���2��jd�9.���j
oa��̸Ҍn��Hg�
�n<�O{��<�����O|�T ��Q���*^������#R��ƷNcb�:��@4�hfLQ���&��*������;SNwu}I���"%;٠'��F���T�$9��M� �y���X{��#b�ϖ=zIy�#ط�:�*n�@�f)B��-D�	�8=��'�.i�ˮ��a�g8C�z!IJ�+�%���d��1���ó8:?��{�[��٘����'O�̹���[e,{�����[�m�:=<�q��(�G?�	,-.cvv�<@A�B��	T�lwE�����롓��e��B��y+��ɑ��ί���Z*�hzV�D��5�:	�l5�a��
L:m׳M��v$i�!�C	�<�}�~�Ǣ;�k���f�3�^����L�`����!N{��5_�]e
E������N��r8�shi�8��ʞ�s/�%��R).zhV�z�R#D��qO�f�Fť+�
�醃H����Q�&���19�����u��jauc�"+e��|I��q@�T���MoF,&�XIGכx�����5��o�� �SQ�p�r���sg��>Aq���/��=g^W륏pN��ޝz�TVZ�̬� c� B��nt�(o ��x�#�����h
A�
�����NW(D��i�8��LP�%�:ݮ�������ruA�(�u�q�oW02>�R��9q�:�u�mG�Z���C��i�-J�}�|�O#�IP��oؾ����B�pH�D9tf���?�lV�����,rqJ8&P*W��g��R�R3<U �������E��D������'>O�1;\8_��{���ֺhv)�b !cN��bڑJ$d�	.�XK��?��ƗH>��`v�,ZHxDE�ֿ��d�%:�=�ڐDi���L�X�Z`oS4�՚�	>3�+����o��1�B6;��W�������8O~jmGq����0aav��:K�;t�f�)��ҿs��D�Һ��Q40=�D<��'p���Q�u�=x������W�R��3�1=}�����6�)�/��V�gs�
��t�'���y�l,i,�Ql8zʐ�Ƽ���9�ڸX5'v�v    IDATE�,tdlT�DjUСSd�9�P8bcz�F7\�,\�З�6M���C��(F���¡�$�%���N��ubbB�Z��d��l��_���������p��>|�#����c����;~Ad|\^]��˗��������'�[��Z\����|��W�K��H�ǰI=����b#����Q0���>���p��;1��r'Q4�e�q4�
.���A�S��%9��ZSDһj����φ�X�I+̄�˖^�JP�޹��2q�=i�u<��?l�mxn���;�������*ā�V @㿚���uq\����D<>7��Zt��bZ4B`l�b�c����Ѫ�1?�G*�E����|�Z+���'�\�r^����%=?���,I��mτm>NS�����<��\9񳹽������E����~.^ƅ�WPkuN���I�P7�@xt}�1����d�c������vSr������0D���]��R���x��ѭmbs�2�:��������㘚���p&G�2�Qk���ʯ����s��9�|�A��Pa�G=./ⓟ��@L��1D�-D'�<��L�TSHk����DJ�P��D���sN*�	�@ύ�С3C_�|U:�]��,�6�6�"��Cg��1'2V�	�@F�aE�,�Rx�㬓�aM��z:t޿.AW��F,�n9q�>�8���`��#�&J�m-p��:�X�=G�Z@B^}�d�
���@r|f��Y�ne?���w��O����~��*���&{2oULX���ý�C�������^|�_���'瘔 |dG#�T�P�,r�F��
5j� �����g3 ���J'5Q�����
uЬn����ib��#�Q��3����QN�����I�{�Z4��F<=�S���2(�*�P jV�EϜ�w�䡦3�;�.�F���������GNC��SS0 !�*7��Ю���,����KۤO��|��$b�Cz�=��]��%׼���K����Jٝ��,l"ܮ��v�y�p��^lo�*�<{��.�L���o��&����4�@M^۾����_[�W�ՅU�K��&X�� =2����>���dP����CwY� S�A)�E��B�xR�R�a���mݺ��u��Tᏹ�D������oر�v��T7�P������-�V�{'0PB04���9v:`?��H�����?r�����U�hX�Z�%1�����	 �h��@H��Y�;u)�M�R84;����p��C�t�4N�z �\�HL"UY�PH���<m��$b!��5"�Rk�̞��b�D�u�%L��XВ�m,�h&�n"3p��m����P�&ӡ��8t3���R4B�VA����#�hU�ѪdL���i�pc}���QqAs��\(
lF6��Hi�8�H�S��*V��U�HZ�ёL���8����{��eF\k��!<�,K3�|g9��4_ʞIT8f#��#��ӡ�ѡ�����z2+��~g���Ҙ��F6�i�OM���Yy�FK�<��F���\�F��@T
�M��;{|Zb�l�s#��g�,_5�pDe&9zo��F0�-�_��ݼgDX�Ans� y�=xF������c���#��r�IJdv������;A^�j+k�TI<�B&�����M���ATJ[VBcO7�q�4�����t�0���a0�J&P�^C6��o��y�p���8�������S�����i~��D����>�)<��B�»>�,�S�{�`�DB�+��,���;t����auuQՎZ���SvIp�f�3���[%��Z��{I�����Z-k�N��#t�C:K��:I~�"Q��Pۛ<�������ŀ�r��D(�8˰�&b�:�.��Z�a��[�^���G?�`rzV��
��c��r��r�3�$mw����'P�6�]�b��|�#YE��9ts�ж6�1�q+%�vU*&P��ʔcAd�Z�)����a�474�-Nye��|�R�b�m�]�0�����Z{`����{�V��w"��	ٱ�>�6�����s�M��r� �Gի��W�<e<���%섶�10� ���]���^��5����eԶ7��~7����Ү�^0(����}�8��������:�BX&7�7|	��)��~��9�R`ˊ�O!����8$���BNS9�~3�{N-�n��8$j�F�Z�tNLKt�������ˣ]��Q)"��"�M�Y���/7?f�7HG��xH�gx��M�P�T
U������X��F�XE4�To�$���9�굦#y��)���1�|𴒗9���ۇz$`%w�H3ɔ�9�N��=��?Ec*�\*��+����BqL�%��;�T*7���mYO��F��\��I
���bcc�vsk��u��Q��cS�'�����uap�Z13����XT�a� )3�2�d@B#��A��uM+'�YV�N�"�H;�����8jR_NK�O��I.��b5=#��a�a�;_��42 F5k�w���ccmS�Yd�A<���Ə<�Y������y+*�ma |�����N�Û��V�I��u�Oz�� 35�������n�p"�
��2I��(�*�<�������C�nsW�6�*k���s�:�>?C�: �$i�w�t:r�����9+2�D`�Ɋ%c�Bc���_�>�z��=�J���NK�8��H��p����"̍���q���Yq�TȌL�С#"?�S��Z ��-�G��Y���]K`(�Ş}7��0p���.\Drr���[,����@�;t��ӡsF��6�G���l��S����F�MYZ�2s,���t>��S����O,Gn�,����=C�r�ow��K�����ݙ��G�س:��č��)�>�W�֡����Ua�C�߫��۟�:�2r��#H[��y}�G�G�4�Ϡ�A�ۣ��a_4A�m9����*���%D�"Qlm����8w�7�W	~�g��@�����:��3K��0ґ��O	jǈɬ�8'ڱ	�X	��U8b�H�TV�;\����ؚJ�P��S�6�h���Kgu����5�A��,2&�cTHk���,y����"�"z�&�R�/5F�ubu
+p�,�tEC!�U輘��C���$�..	G�e���cٕ���\d,��-Fe�ը7k�&T`� ���C'�v ��}4�x&���ulnn!�H#���܍�pr�yISe�8g�t����̀�p���N-�A���ܨݶe�l�v{
���X]^���M���������6������H�����}���,=}�"oGIg�h�t�|��ȱe���߻ѷ�p`>C�ȡ9�IT��uɌG����KC@�7*Kh��U���A[�h�[�3��X�܋~7�����8��I<���k���,���߂��i��U��{�{sGO����M��v����,֥����:zM7v��N�3��5��+���#:t��@@�q��@oEl>[���нC'`�ψ���F�C�C�=aP��+���$[u�U�/Ζ������a&XggL�B��h:��f�UC���X������?�Rt�e<��Illl���#x�ޏ�}��C?�_4o�5������q)^�wPY��������06=�p2�z7���^(:���}��ru��[Cc�sؼ׼�����{�xEݜ�"eX�|�?=#�����e՘��ٱg�s����)�o��t?�X<��-+qU��E0lcv��w���]��o��9"��z�܏R,j-8�Ob9�����/:G��j�+d��H"6�܏ƩNh���N������徶�2�����V}�e�a	3���T�;��\�(�I��c{��3b�bq�cIMg�>\���_~�=�__���v�Aޡ���Zj�N��3�����'�����j����8�&~j�|��G�+�QI���&gI�ʾ)��tm��Hh.�k��QN�,������s0��,�^\��;rn^:7���G����u�a(w�I���Hd��j�C��3ui�����D=yK��sf�ý�a"e���@�����U�R�c��k�E��ΦѬ���`q<jfvZ���"\�x��Hq�D8��^�� K��n$��pf�_q��.~/�X.[)Y�;��ms۬0#t+��9Mpn���a�D�G�_<��:v<��$�.h#!�v�����y������n��` �v�c)���hc�N��O�L���5�}����)�:s�./�ˠJ"7:�Z�ً�jU��JB�&�Π�;;�2�'��1s潣C��w2~���Xrg�Β/��όXa��,���<�*�CHf3Ʀ�sN���w������ͱk�ҡ��H���3�����(�]��d?�������;{N����4�v�7���E�m��đ�;|G�Ο��������+x���Fg�L��cam��I4Zyǡ[!y�:�ܕ��}�k��s㚳�����4�谺
�ͧ1� �&9�6�f~���T�2t��xڞRF��ߡ�p�C���:ײ����q�{���Ts���#��v;���Yua2���_��O>Pgu��C��{߲a
G
މ԰}D�VI@;��ʢ����h�����x>�=�7�K�����f�h@d	י����Qc�t'+�n�hǉE�mD�>m�j��I�q�:�_y���]�����Cokt��#9�j�)��~/�R�,�	���m�T�&�������Г��8�c��V4LIʶP���Jb�'I�fG�;}�ÂY�,Cٍ$]��n(MST2'晡���Ϟ脭�GYW��._(���cf��:y�G��'��g��v��1��OY�b��4�˨��g�L"
@8.�q$��1
)`�#(.z�$���~L�L��JoY]]Aqk[h��o���:us����~s�x��Q��u\�l}ģQ��y��.��G���� s� �5Ə��پ��Y��.�Ԫh5m�Nsﳧ�uC#3�?������͢VX�T.�fa����/~�^:���.*ҿ���j���^}^bd�`R�_����'҉ˋbHT+������C�����5[.2�bP��d����D�X�X���Ls�;�щqAw;t_r'3N�X��v������-�),�brm��;9��9trp'����1��]�T����8qp����4��?{�A���?�O��?�u����ɩ1��+�/�5�z����?�Ǎ7>�?x�W���V3nD��G�D�=�XBY�w�����7�}m/�g�ޡ*���������w�$��JՊ*(���"g
�9㜙R��U�s�W�;`����C��]Nv�����Lm����'�Ǿk|Ͼ���k#j�<��b5��k���=������0��g߾,/��y�j��7C*|�be$Ƙ��s��j��8��K���j �Lc���C)"�^q��X�H}]2@/�Ud?;Lx���!�tV�'q�/�Z�L�I
Ƭ��ʖ�IDU~�*3t��Ʈ3=�~�x�����w�[}m��:�ɱ��e�i=���M����e٫0sN�B���$4l� �mJBrƜ�Hca"u��V�*���´�o�4H��2T�����=шrAr��#���<j{'U����*���B��8]���iw����[�4rc���(�JB^�	�Sob��>�#	��`&	L��T&-����T�4���m�{caY���!>D�n��(x��9�|3��ir��QDK����MLO�+J�B��C�V�� %@9��P1Cak#9�ϡ�R7{i^��υ7�Ԗ6"J,Y;��q�	:Į{��Sȍ� ��2���eF;Ru����v۠�ͫSF4�)�*�^�@/��#�0^q�O�]ZG<���3'q��������z��8n��1X[�������M�'�q��b�1t�1\ZZC������RZu
�DD���z���W/�]����U���c�a9���O�pE���'����ǲGY���8���f-�,$�l�&�72Y�0��uO��*BCX(�i9�q�~o�̱���^2�L��B��ۋ�;��{��g8<�����=M�Y�Q���&���b}s�/_ć?�A���vB63�����1\Z��������Dfr��j�J5��l��gQ��R�Mɡ��Ή���,�k>��Q֦����	�0l�Թ�[��*E�$���k3�흱@o�.�I!����9�(�?�9Έ��k���/_�����L��e7	"SMs';�1]+�W�.h+|���^`W��wD�k���Y�P�d�mI�*w.;��t��~��%�`ϐ��* F !eI�T��yP����ǣn�����?��ū=�jg�IG;ZށM��ر�.��y
��qם	
��1�y�R*�s�gl|�����������|�����z���N@�[oȡ�(���;�"�=���h4������N���-
R\XafE�3��m��M��;ѳ�$�K�N�(K0vp6>@#�4�̜hd݆�#�M���-a'��>x��̟���HjY.Fr\�����V�BA@�0BH%�h���1���Y��ɐ���]��"��������		�Z睭����qdψ�2k+�����٣�K��(;H�AQ�ѲR16���+W/��yiJ�vZr��m�t KHfVπX�P@8��p�܁��H	�fe��X��ҝVI:�7����\�޺��f�ɃO��D�0�[�������JD�y,]a�F��3.o��v��2o:�ů��e�'C8~p�y���/��f����L���O�wމB��7����џx.�T��~|����G��"a�T�[)�é�P\��TU�,m�X�B�c��'����T�,���A��-���)[C}}s����Щ(��R[ ��0�#	n�"(��Hl0�E�$u<�й��<'���Yu!-�[X��!�n�[�B��������H��H'�S|����{��|��w�?�_��8�t��y�韾w�y�t�]���l�q�����w�#ʝ��{U)5z�&`�)З�����0x�z���]�j�~��1g�� ��c�I��HX�[��+�Z���'��|�lf8��cdՌ�C�+����R� zC��,�1�����:L�	b�U7��6 �qvt�C�q��y���W�������;t	ϙ�H��������ar@�T����g;�UW����Z��`���]�:��&�Lp/_į�6�'�}�D��u7��̒?��`O_�Q����=��+�d��*�Ρ��$G�����_������~���oӡ�����!��͍��{X�`�ܓ4�M$�DI{6%˾U�u���?���vV���^��8t.J��H!p:�$.Kh�lX1F����N��c�����;t+�������Ƣ8��&U�����P��4�+:g��	֛߿O���l
�t�.�w@"�7	aܼ��r����
��Aܨ���g�&�p2��:-$v6ǹxj����"����.��Z�,�ّ�Xe6fm9O^�jB�H���n�P@�"\�pF���s�>r���YBp#�R4LpX�@y�*\ϭ��U��0����Q��`��{�ʧ�g�uBf�L{-�]ǋ_�#x��'��O�{Ν~5]�^��#G����.��7�In�[H���]�<�b��@<�V7��#���
�V��(���i�6�]�0�Aǰ4�|�����֚U])n�ډ��U�`�N�N<)R����JE(l� �c�G�nG�'��g&��;_r�#1@�ϟ������w�$�a`?�VU�"��ƣo܋����G�_ř��Em���HA�ว>�������g?��p�whݖ+u�|�,�	�����?�K���3�Oc���X-هk��k�C�-ΖȎ��4����VR��3=$�I\[��ŁO],�������D�+`�����!�Q�J'W-#��J�"�G$�$B����OO�S������u�m�������k���
w���z�zV;�w�F��    IDAT�.�	�H�Z�/0Ti51v��v�}fc���xJ	�t'ȿ6<+ �>�x��!N�T�5?l��N��:�`�_�Ml��t�ՠ�i7v���?o?� .K�,aF8ZJQ*f�D�9��C���zŻ���{�.�V���/��P��;t�}����Ә�8�f�,��c��,�
�W���rԑu ���<La��n����Y6�%nf�h8t�wh���i�#48��h��EFCq����=e�K+hT�W�F� �K����L�X��`Vd�Y�x
�R��.[#k7�qE�Ź���4̐]�=(�_�=IeX�%j}rr�hDz����| �F�tJ#t�Xc�D#A�gW��(��Fa_Ic<���kND���^�2��m"��(hX�z��@r��hs�:�l$�c�������4��`pg�;fCt�T�J&�H�Ө��fb�LpC���s�E����Y��h�"�k��=4Zu$�a�6���g=����D�����g��2�\�{�㕯�5��7����W�A�C?�E:?+��F�$FCI��u4��HnLtiu	�0�5i]YJ�5שԑͩ��ufM���Jg�

�65e�R��=��`ԡ��y�TR�$�<lup��"E�Ö�A^�d�Dctj���Aއޡ/)����M@����]������Qڬ���F�	4�}�{q��C���+¨��U�|�}�~ի��]�|�e<��߇�����7_�F|�k�B(5���,Z������k�����9u�lLk������u{v�(��h���gj1q�"d��y)3`6nBy>��ջ�Va��?� ���5b����w�6^�؅��M�g���	��5���s����ʁK�v�����_��k׉��ۃ*�s���)&UY�F,�#���@��aq�����TU�$�ې�y|�O2E�M����g��$�� 9����^��PE���<��A���{AvY9t���ǯ�z�����9��[�NB�Lq�����D�A��C2��h��BW��0�*+*ǳ�a��;%e���8v��5�zT��� ?�R�4���]	[�%��
�Jh�md�l$��z�h]�$h�҂�����e�4��ӡ��G�1���N��o�pkk���8?��V���}�c8ޡ�Z��S���`.6�WOL�펀#�W.?u�Y[G����r�c�����Mp+
$�Y���H4��܈���%kd��\t��BΛ�:#l��6��B��$���)��h���	�4�C��������m `ee	�FMR��v �/-"�o;9��	OcQ$*�F0�E���gї������3��B&C,���>��gH��XX��J��mf�#�����ٟ�)�_��hr�^�d�	�U0�@��@|u�N�����\YP��l7�vTr���'��{�t�L���͐��X��CH�
���ɹ�����/gbټ��/(�L�l4}�߲VH<3���~I��)�F��P�O�� U�Tݴv�ٓ��RB�R@<��co�����a��|�˟�m�� ��<uZBKB�PQka��y\]�*���48� <s�p��K�/��<�-�"62���[��9P���5e�k%_e�&�U�0���^_�_2é������3bX�`�����+,�Wf5F�V���!� ��/� 	�U+Hg3:~������y����Ys��X�ݥy��f��=�UI�,-(������z���1������v������:,������b�/���=	��c���9Q�ׄ�ɍ��S����I��6���aŎ� �4���Vu>�c�y�й��V�ů��)�1h���J�UL��Z�2�@c�_��N��@��n����6��ʦ��t�d������ֺ�{�B��ZHe�h4�aY��K.l�=2S(Mc�z][Z�Nw;t��͞sHY �x�;��p@:I����#$(��>_(�~��q�'D9�6��+B�sY��� ��H���T,.f�H�Ξ��lj���8p����C����F��DO1�6��]��\%�nW:�t�s���3��|NƉ $��:K ��
 ����p+�K⾞���7��,�	�p.W�4�^�����o�;�%OhT���%�OED���/c�h<�:�ǒ�9%�jM�W����;�jD��C��F�PC�T�'K�9�E#���dy;���X��6�+��[ Das�*"�>ҩ���r����� �&&T�__�T�[X[s�]@";�XzD
k��H� ��N�9?;���itQ*U� г�F7h��JYř������Q�P�
�0�K%Q��)��9�F�)U(�	u����}=��%��m}�V�!���9�߲%��bȪYmf0���;9�~�!�  !lW���k����!,_:�#�g11�C��-r�Lv�Jӳ3��(�
�N^^^��c7�2w�؍X�(�g�/����	br�0�+5��Y����[���n�>�T;�^��֨e�lu9�����8ȃ&�� �/R&��)��1G+���ǂ�O�8�C�*R���'#C�i�s=��n��;�A|�4���`=��ϥ{B_*̧��S��}���n���;\T��ip^V�.�kּaE<'�1�K�3p-gI%>,���T�V126��^k7��~bE.��63~�Dª�������Rf�vF6e�_�1q9�Q�\����:m2�[$}�Ρ���Я��+/�������y:� �,�&3�rw�%w:�4�e���.���y<����������T���̭���.%��k^;ݔ���de���ȧXX&�hI2G	��i0����pVV091�����i��o�Dvd��PmVhH�� 6���|7AR�~[$:�cB�Ǣ=���'�?4�|�q��Ξ��h1���� BD��2��i�-�1|i7` 5n ��D
\Œ$Q��iJ�~��YDH�CTf�F��)Qn�//���*�g��u8����U<����vͺ�c��etl�O4̤።�ha��A#f�e.�j�x�	t�1�t2!�lL%�yQ-�tkx�+~������'�����Q��Q��Q)7�1`
�d3ds���Y�v!��9 �^�D�:v�.��=Y_]r�Kcj��=�ML������1I^���
?&~�j��^?� :X޶��X	V8�Z5��İ��",�)JA�'���w,���W�.��g�2�]�N���!�&�i���,I�,� ���q]��"�F��
��z�Թ�rSwە���8ǡz�m�����8�u:�~��7�C�QB�R����6��S{�&�}a�\
Kˋڧ=�9�ǰo��^��l~����latf�jݴ�w>;��g�
Jve�b�cO����8�>���^)Hlh���t��"�4�JJ�W���8�3>~ԓ��7tDq��j����!ft@�FK��� �X�ұ������yۈ�#��X��O'h���Z��)C�����u�������P�ٵc�|v��7K��j�~#�aPG "���~`��`"ߛ���
��'K'�h�T�jQxOMLK.U�t���
m��Gdi<������1�6lM�������cŒ�A����jď'���gt�x�W��3��U����.B��8�VWWus9%�ᮔ���06�Ư���@���m��o~N>x�����vT�i*���FV4:ol�˿<��a�8����ʑ�A"���Y���1Ұҡ�m�)�ZU�K�x����x��XY������"=���Q�(!�/.�:35-#��E�\��o����.�Q�:�_��?,�	����	�p��9LN�!Ƭ��79􀜥	�Yt�R>�4�Bcξ1#�RY`4q�G"cb��3@��d*�T����f�'�����O�p��R���&�lT����h�4KYF�a�U,OONM-o4�x:��	�_,Ir��]�]A!�p
�x\��7j[h6
���y*~�E��ѫ�������>�` ���m�Ci�����L �A#�����QB{1�fI��t~�~�A�Kkx�����X�Xŗ��%�>s�zc��a����Z�\_���#7(HZ�\C����$���d�3�u>Xu�3���I%�~5K�6ry�؍r�w4"��Z!t�M���!�J��siLNO�u�V�Ʊ�0ׯ�i�:����L�F<����:��:�9��G��P�`�~�I��A�q��r@���$��F��v����G��T�ۮ�	��1?>���Ƹ�m�T�2�[ő��F:t��:|�,, �̢�`}e���գ�*�dK�$�r0î���ֵ"\_ܘ*� b+�� N���>���ſ�(_$���G�Hj��ڽ�f�x��[����}��K�<��O�w?�ɸ�S�Ĺ��wO����I��@���+B�7¬e8���!l%�������N%wv�fW�6�l/k�$����|�ʜ�yԂlR�F�`��J���:�	��=�@����x�)nT��s���Q�C-�����3�ҝ���6��]@b�$O��?���`���(���1�df�t@�G�8:����_y�]��F��o�{R���D:��d&G�<�8��d��7p�cn�/����j��G>|/���!C�G�C�n�)�˺T'#��ކh�D�W/0��k- ���Ƥ`��qRi�E]F���D����IbСzP��$��^�����ш�'?u�W�C ��2�t4*�K�h68��Uk���s���8��������ɧ ��7�7��=���o��~r4�d.�H�FY:���4�;�L�{h�ے&\�tQ���"�I�Y.��py�F���Q-�c,�@asScyĢAT��hTʒ*���x�S��o��u��iسb�H�a��i�j����5��*c�i�<-�s��b����me��TSӳHR�Ԥ�
$�Ȍ"5���{�PR�L�N�^���������W��GƧ?�Y�j��ST��z�t��#c2D�r�J�t@Aε�+7���D��P����r���#�����w~ �y��Ui"?��P�&P�Xߔ-�C����'������x��Q�UNbS\�M�^�T�z=YY�.��vAkF(j7��RYJg���p8�b���1�VW֔���Oc���\<n@.�s9P��F�I��Wߣc�.Z�IB*�Q�D��jU�Z2��l�"�a'4�E&F@h��Fժ����C�'��"�����o�E�A!�6�ɘ�}gǂC�7�@5����Z*Ԇ4-���s�I\��Ø��(�笳��w��!U�c� h�/	糰���''���L���Ds�#��� ��Q#!��^����p�T�w�4R���*`����7ï���"�6��׿�M8y�%��qQ[<l!5G��#)�O�A?~e�C��V�����z�����)kM�P�A�����(�i5�XB�s��ن���$��lc9r:r5B66nƵ���q�O��Hp(���q�� �lu���M�$�����s<�5WVE��lc��
D��ӁU�J��x��d�H��Ɓ#�˞6Ŝ�	^Y5BՎ���bȩ�o��$3:�~�e����z�]/����߬��{h؂����#f�q.O��%ߤpK�l������O8������w����A*3�N��rs�*�Q;�9tƹ���M� nS	'�v��p��{��F����͡3S�j��a��-�5�a8�H�y.p�m�>e:�����s��	����?�E|��_C�F�Ʀo�\k�k"A���P�R*h��%����"��^�\<�_�ʃ�؝�Ǚ3W����o��� d�e�����<�Hy=�4�D��Q�[���(�I��om����~7�4��"]L�&��
�KhP��F���c���C'%�Q-�Y)GK'��X�=�I�04������D�i�e/6
cmcSN�iO&���'����-�t��ø���#��}�V����f+ !��:�;����������Y���8p�j[�j��$�o0� �|�z�D�;�6��>��[2^�(Юl����x�O<��E���~�^���"�cs'G��Y�v�d~ǎ���@���"7��4z\tZtL2vΨш������������˹t>ó�
3�\W~,�[�σ���HD���cf�c�ɴ�M� �r���]��?[��2o�l6t�t�|.:��9X:/���l}6⍟�<���N^}~b��H�5σχF���k�Le"�Ϡ��U��_t8���1gF��5�	��瑠#fK��2o�`�F ��$ێǂՠHH�IVQ(X��`P��fP���|���e�7V|��mU��ٌȔ��+�����\G	r1x=�.��t��Z[Z����R���Oi����ħ>y7���m^P�������ࣈDSU��\�蘭��{����[������(��ē�?�'��a�D���` K,I��)��X�`���U�V<�l7N�ͺ�7����Hyj�L�A��a/ %�n�qe�N� �b����H�`�UAU��G�!8��F&�R�>��\C~4zǙ�`OA�5l���<n(EP�u*���~?�w���K�vf�5t�ʚH��lˡ3��7$����t�@8�G��ūHf�Q���Ɓ@R@*u@��J��hH��e�TN�L���`P��ze`�.�����F]�4PD�"fZ~�E��F�0���	�C���	$�!uK�>�Ͷ1��*�񵺼�J� ��*g���X	i���#I\�zJ�2V �u�}�(T�����#2x,�R�ݰ6Fp R�``p9�\��bG
�c���;{�<��*F3cȧhV6�on���
P~s4���e0�K����?��7�����ѣ��&G�Fq��93�n��K�,���*:tf)T�c��$"��?y�)����O`nϼ��/.o�o��Q�:�y��Ez�����+W/b��C(TJHdrHgG�ੇ�er#j�P��e9��,��V�c%�AڹO6��C�0=�����$�A
�������l�k�9 D��m�np������F<LtG3��(՘u��ƚDvQ��X�eڑQ95�Կ��l���c�u���Ҳt0<3)j�=d����q|��N�N������i�	�c͕��P,��Ӱ�j]���ɾ�S���Ͽ�g�>{F���(��
`��h/h�©�����BF�A���)I�3x~���d@��1�;�8.�38S�j�~[g*��r�aF$ȉ������oasՊ}F�A6��S�S���-HYY^9T1p9
������=eV���p��/^[�^G��uW���=e+�mN��./"?��/��K��'>���_���4._a�G��7i�ޮ��7�B�uL�VO<�G錋�:h-�@O��^=����Ȏ�����ϝ�q0���]YZ��f;�NY��AV4�:.χA���L�	�~_��}UE�����6�Av�e�bxt
�:c�L��;﯂MW�,�6M�	|̩���1�5x�]��V]�Wg�i;<�ߟ���K��ޏg�{7�5�'E�8s��]��@�}뻿��{�.��މ�0F�"`O:�}��²I|j���A�:",�N��h���I��Ud).. {RF'��y�'Gj���?�P��5�&y���,�i!B�rfs��N<f�T���������n�,���8��JV�#k��9B�	�m��6RؑLVי�G��0#f�;39���q����e�\������d6���#��()���9*����{b���ˋKȥ�⏟�����&6ַ1��#�02�B���ᇟ�,�WA6��X:��&�g&�t���Ŀ����u�o���r�ܸ�\_���ЕU��9��ژJ�YU0���8�|�-���$f�����X\�Ɓ�Ɲ��&N�_A �@�~�d��8��	J�R�'���e�Ҭ�ם����ᥪ�ט�-��E�C�h�cv��N!��7߄�o�����g>�9��߾��(�g������ul��㦛n����&��ԑ�P)nH7����v@�    IDATAekq@�i2� x��'��:::���K45�''-�#xM�mD��F��D\A+�u����݂��q����fY�_U����A�OG�g��}iX#WN膙1������>���{	H� C�^�����ê��
��T��c�SA��LCW�\|K�X��c	
[ֺ"������-_` �̝�,�Y��2Qϭ.R��ew����k�sT�`D�Y9�>3���F��i�+Xq���6�
�Y�X���� ������r0d��m=7����Ѭ"�d֞i��:�S����!! ����I��m -@ҿ4�A����Mt��-�G  �J�$���Bì��U�+�.�+�����(�ط���Y�ZI��pU(�\�����m�E�INJ>�Ϥ�R�v߽�g2E�{DN��<��F�F���HZ&��g2�cŁ����9l��h�ī��Pd=aK���+�$�r�n��>�c0��"��6�%M3	��GP��~?�����K�9��f7>˒{�g:�#*[СK�K���I��A&I�@GM��v�f�sL�*�(��'@���q��j{���M7fG��զ���鶐�r��Ju͎9tF�~�+����9'��hhY��d"&b.4��P-�
(3�v�a��f:��A� W�抹���ݳ�c���T����v��N7��߂ѩ1�n���o!�`������;to,��V��Fr
+IWʌ�^kanf���1*u%�(o^�H*�~�$��T2�=3��x�Μ�_-�7����g~t=��"wf-/^'9�%Etx���AVk#�V����m|�3����x�R�l-đ�<�v($��g�n����z��~����6g$I��(*պ���?��"\i����a�*�"��5�*fk�n`z,/��T{�C�Ʀf���)m\θ77�G"��-7Ʒ��,�������,Q��ie�BQ����f>lA���ec�S%�4K�t�t�tD�Cp]13��#S������x�S����{�������ku1��ґ���4��GOc�yʽ�亥�T�ա�5����L'E���H��~�8��r�<<���_x�jј�V:�P��c��ŵ����D^D¦hTƓ{��b��5:c���г�5��?�s���#{�F��t&�Fr(d�f�Ɲ��y�N��������P����M�3w�xY&�ؕk�N\ ���z�4IزI"y�1N���P�}#��5)�M�oT����}��XV����
rĴ��6�?����`p/r}�9�	�	�#v����6�E��-h_k��4
x]
H�\��P�pt�_����U�vf�S�'>�����x|�Љ���9��歖)k��
+����F�Y�	�,-�YǂL&�%�j%�jɻ_f�bf�>���ɉ�#&gHH���h��s��y{�Š�1�iA��(cq���N>�b������O�{~�7���RO����Y[X"�'K{�6�2\���ED��Q�A��YN3P�Z$1F��TDC�Q�mayeA�x#�IT�e�HTh"� "��fۀ>�ye�-�6=#Q�4��!��y�JDc�s�Zht�ʄ�	�Cύ�w�[2��d�L�FXFӁ/h��
�2#����%҈��hD�ݲ|h]��1��ǵ����2VWV$C0�޽{����J�*�NF�p��x��t�����!�o 	�^)li��S�6kX_[�A��&�����
���}�l�СC�����2�*�:��Y���a<p�{��?�r'�Y�5qaa����Ma��E<=�>��������5T�e!�X!�B,np9��0S)�9��!̀h�0jTό�TGxA0:H�O_�@:�,�֌O͠\oav�i`Ӡ�*E���<[����o0�]+(Ü�߃K��Cn-�lnn�P������L���rt�r|�l���7j2X����
��J����S�N���L����t4,�K����y����?ao�t���9�~zļ/�������O�&'.�1^3(��v%g���^�����J�絝s�=k�#βԲ����q2�1�m�u��' c�d����J�l�I�̕�`ӯ���v���'�MVA,;m�I
�I�[7�!�Y'�ʙi2D!1AM�(�LR,	q��X�JU�6��t궎я�Y'�>�ӈD9?E�����	��+" �"'}%.��H1����S���N{ů=���6)���ET4�e�)�k?���������g��H �q��J"ۤ�>����5�@�*���~����)�pRI�:
Z��qN���5Ե�hPʗ�F�x�3����"�7���z膢h�60�FwĮ�dk���ޡ[��KW�/ �2i�}^�:���/���ګ���t�d�Kui�FDe�z�*���r,37F���i����,Z�rA�;>�W��7�'�+)ժȤ���tJɧ06�r�Z�d�h�NQ�c�Is�ѡsp4��%q!x.pC�w����c��ca��2pISV�ȍ�q|�4�5P?#~"����C�]�ͧ�C��d���.&f�"�����"&f�hv���Zʮ�2�Iұ�������{����ss�2��Z��S��ۏ@��^��#'�/�1�K$��sI�z�>왙R�J�����͚I����oq^����Q�:�k`���:n�a��9h:�����|&n��(���ON+�������F_��9lT�hv�$�B�@ґ����F��Qb�@�9jA�G�*v��e��3	�����N������������
�-,� �Ψ|ǌbuy�`#����O��s������X �&I`8aQF����z�!fA��H�1` �R���-�R��q�^����}&�K����\����%
\��Y�v�B:���;t>K��q2�f��ߥ��A՗aeQ�,&ty�J�^^t}��<�[dU�/^�����%Z��X}٘��ǀ��~�#�eʋ܇<^6m�BVט}ҹP�p�Z�M������-G�����������T�Α"�,/k?+�i��"+c�:���#�s��!������-a 8�s�(p��pO(�����af�ܻ�ֵ[}e�M���1�4��  �k)�H����)��X�c`���X� �@�c�gϝ�h>��ft$�{�
���F�ϟmH��"���6�iˀ�LV2��	s���Zѽɤ�X����1�M�!^�/ի����j��@_$�i>�Q��*���|6��1T[����ai}�%T�=�Cq�
��F�+O��G�����Ǣ�����^ ����p^�%w:����/�̷έ��ՏMR�:�nɡǍ0�Э�ʞ[B�w�;U�m����8�Nm%��E������T�"maf*�������4���O��O|��2�0��E�]=�v���a"�K劜�"�^W�D�ڙIV�F%���hG��; yWfC�B���(��:_f^�I�R��ei\it�2��eYR�*"[I��c�����<Z�h ���%!S�ݫd\��6��<�����-f|�sӸz�����޷g��u�7��߂�W����ͯ	���F�)TJ[�g�HD��6�����g��]w�����^��3�HH��IOz��6*78���@>K��	|ޏ����{�7u^$T	��H��E03���]Xܬ�ѥhKl��(Ƒ�Vd��6���G�	�9��p���V鮧)R������mS�<��L�a�ZMR��Ȕ�epBn}+��'h�%խ��q̎�P�^ƕ3 ���v7��#�%^��2{}4�\/t��F�H��Ñ#G�;���yNt����ǹ�i�����,Z���5A�L�˯<��-Q�p��c�T#މ�������2�qX�����g�2+�`���w�7����ٳ�N�3e.��F��x��2���j;�����'��儕��g �2�;�/�	�3����<0����[�;O 9v+N��L�r��q��<ٻ?q�� �%<�F�ػ��X,z�L�V[��?[�9�{��l��1s������޶�=��pŦ�%̔�=fCH��Ns|�@���)3��u��+��\MP�)� �-�:�Ϗ?��ǎ�s���$��,yox��1Uo4{o���Np�\�[[�x��e����:{��J�Ƞ���J�V��xJ����5�|��
j.\� ��u�f[�J�V���߻D(��Ozʓ�y~ˋ+����E�i�G��D8NQ�>�<��Z�nФN9�ħ�Uz'�;�;��9?��*C���;ؔt���.Aqt���_��{/m��ՏNԫuD:�o&(�e���W�� ISiv��s���{���蘘��ЉZ��7���}T�6^�K?�G߾�mO�y���)��M�1�c��(�կgdF0RV���J�dts��<���T�"�#���M#BBjW�Tx�c�Ź���cGo�F3�VTJ���X�H�Fpey�h
+%����P"���5ē��\\F�!���U5�D�ZI��3�E�8��C���؎�� ����U׮ �cf"�Fyc#)�V5!G��������s�p��G-���7#�]t�g������w���|�p#S.��c$�w ���IJ�����]*!����za�ޒ%��j;-�8�M��c-�=ҡ�g�r_Ia*��Bs�,=��U��1�Hg�sa�ǗR�ݒ-!������*R�B���O���~���&GP�\D�]ӱyݬTИ1��⋆���h��Ј��W@K#��ʿQթ�н��"��ip�=�>��fS9lo��%�s �%ׄ�h�=�l���oEX�c{f1���K��<�Q�
���g|v����p��������vog����4B���$��xQ�"W�"T���)	-	M �J%��F��v��N����z���x��gý��e=�~��k�5�;����~�wX��x<D �9���t�bXk3;k�#���\�z��)*�̜��V<C�jٌ<}�����s�W���[@์�1�b�;QY`3#`�tM�8؏1��B�q;/�G��½��/��	�Y��iP���Ҷ>��W���X,���!_O�q��j{��VIЂ������2���o���C�-"@d����k�ڹs��禔�RNh<�R�bF���ujꔶNn1Âuπ�[p^�C�?�yŋ}�}��/���=3�c*2���|8��uLS-B�̳����1�����v:6?�^�'=����[���n�m#��/�H��������g<�6�(���a�� ��ظOd���=��e��[R�ЯZ'�b����K}����PNG`>��%���Ө:_" � d��Q��3^������O�����������[��0��d�e�i�b�-n��Q�ƆE	ĺA��}�:AoU��L�2�Ԭ�!�5ޭP�6X���#O?�������W>G��t��u�_�����4Z�ie�`���Q����pf��83?�=	�d�N=�B�0
A}�%kz��-���˿4/�XLi��c�@�	��C���|�a^,�x.k]��[��ܥ��P+A����E�L���oF%�a����o�:Ҽ��:��H�6��- z�1D��N}U��Ym+i�hA��R���E�:�-/�;o���)]t�j5���x�_g#�qٔ4�ٱ�L�"��{Bcc��# 6�_Q������6>2���jviM�dA���z�����j� �	��i����雲�F(٠nC���?Fi�6�@;��P�����f�G2[[`����H%D���V��p±xWՕE���]���_��Y���F�Z^8ed<̳�Dve�>B��1���OS�ҵ+e@�?ak�9���ȉ�<T����d�ǇF�ϕ*Q/!B��<�6��x�s\��Ɯ��F4D}(��A�D�F$Q�9 ����-w�H��/sD�By�c����f0�hjt�����[�)����PN9<� Q�Ŕ�Q��M��_Y1�bLs�*��N�<8)<��쨑�GP�e���v#��-�a7�^�� '� n�wx^x��a(�-e��`(eꑫ��J�b	{�@()������0}*ZY]��:�#B#�,`�.z͈� ����zc�QVǽ�Nx^��shF^*�x��7�0��1`|�<g��5kCLH��A6�;Z7I�x����Am��ʊ�߯J�qy�l�������t��I���h��
#��<htxX}���y��(~�����P�þ3�1Y�?��l���ҀNL�+��h��T�0��fG�ʈڤ�t�LY�#ߌB�(Qgm�]�#�R@؄�$������S��'�B�l�_��-(�N7;��^U
j�H�S��
ݐ�P��ZV
8(�`[ӻ@-h����= t	a^9p"�R!8���/9�Bn���k^0݌r����I��S�:�n�fau<�D/b9Da��Y�Bf� �BӅ����(ݫ^����׃>h
뵯}�	��o��ʽM=��z��.�P�Yg��s;=OLj��J#����:5��FF"mM54��A
T�!�o%!��؉X�[Q"f^��a)t�����u������:�8���*�`cj��$�������wߥ���U�R���n���cx�^d����͓2�M���U������NNY��/_��:묳t��س���Uс��:2�n
}f���NR�k �ǵ4;����%�����O+t�;��3o�{�S���cǛ'd�y��G��?B#�������Y[Q!�S9+m�S�[�cޣ��NU��fB��9c	������M�!�X!2�����Q���V���P噝����@���8��!�+5Mp��9?�^���w�I��?�&���!hzt@Bńd*���������1�y+`X�u����w��!�d��m��w�!Ӏ��`$3f�Y5����r��-56:l^)��O��TJ'N��j����ޢ��pM��"K<��p�{E)0n�~�cu�h�{�ʕxR#���]שּׁ��d�%FF!~�۸0�x(Y�E�� #��X�R���X� ��⼭%z8`�k�-Z^�ZU����|�����ذ&\9�����PC��� /��Ȋc5XϬ���9�m;l�<��!�s��Uu�A��߳�3V6K�8ꛭ�ur�S�7g�H	���Y*�"3�J��ȸ��W���ِ�c�!,�����F�0:��ђk_\ԙg�m��z�.�*]�S�IBA������Z�O3)�Ri�9�5�4G٩Y�V~Y��H��~Z�O�ܩ�ِn@�=�:!�~�7?ph�]�^f� ;䊪uK6S'��jo<��
0��E����))�������t��Ŭ��Pv��Su}Y[�hyiJ�R�z\��U�-���Km-hy��N���!�X�t>��F;X�lV�9���uJD��c�����v��fsaa~�Ƀeaq��-��=b��_t��������/U+��R=��|��Z���W����Q�l�l�.-��agh(���)46��l��/��ưu��	k�b��DW�d[�|�.����-�y��z�EOQ�YU�N/��)��ڪ���gt˭7kue�j�/���p
��w���ԋ.����;�zр�Nؽ=|�rg�|�+-���C���@����gj����~�n�����Ik��1R��Ҫ	lT���n� ������g��Q��u��jo)�i���� xOЪs��J�Q���eC9XV�C��{�c4�X�W1S���s��jyxL[ǆT]�Q�B�C����􋟮�?��f�=z�*�(��{�~S.¦�l-�#T��2��(Ϲ�fS�|#���9zI��&�P �~����u�=\�<!��r�3a�z�l�=�+�ّ��e0ŗ���̴�f�-� E�1��\rI �)����o��>9���1��P���3r���QH�-Z]3��FS.0�ues����V��3o|����/�0�0�� ��I�C�����t�O��n�lN�7~Þ#�t��O.�a`��L!}�;��ԉ�5��Bh4��W�J/x��ۜ�w��"���1���k�S����fG4�M3t    IDAT������Ę�9jF���$�6���:��}��_��͡���]3�׽�uz�s�c�u��?��%�i��뮻ΎaK0>/	|���ik�cQ��sf�2����{}���g��r.�.c�Ї>d���x�qV�yj�/��7 ���q<���_�N{n�=�x���hԮ3�����3���旭1T:W�&Z$�(]#��ƩL��>�9������Y�1�,i>���IC�SR�$-n<�.�xR)�c�^p��>tp��-eGjkU�5�k�Щ�<u�ա3Al0��)�N@'{��� X���ڭ�T�p���fU��3$�(aɃg��W��M%4PHh�HE��h��5����M��"B�J#����y��r��ow��/��+L��;�� lm�|�W�^�E]x�E���}�h�y��y��ʗ���r#�k��QO�S��-�["�Fh�@^ A%b�P{	C�Y����*a�86�����%�A)M3��K��{*��ڱ�O}EBH1�:qX�<�����=��C٠��g_t������،�w�6����{�'6P�h�533��;δ9����c �X�i�Фv������TUN�x���[��&'�(���m]�֛X�t"(DL �	�.�n�xd����K��!�ijf�����:�|vnYtQ��WØ��)!-B�Q�먱��.��꫺���9vP�'k���V� 1���<3�H�z ��Ba3O|F3��i�>�k�.��o|�	#s����yG�&��Ю��U�#WĚ�wK��sα��(B]7�L���dp�������=��ݜ���rqO̄��+k��[~���� A�}���i�m���>n^��Q�8z�� D���;���|e#��%Ng�}����wY�ɯ����֘�����|D7�x������܄�u��/�>����{,���2�d,m���o����:k�%t�K^��#��Q`n\�nvt��3��ꫯ�=w���(�F���^��ٟ�y�o����A�3���������b��V���)��U��]f�``���,+��v��aڶ�/��=t��k^�]u�U��s͉�m]����կ~�F�:s�G������7�)�Y�4�u�I�׽�+�Z�͉���=�y�^��W����;��9�o��}�oZT��c"�#���|�~���i}0aB�+Dɚf�\y�5;3���Q=��'Z�6ԍ%�A�J��Re�HǨ��u[����|�SOf��ik*B���ݦC$\(��ɓn2�\�h��I�C7���o�C������
=�l��B�:u|C� JD�o�<�ytyh����u:�S����͚:��r�'��� ��n(_Ω٢߲r��PuaZ�3'�T�������BlxfdD�=� 0C���Q��������:��sM��(k�5S脾٘ ^��Y��w��?n�sL�2�镦:ɲ���֝�Wߖ�j���dT��r>�[�B��E�M�ȅ|��5�k�(��r3�S��Y����1���+��k*�����RVՕ%�8zH�S�y���<���\��%U��j6'��c��~:`�3��/^�fӄR:I�*���{��?]�����#�+�����<�UGNNi�o�Z���4��UX� �H������H�z1�S�K���Z���45}L}%���ȑc�;_]�9�����I���D��,��u������$^��	�c-]x�6�����wjJ�V�*����n0�>ք����y{�[�bQ
��ں����}�몫ޤ�'O)�H���:j�Q���a�y��[��ZU��T!�����?�i+�#7O/�_��J��7���z�ޠ�����w{�_:ү}�k������,��;X����^����'��@�^��8�ܳ���o�Zb� �SǞ�u��G?�QC�=v���Ĩ��'>�	�}��A�H*nƝu�IM,i����ϑ�f.�g_��͓�%Q+{���n��VS���?~�պ��7���uB�/}�K���>g��L��7�]��]ܪ�)�����6�q��¢�4���^����ր�SR�N��(D�n|��7�Y��Ϟ{����կ�����r�J�``n0ެ�d"f4�o�ݫt���-�Z���|���_���x���IA8�s���y1Nx��u��-s��g<�Y��?�S���D�o�q��g���[��V3B9��ɍX���q�o&(�����o>`�Ǻ6*Z��_�"]���C���Zo��Tħ>�):x̺0"oZ=��EM��kfnA�bIM�"�:x�_ԥb��LY��p|�*^��\P�F�00k:�W��gﳇ�O*��u��ᡣ��i);�B'�΢*�Boa~�Ѝ$�M�4��C���XF-t3�����֤y�tOkQ��$�Z_�Y�uHX��V��':�+g�QS[+Z�=��G��aK $[��MGÂ���+�՗[)�5�5���k��_�+��e�]�m[&u�?ҥO�8t_��6%C�F�Bx�<;�m|b"����ߩ����oߦ���
�jǳƊF1��Q�vB�+K,W:�u�R!�B���`��A��T;���um�ܪ��ұ�)�K��C��oѱ#�͠�2>�Ǐؼ��Vt�]wjz�)���[&���$.��\����F�{��2�-[��+㡑D���0�ȡ�vg�}���A�.A3����Gz���b�>�W֠���ؘ�ͮҹ�m(�7Vk'jѴ�;F�I�R'fy:�~�ƚVVgu�S����v��l�n��a}�K7jy��N;��jC�gl32
��Q��wr[�F����)��k��h�ݖʙ*B8o�:YZc��������/6�F����y��wgax���4�׿�uz�k_g�Q��/.�[��@���˿�����SS�A1����o�/��/Xn�2�?�0o�[o�M�_w����L�ODg���������<Sc"�@iXJ������=�t�M����Ͼ�K�袋x�@)_0J[������t�-��3����k�7�@!�YC�z�զ(����xY���q�v�w���t�]wm��Hϐ��'Ș7"<�����w�k�ɮ ����^����/j'�1�#��;!w"rD3�S������I�_�)�L��Z�àg�
�@{�fx�k+v<lr�����7���}���\w2`H0va*���ݪѶ7��0��W)��α�$J�5Z�0�`��O�{gx�I�ƃ�ʱ<3��^!�W��xn�!�b���q�Gk���}�ȏ��E�)&���(S�eX; N~C��3n`Ң�AS�ҕ��v�ܥ��?a)�uk$�0��x6c�g�B�
d-��	��Ǖʕ�y/�����ܭ����)t ����N����������w�z���Z�Wi��TO�8�DM�R�R7V��I,�$g��)��ܪ��\W*�Q1W>�6�"=�!h�t��	k�23?�����T�imԩÇt��~�i�amk���⥬l�K�k��Uo� ��Vh�:��җ\a��v���g�aBp��Q{m�%�k֨RɮQ����Ȩ�}Ú[k�7߭��]Z�������)D�0ɘʕ�:I��b���ۤ���Jێ=j��!s�RΗT!��n(�ZU����^��Z_�S_9������.~���b5�K���>���6ʕ�����LpaH��Q$�?�ӯ���<h~�a�_2���x�v��8rƄ��Ƕ��Ǐ�4�M����ubaU��`h�Z<�� ��*���aej=��ti��6����#B �M�^]���)�����~��.�������ݨ�n�S�j�Zf�T#�lݸB��єR�6L��kjW��\_���a%�MM�:�g_r�Jٸ���cF@AHt�9dyh�\����PV�0:޽{�i߾�&�Y?0�`#m�7اm[��2P1��W2�AW=z��-��9��v?d���VLf�PN��9�bP� �@8p����{��ff��X�P<N�A���)��6�9(
�H�焭�A�f/��|�������sȓV-Ε������D&�n�@��qv���f+0�5@�G<�`p]R4��1�0��s ';e����?�\^;�3Jk{`�\ܨ8�K���YLn��'��2��]�xh�"� �#}b��r�}���FGH�93=���wX��gG'6/�[Yeo\eO��6�^�ci�M|�ND���"j� �v��e	߇�x����}[�c%��oT?�kk������&���8����� �R��0�KD�`�é�=Ǹ��r<t|ެ�(���>+��/ �}&�b! ����
xpxDO�s�������N��s��lN�g�U,�Ԡԓ�AVe����pS�R���6Gς\Q�dΪo؃O:�;��|�?ߴ���4�������� ��}�g�a$�,%������ȇP{c}]��j���+�i��NsY������kJŌ�� Iss:x��I�����*�(����GԬWmX�ԟ"��5z�,��k-b��a� �
E��VK�zֳ���߼����%��+��L��o�,s�3���	+7�*��Pk+Y�7��}=���eK�%3�VO��?�cX԰N�3�j�f1�����,֩9�7��h��Spۯkh0���!�5>T��j�\J��:� ���Sk�Kz�G�;�J���`_�!��S�-����!�U#f�;�~�2��9F<��^��U~��a��/�`D�ʠV	O��~x����^kiey]�LY�Bž9��e����"��$==l�-ct%
�ψbZF�ܟ{���W������7��;���[����X*���1�%���e�{m%y�a{u��o^��?�Z�_���ʹ����+u�]��_��}�=p����Ep������s��v4�iR������h��ɴ��Eh�	�ެ��+X�Pπ91-/.�P���O��=j�V!Z���	QD¤--,E�!u��ؽN���^`7�8'���RH�.h�T�?5��zw<+�;�f�f و�āb��X挺5j���t�`��t�� \�x��k�T�1�>�N��`(!�P��e�$˸�>���;�bqaY�#�VҴV������>�<�nG����1 @�ܗu�"�a=��1�����>���9��q@ ��T>�I����6���y�;��H�v%T2p��R���K��|/��R<�y����0﫫+F��������@R-QC����^	�/�/�/7>�>Y�Z��r�?��]�&��Б����>U�J�O"֖�Pֳt;���-X�t^�dF�L޼�.�����M�h`L�O:�o>��7�9��'�Nyl����C�,`qz�6�mjX�@�@o���I�#�P{.J��ꬮ����?�R����:���+����Z�N��?y��	YB�P9>���u�F�j��,T��@���ؔ����� ����IPT�F�O��g���LPvX����-gS�*���KIK��VK1O�P�oD���)�)�40�z��*�k{H?��e���1rcԱ��N�'%i4��$��J+ե�M�h��]�[�� ��)_H����J_V�'Gu��ǭ�<�(�I��XU������)����q:�%�.���7N�k[�,�G�������4�Ɂ��.-��#��4�_<UԹO{���LO�� ��ߪG~\��:ݤ��@�����u:f4��V�<-:e7!���q��wʌ.r�xp���ʚ�|Q}C�j��:�k)�V�J�NW�^M����T]��|�f������߹I�=t�^�����ҭ?���5P�Zl�B-7���?8��������V���B�F���!����(��,�m:ه���RWH.9�����O+K��+��:�m>��)�Pp����!Y�,	��S(���lϑ�^v��̑n\@�k5�Q�=���/r��1g�Z�P��~wc�{�㚼o��h��0rC��8�����WH��ٟ�%���h�bv��#����Z���?��_���s�<7��(�6gN������p��s�Z�o[7�uq��G@�ߪ}��	&��ĽL��טCOe���y�:�ܺA�b�F� �*�Ȑ�xVK�MEL}�:C��g�t/����ܶC�N�hϞ�Z�7�V�r5����p ���*��㮵��(�Ș@�O���R�5����N�i�z��S���Þc���VL��zP,h`�dbaj�BG��MD�Q�+%�ڱ��S��H������k��|寫R�il��B�\��R��p����he)(����K_�����F��\2Fx���`Ųa�:g�����
M(�%����R�R/ܥcYɄqXpx�놪����A�YDZ�b)((�����)�(�2�E�LޔK�[W��w*�ho[���NM�P����0����`Yw'�M���̩�<`��l���eW��<k�PA'�2 �P�����T_[R����ʲ�� F�H.�<#s���<,�GPA�S��Y��ڽ�Vk3�J�#*�G4<2�\Ͼ�ť9�MO�Q��z�g�&t5��I�"�Av������ga���O���5)c�����T�^[(fM�7��;��B��������v�W�]��s4X�����'��o����99t��<���T�:�[��.R���_W�T#�B�e,g�^��#]���q�s�+a�o���ެt6+]�S�����9hW��/��JϿ�J�C���0>�v��vcÿ���s��T���k��^} �Bd�x��u
����V>��ٱ>���Ct������(j�&>WB��z��:�a�"fR[O'�i>�6�4���C7���v.t�W7|�����݋>�Pü!;�g��U�yZ)W��S���Ai�+��Bd#�m6H=}@��71��7c"j�ΟV��.|�O���L��~�F�[�jh�3��ϱ�	��y���L�/��L��T^��;qZ�[N�n$3!�ڋ�M~���BS֖Q"W�:(�t2��S蔭�����ǎ�ࡏ�������0x�Ч��k�^��RG�1�9:?(�9�lJ�em�����/��+W�T̨� ��E��4(hk:�N�Rf��+����{d�G�If<Fm�+t������CI���Q
,�j�~&��T-b�B.X�5qiyy�L��4Mb*��Q�Z��jkeyM�^��UWB�+��${�6���8h����{����8���&�4i�Q
�[�M��	*X�������٬�fT(b�J
��GH��R1g�T1�9���S�+�u��O�~ �D�9��x���E]Rԉ�d�U��Q�hE�d�9�#�5*0vF�LMy�du��~]v��[U��G����T�%4�PS*ӧ��I�C�Z53v)�A`�3&A�qiSKIb6����FC"'�O�\�X����[��C/}�B��������N���W���b����5������_�/Whr|HǏ�z o<N��`Y]	}�]�P��!mr�s��n���@��9a�9OKSE?�=����=��^+�q/��{�(3����k�=��Q+����Y���r�h�cf|�<���ýxϣ�"q�������vD��¼�ܿ���01y?~��1� �� �b�+�X�ʂ�1���9�g�!o+��Yq��OEx�'W�f�����$t�
uC��oP%��\�����8����#s���}T�)d��ح��)��w��b?�f#�Z�l}t�c�ȍ�1��������j!E���A��+�#�
�;����x~n�����!�i��xh���n���x�����Q����/��B_ t�x&T-�ЙG�a�G�
J��	Q&s�(k#�w��^پ!+�1<6����������w�|��ڟvz}c(t5�M����8�l$)�� �h}1�Tm{��
���Z`�B�	�W�e]�kR�����ҋ�P�N�yO�D��l,��C};`ue�?����������	"���]�m���t{~9��    IDAT�I)�6���	Y�cU�M�n��t� N(Wjap��8@Q��P2Z�g	������ʐ���r�A5�I�ќ��텤z	.����03B�(���E+��@u�}�C���Y�K�+VRD�7��ۜ�
/t�X�O�xb�쬯T2�/q�N�!��4Aw }*�IE�O�k �G�s��ڔz(0��5[��M*��B|)��~���j���m}��ާ��ff{�򗾡[n٭���R�~�O�T"�����Z݆���ܬ�
o4��N��J)~xC¼�NL+��(�+��_����8
�M">�T
O�hO���~���c��{� /@п�#5z��?W�nM_�������g\�{��(-����)���Ʀ+@Sr�<���&�#�2��v�����v��:E�yHҏqo�Cś=�͆�{�ӛ#�"�Ϙ���u%잔�?���B�D+��̽��޹�>~/��{���6��H-6�<mPd!b�څBG!�³� 
�ܩj]�,*g�uh�9� ��?7�87�+���(��p���x��#3�ڹ���Sk$�w�>QA7F�'��z��l�!<=��13���z@l�͹?����ݮ���O]�=xP��P(w�+�xr���
9w�&o @r��$��G�����}M�z�HǻA�{��0z�@h�d/�CqaPUa\����b`hH��9�f~�	S��X�<��U��� ��)�!b~�'3��2R2m!���X�st�I���h�W��g�����\w�70^]o��ڂ���@���n( +�(NL�9AU蟰��U	�[k]�X[�Ы�x��;g\t=-�Ci��^$��<�,#W������ǭyc��O��N[�l�����Y�_ͅ�(t�u{�Y����*,kC��s�y��\Z]S&����ZOk����nֹ,�/���Z]�նr�e�}��$쩛�B�����n$�b 0B'1c�]�P�,|64���Y����>l�yxp@�4-(��4�ק�m�� uPsφ�Pd.l�m���Me�	��`-��M�ðG����K���B�$�TL���:9�_^�S��ߓ푄��/ܮ�~�_���R"UQe`L=H$� �6��Ž	�.���S_Y^V��T_�d°ըYY<�3S�����U�z�nM�xOM�?�г�b}����������5�ׯ����z�����_x��r�ٺ�޻491adA����� �˴���ҌD#
���Q(�T���]�B����R���+CW2?����.X��D|(t��{�\�Sq��Q��
�����. �g��{�~}�����f���{�s�{��N{-P�FԹ��m�C87���?S�Q�x�����f�sG[��n���w%�a�r��E�QK��fC������o#��xk_���"�q��y? wCh~��m�����������>�����C(۟5��S�k ��{���S>����9:�k�4�-.n�x�k�:��_�`\�׶?�$����\���9A07�vl�c��g�{����z�}Z\]W2�5�� �UQ%qa˩R3k��0�cz�<t�8�� ݳ6?O:b�Ggz��3
}��nopK��1���2��H��O-�B��`�����F;Ԩ3i,9�K��b��3�+z�k_�ɉ��L�)8
tg�|��@�,�[2�&�\s�q>�,����+�X��o�,n���A�A�4�!�ټp���(�Vt-��Ņ�Y�d��pM8�)}�QϘS�Ht����2�Q��1�detBM��؉���A�����B�l�6��\.ivf��T�$�$�1�6�-�:r��͒��t�p(u�Ž��B��u��m����
��o4�"��"��,k�2Bc43`Lf�l&gт����~��$|�+�cz����e������7���nݭ��_}��ު��@���ڼ5�1Ao��	C�w[��;�b����%ujuU��-����Ջ���1�I"����ſ�'>v���oilh�z:��?�M/|�3u���t�}?6�xx���`gk�Z5��Q�Z��0��i���b>c��J�m^ �sl�f�D�fW8�=@W�`��{��p��d�^�\�q�x>�=/�oV�.��R?�z8�kpNC!G�{dD�~V�����̕I�ЙgJ�P��q���;����a����� �2���#��Z~ώ�	ϭ�4��i�Y�\���\��s#.̩�����U,!�o)�(d��1�ޮ�=W�O��s�ȁ������'�%�5]�2.��c�k2�<���(��y��$_;~.7v�_�~�f�FUq1�UQ��=Z�*���@f�
P�t�~�yO1���ji�j
T{�Dv]�n�P:�[	��7�;G�Ǔ�C��K�e��g2O>�N����~�=v|�]�^�$
���E��B>��O+t��2��d�l��ZƩM��ÔM�9ѧw��J�ZK��2`��ҐNt��@b�P<Ԅ"c�paj�����P�c-���ѽ5d [O�Q��l�hs�EEc6	�8��sv��{����Nlы/��"�o����ܯ;�ۼt�q���w`1� -l�����K*�hn���Ū�#���IdR` �vW�������|�q65��y=z8䪠�{@�I��Gbh�fK�T���n��s٠SS3v<��|Q[�]@nAq�'c���5v���; �F�Z�Z/�(����[0{�ܣl�@(��&R��e�^��`A�+���i�s�kJ�˖C�>�m�e5��T݀����|�y|��^�& ��L^Y��:g�l��U�0"���x/DE��mkLy�Л����|����u_Q�P֮[��8���?�����u�E���@��FU��S�I�\�Ѽ�z#�prVA�/�s�geލ`$����
���a��B��=S�@B6(t��$����s<S��{�/�r��µ��^�;�KQΞߎz�\N�7�K 2�9�{_�ύF��0�����e�\ÿ����aa��E}�+J7�1
�&&���;��r�G��]�U�P9Q@�y�D��o���V���?�7{�1��+���5�{����<��Q1�^��c��3�HS �����c�@���@�9��x�/�1�Kw|.<j�Lp��a�2.ƈ|fn �q��SF�6 ���Í3_���/�y��ό�x ���H���B_\����5P\"�1>w�\��a1��q�tb��/�6�;m�[鼔��\"?�T(w��}��ÿ��7���j5��M�����k��.��\8��X7�0���{e�%��:���1��nաC'͋��:J4�u�����׿�8��*)Q��)ш��p\X��[������AY#�	��7��[����s(M�_X��l`|�N(�����~劗�|��v�E�÷�� 7�<�W?��Rt*�~�NMNn3����	�v<�D���3����CO����������	��K#ZYZS![0�Y�Q�23@s��;ݮQwҔfb��/.��67��n[3���M�@�B���c��RZg}�A�3UD)iy��wxga^������bcۦ0�K�љ����Κ�����/?
�o�%x!tI����m�y���e_�iqeY����.k������oC�#X���54h^��&3'���3����e��E�0D��y�zCC��>s������M�����ֱI�}�V͞<�}��g
}����d�y�4A�Z�����7����C��.y�`��{h�͹��9o7�\Y��ܬ�]Qq=�i�M���5н:W��7pQJb��*�h=��9\���C.ؕ��Ϛa���Z�%R�\���.{�RQ�7$��
��Ǎo�B`O�`���5�?�2�n���;�7ƽ�/F�S~����Fډ�wJs#��R��Q�����2�ߞ�R�t(�g����ϛ}���9��w|�r-��)�����şO�y�(��3n/F�Gx��|�{c>��<��u�!�����3��]v�̼*�V�%���elE�p�
���{d\�k.%���7��znD �aۣ�ϡ�0�m�G a@q���{ʅ�����������m���P5��@C�blb����s�Jgʗ��K��Ζ�2�{g�O*������Yz��o��5K+��c���K��BN�B�w{j-�i�h�fN��@^;wn����ވ�<@�~J�^S��)=��I��_��rB���o� _��v��<�|������u�!�� [��L�V��7t������V	���k-V��i�֍/��ڿ���?Z2�.��)��J��01�Ug�8�<n+�H�Պ%���N,��B�wxF�p��R�1����fq~Q�L�J#�N�ծ+��)��Z��
��}�:95m@�銕(�)�铧B�H:��R^Ǐ��C�U������{^-<)�C�ó���C���7��#/�z��ME
���`FeK�'L]���,պ�!��ToJ�1�S�����s��F"��֛���Ȇ�@b�5c	��m�R�XU �$�
e��3VC:44�B)oh]lK��E
=x-R蟽�}�ǯ|U�����׹��k��A=��^]q�t��	�}l�͑7�1A�Mox��k�c��Պ�P��el6/Q	�{�� �mV���"�7�M(������Ay��	B0t�������z����)��u���#�����滞����5����m�.��7��ρY\��1|^}��l�X�g�Q�cQ��x�e`�#�u}f����Mh�f=��J�q{$�c="�3�^9b	���3��5�X�����<���H�����9x�g� �I��u��k?����E[��6��1-�+�=�����Z����i����}��<�䩎`��L�V��C�J�4s@��`�%����{ꬩ��'��+�V�7C�Ӳ{^��σ�[o�u�]X��(���B�d���ʊ~�u���������?�Q-�VU,���̩�)�Bg�OF����kϿ�����������X[Tm}�<t<�ٓK��z��`.���)�g�_~��t������s���5�\W&�W9�Vc��vm�[��-�dT)d�MŭQ9x�c!�Bo��������M��&+�V�{[6gǵڡ;�[�������p��;E�X��J��e/~�v�:� !W�Tq�Ո#{snq1�bY�,�N<e��Ԓ�q�j��yU��*F(paRu�_P�޲�>�x���ZͪN�<n�cCC#�j�Z�����͒���y�ݶP��W���y;|�@aP'҇x�B����²ż֬7wh���P�`���<���Ȋ��S5`�U8�3��^:���z�S��HN&Lh`tH�XK�݆�3N"BX�<��E�C,c��-n�aC�����L!�������o
}����y��x������!S觎�7b�ѡ�榧�B�ʸ	c�GL�Ľ.֝�#-��7���Kw��B���~����$k�Ƃ�{#B�G}\��$���fA�Mӛ�!������|��|'��Z�vwCPb�4�������Q��������W�@=�X���	��P��9��^Vű�p��,fx����q�=糏=��@D� 7ܠ�{�~=��υ�L�Dt���漶�r]��B��1J�O�)��� +(�bf�>N:䘀�y8�?�Ә��B���� �лGQXG�G0�B������cB�@��Ζ�B�>\bD@��}A�;���>�����\�+R�����d���B����25=m:u�t]��=��v�JS����s�a5!Yx���C����y����;��n:vR}C�Z�6/)E7�t
��^/u�퇯������Z��^7�nu�M����Ԣb�H���*�:]��+�x�^���48"���o?�}�|�]��Rھe\�ڴ���֫~C��EsI�	�C 	<~Q�ez���ɇE��}�B�8�<p.����"L�0�1�h�d�����*fs9�_��W�t�#�s6u�,�{���<s>8%s���оc��7���妊Ó��J�wZ�w�F���k�UU�fLQ:�O[����sv��J����f�-�47��t!�-����M;��O�:�,-���Z�S�P��B`�9qZզCI 4�6��t�J0��Y�

=lSB�27���P��VB�>��t�i�aуK ���\)��� ����qp���ǈ�B15YZ��  ����9�WW�}���o�_ӳ���M�(�.$�\�[���}������WoR![Ԯ��Q�}�^���irlD'�6�7��ny�N -�<��<6�D��=`�.<]����a����֔���x®�s��g➾��?�t��R'QY����r?���������?�zH��f�cƅ<�9Ɓgu�x=��ʓqp<�4��Hf(a?�7�Y0
&����^9���>4���>E�Q�ڔ���b��G�G���\~ots�8o��e�Q��S҈��s�s&18HmqO܃{�Y ͳ�8�y<�2�W'�� ��ȳe�8.���+/GΛa�
�u�V��) �,�uI����/��c2� )�������sa�D]<=���S�9�Žr�n�r-�ml�Q�?�zի_m!����S� �\%�22bLq���r�cJfs����B�J׿g=�R�q�#�o�y� ��'U�	������߀X�o����}`�����m�����S
}���!�B�%DmQ?e������&'��Sҧ��I7�~�ҙ�ƆL����_o��46�W.�@3����%r�,Ґ��"��'�5��	N@t,�fP�fљ7˂�Ń�^�N�h�K͒���B�l�e���A���,46�:-q�[n��:�3ZPx���~�#��?~W�^�����U��c=���Zԛ&�b��,5]�����_ܪC����43���jC'����v�RQ.O��^����O(Q����������j&=zLM�ݶ!�iSi9�x���D$��"O�m ����A��as�斃���L��C�G�;Ke��LF���m��H�-$���R�֤�§�5� N���@�Cg,��� ��=4 YW<�4}`hP�33v�F����P���-S�ܧQ���_��2ɬ��6�ř�:��#z�󟡳�M���C٨C��CG(!�<���D�p���^���+yW⛽�`���� 
!��^rmr�A��a��"���=R_�;�koV��g��3���x���}�ၒ� �ߌ�s���E�1���<��91��[`<l���s��'|)<R�<���ӭ��j9�˹� ��"�!bOcLx��=KOy�8߿��K��^.�!�=&�X�����Mr��'� C�Nt
b�$
�1;vܞ�2��=X�$:xqNc�o�,��YhÍ��)CR��p4��]�L,���&3)�X0��F��#!A��HkƣQ́G3H�a�������j��w����F� �ӣ�Y��S%\���>�y���민������g�07(z#p3�8�6nٺ]sK�V�^oS�Li\�����Љ�q-��^x���zt��o��i�R*?ys蔭���_}˱��[鱉ե�:��:e�Ԣ���B�Ĕ�k��q�M=���i9�'��G�[mv�c{M5���Y�Ի��,&��@�f@M9M�/���Wr�|F������9l��)͂s�W��+
�CT́)���%[d��Z�~m,Z�~�/�T�^z�@ײ���ِ,rB�,��q���Ǭ���;l��֚��+�������O5�%�l=GUW@�� �RU��W���铦��ܱEW���i�"��I7�`Q��SZYoi��R<Ū,]@g&�jJ�N?zO�+���A�X�9S�t1�� DtP�}���l�ը���Q�(}�O�,k 7�fϝwZ��))�x"#YT�c���(Ƴ�Z���ι�Q�Ɉ,�,t��fX�H8	���2#�{����̆�3���9�u �!�����4\N�s��s]���t�?��J���G�����������3R�    IDAT=���G42:j��*�/�	�ҁUn��\�Y��t:�B��˽��Fk�C��y��� ��p�ys�����x�ω�7�c5/>Jx���ɜ�R�3!�@g����}j�=�c�����lw��eԹ�{��v�=�ؽ���!�6�B����۲e�x�6?�w�6�D�u��g��s�a?���|/:�`X06ΏG�r�^Q�	(���.0E�<s��Õ/��;��=<���5�ϖ���_�P�����5��0.��)�b>h�j�\2f�c߳j���￹�W85.�!#�9�&82�3��p�7���ߎ x�T��/��3���� u�0>�����
ȍ�Q"(�sϞ=�I���uP����q,�9�Ƣ��"��6��!mGw���am�~�V���#?Q���{Jn �an�5�/�/�?�aiaE�LN�r�9b)0谾��٬5��}���CG���/���o�A,92^]m�]]��:l=�<�Э��P2�檲�e�[�*��N���)S2��N����I�ܥg����I�	e��}�|��	���<!���v���{�>������֎:���Қ�έVБ,B��L&���b� 3��ir˸�?�lU�W�XkK9=L����v�x�T��I���3w��Z���^B�?z@��۷k������ڒ(8��l[y�@9�k3W�dOoy��EO��t������_[w��}�kvnA��[�0�p���n�B���P1S���>p��!�Ŭ�}%#�i�`
�m��a�xC�Z��u��)��ݰ�c�<F�j�r�^yH�X+��u�������B+X4����D�H�@,�t�"�e$���wcJUc����y��C��Џ�<ZH�c��]�gHW�by@�>i�Ϸ��n[�ZK#�����{��k�����z���4{B���ſ�,]x�.=��ǡ����&l��_��́�O�$u`��\~#&�!w�yoV��Q���Jz� D���� Թ�U#�N��q�*�\��p���e�^�! ls�e���F({�׽G��cxЌ��*���Jj̣\�c9J��a;�E�}��m�7D�Jf�#�QЬ[G_��BIEC��|=���E�����C��]��ܫ��s�xnxќ��a��;��{p�=B倷P����0�������ఈU�e�g��� �a}>��c��؉ �#��x ��9/\\�޽E\"���t�	}�qg,ڈ�����#������C�n \��p�L�t�g�1�}x@�(���Glp�a������!T4�����DҞ��1C-t����ڶc��͎|�q�Z p�j9�R����f�nitb��]�Yo�*=��zM��1���ς�Ji˖�'�B��M�}��#�nu+�FO�ڪ��@����u贀D���*�SZ�;���:���:�����,<��H���3������lL=r>���(���^^�F;ϻ���>�����S-!Axӈ`�:pJ*@�#������gfz�W��-7�urBoy�U�����yįy�kl�������(Ӷ1�7�P��1/<�W��c���ܭc��޲�:�c�մ�?���&����֖�tƎ	U�TK��瑽*��5���V;�yḆ��8�Lc�3���+��y���>S��Q�ݮr��*�ecO�
�G��ܯ����z�V�Ox�E)^�PT2��F�<p���^�eN��5��j�=�n;C >�NS�$
/��M��n'P�6�`b�Q���V�X�F�R�����BO��]���>`�?=3g7�r�r�~�c9u5:�ı�[�j4m����蚏F_��?茳�V_)��SG�4w�����1�=�<d��Ľ��6�I�v�i:��X�X��H��g��y�%������59ƅ���2¹��}��5��2�7����!}��r#��z! �B�À}�7/+
:4�@PUq���\��PQX^�t�%��Bu��wsNE�R߱������εH	��r�
O��0.����zE �]c<>�s�%�3F!sG��H��_l�}�w�9Qƌ�(�I���V^(H�炏�7���\y$��s�`��M�Ƌ��c�����d
MKx^��wμ�<��@(��H@�#��֕FO���
����C�K@�;�##�� �c.,��r�χC����?k�k1/�yx*�#���@34�k�c��OMp`�d�������3ͳ��z��+�=p��WT�5c�v�W�3Z[o�����!��(�@�������r�ޣ��h�8f
�����_C/a@q&7��jWq��I:�$�¸m<1��R�Y5�ft�	�ş��*Y�s�s5����c'��MY�n«�TN��ߣ}��^\Z^P�T� V�F(Ai�Xݪ4aV*Z3�Q���ZU�++���@�^rً�O߸ш+(���
���'Hs�V��t�q �}��6����p���zɬ���;i����.�Um6�Z��y���)/*@��R:������Yx���mZ�F''8���3B��T��fbx4 ����Z}-x3���p�Y��:�ٓ�t�S��׿�պ�s��8���E�Í_Ӄ{�ʳ\S*[��L@�ֈ�t�.N+�骘��]���Q�(��k`�b��pZ�X�JO ��|L�~3\h;K�Y}u]�l��~}41I���fBn�[W���©��]��}��+_��۫{�W�lF��z%�:vtF���S;��~��S��q$;���������?����]x�.�M��ܥW��E�/����f�sC8Y؛r���Ҽv[�!T��)���5Pϡ���P<��߄p]@:��X�Q	f�?�y�^8��+�r!�x8=���˨�Sv�ہ���yݛw �!n��x7����3�)ap^�\�`wc��|�
��!D�z�v�
�NH#�p7�3^��x�������Z��
·�X�x�I�Ox�{���=Gƀ>~�)8�K�ayq����� [|%Ž�S)� <��϶H���}r(4R��b�020&�gݶ�qO��
�������<x�!ee�$�hS��n ���^2cF�{5���'�(��I��F�1r���s���?kK�D\��W��Q@�m8���=���^%a����f�rg��Ƙ1�5��N����Թ�urf�z9��i��cFc�����r�\�Z ���9k�p�LZ�R���"��Ir|�W����U{O-�q�WChw�0�-ip`�&˨_�J�:LV�<&WK��J(��*�Zՙ[���߿R[����܉4#B��`��n�Ls�&�����~}��3!D��\<*�ht��V�)Af�Hf�!7�oT����:-aW58C�B�XҼO���#�Kk*U�O��3�|�_�R�:��pI��&b�e`�P�T�tAK�5�֫�Zԡf��P�XL��YlqX�p�h7KyXW��V�лٔƶL(�I��ba�8~��ֺ��&FP�Y8t���xY����9��9��wL�o��m���M=t��u��ipl\�;w�?��n�m�2�՚�@��7o�������*ro}}���%�Ծ��48ܯ�撒�X�z6v�+^kp`����1�jm�n� �a( 4����Mj�Jݺʦ�z����o��K5P�~��;t�7ꜧ\���Zq�r�Z�Ŕ�WCi�	�1Iƌ� ٪���?����Ǯѿ�t�)����KS��i����y�~��;��8v�?�!��<,z�G]�,��\qz>���ۡ��ߛ��7{�v����#��`�!�\�"������G6�=�Y-��L��T��v���G��y�﹑�1.��Qx���� g|�G�2Gq�bXr���Y����Fٔ!n��	w�w��8���t��ω��lC7���<������H�����)���-��y9��P �˵����d�Z5 �[�t��8�ύ0>gx�|Ǎ=������3GF1N�_H;����S#��M<��
��E
F��	�>���n�F��#�50$87c�~�87��0^^<g�ude�V�J�<��µ݈t��������K-eE;Tr��ˡ���2.�g<�9:5�`(w�e�0�"���2'�IV��;A����Lf��!-�dV�w����|�_o�ɥ�uz���
}�z�M
�G��-�OzQS�yT)�3���/#]z��z��@!�b.�D�j�k�d��;gA�Sp�� ����{v��-�Z��t����q��4�ڳ�X��:�
)C
`��G������)��	��ZX^S�<����F�K��R�QO�
�Ml��.䩢�����M�6Z����W���R?;:4"0 �,\��1��2B\�[&̃�{B@�8a
��lk|dT�|F��r���"�N��|l�)��+.����Z�nj��O�2?�;~t�����ӥ��y���?�;�ݣD��z��2��41R�[��Zm����=��?���9=���v�G��n]:���0D*<��W��O��C�N���%��+�]9�˹��ݒZY H"y��&y0&9`��klcc� �c�Ɉ [�$��S+t���z�������_�?�?�V�Z�^�WU��{�ga�ˎb8zl���`4�{|��(*^���i�L����*����X^t���R�\x1��Q�V��B��nB�{��c3���H���4����4�\�m�3X[:�ZaO�p7� 5��и`��N���Ky�,�
���f���q��,�� 7-n�A~Na�GyľC�74	�pc��H�r���Jotn�
�SxD���Sސ6�.W�^eqF��_��@]ǑA��%��1r��]>���Dx�C�b�s|�a[�����uC �qy|z��.��y�u�$lyyi�H�q����yz��.�J�������y$?�7��|f��Y��w
X)o��Z 䃤�U%U˱�<�~���y]q2�J-�$��
E[��+u��i����1e J@i�#�F��T�շk���	�V��_��L�� ��k��na�_�е�U�^޽Ҟ2�d�p>�`�y�VV�Q��ݣj͑�Lg�xƥ�[�M7݊X�$g�y@���ͨ���D�C�!����S�C�/���K7�m�r��;��$[��C�UJ?��ͪ�\��e�t<#l�܋����M��}�a$��X�r�^��x�I�u<Wgɒ���c��|�=���?�ϾH���l�v�LX�e_\��^$�B��md]�x�9%��z������`�k���c/�p#��(�j����bش�t�L��b��i�|,tl��[�n�n�X�A_�шa��]�;�F.|@��ټ� ���B�#���5"����E#����ԛ5��1�62�B������ٸ��]�2������0n�������1��|���Vm#���6G̉��)\��o�Hȝp�R.��\����8�o?�ZM֡;/���$�qsc��Y�zv�:����z�G���߄{����8㜋�����J�2�V�ᒧ��7��C��^�U4j%#D��h�3�!H��B	�[�@�E�����������W}䓸�C&����cu� VO<��lg��fMl�aH,l�:����m�'Da#�/z,�2�yM�abu�=���ٓ���6�7͹�.�'�%e.����w
��k��-� s���U̍R��1���H7({�1��X�<���+�+`���Qh��B����1�SV� 	�/b�Ho�|�9^�8�e�>���9?�"�|O�v?�R ��(mFW�uj�g�y%���.�ݲ�����Nb<���0�9xM�K�x��Si����K��e���ҵ�H����0�V�ۖ����1�(;OD4���W�a#��GF*�9��y'_@�ևB�"Ur��4�ymJmp�i�{�O^�����q|}���9��c���Y��$���p���[��c�B4�����$�V��Q�&�g=��Ѓ����r!w�G�t��]��Q���h��!�'{����A\	��y L�:-�`�X��g�v�������^�r+�G��ZȤ����R){��	+��������9���ق���ب����R��Y���du�b���5��f��C?f���4��*Bስ�KeG14<���("�ZF������'�i���$�Ћ��FM�D9OBm���CwY���7�y��P���4=c���c����2հbIc�3�O�ql�j���g�N�A$�����W�R\r�L$�˦�,�������cC��:x��<��QL�n�� &�b��?�C�C=4�NS�֨��8ݢ!W��
,Ο@�^u��k)�
�?�o��u���d�pl~�ӳfQOoڊC��a��#��(��R%e��Jy��A����������\~���q�C�bz�t���HNoG�5��������/�->v�?ᚫo����ٵ+�q����8w�.�q�p#��87�g(�h�/��;h�G��7s����=��f(�(�yy�������z�p��k]9��ܧ�o�	����T��󧀁������A���t�jpn|�sJ���7d�ϱ(����y��s��~X�8#��	��z��K�E���sE�? ��Wy�J{褟.^ �����[Z�V�H�h�ؓ�Bv��.���fȹǘ�/�:�,���w���Q�]� ڂ2�\��E��\q��L�u{#�E���r�R(2B�\C��8#�
�N��%�pp��{<��@Exh��,Q����/Ej��йy_%BT��˝��r�dU4��q�gU�e�W��Z���h������`ȝ|%��C�� �!�~$ʆ���`��������t�r����8�ת�;9t%�ȟ@�eh!B�qa`���
:h�sx�3/�[~��(�.��{p��!!9�0�F�eĕ�w��ҥ��G�IG��xw�}�u
��kM��C��.W	|�s��sC��a.�d"m��X�G1��i�6$�i's�T��湓GնF����-�$�X/U������A�I�Y$3��G�h��9k���1���YB0FwϚ���OL
��J�N���y̡3�N@�b��b�����8h��l����G�P+�����'��Z��e��ҁ���4�DƱ��ø�w��R^|�MH��a�^�P2�׽��DH�\A�TD����vnA(����>������l5mw�G,�a�����ȸ):�m9�R�}���ܧ\�b��;�����H�nF���!~_�����9|�d�1����o�>��kϋ"><���f����7S��za��#��>��O��OC�a�ڶ��q��O�<���>�k�v�UP�V!s�T��r|~}�4��~��f�¢�����]��n�sc���r��;���t��{V9�ꑝ7@���*e�x����r�"�i��]���`xV�Y��5������9>I�*�j��HĮ�ת��@���g��OҤ�C�s�k���G� ��2e!/V���2���z�O� �����Tp��l�t��Q��j%�~��e��GA���)�y,�@�Kn�ƒ�D�U�>�Gs�"ǃ`�Rqh��%��C�ºP��*��`�$D���t�yE��R���y&�$E����S�E�*.:��V^Ǖ���x��]?�� �06f�U�/��Xl��hɖek�@�v����ia���FWN)@��������VJ�O@g���5�GGƍX���7���Aup!��)�EI�z�����ҋ�Gǫ����P�H5��`���b	M��l�A[�P&���CXX<j!���C63f5Ձ^��+w�E9Mn���35IU&2�]n(��[~��Q�'���d�m��D�Z���v�q&����;�G���f�8���z��(��,<D�%,��:�څ���&3`�=��9�肿r.�������O� �5��'}jb�<������ab|�"^#�Z�>�?�E;�1��B��5P�o��c���'���    IDAT���*ֺ	�� ���U(�8z �T�m*�D��P��|n�x�F��F�Y]<n5��X��͞�_U������q��x��_�]���g�����X���pC	]� ��B41���ҙ02�&���!X_Ca�(�!`�T��w܃r+���k��z6Z�	�")�Qt�ģ���_���ᓟ�<>�_���4�;�4*�8���8��mNceei��Y�Q��.�=Z���*������iʐ4�������$��yפ"7<�`N���X��dՠ�������AGb�Ե�˳��! ��e������Ǔ���3|	�酩F���wM���!ο�w�m5/�'�A�%h 7@ȿ�X���xu][.�f�S7���N������w�_+L=4�1��6��z��N�t���6����zU��xE\������{�6���P���q?�A'Vk��q�u9���+}@�2�N�>4W�� �y�N�]�rV�p�*�Z��!����?V�l���~��"Ez.8_��Ǭ����ly	4?6o�3)'�C�j"aZ��C�޳���>�=+���vR4f|<�9�;r�G@��N@G<e:�}J�����/�.U����� ���F��M@7�� t�,��*�c��	��P� N;��l�d�
{��M���
).�"
"� ���&v����Q<Fϐ�N�Q�#Y#Kg��v��䘝�0����!���mTv�Bd	�en��_�������7�)?��N�&[Gf�m�������b�z��FF�vw?�w����"�Qx� J͊[R��A�1� �LՐ3��&gN:%Y��o4P�=���Y��P�h�B���؄-�����\#�86�nF1�C8�B���{��V\x����h��D:���On��
p���Y�a��!�b(;��� �n�hӣ�U�ؼmw�s�:w+B�.�W\k\�\=ɛ`u%�H<�c����C7���[\�J�DȌ����bxj+�� �:04:�V5�J��Gߍ����Ǐ �Hu{��ý=�P$�PxH��ʠ�"MY-F@��}�e�g?�^|�3W�ӟ�
&�&�s����<���c(M�j�%G���qz�ʃ���5�p�y~�K���)�\{�����u�~ t�&sz,���9לj���A�5p�!�±:.�/���0�2�Y�=/�?=U^���yS
i�o��͚c��	,
e��_�'ߓ��Q�6}��US.��c��J�qV���䵹�`�_�3�����"ּ�DOv��v�4��;��+<;���7#�os��;�NA�F@��9�[��|�Q%�y��S�ԱNDDΙ�Wiv��u�k��0x��w�^��4t�_�Ĺ�MF�"*��T��_�N9\�
]{�f���Je�p��8^��~)oM�n8;d@���G\EŸ3����լ��wރv;�Z�������9:Y��� ݽ� �:Y�O�S�C��_�ˣE�͍Vl��h��5Ѭ�w0scQ��hR:�tz�X��^A{ϼO֫[��>	j��������!v�<�f3)lߴ!�P)/bl$�J�8��[s��A*6b�8=�E�@3h���6>{��p&=d�I�N����$^���]��w>d���qg���~�s]=f���ب5ya?o�lC�z���7ⶻ���vT� Z�$�2<*�1��Ԅ��p:eZ��FA�7؝�R5O{jf� �]ی�u��)��C![w�4��N�n(=���it�z�2��E���/}�ٸ����Ѱ�~��z����W�����|��#�-�ʹD��nJj��7��矍��byq����|���@V�N`jz�ھ�HD4��,
�yd3�`nlu�����_F'Ŧg!5<�|�I�&�MΠ�`-_��-g��N&�V���'o�򁇰p�Qt�u����}x���f|d�����7��"���&�`����h
_��{�w�
��F���#��������K��0�( l�s& p#�%����e8b�#�z�
5�	�_�'_����A�%㖿�P&0�w�~���)�Q���(w�MU�)7R��),���胹eG�W^������B%U9v�0h���@�`8�%�O��q,��8uL���)��E���=�w-�d}��QM�<Q���� P ��>�ؔץV�rּ&��Ivtw�?�k����L2�V���/6��3#E(�����"��<���wd$h{՚��w�e�(
�9��d�p�Ůw^����������n���ϫ���%���ַ�s�{-b��2>-;вUQ����>C��<=t��M�眡84du��>��4|�K_���:�'�̑ Q�����Lإ�~��P��M'�J%P�>C(�53�����_�����h����k�r����b��>HGx��{� 7�>�*�`�u�Y��J�Ȥ☛��W��Q�!�o����{�E�.F�k���ajt���`uє�ȵظ�>T���n]Լ��ُ��/~	��y����i�����]z� ���6���&�K�a:7�J����VkA\�͛���eD����Xv�IY蝞�1
��@w�s#�z�rAvzhV�F�s�����63!k$�5bq��$��G���nC� ���ћ^��>{7�����ׁV���+E$G���~��k�%'����Z%o鑏�o��OC���=�r�D{����k����)�Y�nv��ΐ;�S� ��2J�*�m31"	D��Ǉ�DM�@�%Og,�Q'c�㘻��kȄj��_�����ǵ�M&����C�Xc��n^8���,Z���4"Q��t�D�k������>����_�	��0N��F���ؾe�f'f��v�J��'��-2W׭r�im�"�ɫQ'/�J���B�bsCb�H�g�g�=q��Oc�����b�s�
���鋔��"Q���A����Ks��)��͛�KLn^7�0�>C���2<ˍ� ��h�50:B�<���e8����P<��X9b�[��O	��'�L�'�S%zJOp>M�>����i�q\<S{������}�F�O� ��	|�}R�<h���ދ�h��V���dPh͸P��"!�ᒃE��S�S)K]�,w�������С�Η>gy�bq�����#��ce���a��x����oJO������S���q���̓��s��� �"C�º�`C&��Q)���O�K�z@��B2��2]��A���t�?�vyd�l:�P��~��8Z�~Wz���O=t���YP'��uEӋu�u�P6q��d"�P�C���^�F�X��m��p��Q�s��j�W�R��m���N�N��Ұ\����f���]��l�R���|9F�G13�:!�A�4;�!��/�Neq�Ӟb1�����q��N�C+��a��z��H�nB;C�M�	�F]�~����������u{�*Uc���Ǣf�Rnw��!��f����=��{��V���3q���E���W�czj�}p�u���M����h�0��4$)�V����{���vcm��Bn�RO}��ȭ-�O��۰0إ��|7A�d�Ͻ���Xn�L���b�Qct�q�j�:A���b��3��fM� �2��=�=wބ���!�Nq��x�z��E�@|dk�ť!3>�Dj�����7��F�z?>z���u?�Pf������&l�C:�i�o����m$(yw\K"������ɔmb����'�q�RH�����67F�뵉*GI��F"A����_��|�;�����8y�
g�|���*|=�S�6v<���u3���SF��M��@���
W/l�h8���p��|��A@:��aȞ�j�Q��	�
G+t�<=G��RF�t���4�v��F�ב�!T*%#eQ+�F�Ͳ��.�̚�p����>0��=`n�fPO��'�<p,~ͣ{�P1��$]�H��S<��4E��;�
ϡ��C��l��6N1]�%�Kz�|_5��j��E�\����}����9J�DϚWU*���*50��Oa�y�ܜ��KY<���v��	��US�[X��رT����`S������lͮ�t3TL%/���L\&Db {��L�m��S�C����G��[�^|���mb�q�wzxC��uTs)_�~c�Vɣ�f�2�2�z^�nc���Z�h5s����1�S������XI*<���7�pQ��9t;ƒ���?\t&��`�Z�5��͠d5��\����[m#�47�յ5�ڹ�V��4�����;���%�)��A�G���[����*H,r�y�:����z�����F��@�ga��Ih�d��~�TҢ�j�k���k��q�߽���ݸ�K�����x�kd�[n��|���H��^|���>U+k���'o�M\��q��<r��XZ]���]�X���~��8�o�q)Z��F�h��ѣ�r��V��$��E��0�"ec���:�0"�ʵ��&�RA�+�x��G��Cm����'���y����@le�����fؤ��D��jU�Nf���}W~�J|㺛0��eO�����؃�b��s���ȭ�Z���#���z�A�7J�r�b�>y7ƫ�K���3���Xǖ��9�Io��%h��U��h���t%���X!~�]P���˘�+� �ߕ�+��qT^%�P�^9]��T�� �g�r0n�����ש�l�rI`��x��3^?�A#��C�  �s��wd9���kU���}��*����qs�f�9'8Ѡ�|sS�񾰰�_��_�]w�eF��ϼܔ���!�1m�<�t��e|���4����V�hQ���M��.o�W~\������pEB8�|_����`>\޾3�ܩT���4H��e������w�}���H!��l�1H��/�\{��ok*������O�5�t#�}��n��6l۾�vۺ�����Ë��̯�M}��v�%��#H��0��0��$��.�?R쏼����ˣ��[���H���B�~��>��Z�2���!k�e�X��� =�InWQ������^������	�w÷139b^z���zm�n1~�cȦkݲ���0Z����?�sqq�V�}�P?�"\�sp�Sγ�5d>��
�����K���l6���M7�/z1&f��ZپC���o�J��^8�b������
a�Cg�6�>���t��i�0�^�).���9�-�����c�)PӔ�6�I;�@��"Ca���6�)�=��C<�m��D�ě�����Q��?�.�0:w:b�1�KE-4+k��#�!�blx+�Tk%ē�MO`����IU�PyB
u�@f�c�H����6T��c�!bqĳcƳFtk���@s���t�����ID0>3��䧸�_�E�B�Bvr3���B	��9�j��m������������k��H0��?�R���܁�����_}��^� �{n��x��\ޫ��k��k�&V,;���q.����;[�`���e9}kzH��|�(�)m�V����8^���1�{���ƾ�<� ]5����j��MZ�m2*�|���1��!��^���3�e��z�^��A��a��0OO�@,<6��ҥ��ss\
Ws�����g?�3��ca�w�`l۾�ِ=����,J±�/��o�w�w���4gߩ�Z�қ�3��{!v��W�qGT��LU0-}�ע+���5��i_ss���p�ClwF,�Z�zN5O�+�)�g8�4J���k�:�j������ .-~�������\���x 2r�ٶ�]�h���B�]Y]Ŧ-[LXfߡ�8pฅ�	�L]����}|�������Zr�t6j��N@F��f��R������G�ޛ�^d�?Ρ�O��� �?ђ�=��dm����W,!�ct4�׾����睋�p��>��=c�0��*��2�5+y�gJ��U��ι�he��^�gi���<��qj����=�̡��%/D�V�E�6�-&������]w��!�I�8~�*������D"_��4���-](#3���D��]�Nǲd�sE����&����k�;=4JeT+�SSV�֦�
a��<¾pB$H�� �Ѱ1D#�����E�i��Goy=���D�J���Qo5q�`�\�R��;�9`=܃�4�u��gz�^�z��3��"�r�ض}睳��c^*7�����s�!�����T���+ijd����+����#� �C�b�7ahd�1~�U������-�97��0��pC�ø��[�� N E�F����qk�h�_j�J8��������������� �h�<�}�݇�ݍ���ⅿ�Kط�	�kzm�J�[�8=��sM|�,-�*+�nP�M*��[��_Lcn���ˎ�I���`UB�2/y7��kSW�\��<��.$���N�[�a<�E|���y����2&t��w�v�^��8/��1�M;�.�[�����!�]�^���y?������|��-6Hr�r�2*�s��sA���g �LXİZ���$�/-���x��x=����b����K�xm��2 y�SJs����J����pye'�#��{�rJ1����p�����\?��K��9��W����?�*G�E�����_��5%i�5$��o�_6����#��?�`[�����M�ࢧ�?�!�>���-��jw6t<lO5r�+[$�9���:=�^<a�)I��o�?���~�]Ǌ��nx�,=t�[�N�g*GN�3��n����	��<d����i�,��ǖ-Y��ͯ�3���$a�x������F&�D���J�:^�Nk&�D�d0�B�.�f�!lz&l���q��b?s�4.@Ww>�׽�u��_��}{�������ãXXZB�M�~�ʥئ�u�dUr��N-`���1�To�g�����IM��l#�����m�F�f�x�����+[sD��I@giN��T<���)x,+a� ��|@�M��� [�v�܄t���H%�����ۯy����"�b1=;�}Gcd�������%�㣦��c���Cx����I?��V;���&ǳ��ģ(��0�ɢR���4Y�W�0Ɔ^�r�����M8����&�7#g���廇ǧq�O�@85�~0cVv�]��Ho��������[f�p�����Ǐo����B!����U�\!��׋X�޳H(���2�ݽ�����}���1��3�z�n;x?�ڵ�����{����/�1�����ZB+n4\G�¹q�y�\oI���!I�D�d��Ir��y�7�<�~�;�:�W�Y�����k"hr3U�φ��1q��������<}~���M\�w���[y~z�|q��I�%9[�����IΧɎr>8?�?�5�{"�9`s� S�-�eи��P���F�Pl�۾p����Ӱ�s��Gܻ��Cg���slg�w���7o�b�����x��T�M���J�\��J�2���D���z�"�1J)ֿx@�8�^�\�^觼��9�u�\C2DźW�%y���(�V�Q��rӻ9n05����Xy	�"�^��3�Mgl-��
�Ų@
ˌ�M������X�M�=�J�{�cf�G��N�n5��;=�S>���r��_����E�u/���[���ekYDBQ�׊Vk���]��\��ɒ����çϲ{(�E�'��j�cnv�~�3Q��q�O�E��-E�.C���~�L���Ix����~�Mձx݂cܗ\�:O�B1��
�6d𒗾_��7-����MV����Z��:8�̳0<>��ܺ-�F��Z��H"�X:�ɹ���'J�����u�F�Rܰ C
�JN�K�|Q�=@��v�E{H-�GV�����q���C�FBֻ�Rv=��B*��������l���m��EϷJ�=�>�b��W��7���}���7��K"94���f睳���#�a�^���Ǚ+\���(#��>    IDAT����J(����lQh��K������Vӳ[05�وp�U��Hē�2�ѭ�cr�td���f�����o{>����]-��sva5���<�Z��-�w���5O� ��R��p,��������H'����������g>��|��/~�HϺ��XZ8��{���ho��7��;o��cHUb+�1p"hs���j{�sg��ֳ���=�������dܠ�W~��� �Z�E\�4Nr܀Ur4��9��x)��cs<֞���}���X5�򤌃��`�)
@&�]�ay��'���9Ny��F^�c�K":F(�>�μ9����3bMk<
Gs�֣�O!�d�h\|�yL�>=i�+	p�W.������N���Έ C����]={�tw�>�t�c��Y�����.��bK��:��|s.�n,̓3���G����(ͫ�;���-��)9*��b�d�W� ��<J��^s=����X��������7�uNIb���T���)F�Z�w��r����彑��y��ß�w&�u)��I��=35�mo�!�p��N@���šc'P*�0�����9ˌ��v�?Y��d�g5���>�9�����9�{V��W~�[�=�����	��͞F�V�p6m�������ћa��fbiR���L
}��������s��mK�N'�@�u�	\-�!m7�l�Q��[��Ǻg��ۈ�	ڮ�c�J�±M����xN����x�X���Uˡ�&GS	c�S�f}y��A�`Ӷ����8���"
��L���׼�)Q��a{m�|�����ex����iүd�V�(��!�۴����დ[Y���k���:g=�{�eOӀ���V�Hg�>�׿�%����#��ٗ?�ο2�+>�|�?�U��F'��Iصz�u[��U���(�ȷ��+ȯ��x����{E4F82�@�욲\*����^��W`q9�#�����2>���USڣ���D��.u})�Q�-a4�_���#��'?�76�5�h�P�s��BT�]�w����@�Z������#�(��[]��>z��cW�#�>y��L���s�D!�����G4�����e&������Fp���t��hd�h�"P��J�x�yi�I��y���)N�7s�yΫ�Z�!
d]�թ���_�|m0'���ğ���
�˃w%U.�.Ä�T�h51�(�������A/��^�"��A�r�N�@�腓��ۜ(r!��S�w�pQ~�6"e�����@��9t
�����mIi��(�g	��?�4Y�����PXǉ�ƂgZiii�>/e?��)*���~��h����z����"�2�4�2b�\�yۚ1�9ʹ�=]#��օ���""K�A��z��]�TMa�O��%��h��-��k�1u�c@ 	S\�C
��~�F�YaOF��0�?X�F-���"V�H%��uǗ�O�W�E?��.!B��/�d���N/=�F0�B�������_�����^S�t��Wo`4�a'O�ry�+M��o�b���[n��$[i���T�15��a#z�?�Q		ud�yA�PcZ�lb���n�:\��@�k����l�̒c�=��G��(2�P�ٽ��Ƈ23<�a��l��y��1D�I�9�0�M���J�N����4�d\��ȎO�����x���Z�$�p�q�T�B�ϩMnc�ѓ�Xr$R��^C)�C4�ܑ�'�����]���4���g^r83>�S)̳�㢳v�Mox�Uԫ%�;x -��s/|*��a��u�E;Gf|�r��ֹq��������e�-���������'���-���EHRk؃�	�̲����XYYá#��q�nԛm�╿���w�����÷~x��I6Yڦ�C��ࢋ��W��=��~r��n�s��(Z���>�b��-[wb~qC#C��=������/��\�����[7܀k��I��/��-?�톇�v�B�]�c�ݍh���.}�#܄xm�ZyCYL�6��ʣ���eҤ�ʖ<οu;/D�7<�Ε��g��{P�E9`y��>�Eώ�b�\�偮\�f⊜<����
��3����@$�Q��s�x������5�y�1 Pn��c��I��yz�Y�5
��P�+�S�Y��V���1hp�]�]���A½ǁ�3�e��&�7�uJ����̌�=�E��1�9F���sL�[d2C����Zn�(I�T�=�N�1����k�p�b�ʕ�����h�����(��y�K~N�t�)3J�0���H����}�OgT�6T����xO�փ��Α��<h�|Vx/�O�x�\�2`��X�>���������kL���wb~a�+��t7��=�N0�P4�~4�@2k���SNX�����|���5^U�Fbu��n;�9	�Eg�3��!��5�.;.nv���a��l����+�"h34+8�a��j���i=�QH��^�Tj�?v6�6pg�s˫Z?r*�9ˬgF�3�a=���X�4�N���Z'8*A5Z�u�a?�&��,�@��<��wo:�4S��/9�^�L5bs�Q�Z:n�Ԣat~O�+��lT8�t��}�=P6/��6�F����+�i;�N��e3zl\���	+�����A���N��)WN�i睍�|���k��������On�mwއ-;�ž#�f��sox�e�Ic<F�k����6�k�+���h����Ӯ"�p�)7��y�O��@��ۊ��i�s��dabr�^��~p��8}���82D���=�g\�4<��M���޽���X���vl�v&��!x��/ R���.��i�y��7b$��?p���q�羈����M�T\E��ǁ'�����=07%�M��`ܮA�en,
r�W�<ܶ�A���VuD����ڴOzI��9���ǵ�E�o�?;��]����67m���N@QZen|_F�lKm��3$��"E��
�+l������� �p�n �ʯ8NJ9�yu�´\g�*��sDT����Ǳ)�����~E/���,ǥ��As�9��<㌝v���/�*�����4Ǥ�	���]E��@9&44�?O/��!C�g��(R��?���9FUb���8��n����}�g�:�<E{y �����urr^\���(���D�vWٜ֊�娦��q�.[����Ӯ�
�d�e�_\��j˹������'A�̩��[���7>4_h��ލD���z1W��	��^�D�J�����I�0����h������0̍t��s�@7��/�sMLx~���GB}�������"Ïz}z��Ō�JD�y�]I8
��^C�$�O�@"E�V���v �����b���G��Em�Ds۶��|'S�1ی:ݾ1�i噐Lߕ��ܫR�<l���xa�����E=��_�RX��m�4��.=�k�;]��Э{[����� �H�ڨU+H��8k���bz4��;�v˚�����qǝ��.��2Sؼc'�VPc��U�p4��u@h�^.#�(�WG2��(��6�p��ɬ��ֶ�k���sg�O(6�W�@!W Ba�3�hV��cj�n���0�5�����5����X�R�#C�z4Ø��҉���[�Z����f���M���xe���,�����q�W��V���>�g&�ӟބ@�ë��+���j��C�F��s�_dŁ�0�:il�P��_�$?Ǎ��(�D5�!c��n��X�!���<)��Mǔ'�U�17u��	�dTXdŗ��X��{Z�<֓��PxW�*@W�����	qц�ݻ���h��x��!�ϱ���x�`TN�3�5���'�Tޱ��(	����9/��Q^$�#���x<�P����
�ø�DE4�-u*d�'���3�1h�=�����}�L���y�����cSJ��c�D�u����ľ������N>�,q<�&<����RN������'�9Ǉ��{j�v����ΐ��q�I|�W=tz?������߽�����^{剒��z/�5;�Z�D)_pGg��Յ��J���ų�}~����߂tv�^�^�N�tO�|�qζBj�����ZN#Ɋ�h_].$p�D��e�~�vˀ�i�^�ら�D�t	N�$�!����m��p���@��Ǐn��pM��"�������-�Je#o�n݊A>����I�v<�R��5ԙ�c�d�<e���BӃ�"L/�m�1���mr�Ѭ�Q-�#�b��9�����ı��l��1�`��}�x�!c��c{�����yj^�`�KF]��!��1��O�Pm��q�S���J�r	�j	�d�r�JcɌ�R�����լ���<���09���ʊ��ܧ��Iی*nҼ'�X�fӄf��ch��HgFl��H��Y�	,-�[��T6�7	����Y�}<��g3�D�y�J��b��z�a�t�N?�jC�,�k��*
�گ|�^s=n���HD¸��p߽w����&b��a���(�;�Qʋ���k+�,@�����e��J�"�#�T�����;�N�6� =�!0s!m��Цi�_�L`�\��<����څQ��*T+�A�Q������s��.�?e��:lc�B�߰�s!��yOn����;c����"F�� �f7���ƒ�'y�k�?y݌v�3"�� 0����ܹ��I��ǖ1���s��OP�������A��1w*��]�#N攝���E�J�A�<[C��2�Dp����<�kJio�~#qE�7�*1��x��t�י��9��קT�ຳ��3�sdc�}J��)Ne~���M�0�ș���ɱ�~A=� �r�8�	�F3��3N�)�w�J��|��].�^�@�`�z�!�tn�v��RQ�\Z�ٻw���;ز8~��C�Ԅ��u��tC������@����ΐ�m����9�ޖkg���X��ud�v�e�b�ayF����}����z^��J<�����;�ׇ��[����a*�˧�B��^b��$���i�_g'�D�p��%}˟�=F�0q^��<s-��痦[��T�-�@�ը�Z�!s!w����9浕Ut���Ѹ�DГ�.z�҉���m!� �azl�$v9w&Y*ddj�	T;]�=v����Ma����U�kc��6��M��Q�W��p|�	���Ex����9�����0Jf�_��} 34�f���Ms8<���ci�bI�D��--�@8Է��^����D��(M�p�T
�U����C@/�x��#k�o�}\��H�8��y対Ǐ���a���/��A��҃^�`x|p��(�d�?�߷�l�����A?�H@W�U^��Kb��[vac���f+��^�4�h37D������?;�u�i:̛�:��U��?Ǡ�+�)��ǧ�kyo���N&�ɐ
4��U���BW��c���]ˋ�\�iQ!`�����F��3X\HZ�d�Ô��wynΕk��矄E�8��謆�="��0:�[v�v5V��� ���`4D���t�/����62��;ﻈ�"�ɳ��4.����ɠ.cM�4e�g5N�Z��Ω����9#R���tI�f��WsH%G,�i�����9�ˡ�6 ��C=�S
�o_��������6{�@�ٵ.{��f(^Di=g��=�=z�=����K�g�*X� ��|����I}v�Sp��0Ӡ���!��9���;��X�N���'��E[��o&��=��Ҍt�M�Qɯ"��`ۦi\u���1'_��V|�S_F�ME"#�u�L�kvP-�l�'9��>�l�M��c{ט�z�ф`M��XjB�	�]pD?��1���S�#����.Zuz�x��(-jz$n9�~�mz:r�tE;ˣ��cTv�G�����'��c�D�����̖�q|��~<�J�E,D��C��C4��Ms��H$�(����lձ�p��YLOc��	x�Z��mt4Q��M����Qo�e#�P�P!�O��ѓ���{121���1�W�N�$�������љ^i�\s�d2�6��D�Y�Vꨖۘ��A��1��@��ё ��N�<����8{�N��]8>��:~�^�n�՛�U)7\�Zw]�h���6xy��Kjs��*�Yya��)y�px�Muك�T�X�$`U�]
o�h˺�I��R�j�����X�)��>+/O�L�\IQ� 8)Ԭ�O��U�{9AgЫ��(���<��y4����\��������6: wZ0���L��T�/��@�)3+T�#p�[aq��<��lԣ�@��X�y��]����w)��o<�~�{��p�(�"0�8���#4>�m�+��7�RY�`$�s��Ґ��x�ϵI���$��3�����y}ay�Hq��.�.@7�F���I�`�;�{4��:��u[���o��d\p��	�+���������f3�C�Y.�KgȽW7&���0�:���E/���o6E�v/�n/�n�eZΊ6"���ϭ��M�0s�	�N�����/��U�:+ۤ��V^Ǳ�p`ȝA�H��@��g_~	~����j	����x�CV�Fb\�l��m�ԛ&�s�潒@ǐz~�d,}���b)$�CX�Jۂ	Z�Ǽ��刬'-{����{�Z�X�X@81@wd&G�akYz� �*3c��qڌ\x���E1:HD�z�ݨ� �I�3ع�Lx�-�^m!5>��b�F�@��8f&'164�cǗP�xhv�,u"��n�3��,-���sתe�>0mB;��&�aC����Ǣq�ҹ��0#���ߪ�E0�
��%$ba�{J��y��d"Q�a0j��@7E��Pf�O,ct$�P���C2����<�J�C)Lf3S�w}��
^�ꗠQ+�R	����&]��70�	�s�p%00�ȗ4xMγ&��V��|7�g^��"77�S17+�`ޗ��u�x�(��[�]�y�@�He���x~O�)�7X�67��m����`�@Ӻ�U��+?+ ��s��ynI��Z%23
)K�@՞snu?X(>��B�������j�ȊR2c���۾#cX��1���I��`p���I�q)�%�g�}PA^��2��9�2~4����
�#><������/����`�Z��*�Ces�*�lPZ����j��up>U�?��q<<�I�����Xlcl*W+��ۚ��ޅ���6<��u,�䱸���}����YqD@��6p?r��w�mN9@�k����?���./�z�@8�A�P���a���X8q�H�<�p�m�(��p]��B$�2��H����8ˉ^�-z�ldQ�&��3�s<�ڸ�J2���An�RS�<h<EkL�<���~��x8�h�2�$���g��:��T^K�$i�x�*:ͦ��Q�9���\�a�Ă�omٴ��r�)��,Gf Y���[��6��JAhd8Pp�s�]_�D�6��N�Fu�]!�?8����ܗ�D�uLE.b�p�`CrM*IQA�17;��|��ce�(���|q�'�\x�E6��?/�"��W��\��O��<�f�01��4E�����	Z�7Q2hbtF����;�XF��p^=���ZmW��u�� �h��7��0����m��ŋ��Kرy3�N�[Z��������������,��q��V��+���&��������K���8��8����z�S�o���P-l�v^%G��$;��ԁ�S���-����@��Y��Z��`�l��+77i����&��(7C_ʯ�sb�S�C�v�Ք3��1:#��pWG���ug�l0�N�����XDZS���;��T��3�.[boK�D�v2*���Wy�@������	�	}�H�F���~��%0��T�@e:~��"�����[��J§@�c��Z,���\��<`]�"����^Ɠ@Y�γ<X�Gea���j��F�w�_�n�3~��U��P�    IDAT_�S�1�S�s)�s�kUjH�^��߹Ɣ�44��a��Ȉ�����e����7��$�� ��G�03��Z{�F�\C8�@��%��l�b��v���$�Iz�$�@�ҧڧ�ru�wi���W_��b�V/��+ru�q�H�r5�A+	cٚ�la��_1�F�D�QiT�'8sڦ�B����!'��a��I�c��yݬe���%a�4c��őQo�z:C�$�����Q��`u�lOJMx��B�k�Lk8�quHd��v�ځ+(�*������0;��'����A�A"\Xu�cc	S��ȅ�̀�աl�~�@��s�I�k�X��ʗ�:���m� ֖��R�h%��p����� 8@ǿ?X�C�><��}:��ηcn:�Օ"�
2��Ϯ�����g���c�|���W��ZBzt�V;�؁�L�V��ٙVh�l������ay��2����\��k�C�矆�~Yը�a?22d�@�xM�VW�}^��"���	e��������؁�����L"=4��@fd�P�r�@ّ�U30Bѩ�h4p��Y,ޏ`��raoy��Q*�l�!0�4���6c�T>Z�@O�6~�[�ꌹ)s�Rm5��	$|_^�͗_�r*�6`���8=v3���6�a�J�.��¨4$�*�2O����:7�2*X�(u\�S�o�k���������X����Y`) �y��+5�sX������+�+'+���(�  ��'O_Q04ry�v�L���=+��xΖ����(D��h��z��LU��MM�]�`�A��d�2�8ni��3�k�{�0�B�ڏ�>ӽ�1����WD�ȃ)��ׇT!b�ɜ�������� �CC��}:3d�^k�q��<*�JZT���~���������;wn�%quPBg����~���?�ׯ(V�算��"�U(�B���R��HP��iD��H� �P˼\��]�Gϗ1S�q��}@��o���
i>Y����9�P�'��&�L��_��+�ny)z�ѐ�{7U��GG�Dj1�G"�@�тG�z�^��WA�D��fL�Mcimňjg��/x�0;1�J����$j�����R1�ˎ\4xh܄#�!W��㦭B�<[�~C�4������%��T�R�,���K�h�+���d8�l�ߡ�N��� ��6z�v�܌���]�D�xྻP���a�Zv�w��щM8�����p
��Óؾ�,3�Z^��*����`}���wY7�J��3w����Pr��H8d^6�L,@�sK�n��%��w��ĢX<v�����w�e��T��XZ8�d"a-k������t�y��{�ŭ�݇��4&��c����!6�A?�C�Z�\{�\A��רᴙI������x�zן���}6'��X[l]��`�[?��=��+����s�tej.$�75>K<�_Ոu|���8�5)�̶�j��at��xn�
�+�gJ�''Y3ꚴ�;4��o�����*ϩ��$j�=E�!8�@���'�cKmO ����p�}2��#��6��)#����#<�$M����?ߓA�k����|v��%��ny}֐�G����Jp����[F� X�9v�B΋R?��v��眿K�)����9ߊ�(7�5�c�ZyO�����C�
�sli��S����)�����{}^ڠ�"�WZ��f/�p���G����k�ei����-�>3��zO�=�R�C$���N�%�6Ӿ��G��~�f���:���␇������ P�`�ժ�7���2�p(f&5��z�Y����^0�kA��z�@��
�j���%����P|>W����\����O<�Tk!�"��w@0g��Z��<�v�<5k���I�%_,+�CW�TP���-G�f^�eaJ�����m�AO "~�5,p!j�h�귝A�׶Z��̰�4Y��m��naj|g���*�Jz���3�R\Бby`6�K�u��S�&oJe���f�f�1I���БU4��y�H�X�x�����<:k�5&n����an��U�1�C����D�<��V�ѩU�����Iĭ���@(L��L<�kl2����G�w�M��]�v�,�#�<d��ҭ�M��k��G�����R��dr��P�x�r�do[V	������Sw,w}f�m��M��Qt��w귭�.�b���*�Z���[E*D*������s�f���ż	e��p�wa���1^yWiPu�at{�ˈ��Xg��Ӱ�G0A:����_oëֱ}f��Et�X[=���篰o��f8Q���dn�4������qT�i�t,]W��w�K��
�&Gc�s�ߝԪ+ˊ'\N��޷�_��(Λ�sS*9mw�g9&�y����x�7���_�B���8�Aje2�xl�8�k��;��kS����� �ʀ������ѣV^��Xغ^�?v ���v����3�{�����%�*&�B�/�G������wQ�����?�'�),o��/6���&s*�1��օΥk%+�Phj����c�ҵ�p�8�|i��9�4���"-^]�6�&yE$�w�0��8E,�5c͑X����(R��ս���t_�<��Ѣ$�����)H�o��*�`�}n�V�M�ٳ�J�X�y�|�,����8�q����OC��~?[�z�����~��v�}F�՚��z��{���4�F
}7+����l!�/��=�ᡇ�]����K�|��/��o~Y$��H�3��56:a�-�e���Z�E��j*�10%�s�lݲ�B�6�r�l7�J����s�2�N0 �?u��$0v�T�*��%}Z��m���B�v�?6��'��Fլ��o�����{@YVV����T���s�i�D@���b�qt#�g0T�Y1������H���r�u�n���=�ٷN7�3����굾�V�[u��s�y���{�g?�٭E��١��H�#}����<����@R���R}��p�"�M���G��T����a�#��,-]h��7M��GR�^�˩OCϩΛi�q�����y���j�ШOZ:Q��mգ��5gy��5�������>�=���7���m�i����%˗����_]�E^�����;��Ѫu�,��Y���L猾�C#c���m���J"cu�tXD�IUԫ!��N�.\�|8kXub�2V�y�Su�O�؂��K'mlxH^e�Olx���tڂ��l�cZ)�	H�4<X�E��m߾C=��J�mɂ�R���l�d;�%QSE�
٢MO��x��6�s��m��Ġ��ԓmr��蜈�ˏ�y�|����N���H��N�DN~�]��b�B�R�-�=+ț9�Z��t�w=o�/��+�<zdn`�<'��Gx!�M4	�`z'��[�s�h�P�$"]F�g��=�v4ɍ�G� |?�2���p<�w�7n,��&?8C�W�*IŸq༝U�cGt��P�$7����ҝ�_�ip�=�]��~9Z��厀窹��\���t ��px���C�޽/�4L��x(�����^�c�2As��9�>fqă�plG���#��)�38N�4�=uG�� �xxd��qH����p8#���#A�9 w5�ID��{Xb���*��g�)OںuO�9�.Z�/�j�J�Nrg=��S���yK������A�ۿP(��og�i�\ny>�os
V�oA<a�gy���11=0T�����v��~������Y�t��{�젱<Y�}��+���Q���\�1`r��W�[Ʋ*�5ʕ;Q� �32�*^�0ye<�] ��L�����O�J�6u��#��ֹ�l�>�h��4{ȍ1��熹����X�(HFa&��yc�ł$�D��.$m[[l
�vu�r������̳��1���u�[�*r����X"[��=���Y2�_<���4��U&(-���Od�'7�A��ר�-cSַc���6���r�M���z��1�O����謕��6���p�����Wy��/Y�Ng�Z��"�bK��MU)��k���M��f��%?��_.��Ӂihz�8�4U5�'���)KOW,U��<7nB�LY	���fwwX����|�����,�~�:���w(z���!�I�ct�b=s��Xy���v���~[�n���vYK�])�d=a+�.��;�X�&K%jv�qG�S��+d'�
k�^(�J4����fh4D��S7�ى"ڰ��:f6G�����زq!N�ѯ��<Zu�6�К�#k7��|�?'��Q+��SfA�mȭ��4o���sq��9o�,=� {d���FŕƜ,����GFBj¡sH�qh�c�5
nn+5�؊��yZ��I[�=n�8?�AOA�R���N,�:���^��Bd�4�7T��8���Ѥ���78V8H�-���k�{�b9>��1�9�=��<����;�q΄��+�<�qn��8<#��A���S-|��U��}�ݧc9Z�{\@F�7��?o�˞C'5wh�n�ǹr�Gq�l�����5�@��w��{6O���[ڭ<U���1�>�n��8����=�~�<������������O�k�C2���T*����h:�"v��ٶ3zo"ak�\o��_�DL�t*DC�C���?\�<�En�9Q<��ʘ�s��Ӹ�`I'��NSn6�?+SK�0ɯc��=�Q҆���ZQ���G=�tE�F� q"$Kn� �X��2�/T�r������A�$�e3�&������������=^.ےEKm�\�-��Z}��]�0V��'��3�̒K�[$��� MZ��N0�k��D�j��S62<hV�ɠק+6ݘ�B����y��x�J^����R!��;lἹVj�ۊ�mŊ6g�|ۺe�����t����Q�LhP3k�<u�۶c�z��&�%�6�o�z�C�J���$�}���2�+S��"�)�� ����V+�tu���Q�O[6A�!#�������뱅K���m�>i��,������0O&&����|R�'<&�j60<bO?��,X����S�w������H4DË-���m66�o�lݎx�a����َ�;�R�l���R�5�͞�*���n6��J���c���V�Az3�b��~��1�Iȉ�Ɖ"U5/ߢ��� ��>97����oS4��nti�B�qժU>��4����{��!D��p�_%��W�QT�y��a|^s����(����c���>㑧�U8*8���*d>7��#�<���w�f3�l. D�g��y���n��x^�}�R����O��I�n�&'B�6��p��ktG��9���UF�}	*�Tk��`L��~�)�8��{���wْ%K,��I[26�n��/��Bw����Vy��߯�O;�9	����ؘ]x�rt<���y��3�hvN���R���׾f<�����������:+�
���c�����/�Ҝ�\��k������Ur(�2Bk�ڰ�����_�*~ZoՐ	Oɠ7txl�iJ�����`�/������׿�b.��b�R��	��w�� ���c8�=���Wƭ��*A�w������˪�'�ڴ�a0�le81穜����r�4�'r�t¦j����C${�|�`84)�r�~��;��rҜo|>9i�A�7ϟ��C�j��І��&bc�3"A� ���I{�v�i�`�qĒ��!�)� /_�B0�3O>��y��TV%k��{�jtd#���Z���6ɧ&Rt>�4�l��+Ԍð'p-��������*��T�����Y9k�N[e|�*�#6�c��Z��-[��ҩ�X�S޺:���OLXoo����[�q��[����lgߠ�}�I���,[�[�T�bkQ�+�*ض�1K�,��cI�z:�
�<ڬ���M�ӮM�,�+Z:W�u}�jS�6�+o]�I���[�<lC��mv{�V,[lG~�-X8ϖ����ܿlRb���ў���c��_�L؎��홧�Խ���;��{���N������/���oЏ��AKY޲����鱑1���-���b*��q���G}����TӘ�1Ƴ���!J���o軙�k��<�Iڥ�\fS�P� ��Z�ys�jLC~;ag�}��:)�uy~�K^b�y�{�����V��4]�T�_�R+��	{��ߦ�:�8�2�[����Fm���������!B�!}����5�:��õ������FF����[go{���0���+����g����?�oCC�\�l�HE03̈́����hxp��E]d�w�Y�A��MZ�.m����鱟_y����Oh/"�ó�1�'�t��X7@���[2-�c���7��}c�R�8q~���/�YӞ��>���hXB͞J�-��3ϲ_\�K yz;������������/��T����e4����׿���^9�^a�h_��/Y�sԝ'�Z�T���~����J������W`���6gv�*X���ݝ:ϵ3�>��	q�Jƈ���=�.��+җ`�dO̤2��g�<��dì������V��|ݎ����c6o�|��~�,w�Z#H�ܯ�~������Q�
�}��BD�<�a��S�t([�s�J���N;lr�{5B���{��~-���;11�po4�-�d�?L`g��H�M�����O=i�c���8�/[�M�������:˴�7��u"C��^�ˤ�t �@pcs\�`����j�:�"�%�cL��0���]
��=�y��0��"v�iT�D��*���P��v�������D`D{�e���H��=Q��x��kY��ɀ��EӰgĨ���,W,)w>��Ix��v��Y�\���ꢉ^;:�V��[r�t�떨���Ԙ�tw�a/|��ң��~3D-\c�Ȍ���&5�=�&��6:2f��C6^�ج9=��Ï�c��Z��Y��+��Tض�����:�
-ݖJ�����6+�ٜ�]�o�����o�~����\������w��Ƕ�>K;mz���!+��V���N>��v�����M�m8W"k����ަ0,ry��A�æ�?2*���'��M[6y����µ3p<v"W<Y�=D�f�*Gĸ�ܾŞs�A��ם����o�َ=�X��> ��iE�	��;�-oy�"���� 0�!��n_�����r�ixb|���a>1�0ڷ�~�%�!-����j_��W��AX9#�c�Vj�s6��d��
���7�N�=80l����1�c����(b�;�ܝ����`3e�6�è�w�y�3��9��#i���þ����Q�Q�T�UN�	'�����U�i3�t�-��?���v�?�ȀF}�9����������Ο���T]��M"�3>�ׯ��o��U�Oe262<dm�a��) )`/a�	,�0�S�&c�����[o���`0V�ߕ+Wj<����\L)-Z�&��?���om��w) B��%�s�ى�~�-_�Ԇ�Fm2jF��Ɵ���;���o��_�x<�y�3�l^�1�^x��!0�$S�s����^۴u�u��Y���J��Z��*{�_����0Q/s'�y�%c�zضmK�qT��`�.Q*��c'UD�G�˓� ��Iڣ=�u�,5� 
l���B{�ˎ]�@T�{�I�����j8∣l�A��w�m���`��sm� m:)�+<//z֞A?���W2Tь�zJ��rꋞ���Y>��Ͻ��o�(���<rT��	E䮷¤����t`�rs���=��#��Lt�;w��榣Z&h�9S��0�󐛟y����3Y�K���EDl|-��"���$�cc|�����dX`��d@�r��N�u�w�Y�u���'y+��L���h�<U*�nJ!/�}�} ���,�tF���p�L$�I�2��4͋"�m:Y��q��ڕ�跉�!���a�YK&�IY.]�jeج1aGy�������'K����s���u(Îw�x2���l�'���Mv��j�㟮�|���;�,��f#�S���~��ۭ¤��    IDAT�:�ҙk�c��I�a����v�q�m|�l͚mv�E���[&�p��A�ӝ���qء�����f��n��8�%x�i��<�.�7-j)���=c�����rP�\��۾�W-d)�?o���Ҹl�K�,�[n�E������Ѐ-]��V���x�>�%�݈������택�f��V�ͯg��)G�9d��x���5���U��w9!������z�z-�Fr�'pvҖ.]n�|��r�P:$�c���R	e�8m�R���W�P�&��Xy�"�s��w�~60اTd��JU덊8%8��C���Ï	�R  �([U��_p�R��*�(]�>��|t���!P�§�*e;��� ��#�?�*d���f�=Vj#���6cɸzi�7_�4��ȹ������P��\� ��r�?�F�3�M�4:>�n����.����oO=vuv��'Rؔ�bE��N=KZ�T��;�p�[l���6��GC�Vj�j�f5D�����d8ps��~�&쵤�@ �X�$8��3h$܍����Fʣ���A.�[Tjk�jeJ=:Zۭ��B"a���o�X�ag-��0�!�2# t��M4η;uBy�)9�n�IyҤ�fR�%�"}r�@��"�8r���K�i� ���D���K�I�s��ۃ����xX�9{q��b��̐�ºBE:��/iV��t�@"�����?�����������SMp�r&�WJD�,�;�f�d0���������
e/����kR|2�QI�k7����ϜGܰs<7�Zl������7�q��#��#�W��ǐӏs�ݟ���F~�U��#����j�-*)z�DT*j�P#�,��YN@�"JO+�~КG/#�\��j�B�5�2>x�\�2�i۶�i�f�Ҟ���&ldp��z;�-������)���D���,>ƮH瑪��gSd�"���m[�ٵ��6ו��g<������LY�r��?f�D�f�,6K�go1�*�9�m��h����5�����YWgɺ�3�uӣ��{��o�#;��h}7mV���Υ�\	�Z�Qo��0F�ǚp���Hk�YhMu�5Q�<��_ߠ�U����u*'|���ڷ�����T_��y���&�e�&���A2��&"�1�fI^Ƥ^������*�:kVWS�F�]�yx�{Ф�Z�{�L���<H��ym�}}���w��!Ig ���j-�VA�h�#΄��R�6���1mȡب@gg����o^��
Ip���ـ)��[W}��V.s�*z��9��c�o��SA���o��mB����M6j�CKc����ުSHX�+r��b�X
�T�gBN-η�y0l��>��-΁fB�<@$٭;�jB���A�w<-�ga-�m�pV:p,0Tp���CՆ[P>�Z&��:�V��P)o�;���R�^g�l�DO��:�5�e@ü��c�S�f9EA��QB'�F�6m��PL�"J���F����O/rc�6x��&׫|����a��\$'�[���:5�
"a�tV�-����MUH9��V�֦��J��j6��e�dY0��E۾m��4�:]�f�̳���ƭ��G׉��ݤ�T�R�31-9�r~��h(���ݠٌY
t4k�Z���5R�|���n��K�|n�0�?�G��!n��M@�DΠ��;���8��7<�N�8����9�#h]�ƣ�6���7W�+�E����H��aȌ����x�(=w#�����įsOH���;�`�eX1��c0������Z�e���^2�c��ʩ�3�<x�ne�L�����蝎d4�!b̧�}�F�u��w��e�{�ˏ�w���l~�խf�ccҫo)�:� \v��z�'$~���o(i��w��)F��Vľy�6Aa�n���s-�i�����l������!ڨ֔�{�k_+���O
2,O���X��2U{��V�kN:Ύ=�0(�66T�驆�9i��5�y���Qs�;>�0蚓4�!%ӻ��$r_6o�j��v��{����'&'��3�D��
���+mdd���Z�?*'����{�����؇�f%0��vv*�n-����xS�Cd<����"�rw�Z&��Z O���dRH��3��m�3OdCSr����!���8:GWo⅋�Z/[[g�xW�_�8���I�/7`���.�m�ҥ���G(�;��k*M���ӵ��c�jՐ?N�t����@�s��|��D4��P�򰀠��r�q������C�[��8Y�2&/�z��^'�����^�uI��R�&��7���=�kڤz.]�Q:��0@ή��qb��`.��a�x�M���(�#��ҧBkUwʕ�Br;rd�W�;J�\�uΛ�C���ʱ�{��/=#�.��:�Ϥm�0��Q	���a���q�*Ý"'c�z�:<%��=P�b*�F��v�Aϵ�j͆��l����'�W*N����R�n6�jX.�ٚ�x��'�u��Hg��-�Z#E�^6��u�玽����dVS��e$yj!�3I+�zd2�Aפ��l������'�������,f�	|#�O߰�k�?6�J��A�~l�1�fc	�흭����\���ռ�I��������f$A�އ�i�#f/MD�f��`*&�Jeظ��{0�L80��|�4�)�?jҽ�ʄ�_y.��F�l�t�:�KV*�mx�������;��V+d̶o�j��E�P�9�f1�8^�<���Ę0��~g�$_�b�)�v�z۸�ia�r0��\�ML6lpd�Rɜ�
K��������[m��mvO���)ٖ-����ڇ?t�=g�J�<�H����>+�5R��Y%F��r���4��\4ȵ�M�eJ���7w��[�e���Ӷ�� `���٠aS�������~�~٨\�˂X/8��:��9<���:S#�Q!��艏5����,)��MLM��=�J������E<$��+���s c�\�D8!�X�|0P@��N��$1(�'�5��;Q�7��s_���kQ�$ 	�Pn����`:� w�~���-r�x�Ѧ���-��0�	�����:�6o9�pz����gy>��Бv����]�nh�ߊ�B��fBjG$��c\H�8�2�Pf��Ip^����07=bn�Q�T4��|}?�X�f��sF���h��w>��)j�!�^����k~ϕ�������k��Qb�kk������v�;�8���	()`��ݹR+4%�=k�ۼu��OLV{d7+�VDQ���Z߅>��%�5YQ�t��W�|��Y�ت<�^��Q���������^�J�V��
pP�@�b�b`=��A��!����}�	K�ܠ�o�v�CN^^p?O�Lg��
5bn�,�cnt�ДE�B}�{k�(ϿT�'�8�������A�#�n�����E)
�}�@��58rx
-Fu�
=��}�A�����J�Z��:zU�S�.&mV�w�,���j�m%�S״O<��8�߭�����~��խ����A�v|g��p���_�K���� ���C:��7>c�7o�|���>+OL��7��dJ���#C�mۀ�u���%�WX!�fmm�62�k��ڝ�l�\�Ĺgۢ��>LW!� 7��Cޮ<9A�����/�ih�F
�~.Ay��v0W�U��~ɫ_��?�SO=�tQh':!�2s������;�����q^&�!ʦ���F$߿�O9k�	�5Р�]7��R&���Q���k��3RM��� c@�97\�GV!��%����6M	l ����u�׼�Sb��A�\�3s����אG�n��sHH�5�&�$�9��fpBpbú�5>�=R�*#��2���z�S{,	{���~d��4�����G���]ʔ������ż�!@�����-#_C�7���Wia�v�9��L��q�/D�Y�9o�Ü"r�\���l���Mg!
��1�aL���}�n:�1�^��Qr�bW"E��U�D��+\���=�〳���w:q�m�;A��q$���ڏ�/�G�������_��6e�A5���4P��1�Ц���1�/�c��hF�p�6BT&_�D�m��O~򳯸�뿘��W�^ͦ�*CaCp~��K��(���0֮_g��`�8s�Y�����q�Xt3�{a1����s��,� ��"HAq���:��pMN�E��7����l�3��0�
UbG>:V��B3L@:��|h��bTW996�X	i�ŋԵ��%&�Ԧf���<�8�r?�ڔ�ѓ/[>k��>KT�?6�o�{��y�-�O��Er���≄`�9=�BA��� R8��'��k�[	šL�Z�m2T@����=�����u�Rο����u����Y�2�=k�eS����ł����}���n�9�նi�F[�p�f
%g�d��G��R-kx4���Q��>��@�h��z��?��>�+�;ٚ�����y��frp2*������ x� Ϟ=G���op����''HY��ggttt)��p�s9�rJ�쀖E�>�(�I�2J�п�E\��zJL�C��,ɡ;%`�JE}�A��dLo�t�>"t�Ux_���qr�t�*���>����Q���g�A�"�pò*�׆xSww�I���b�)���T����Q U��-㜀8�`UN��܀�:��"�!Q���0.�.#V�7�PK��C� k14p�!2N7;��)�ReR���x�����y���b�1v'�p��������:���������xnd�7JR#8|���nw��\v�Fmm�nZ��5�������J��$�bA�>v<�#]�`q`"'��^�����q�>\S؏ܩ��➤3!M12jT�QYŜ�G�'�&P\D�#��g�}fKuB@�u t�^l?�Tq��ں�Xy:-��5�Wr�D�8�S/��֛���޾*U�@vb����V����C/�c^�#�=��Ơ{��p7�)��1�39���65�#�FpW����|#����:����#��~C�Qx<:�=R�'	��0=���7��!_�� �In��AM�rSH�����u6�@�<F��!�iLU�T�����"��	A����׬P���V�R"�i�X�TY�1U����w$C�,j��a@8O����Ժ��g���ںm����-۶َ���?���X���4�9�T�Z`�������m������_��X��T�F��r�B����2Em������s�,z�܇ 6T�� ��D�䓽-f W�tHu*lbO<���p�v��7)7α��4�Lh!�a�m�}Z�d� V�uVkJ%�� Ёj��կ�7����o~m���U���v�#l�D�l�aQ��x�u��,���z�%I�u;���:�0��o�2u�u`w�����jL�I���+��w�R��'�����ϤlldL��ԵCb�D��)S�u�8���.z�|��@1ʐ�7¸� �x��&Z�^H� A)�BP���L(Y�㣍�Ȭ�Y#�՚�
E�OU�s5�VVA�_ZN��mn4�OZ���H�tth.y����%t$�F0�S���
&����&ً�r2 %N�,�MIϙ�"(�i�#�<Y�d#a�R�Z�%�A�	m�A+�b�$�]��_Z��G��:�HX}lB{�ip)pU�:�q&*�I�gH���r7iuD1n,-'i/���4+���2�i�|aƑ��(�Y���EU�,��w�X'ڋ8�d0��-�#����	�Ad��#%���$�&3�������͟#�M��p�Z��b�9U������}�~�9�8���o�B.�]%/�Jy�x�N'�\�v.���GC�R_��.أ^>ñ<�ozlʇ�`&B����XH�#��i�Ct�=7���<�þKT|�\f�`sD�7�qoW�����r$�/(-<����;Ԡ�o�?-��MTW�Ag�QϝL�"@��/���h �'��56��deT��)ki�Zmjܾ����q/?Zb1x���	��3�p��rEH9�r�8'6#���G�э#�EQl��dh�Q��#�AI�n� ēO?�2���|�l��vE����p뚽�n��۱e��͙c��	�����=�����W��E����Ȑ��| �W���8�?�O�SO=a(�-��@�T�TBf���p���5��AP�Jg�����9�T�"���G?�'�|R�H7U��h�*�P��3
���R��3g�mX��<p��񏿷��;lV�,{�O��|P��x���w��˝��|���)Q� P��XZ$��h�ލ�|oԒ��ǉ2�=={9��r"���\6���B��͏�߻_�t*B�FG�l��e����~��J��갣�:Ҟذ���6km)ʠ�1Md�I�\6�/�?l�S�Qw?Z���ș�	ׂ�!�K�u��%���1������s=<��������X�*W��(��"Db��V9�$H]�s��	e�����_�2��7��S:#��`�������	ֺ�c��C���I�ҧ��lmR��DdJ)M�	D��8�z4-<������TCd��ך�=���~fұ(�9�+|��/�ݛW�,/"3NQ�� �c*�?�za���rZ%���w�a�[WO�m��o�\ɦ�mR�d�V��8��s_~�Mw\�Aw&�,�ա=��=��j����ckk�/LgQbН(G�--�ߎ���EӉ��I9D4�z0�@�Uʰ�Vj�{~�߳�M��Y7����͏���2��?t*��#ڐ�H퍒�f�Hq���?����4#��')�C�cP��#���Q��H�9I{K�&+#�Ϙ���W�9�e�]�!����T�{o�A��T�/�A�i1���Ο?_����K� �D�ZzW�˖�pn�^�Ɲ};�,nuJ�5wڶm;l��(לLf���Mo����b���F;��#,���!�_eg����v�r��m�vE΅b��9����r�:|=����x���d���f5��ܙ��R�omm��g�ŎM(��fB��5���h
.ɩ Ǜ
d%�*��p0��jHw0�)�\��~��/}��̝m##Cv�i����<�$&q�`���#c����6hI���{�;���|)#���98
��P�����g�ϩ#�6�`���*f���=��9�\���#�ZY�l���y���m���X:Y��}�=��C�u�Ӗ�W5�!
_�d����	N�L֬�g�-X��͞;׾r��m`d̆�&�Z#j�26A�Y��qܠ̤h�����!�HU�c[�=��ݐ�I�;���V|s�S����w��p�0�p'�%I.Xޤ� �ɱ���Xώ�F:{��q���!�q�|_ �b\Ik8"�`�`,�C�,zRO�4t�j��G��~��):n/<�Q/�	l�����#">
 ��Io�&�A?A��-T?�~�-[b۶o�[��n���WZ�X�}CVGų��ҹ�hй�s�9縛o��+�НA��7r���χC�j~���6�k�`�snН$�{<*�^��g�n�Xd���-�i1�������č�G)��L�Z<�ѭ�u]�}��S)�퓂�ߏ�1輟��c�)Ny3�t.���d"^i����4>�A�797Q���	k-d��3�������ll|�ZJt�
�+~y/e�i�v0�3�?%��y	*ߺU���">D��L�����hC�����&c��w�ޏD�7�h�>���v�q��_d�;��7��{l��s���p[���S����˥�6<��ڂ�G����*ET���%�9b���o����.���;�:poy�[��^*34_y��)��>�;�A#�`xtD��㏯�v4��@c��&-xm���!ң'BE�?�����Ȱ���9�(�я�=��#�sE$Ш��"��04W�b�+%�;�'��a^�<t0��>��Nd��y�����E�!RQ�� �o�R>g�L�N8�h�ٻ�
y�v��U��}�X�-��pv���d]�lGo�-X��Vp���s�������w����ќ)pz�Gʕ��G�@�aQ
M��B�h��G���E�w��<"�7W��    IDAT�r��A��!�]"Ԙu�=�S���/���ݐ�1L]o*ڹ���4葡��|J�\=�M��e�AK @�I��4��C}�l�輧]%�\\B;8*3���%0����m"!1��t�*N@���`��q��I�"��#��2�pz�;5�zw�k��y���6[�F�����ދ�#�~��7���|>��	 6�O�x^5�s3�g����X߄����0q�l������l��rw�=1#F��3���ڍ�O�g-��㩀ݣ������/��#����Ь&t�c�c�1p�����[�'�or~8"Lɳ���i#^/�F�Kk�h��9Ϙ�p����K� x����C���(�*�>���4X����#*�;�C;�V7u��,	ģ��[�.� X@��~��P�J)a__�m߶E�����v�=�q�=��c��Ҫ�x�O���m�[o��^���?����Gϴ���$�w�m��'����1_a��DB��W\!�: ��:H�50└1ƌ���XӠ��I�~g�J`�o����,ۯ~�+�����D�N�eG��#��@��`������Tb�2{r����HTI�MِTC�SX�!B�7lx���a]�E�@��|r&"�HY����cJm!������}�5��J�P��9m��f�H0SX,H�^�����߶~�#v�=wڡ�bK-�����k���y�.�̡���n���7`�j�v���}V���U���%���4+������P!�B1�?�!��)��6�Ȱ���p�"�h �H)�)��l�<(j��{�Z�M-����8j�G���?c�B�?�}�=�Hd'
�|Od� �Ŝ
�h�B�.Tn:�P�)��+EêL�?R� ������H������S9	 +�@��}���<S^QE�N$g�G� E]�"�Q0tP��TH!�MU�K)�-X�Ш�9JY�ԡ�Di/�C?�s���[/���=�j��t���'�\nTV��xk�3ɡ���C)�k8�N��;��ll�e,;%w*�|w�4��dO���#���<�@��G�pk�P����@�;���S��D�2��A'�.�Od	''Ր�\,c`��OM��^,��>�Qb"_u�b�4��iR��{D��A�U+���\n�8�ejBR,�{� �����81�C�C���*��NQc�e5v "���_x�΃��8��f�-?��s��[���m�4끝���'��[oY#E��s��)��fk�>f���;��c����Z1#��g^����a����D����ۥ}��_�Z,�V��C_�°y傐��< ��  �J�	r�[�n����7Xa!��Q�6k��t�M���H��b�ר�E
Tڔ�YK(?�w��.H�.i��s��>��K>5��Q�*M��M�En,������w�]�G�('G������L��3�aOس,���szvy���5����i{C��.ٔ�++�ۗ��y+��v�9���JĹ�a��+�N�����r�/��A�����Z	�jݶ��K����Xѐ�t�Bbw�ĉ��&GG�:pܐ�z����!�Ǵ���aP�l�o1�7�i������p��	�7�ܮFj&X	��N�U����cx�PȰ~�,24��U�9n�=B�A�CʋH�Qd����Q��=�l�͓�=%
&"��K���ߤ�ݠ{�b��,BT�H�R�3��|e���{��l<
Z-ͥм(A��NL�`��6��A(�[9t.���{��7�ri6�;��5$�``C�� ��$c95u���A�|y�Б��=*WH��מ��:�u���C�>��	��Qozd1Hl�h<>���l|����=��;	���{�]IK���d��4�IFz[{�r�2�Ţ����M��&���6]���ļ}�;wR����b�#��R��o~�3�w���N�n2ec�L
�(��� �#��A)��gm y���Ԗ-[�T͜IT�e �
"(AG$@�3�t�)�3�cc��3O
�^��	��o�Q���h�r���z�[m�k������}��7��[�x�Tj��/+�C�;����x�F���1�+���Ƹ,�Ҫ�tϒ���߫����7o���=��0��������< �Cf��K��G՜Q* �@�@ZD��HF0��6U%U��Q�&KCu $"�B��T�I6V߈f�%\���vs]��g;�3���􈯋ݍr$�w�.m���I���!�U�3���-�ۚ5wXg{Isi��N[�h�-Y�جV!��Zz��xc��ٸy��wu�hyB�p�Ԗ��Q1D¦4��DV9��HF\)�E��r̼_^���NЊ"���Ȩ�S9��A�G(����Q��Ս|:*v�:w)Úi7�
"�h�i��#��ϣ:�{98�in��aj
%�R��Pܠ���m�5Ƣ!�A�p&��m�#��.�%ʣ�)���;��en�Ȝ0�i׾�[%���`�9����P��H�)��b�M#��/YM�� �
)��:�쳏����/���:����%D�Fǻ��5LT/��[�~]T�>6A6~&<��\Q�{.:ܴ1������51�5�ͫ�}��("���	���=�o��?��O��D��ݺu��ҿ�rg	�HowV�lN�$A�ʂ�{f�����3��u���ښ�j��7k�	�kҎ�o�r�ڥ_��Xf����3� �J�-f /�k��J%�� G�=c�a�0���c���#��FQL ����iaA6�!�ܭ[�x�ي��7��w�i[�lS=�qǾ�FƇ��;�����Z��;�z,�$/U��Ĉ�ܹ�.���l��v��'�!�<_��G��bZJ*?��_�b�J���v�u�YgG��#�ȇ�O���~���|��U3�6n��leɵ3.������f�����T^6U���׷�)h�"t�� ,Dޖ~�D��Hl>����D,D2�H�NL��Y�W���T��K�l�nD��ƝҦ�TĊ>�*�˾�=�6m�{H3�9����������.�Zm\+rT�[�i�	E�Y6�ʄ�P���Hy�ZZۚ%e8yT,lx�	E��RQ�Fy?DP#�V���B5�A
�uz�^[_@6p�@D(�A��#"��h��ꑈO=�"% �P~�eW�嘁v'���se�A�sfN�#��)�m�n5	�;�Uf�н��L�r�@�.��]٤H#ڪO�0d����Qyrd�)s=�g�cӜ�Ў��4��3��7�l�
%� Jk ���>'#��fv�e ���B[o]s$��G��B��~��FҲ�9� ?�|�2����v��������/�{�G�r˭��r��`i�A�\'����;Z��1W	V�xni))���W1��h����
�67�~�8��:�1�����[��!�jVYV�"��;����=�]��Dܠ3���M��Og.DA�#�SY��ɢ�zۅ�͝?OD( n"�r��.{���H����o	�ߥ�9" �=dG#�-L�L>c}��p�;`�J�����+���и%�^[�~��e�,�!�0CJ��Y�0�i	]u����z�[r�Gu��_}�ua��SO�B�ݜ�5z�<o-�1%GO_d�ٍ7�lW_�A���W�ƶn�l�����SO�|��A�B�ϒ/ok)ػ��.{����V��w��^����3}ϙ�D��Їԧ����5'�'��^}�ډ�����~�/Pچ���A��q�3��a�<��!Y�ӟ�d�+2�R����C��fF��:?�ß��Ĥڻu�u	v(���P���� ��ڪ�B����FDe@�_M��H*9�(�(�����B������݄9�&n��<w���£Jr�@/%��Q���Q���H�p�9Ѣ2�l�$�k����BӐ�	9e}��I��q<gJ����X�3�g�b�QÙ�*�:82nĢ��:�g-�
F��A��U��z��8c���=�3Bo
n��f/w��d�q�HI8���7�����k�N�
7���)S�Y��G^s^DppW��Q�Ce�8�S����O���h���DN,i7���0����rŢ��s�J�"���EI*�m��"���Fjz:��9	�T�I�b�&���o�ZlO(M��zP����Yg�}�;�\V�VW�h:bFu�L��y�[�I&���ԈTi݇��Am0��J
6z��O�d���M�>�.j9H2��Bssu��-	݈�K�q �c�����ϻ ��
��ĉ"�E�H��������PYH#{�V�đtv<�����;�5�[��9=s9?��f{�ɧv�ޤ����J��j4�կ<�>�gآ�s�@W�D�|^s����]"���S�l�w������d�ÔS]��_�e�]&x�?��?d�?����g>�	�\|��v��G7#y��Ѐ�+�'2�;�� '����%�|�6n�l��-�#�8�}�1�����O��ș��ɨ��v"��O>�N|�Ծ���>�tF�k�w��u�Gy�}�#�����A�y�f{ӛ�d_�������?�#�8��p��A$ Б;��sp`HML�����/�F3�G�Lэx`�+�ěR�$s�J�:�T"��=�΄nN���(u4mƩ��F/�# �����2� +�|W�t�M�L�ܜ9rX�֐:ŕ��WR��;
:�ȕ���:�*�j>�6�Y���$G�jET2цXHHE�Í�p��C��7lR���r� a�"�]]$��F�n��R(�濺�)�����1˶����� Uk)�΋Ac!ŪSA�(�I���XP[���dĢ�wY ���J�ҘH���H�D�]�����>-@��� ��!�i��F��j��jMd/�Ix3"�
�IWG����(�P�[Z�"��<�}N�M��.ΐY�l���h~�MP�d
�`��t_1�㣣��٩{H�a�����m��mo�Y�ݶ���R,��Y:���ܜ!~��T�ΨM0{�*l�62��L��O	k�m#4<ꚭrR	w!e�3�0ٰ��t�Z�MUR�d��0��d9k��t:�,�ꉒ%��L�X���gqz�?�Ú+�	8�t���dp�5����g�y����q�e�db9�w	D����B�%_�'�̗l���|0����d����Ρ�2������μf��ݎxN���{�:����u6iw��3�(n2�R�y�$^�����p�ٳ�3&�P�֙����e9sY^u#(v�I�^5�4;�:�QO��аMV��T��@t�}#�*�c��1�/Y��לt����T/Mkj�I�Qn�������_��7����ى'��h���s�����?���=�\{��o'�x�Z~���W��SN9�>���i� gl�;��VWG���s��t�JƋv�\���o�^z�"�ŋ�ؑGe�<��q�mv�����?[�'^<}�i4½���7彿�ŋ�Ӿꪫ�(\�׿�h��������Dd�Gy�>��O����OZ�f|/Ft��_���qU��1��c�	�F2� ������{���\p=4�	�Z�֋"��Awt)��Md$$�~OѸ'ڬs9�� �Yk�Z#t�S�0GFe�D��8"�5E��,�����.E�9��R,��Ҝ����o�k��C|Oq���j�]�գW7p�_�Q�����e��K� 
P�c��K�w2��WĔ��7i4�\������۹>A�	�����������ԐK#�#ڨY��)�Ѵ�x��Ѓ�Z>ע��Q�;Q1���nu��Y�;�s��D0�Mf{mR�:m�V,)=��w������a�_�q]�k��yYb��~%uF��y����Q<�E�B>���lYmX!��Y��-�S
Y�)��z������F*�s�U��U���^���u�� �RnukV�`�c�d�-^`#C�
X��!o�\�r��jr�ptK����! �1U�Z��F:���k�H����������e�0�����m��Ŷ�{�p@獳<Q�v��l���H��{����T��z���}������d"3:<6�oht��X}�j���5K��R���T:	
](�$zH�J�8�:�&{�^1���������.-������˳G�M�f:��!7��D_�6�н�����W%k��$�EgS������>9�.RR���GP!�U�a�Z�;����N�إQYP�^�����3�\��ל(�sL����߶ozMX3���:|'c���p��6��ˠ	�M�Վ�D� >�i#��)2訹I԰ְ�_u����l�K-�Ȣls�ϳ{���9�l��o��������6%ʩ�9��6w�|{�[ߪNbD�D����'U�d��OVc��]�i�f9],|6<��u����elp`X�z������v�z[�t�����;�C���϶jT�����)�!́3A-��g~T�t�rm��q�	�6*�kzJ�/�x�;t��x�+D����[u�ѹ��CH�ײ����.�dt$��`�q�z08
�4?w�ݣW�be��2�2�IP�d�G��E�*]�)�0��J\�'ʇ$�R�&B��j k}�̳d�|�p��+ ��	eo��U˽��3&]�%��*� Ș�R�����{�(�T\68+H�����ǡ��⺅�C���q�)W6��'�[Z��
)��yH86X���9k�'HRkG��I,	�T���Yg�l��9h�^�u����mb��N;A��Q�[���a3z��\D"*�᡻r�>�X������G?��+�۶-�Vjm�R��8 �F��|��g`sGfH�i� ��5!r-��C�es���)�n5�h�S��,`.@������l$4���:\�dG��:���Ȱ͙7O��A�0��o����a[�h��رSץ=9r$�����R��*�\���]�����G��Ouq~�ϬY=��FykU-�7n�i���mW\�7;דּl��+'w�n-[}r[:���XH���ӭ/y�Q�_y��QG%"&T�翻���7>�}�C�/���Oɦ�ǌN���wu�n�D���v����H�I٫���q��}�%�\n?"�d��=��Dn����z:,��Q�y ƅH=@�rQ���������=Ro�����)K0�ΪG4D�.��m�rJ ��X'*)!��"�Ot��}d�a�;��%M䚹�m[w�����O�Bn�q!�A'����z[�;����ҩ��2�CC�R�MBw;���CH�S�"������'�l�,_��^���'7��"���>'�%X�l�6>�I��ήvm�0�1��Q����2������x{�g䌨�,����ڸ�t�b�|�@(q�_6f�h>s�]��w����`Џ:�X{���d��9��v��Gex�nR@�Cڔ��ݳu����huGs̏�{��CJ!D�I��8��XpF�l�w��k�	Oj$��iSĠ3n?�(�R"U	��ƀG�l����ܧ(�7�WJo0�Zl�R=i����;���P��Es5���XG�\g�����15����H�L��`�dD�2��Dnô"|����]����AJ4�c*u,
�w1���a3Нg�A87�����^C��x�j��Ü*79����x��i���0��'$"�mپE�.�wߠuu��x�-V��5��-v5(����Ҩ�)���/����q��"��"BoSʾ˖ے%�lld\)�<*'�4郃�Ƒy�K����{h�����+QzN4�#v���v2�qe��Q��� ��zs��Ozz�'�����t�snWt�w�@G���&��Hߛ|q�;�:Dz���Ino��q�B�,<�M��R�ȃ:�(@:�RNj�K�j&�f��P�5�*����n�+~�S۶}k-������u��;~����׾�O���������?^x�7u�}����{�!����Fʦ(�-�-ZK>�����>��5�^�H$�s��9r�:^��=��Z�L���wh�a�8�C��b�Gr����    IDAT�m��Q���g�!3#'�x��>����ql���^���$\�;'�)��n5���w&�q���a؄��;��7O��W��zab؁;�~#��+O:Q���~�s���1ai�P8Ǩ�G=Q�VW�k72�{����'oKϷRVu��/Zh��;m�]w�����uutkÃiJ)��X���Cy�Ϲ�ʠ]3�\����hT��*�Q�)�aT�#�|��۔�ƩY�p���W(B���5v�Y�!�J��&݋ �Nkc����8&����l����g�����T|���{�v�iB���8��:��?��?�����Z�d�>ØSg�w�7�0<���{�Sj���b���A��`E��]b�Aǈ�$ep R�Ȥ��g���J�Q�`dt�����L���?��	�WW��\6o��������C��]�>7�M%��,��	�tAy��H�����ƅ���)U!ʋ�:�%���f.�XKg���kr�X�Ir��M���@��?"�48<lm�-6D��5�@�TKLOArʫ��:�!�r.������f�L���[K2t8�LV	�f"�-��EFLD�640(��jh���Mӵ+�A��(�}�4�b����Q�Ż.:/�0�\MOU�� ��y��A�Dklg/�"�9;�6���|�I�sV��h��_�<l�Ã6{�����FkJ|�+��D��=�[@p�(�lXk�E������_��V�L��3���Do�~r}�L�t��Ĕ͚3����Z�P�R[+�k�:Y~�Q�|�������}�����W_}Ǖ��v��7�rf���ŕdv��tڲ�NK�l*��^5�k��r3�Ag���pyvQ�9967���ha��q�&E�Y#}w��ȍ�<.�����(ݽ�]8�e�6�x$��bg2�H����o��ҍ�nJA���l�l.�B������?4���Ƞ�GD�,�!�u��׿�m�(&�Tǀ�O$$pȡk�:�q�/�"9�W��{�O��{����=xr����S�~�ӟ�s�s��'1�\��~�3A�?D�tLc�Bx�ǵc���w_�� ==��z^]��Pj��9r�V�������Ï�G~�x�>{���&cI_t�B�s��Pi&d�1��މ�pF0،����>���=>C4!�c���~��J)�Y�F� C�u�����/|�6	�yt�}bD�#�c��@���)EE-����O����w��=� w��5Ł�Al	��=m�4�IH�C*h�����TeR�?�*P��SW�m�#�6w�������N�Azc��8�r��!E��.��ς�݆�b*���>1�#�8�q���3oC{�9P 1Y���d����Er�{c���M�X�����uvv�Tm�jպ�'sfϱ�;vX:���Y]�����h�"���l!k����E���!��γd;!n��g:iS�r�*{����ϧm��qR ^X����1vt5$����+�y��W��"%�*�I[H���C��"�,�9�2g��ɡ�f@��2�H�\_�}
��t������~��������ۂ��^6�P���`�K��je�J-�'�Րu�SԿ�/�j*m|r��u��J5 /�[7[[w��s�a�4utS=?�24���'Ӣ��-�T��m��&�c�!m5V�A��u��yN������;>1&�Ṱ���׼�������N�_X��n�T����_����j��_���:^C�
~E0�r��ɡ���8����4�ɬ���^��ݠs�պA��s&�c�=���ĉ��p��p���h�F]�<o$�8*=�G�|��i>�f�ם9�5/��8'�x���q-ND�G�oXq4��ϣ6!w:xCŹhq������{͌�;��Ë�Ԑ������ D��d'������;����iˤS֘��/>����ۢ�󬣵�� Þ����_�M�1!B/�Mb'����g��w��.��BA�41�ꪫ4�_����?��~��_�O�����'�}C�u�ю���a,O:�P�U�6��;v��!�aйGs�γ�>�֮['������K.���͛��c��p��)��>�1E����O��+��B��y��p���^H��`�cؽ��{��^�k��#<����e2�>߸���P����3߁�ߖ.��Aۂ��״N+�r�hه����Fj[���������ẉl���2Z�8��o �H�ٝ*��G�HRi�A"�N5��)��l�2w'X�rM�'������2�kZ�.CQ�Pe½ŉ<�c���$� ��֕W�T��^�*��Y�8�7�t������U�W��d�N�Vɥ�����Ν�v䑇[!WT�b�h�LF�g���p���ب]��_�u���
�mbwi�������������Z��))����G���R�X���%N2!�H�wk��F���8��@�J�a���V��47b)�AX�*	̀���=�pkEh*Ry��Z'�$:d���o/|��l��+��_�B{޼�s��9�::[�nٸI����J����z�G0�o~��^���q�io��?^��w���]���y�(�E{��/��;L�w��۲e���sy��zʛUـ����9�ß�Lz�=s��z���r���g���M����s����\&%�(Ɲ�K�,�SNy�-\�خ���v�5��i�.��jet���ƃ��w�����v�����]���+�>���ή�v<�@4o�B2��A?�3��������Һr|<��94g�����������0�^㰙H0�b3��̉ĺ���tҌG�>�n@���d�'�91�s���0;�E�è�Q^� � �F�`�n��i��"�t�q
��d�]��oj�W��K2Ec	k�x�~��a���/)gt���A	U�V�3|��!j����Ӣ�R�<� �緼ٖ.Y(�.�u������yJ�0��`z��J�x�t�Ia,1|�#����)�Ⳝ7�`i�(ca�sf�Q��b�8Y����m;dЁ�1�|en���O�;����Vڏ�#mҒ��&�@�� 'ǁ����e�9B2]t��r6� �Yg��(���/;�H'�a��D,���0y�|��T}�;������W_�R����*��Z�F�jQ钬WDZ�uf��&@�Q�\nS�`#ZA_o�:R�ɑK�� �å�P�Sā	�8 ��	T	T�hI4E�-�(�=���m*�1�jͫ�����5*�3��g�Y�� R)Ss���a�ONJ���}�~�]�_���/s��O~�#ݗ�����O^l��{�P��N;�>���ҥK�5@����~�#��e�_.��U'���%9\��G?�Q[�~�]�۫e�~�!v�s�k?����?^����N�5�EhF:m�����m��裏����V*!T����/604�ySOD:鴈����j���vk��$���G$px"ޘ1�����9�/d%@D��k�1�m�<��=�����Q����=����c��ן���������Y�4�㒯~�֬�˾��/��B����W�z��_�L��җ��>���{���ؕW\iK���\|����R:��;����~�[u�O}�9�T��е�uٿ��]j|�=g���)���j9f�W�g������y=���.���^���)0�����~�.��[��>�ڷ��}���~.�%�#Y(�7զF����ν���N�?5�|���}{�O���S�Gk�ʴ�j�%
�����3?~�m��~Y.��O�"'���/j��%l�*G�~6l��d���<B�=���)ʌo��f��s���g�����wэ��D��pa�E��<�A������;�Ht�p8�ʏdj�_m,c��A�;��A�5�^�!O��sζ;Y<_�غ:{D�
��GA�ٕD�'C7!]k.�\��j�b�{�)����z�:�ޘ���6E0R��1�����YY�t���=�Q9��3�LN�c���G������1h�s�e��������@BU���`�{E��PAAP���
�]�+��`�(�H/��dz���;Y���=�=>�9����)�s_�,��ޭ�T��*��+�=�9�͙/_s���l"���ZV^!��}��H�~ܸ��KJ
���$�]vtǆA��1��3A�Ю=�Ν+I�#7t�#+}="�1���K-Hy��mu"����(0U$�kv����u�y{aQ��	�_Q���������5��Y��PJ��ZDx"���"�%Y���@�h"�P����%=����`"*8���ziR��0T򢾶AQ��
K����j��:� .�ﬡ���h��J�w��I|��hg�q�4��j�3������	��ط`�7�k�9�\��9
����m۠q�^L�1m��$�:�\p�r?��,|�]I�֮[+���uLD�?�x�8�f� Fd˖-":4��+ɟN$D���̕����h-*���~=:�6lB��2��)*KYU�+Ľ��!k��}���/-�i��e&�c�
�����t)R�1e�Bœ)�1��hv��uײ�j��1� �J��H�����b�#�E]�7��2��2��i g�7�V���#��q�n���n�ʯ���ŋ���ob�o��C?s�t��5���+e�VW��AÍW^oq����}���fc������^��7^��'�UE�y���q�q'`ƃc�u�c�}(.m��F�$]+;c��w�h��F\��3g��a�ʘ�Ӈ��1�q�Y����W+fPR1�ҙhƈ��^=;ݹ��ז�7�9?㻭[�z��u��ݙ��+�n���nk����Z-qc9��uu�۔��g.^>@���TۧJE������]e]�����Z��\�Z�L]�H5xO���q�E���|Aa�E��!�0�C�M�|��l��骓��,=	��*L��q�\��]����Fca�s.Οg��dɗ�9�)Q�����{>V�2C�+��~Щ�^ֱ=|�u�:�?�t�V�<�n�&+��V 1�rz�G���R��!e�C����7˦u�q'H� � �ky�Ygaٲe� ��q�TJ����<�Y��5ջ��+@]����}���
Cr����>��6�>�A�˓�{:+���%�=+w�j��X�kJ��
�\8Z��g�'�ئ&9G���3i%�J�M�?���$B��9����Ҋd��x��������� �;O�.�o�3�$/9�&#�	�-Ҽ&Ǚ�1I�DXE��H'���Y�(�TO^~�~�T�w���+��f"j9�48b ���]���2a���ZI��=����צ4�u��D���2�*�H��p^�}�C)��Z45��Ǩ�#��3�I'бC\��2��ޥ2�W�|}�.��[�Fޝ���|G\ ɸ`�ƠĠʎ!��K��.�S��7_�.^o^>^��WW�̳��ò;��
h���d���+v1�p^������G1Ｓ +W��D�sq�;�J�[��t�DL��Xk��ʜ�k�p&rY�*�G*�t~[�ja@�X�P�t7&���׊�������}0Ќ��=g�u&��f���v����~��>|�k�ph��H}�љ2�z��Gѹ�B�x~^�����_��Eb�֭�6m�xP����`��A�ɬ����T���M��9/c�9�ԹR�ݺc�o[䙡3^QI��r�!�"�	���� ӧ�-�+�h�v��̳Ͻ�޽���SNǹ�]�=�;J�#�D��믾h�C��n�ot~�u3����꟟k�em�Ft��RܤI��^����k/"�u�ՁMs����ۚ��^ �7���aKZs���tk\�r�s�� V:��9���Lt)�[�<^=���芚�/�΀(�Y�8~O��������5J���y�w������"J��}Ὼ���Z}��v�|��Νg��-z�_���@:=����F�2&dL��20-����/�QG��N@�,����\XU���^8����-�8 �� z�����İ��H!o�J�o���C�6Xy=D��h���}�I��1;g��96�:��*���C�s��,'�C?\�y4��g��{X_['`V
�W��	����~~O3 x�x��<g��ֻ���`�����Z��=ד���-�݉k��A��e˖K�!�GQ�f���BUuL�.7:v(~8[�R-HwR'��l.DH�2)Z'���R�<�b�)Q);��c0h�<:��N�y��!�t1�5�(a�*!;��R� ee`�M^�_K^���j��R��D	��2�lCi+��J���]$�y�[L^���ЕJ(�S"��w�GS�^QR�Z�E��9X��+���<�ȃ�\����+��~�T��$��.�a�;}2Ra`�8�s�ƦzL�s�8�qn��{b͚52�)i�+�]��O=�~�9�^�.��#����V֜���!k���H��4L1����&)�j�X�Y�6�	G?�D4*�7�'ـ�{�{m$R�v�T$�!�&X�7� �r��f:+v�7���n
��=M�
�Pd�bFsM��q<.j����\�	��ŏ����1�
(�����_,��O?/���6����=�N<Q:tL�n;M�;f����_ ݷkG]��}�`������u9r��^&�8k������9x��1祗е{O9x����]X��[�c)��"x�<�Ӊ8�>G�SO<A��˗���oĨ+�De�����V���+F]������N�>C&��s�θ��S���o�Y�~Y9{��/V��f�N���k�6s�����U�|���b魜�T�FW��AOK�� �+l����?���X���
�7Pϭu�[���־Z�z>�[N�st0֋57�П��򹕷���uB�g�:H�&�=�znGA�V*��\J'��.��9`�օ�69��!*�q�#�����|k.|��"���R}5��<%����;���,ݨ�!5�v�����t�T��o�e���:���GN�_���-���vvuu���q6�`+�f~�$���2����G_�T.��4\������9��ի��/�z�p�r->X��l�s�'ʚ�pW]5�f=����V�8��"��ب�l���<?~�����geşgK^��[dx���"uόh,"ׇA����~�����x)�7sS�o%7��Z#1����Ͷ��#�ȟ�8E/l�w�{��;���Ċ��%�)1�H���z��sp����?!V��M0׊oV�SP(�J�X&Or��L���ʚ��-�q-�p(w1̓�Ϧ
誒�{�-������%'hM���YL`��̸2R���tF�xn���c!�{�L�����~�2V�f�8i�$Y7�Μ)L���;G���_��n����"z��_6B ����Թ3���#|��b�u�D����hס=n��f�<y0���hBF��WϻQ���ZT�JP(A�GA�S>���p-��ȈO���?��ͰBW#vm���*�r�wDM��7��f�[*tV�|���F��\�O�x$��6��z��hWR���|8�f�}y6�}�)L�1�;���Ũ�W�s����G��O�)Sp���H��g��������Γg���ݨ��:
�_p�6�q�[U�~L�>M�p���}}��gpޅ��!�c_]n;�XUuu��ۄj��D0��q�����KQѩ\Fv��v�\���
<^7��؋�wLB(JeLbKbH'#MCt���_�p�.�b��^/�S����L]0sR4a��?ЧY�j�&���V����@�.j���0nn��4׬�A2e>x}�&���`�������V�7A�fp��t����xt"׭W�?�2�Q'L�Y�+����s}�脃���M9C�$j��f��@��(YF���о}[�����࣏�WP$����Eu}<��l�ՙ.�����8�Xn[\_}=��ܸ��k �`��غ}�2	�J�r���x%Xk ϟ�k&f�֭�8�+ϓA��(Ap��s���h    IDAT�*Z�˩����Z���J2D��u?�F<��
h�xƬ@�	��L[-�?_f䜗2��ضM*k�(�e�E�<��{��+�^k@����w���@f�N�2��"¹���`��ɧ�K�׎�[Ye(c�j�Sn�&8]D����G��MB�V�L�2l����`�<�TQ#�moS�>��1t���H�	����/���m�)B0FW=#)��/5z�~��NYX�ڤ�KdR�h��6щ���]=���UKX���yk���.#1�e�
cF4�V�ԡ��ԓNĸ�7�M�Bp����?�r�f�7`� ̞���n|��8��S0w�c�>�9�}�e̟?_�2������5W]-�(����/||�1�O���}{����/�`��WH%�[q�(ͫ�-��6;��s�:�vB���d�y�й�Z��ib�%9A��0���Wv���["Q�Z� )@ֿXV����l�3Η:�j�R�c� G��]�7t1SR��u$.��B,�b�\{�CW�ك�G����Ʊ'���n���v��O�)������g�~��<o���s1a���h�|�%��ݍ�/�޶m�޻���`աg	H� ��C��ُ�^GE�N�|_����㏘��#���K0f�X��7�u�أ'�%�[ZR���j�3q"��CO=^��~�5F\~-v�ޅ+F��U�\��[����F�I��r��L�W�o����s�ճ��[�_�o���Ӄ��x�5�������[+�ɓ���o^0}X%p1pȥ�� *��Y�����0y���{�شB�~7W�*`렭��:Y�U���=��s+~��?�s��r��ue��n�k ��Xe�P�@f?���Dn�Ǯ�凭�~ u5�/��"�D66��0�:����K>���}���
�WT*3�]���fsJOP�9��
��Bi��B2�1��ŐF�>�,�ɧ��k~���fU��j�V8�xN��h�P�?�*G(���͋�=�����cT��Y0w����5�]+�.�ƍ��'ϛ���t���'��l��4�;D��ggz~��?]��1"�RZ��QS���xL<6qI��<�=g�ɯ�O�o��ن������A��g�2����W]u��9��9
h��=� J��� ���6j��6L\ںt���b�;��GzM��3��V�W��P�_TX3��,�� ��]�x�g�:�;\0�m���˦m+mg�
��̂�G�6)n&��J��U��JVV�I�CWk�5��v����*��t�E�]�ٍ�$�2V�8�h��p�����SG<��â���d?a;����3���\��s����� 6�m2d���	�����p������ċ����&a��{e��-m']��R���,|�=쯭Ʊ'��Iw݅3�8S�]�T��i],{
$��b�IMs�hOAM͠o�ūx�4l@�v��"�9� R>��,N&��УHP�n��aǄ9�*VTB��9�a�aE�N"/�@��A?UY���K��(|v
����Ǻ���?Ɔ�V#�|��rt�섊����kx���0��s����c�m�Ģ��+���Oє��oźu{%Q1�|����`�P��z��M7M�I'���;˖��I'�_6�.�Ε�;�.D�������vq�磩��=z����wv����p��`�ͣH�ނ�s{0r�yX�z&N��ӆ��zS��K��F��UÚT�W趼:獧�9���B������3���PV�������6g9p>��ڬ�t+[�ƹa����_6H��2���ZW=7��Ur��Ź�N����Z ���C�ѝ]��d"��g�U5�9�$A�4_^'��y�q�~��{�=����**YY}g�M���oݿ?�~IY�rv7�*�b�νh����y�X
�7�7���U@��YmF�8�u��7!��㱇f�sE��{��JQ��e�b`s;�Ч�j��X�+����۷�(8�Am�X�y-��T���z܊������G=�H\:�2�𙱋HOL�ω���(Z�6���M:>D*3��֥��=9�g�ۧW/�3F�9���%`3��sy<?���PW��:Ya�ª_@l	�	
�-Z�yy9W����W��8�7�e�
��TNkY��t�(ݍ�����͛D7�IT��=Чw_̜�2i��|��#Ɍ �2������v4����B�=q��E`�|i��u��Rս��bX)p���$��v�����U�.�h��M�3/A$ӊ~��U=g�Hk�i�X����JdU"r`@�xJ~
�4	����ϼ���x�u������sg�p��D4�D��k�)�ֻ0h�$w�PPč�vr�ԡ� �H�㫄\U�b��*쩪J`ܻ���N��xP0C���u��HNv�i9>ۢ�B���	���N���1�h���M���̿�Q	褐r4��� �/�䖋�P��&��f@Ϥ��GA�4B�#Ȓ.s�wѐ7#�N���M1��vmJ���՘��x����6�С�#�n~�m3^����O)�/�H�7zL�6M�K�O6o�U�g߾}d�V^����E8j��e�`�TC��^���t�Q;�GO\v�e�X��kt,/Ã�>�R(��h2���&I@y��?����"�\X��stl����w��+����߭�����d�W+`q8KQ>��)2�_z�޻�u�2��/���li��^}����yl i4��}ڴ�\�b%���p�r!��5>сKg��z���*�lC�r�ݻ�E�T(�v�����ٿ
���-�ߓJ��*x���5W�9)HKE�`��D]s��\�)R��� 5��y7oTe��<�UJCm��4���Q��rBYʐQ�zY����ओO��A$�%Kp�e�f�wR�q>�JtPs^-(�,KK�f�I�-Fx�6�ݳS����}�~�3f�/�:�H4�JK��ܢ^�*FW��1�a����o�z%�N��L)�)V���:M8{�V (v����N*[��F�:0}��r�ާOI$�f���i��*b1<������v#�[�p$�;OZ���������EҖ3i�*�@���%�2{���*ry66�Ċ�D�U 5�uF�Q�8k�p��~�j�2��+1�l+6B�2�^_G%<�l�}9DZ�_~�N<�D���G��1qf����b�7=�#Z�f4#�i�����aäMIu>�m2 ��5��g���� S~1L��A����,I��8�����,ۻlϧ���U��Ox�������-�p9��,�M��ZR�s��r�-Ⱥ ���9���m1M<�(,)��/�\N�����C�PpO� 	����5�.5�a۞��������ed#�bJLA��N0Xl�:]�[���TQ㬝k��ky��1�3��^G�!W���ԉ�)c)P���@��0	��B�#�5ˠ�.Z�rM	Ő�&I�Y���VI<Y��U��B~A�v����L
02��&�"�uQvF2�(��G��(/+�gI��v�.�G���>I�#^W#��
`從L���Z��y`�^��f8�ά��E �\OT~��r�c2�u��k�.$�Ē8E�-,D�b8�`obl�N����\�$�;�4���c#�E�|iBm�^I�ڕu��r��Vx�Ѡ�j�}n3���[�K�\>f�k�����33�����l˽�!}��8���_��)��~0-�&�f��^��T�����T�V�(1UU�S��Y�9�P���k�]%n!s��[��V���Mh}_m�R��5/�IS���ӴAP��߹�J:M�oe���լ��u���MCU�����&#rN�����@9BV��"��%_`��j��"��-3�.e�3)�������G�����&�y�{�HRt"��l����p�=S��'�PDǎ��E�����`�����F �<%�x�y���N�ͷ�Ə������I  � ݭ��REmߵSڞ����)S�Ȭq��[�kl��Zq�Ig%k��{mu56o�$nj��9;�9i���E�_ b7��O�2	�o�C����J�O���j%�ѯ�3S���-r�$ȉ�,i9C�A6�Dm۵P]CS���h��w�^�	<�p���W,��3	�|�	l��E}��!���k�J��U����8�裤J'ņ��YO>!UɝwMƌ�?F^a1�Km�:ڐ6"O"O�a��MQ!�>ݺW⾻&b�k�����N���LE^a!n7��b�N��m�ǝ���B����*D�"�.�)�)X ��DV�LP �\{��9�շ�uyM�)��t�v����:������YmMi���hWR�@]�$)\s��4�m�2M��ʊS�(�a��Y�u��SQQ)��{��c�2��׉*�^��c�?r�?����{G��<ʓ�˅H�|}{V��]�f��^�D`b� � �u`�,j�Ի�E���e�htkc�`.g�4�$��=PW/I:�6��$I�44�۶���21�&z�� �]X�2G-�Ѡ�hi��}��̰Y���*Mt�{J�({yēhWR� A���0��;"����NgD;`5�� �Jȵ�Ю#�����'�HRI��V��7�R���u�u�Zk������y
D�b�J�z0����{�ȳZ֮�h��Uҩ�"����k,+XD����w�{8)��f����O�_�R�'�F�u��ұp�lH�Z9��ُ.�o�5����>��uk����Ρ���:�o�O=z��?��n�֘��
�7����.^��lYs������>�ʯXq�U�J��x!��C�ϳ����A_W�j��k�x�	:�?��O�i���~O��5�@��uW���.�ȝ�����T Tl�N�މ�%���_�jC|��D��ђ��d����t�4����p9����a'�Ո��*�1�v\{�5�'�Xֻ���7�9Z��-F�����/#�2�P'���v"Zym8�mӶD�e����(�&���+*+�U�y������z���'0�cO��-�D����eK%h���kh}v�X�O�|V�\.#���}Q�t�K�/-�4
�l�����a�Ɩ0]9B ��x�U�X���uP�b*���6���\b��l�gu�p�QG�5cׁ -��+йKW���<4�"��] 	�b�;c��`�!��,�I'����y���ɧf��5?�^¤���􍷌��[��������p���51��'�7�`�=�'6��֯߈Ɔ 
�;��,@��P�Mi�K"�]iL2�M�EjRI8�!e��o��*�a�Y��4�H�i1#h��Yf����j�#�z�;���0�-�;j�s_��B���y(�n={�T�)�]���P@-�@Ɍ¨H!��� �3t!�/�`���]��.���WW%��v�s�cI����sLR��p���3(��TP7*5ǌ!%A���_K�E&C8�@�YC�={�!��SX X� G#f+�|�Е��ό#��H�a,AwɈ|�	L��I&+l&�86�#!�wĨ� Gϕo����x�ba��.v,k��wn��&���C�\Z�ND����+���h�� >Z�FC���xmb�D��핮%^W&/��eG����k��d��Ⴏ��hm��!��!���Az }at����2p�s#����]�=KJF�5��I��俠�D�Y�����8,��scά��}zx�������,0����e�G�LNg.d����O�>n܄3֮�y��j�Ζ;7:�u��niKk*k���������B���`6���s���*�ʝ��e���#�k��Q)Ĺ�����5�zn�A����3�Υ�x^���V42�漘�(9��(%���LT��8k��bT$�*�}�AW)�]�LD�v{&)2�l��J�k�$ۘ=�i�ҏY[�r>�y2��U9�q�T�b�Ç���c�Z55)0�"�"�uʭ^t�e�J&h����J�v(�;-U�8�(��M*�#��E�-���U�ˇ�3���,�.�f�Ģ����ɱ�3��I�|v��9���yՁRNpB�"Z>H����b,��e2��u���b�'����M\�a��g���)>Gl�ةdF�)?L~���	(�'�}Axϼ���E�3W�-|Β�tM�G�J�p�U0�?����~~a1"�V�#^xy��t�04���p�<<c@�ƛqư0��ѱ��ޘ��x{��h��a)l+U�¶�۳���R�� Q66��&"��T�	v� Ϛ<ь$��VyLޗ�Q�u㮱��W��h�ދM[�b�w�bޛ��C���ȚD��lnF,܌��I�O@7�޽�n֚5?	��neF3�if�9�P+���1l2���=�!����CU��i���2G���-c����J"����M�|�^&s���V[U�F��g`7�X[#�$��i{�5M�Cs}=ʺtG�dF�9F2�Et����D��`�hP�o|F����˓bgvJb�E``"�LO����ܙ�}	����j�ui�"�p�}�68\�h۾͑�� ��`B���"X(HDn;�Q������b!���#5���;�Ս>� !�>#Enl� M纠_��m��������ѶkO��hh��!��pP:/;2	8f	�ڵŮ��:DF6M���q_�o��d�i��'>�͙�?������?m-y��%#Vm�ut�&`sfn�8l`��'��y�]����秬VkwΆ�
W��50�t0��6U�\_	V&���![�+�����}���~����B?0��ռ��k/t@���K�l^��(K9�����<�W�Xw&��hz����߭^�%���mf�I0[���"�fT���l�Q��&K|5[R�{�r�J K�S׌}��H|ڬ��#�f�vZe��F0~�8�r)�J�������Bt63A(☗UT�\V.<�I�W����߫Q��pD�X�i�Lqҍ������x�b	�ܘ�3�>UQyp��p2��}��j�P�v��N;���Ҙh0P��U�y�ڽ��[E�}����}��Sئ��ZޫMyx�������A:��|�e�$b��н[O�����+�p��c9J��d����4-�����Pt�󋊥�u�op�r��_LV(�s��Ov��oIm���F&��8�f`d@/.ȗv�5�F`���f�A��z�o��Ǟ@��r�.f0��\���i3�Vܤ��S'�PX�F���0�a����x?o�O>�2��X���4�ҕ:�2�I�Ł��S�B��q
���`F�j=fpE<�G�=��b�ۯ	�w�Cq�Eg�w��_����'[�|��4�n;�����;���B+v5V�ًo����xP��P����$���,D�6���M���� ���L8Ԭ���J$(�i�F�mN�գ�[x�W�EZ�j��v�LJ�F�����ET���WW���eE�� G%ѤfΖ�n�	f��(T�.H��`P��ť�2桔3�ڿz��}m�[ś�~|��@ �; ��G]����wj/���=�I9o�3V+��Բ�K&`�`N:�H��!��*��b�l��@�;���m���as(�^&�@2���i3�� ����0_� �ITv9�]���������J�����Z��#�E�H'c�T�A_�|��ƈg)(AMm���8�6DC�M�Lp�u�^4y��Wl�_��?����Z��K���b�#��-eq"�$��H������q��X��O��VKw*�P�xc���1��4��Du֧����4����]���H]�ZK������	ZV�:��iV��>v��x:�3�kl�n�� �'�CW����d���{�s�~๹��	�g,-��)F�R%�
u`@���tA�漲�:�I�j���x8��O��^__'Tj����{����eK�4��Sl���C`Z\dM�"���?��6*���p�V%U�X=�j���fJ����/J�r����� 0�ה_c���9�    IDAT��N��]{Dq����>KP�8m]2{�*�-VVv=h������d[��e�����̞@��<��3�"���q�TJ�f�{�$L�����%��C:L" BQ ��T@���Q�;� ϘqcE�4��4,iz� '(nΜ9�Dq����X��W�"��2ҦL�H�H�Af
������q�ЭKgL{.��<\t�Ew�L�g*.�d���4%]�"n� .}��B��o�)��4�mI!�u��7܊����aK��1u����
]�0�X��fa^���f#�2��0�ˉ��ţ�nx*3ω3)�������=�4�zlX�=��=��#�t�t��U`���(aV��DRf�l1��v�))D:��co����-������e����(F�yk��"�.��d����y&)�{2��(ʘ e�5�#	+WF�M[ �D"�Y4��ʇ�O`?�k�	~=���������O!��bH��s�^p..��\|pO9�������o�������"�1��?��^�K�xb!��2K$SJE1c@ii;�V75�d3�X�4��wI��0��v��+q���]�"|���0���`0Y1p�1h��y�N�إ0��Ɂh$ �ÆX�n�����-]?>�Ԙ�s����>��p
�;����:_�dn�N+�k�B��
H�PԮ_3��y>N;}8���8=Ű�
`49Ė�ϜP��A�j���m��a��6�{e.��<q׫on��j�G�/�{�}�-O�_�*�>�������۠�f۶��?l����_N��h�/)����/A�` 3��������w�i��3�k7fyz��/�d�Ye.Xsy�|/,U����_U���[�ŵ86e��,�����\��:�9�它�n��d&�z��$�>�>Y^:ϕ�9��}`Po�����A]s���%(44	��l�ɃD�"%	��������� �
�dV�~f�>�6B�<Ĝ5\��U�߻w� ������Xl����ү�����`EPXAA��BO��=k�6mJd��ʝB��D4<)r<��
f��
O�Z�T-�Y����:�l�$jj�a�&:�\�1kHÊ*�s&#P�#G]!����
��q�:	�쎰j'������h]M�#5��3�6���V��@����͓�S�E��r#d2����?���k�nq�:m�i�E�~�m�J���KWb�}o��y=���px���aiS2�[�9#X!Y�47`���[E&��o�|'�t�9���f���;.�h�t�(�Hy��
LŢ��p9��vP9.���pT?�VS�����6l����$�@�Y��Lf ���#�LZ6bv?J۵Gc("kc��A��$�d�ԾO=<��~_� ��������A}�[nG�dG4�J �9�	�GVc��j<�ģظ~-�xhʺw�5@��|�9o.�[ޓ�)+}v}�͓�D����A(+�(�x>'���`(�ͅ�v���d̊][����׺/)Ъ֪B�mw5?7!�Մ�m[pɈ�1~�H���&,_�n��R�ݻ�}>[�5��q��C<A�GX��PcB�h0H�M����z��q���Ear�ϤMP��x��� &����6m��/�ڌ��L��<��S�o
�YϠ�mGI�T-�<��u�1c�d��wO�(��K/>���ʏ��{ޚ�-f=3AJ�效�x$��� i��eB�ne��3(��mkA^N:��m�Ihg�������S-k��C�%��:�x��X����={���oø����k/�g���?���Ç��[.u�m�/U���@,�Ӟ�n3&>9��Þ��̉�0��^���_���x��?m�:rGuӠ��S�(l�}u~�ld�G���oi�g2�	�oX��6��yê%��/7�����(7V�t$�Dt����i�V�ro�`�U���<7��3�����$�N�_kI���۪���h��7��r���׳wn#�������>r�m]� 4,~�9P�[�V'X�35��H�!�X�s��g[�Y�gnB��,3��i�tcgv&��s3�^��t*��ݵ9r�pKO9�T�e�/hh���- 
H�D&+�B��Ӭ��σmx�m�c�<���/�*��x�<9S��p���LUO��/�p8q���r�7�i�Z9b�p�_�3[�.��qsg%A�q� �sy��X�vءb�z��YJS��M"�9��v�Y�#��p�M����f�Z�۰^ާ2d�DM*�e���~�Zl���*߸��l�"����'�}��[�`�9�`���5^��J�N��?[����01�{Md��IO3�I"�M��q�)��A��������Y��T�W`���0g�p��#�6#n���FA�ǐ���I�q��p�e�ổ����[�ن`(�T��H�\�	Q��⬦hg�3���������K��P�͜��F�[��MQG��P���ߌ����y��=����f�zL{�q��6D"q$ci8]y�bhȰ2 n³O�D���q�:IdvO�����o`�{�F���x�3�لPc�N���*��w����n�_���u>����%YI%3!ζsv����|��C�9�� �d7jm�[4�ہ��>Ķ߷�kF�n3I@o�7�=��3q��q嵣�k_�JD�j}D��ba$���X(��y ;9�Ri���0���F�bB"����`��p��0�ޱ�o�X��b<��t=��5�A,Z�f>��+�|�K�&`/�+�x�!S5{p�9�/��eб�_|�	��1�{v㚱�0��+����/�K��l�M�)
���7�¨�N�k�a�f��ph�~0�I���J�Ǟ��;��\:I8q&�-e�0�kqx�>����X������՘8y"l.
ږ������xt�s(*l�P0& a�)�6 ��h���֭��ag��a@�~M�"����������S��O�n�QuFcs� �����4��0�T��J�c�T�����d̷�~�9�oz��t�tɦ�լ�1�LT��Uk��5�H��F͗�\��
��wɃ�u�@���Ճ�-C��wfƬ����!�=�R�Ǯ~�-�����;7-L�?y-d��U�;0	��A�1�
_"*� ��舻�׮fNV�l��l��Ue0W�Y�Z.N%_����nFa� ����m�`���*I���h��B�xΏ�l/��%7�%P����F���z�q&��#��%�+����.��?� �˙�n�2���*��H[ň`4Ғ�p^,�������������y�b1t�2����n��<Y��Α�:�H��P��#y���}�p���ٻ�&�̷x<pZ8DJ�?�u��/3���V-{&�q.��
� p����fW}�Z���xM�h������9��[[��	�x����ٌ89��AA4m��L�3+1!�S()�,��{'�{�
�Y���.]���ISp�mcQ����q�	��\�R�Z�~��{�H$BX��RL�s8�`̜����@ƞ��x���8�Q3�4���K.F�׍o��5?�(��]��Uu���/��n�p��I*�f���=�4�q�.C�W%�	M�a����n�oxe��H-R)��v�]��O43RQ	(��k��!�`��������"x����u�/n�&H�v�[�>�77����#3�A���^��"���|y��YX���h_���8�i��S�W����G1g�f­�u���V(������I���*�~�y|��BthW�ں��8�����������^8�mߋT�$ M� ��c���8��cQY�I֬��G<�D~a��6mނE�{� FjI~�!\[�Y�A��]p�9Ñ���_���q�p�'�ۦ�O��H]x�W`�x�DQڶ�}��b��L���4���w����9a����z�-��-EMC=f�{_�X��_}-L�|	j#��]i|��p�8�oOL�g
��ۅ�n�a���sν\:
fg!")��|��.0Y���8P�o�n��r���#�?_�X��?�M�~E���҈{�8pݍ�P\���*D�u��2�-u���w�ɰ�}���u(_߱������Xܐ�6�6��w�����|�����
�������N��8ƕ'���st@8��_[ ��!��웬�'N�2l��+�X,]sYnp�l]������C�}b�a�K`�����W������״����S����Z����Nrix��C?���뀬����V��\�[mb�}]��^K�a@�/�J{����FD':Ac���Hs���m�ۨ�{vV��r��zFi����=d� ����Jd��
�U��$�2�^$R�a���W��#����jz:����LК2�I���\�������q��dV��D���[�3������;T�x��]+:cԕ#���:W�?�Q$(�WM�h���|-�V<ܔh"�*��SO`�1iҽ�����h�t��a�:�o�Q�A�.|OF}����Q�#E�R N��D�p%��n5��y0[��X��ki����s�;O6j�R���N�S�����X��Z�w�?�������c�XBP�^���޽�a���h��F�N��M�g�}�9��� �ʺ��@C|Bs�=6|��a��V�`����3��nD�`­�`O])�]�62)�-Rݍ�<���jkpť�χ���1 ��	���`u��u#��H���h,	��@P
]&<���_�����a��m��L���c�Kb��W"�ǜ�s��v�a3�1���p�yg ���D�PT�:�Ǹ�����PԦ�t;B�$�v���1�EI��GQ��B2Ҍ�G]���o����5!�2"���$'��D�r7E���C$�����X&���[4��A,�����0�pY�%�ųO<�n�e;�:TW�B���Em�1��Q^yοd$�؎SF
4�	�1쌓��c����^h�!����1��Eϙ_ �1%}�&�~�^\v�y���0���y�F��w�t�b&N9��7��������оc7"IQ�c'�B�t�=9��Z\}ɥ�?�pI��j��𡠸��_�yo��O�,C�bE�~yy���hn�Gۢ|4��G��];wƴ��F��T������������f��'
8�@��B��ކ�7\��/;O=�*�uV,���)s%em��ܗ���1��Wѱ� ��t��HB�O��f$�#Q�Qs~S&L��qNi2�8���`*��N&��x�o�qL�i��(
KK`0Q�X�(�r����>eʔ�K�Z�8��BZ)k�AMU�hB�q8Z�ٹ!�k�¡�tm�ɟa��0��*;kf�W-����K��������<0@K+5뜦���n�[rn�-{=j�q)���QEn?�8trDQʗ��͙�0m8Ѕ=jT�n��pE�)�*��Th�Ŗc%�j���^�I{t�x�B+#@<��Rg�V*]���9#_BI&EK������F�N��h�"ټx�Ts�3�ev� �-]���>��M7��eN������(�"��QJ�۷��4�SEe'D"a�S@�2�G���͔R�"˩��D��*{�V�\!�[���EP�����}Ol�����$U���{edС}'A���ˮ��-/������ݤ�ŕ��&�C���9u��۾��v��8��c1�G��\p��~����ʫ��K@�͛v�e"�L߄h\6A�ـaCO��G�uW^�Q�_�����Y�e��5����)G��@T��&��]3�J
ݘ�`6�Y�=�U
���1�ХWo��p>��x+܄���/�qfN�SQ�y��G�V�!}���>X�W��@��!?;!"��#��,�(�)?ґ}8��S1���(.)Ͼ���X���%����TR�-�JY�	ģ��(+�QCŦ_��'��s�:]�k�,��DS$.(�$)�F��X��Z#��H��EA���;�ބK.<��(�y�͉oX�p(j�	�hqX��5erY��I�#b�OP2#6�-����A��ګ��&�V+�#2Tūه�<&�������@4����������q��G���ՋfH�fd�X�I4��Ǎ�]����7�$�ﮝ�EU�b��@^a)j�|0�]��gb�Q\�ˆT8�;Ǎ��qפ'��G*��s�6L�~/.1s�}�Y��AAI'A���fB汛i�õ���!ìGE�6m��1��/��c���QS�f�&x��D<�� 鳁�t*� ��a_�T�t_���+0��s���ݸt��o�	���0ռ0ZmHѥ�x�f �G�co�G�!c���c��[`Ϸ���#��ካ�E4aE8���^$���P���a7Y�=dp$����PpGB���Su�d]�Mf�Y6�I��P�����`�j��qG��[��ɓO_���'�Y����ټq��ik٘��
78��T@W�8=W��8�Ti��~` ��`��Js�OI����}K�j�m���s������N4���Sc
%h�zk����f����j�_gK�(���9�U�cң�R�ь��s"�UoUړ��`�V�l�f%:������b����Ɏ�:��LN'���+��j���sE\y�8�3��&��wu�8��I$�}(	7saP*�<�sV K�4ȯk��ʎ���r	X@�R�����`��Q3���j!��ILHӋ�x��:���KeA�=U�hRXP���j�5i2�;�a�}�7�Ā@'&�9�r���Vf��7�"	b+8չ�~ݨ1Ta��i\:�R��>=k&�+*�{�o8h�`<��su�u�����할a�m��&o�H;#��K/B�6�g�|��2^9�
���B���N<4�iX� 6����2��<BI���:��Z��k�c�t��|���8�,^�#RFŵ���0����!$C~�j��d3�-o�~�p��1���R���p1|��Ddg{2+lVdL��oB,P�S�93�N�o�7�����#e��K�8�묈ǸN-��f�?���pvs;7��QW���� .�~^�	g��"Ē��4�!��$ד�i,�C*@�.��$��۳S���}�RAڝ6�}���|�*���)�ij���U��Oh�"b�Y�d:)�x	蜹s�ZDD�밢��
�:�-FXG�>=еs9:wꀚ�쭮�7?�E�?�����6J��"�+��7��0I����̝jhw�k��.D~I;�b)��8Pk��o��$Z ��:i�7��j�
���W���}?�N46G��[���i����t�#�oD�ׅL<�����h��tb�[�~����cæ-X����/m�ÅXB��)�����D��F�H��{3�"��nS�ʃ�O�.l�&T���k�v��5#�����ڔ�ke45���`�Xp�S����e�/hW���8�Ne,�ǥܧ�9���ƢrV�E��+F��י�6$�p�ꑂ�rQ�քD2���,��ڛ����膻����˗>a�X�����F��g72Щ��Z�{�9g�v��.�K��tbN0ϭ�u�>�����L�t�������f=�W�����;.	F�y����:Ӓ��sxu��ߥ�pL �����V�Q*trGIw&��<t��AB��ơ�0����-�I��u(?��'i�Oə����T)e+#
�ĩB����r^���7���&4/����M���;HCZ���|Qg�v�	N+*��*���t��.	b�] �8�q$��ly��t�2)�1� x�x�	d˝�^i�Ǣt:�_I�x�d�#�׆��q���ә��.{�U�$�]	hL��N�=�z�g�.Q��H�$��RZ��x���JF���[�W�����za��	�C�������Cs (r�D���d5JBU��'Ԟ��������~M<�׭_/nm7�r+6���L�kA{��yHʘˤͨL�(υ!G�}�v�z�N���~�y쪩��YO#�����dϤ���o<Ԍh�	e�y���L��c    IDATsq±G�]��v����K��P� �2��!��f���jS�sfSƔ�M�3��0���3�lۉN]zc���d�wГ)bQ���$������N�о�7�0��߮�/�����m�DVT���p����@�ċ�eA�a��D2�g,��ON�v<�v<^`��g���_�S�Q�I��d	��#A�ԇ�=�ʹ�l�u�J!(%<C�3&���Lʜ]dR�۳^�Y����.�ٹ��}0y��s� \x�Ht���?������!1�e� ��aNb���()*�?�����]q���1�����*(���ן��T4(���}�еK��cH1�ѳW%Nv&��q6����f$ɘH ��D�ӊh�'X&z����׀��{�s� ��?�®�m4��
�N	�6���I��hTX���H'�ع�Wt����s/Fy�^x�9��L
(�H�}
|�h__�>�a >@��9�H�	�MK����>zᘓ��)���3/���KW����8�P��.�3L��H�7��(���%�I�ƽ����N�JG��Y�u�J��zs��ϼx�U�-}��ɧ-[��I	�Y*����G�+5�4���h>�2aQ��F��5^W��\�-���pps��������+c�tK]oº��g ���U�~jn���ǪZ�ɁBǧd��YVnW@���7_w+4E��l���v"%�쓳CtV�T�u��R�k�BU/������c�`E�>V�<fq�C��UҘB�!�Y���6'[��U�j�K��	�K�P���� 5��:� թ���*6���bTR�: �&���N0	��n5�LJ2"`(�X���� ��p���
TZ���ʙeRm�4�P	h�M4:��I��䢡�N$"�{m5���1�D�����Hk�F�5��;-��x\D`�T��e�'p��s����Orm]|t&�a�0Y�"�"����#CM�`.j[;,��(��17�l1(��TR*���:,]����[d�4g#Q0,5C��:7t�Q��j�kл�!8d��x������)�S8���<�T�R����d8�w�zu�҆lh��-�/B����"X,.�,9�P$%Q�~�x��h_�@*D�n��&����Ͼ»�~�ɉt��3��m*�0��F8P��Oęg���=~�-ek�Ÿ� �������0����7���g=������w�}�]�٥�=t�v+y���X���i���)�)�S4�%�F\M�����Q�bDqg)��
ɩ6y�k���4X[#�j�E��mP�q7��c��I����.�m�`�G_b�k`s���:�dEyV4V�D�_�<���WDg��2�� ����d�RQ
�GhB�Deej��"�\C:�!������p��A(�P�O9��9 ��i�xh&~۱U��R�C<i@��PFxT�k�ُt,�L2$상��^��I���Æ���b�������N��7�T�c��F�׉����5�ܽ��e�5�N�}�$3�I%��JIb��)(EJ� �H�HP����  ��N����$$�M��dz9���]�>�yy�>}�~�˹�\i3�<�y���{���Z����t�����~Ь�0;�X��w��3D2E�a��I�Ew�N+�C�H`t]5�^�Ǵ��o.G뤱H��x}�j<����3���_�ފ�0�m�z�n�������$�B������&5�t��TB@f?�c�9�C�GgzϤ	�n��m>�o	��W���G w�TY��xP5��+W��,�*tM����6��%�l�g~�*}�U����|�J����o���w��?��F��=��'��?��cp㿑?@���שs�
z׮��.����C���<t��JMw�g�(ĩ~:��ҘV��s�#�T��8X��$+�?K���U~��,���ZI�J�ܨɳ2iK�(���U'׮��0�e��@�Ñ�[��4�)T�8�W��/�9{�g�x&�2d�Ns]If�5n_S�*L&��>H���$2=R���UI
�9kN������F� �BMQ$;�]��lp|�b~#�[$�唒DC��[����tVX����X<��J9D$)����X�d	�z+>�h�5�R�ДD1�� )Ψ�K�D �ہ�|y),\���l��O>���&�̳���<���~���M�R*�4�GbhX��b1�ɓ�I�D��ν{q�)_�m������[���d���dqO{S#�H�BH��0*���G��k/�Q<̿u�w`wY�a��t���хڦ�h�iB:U@$���)��G>5������2|�+_�I'��3�~:�t��;�Î�	���h*�� g(����a+�l��S�ǘ�Q�����sσ�W�_=����C�ndrE�i8�!��,	!iº��]8������o��Mm�����-��D�QB��r�N%�sİD���tVI+3A����p��k���y��+�-'dܯ�C�ߋ=�#�c�\�/͝���M5�~��{��O~�T� �-�<,�a��AݘQ(d�H�1uR3�.>K��ÈD��x2���q�$TF�K��o�T���l�~'�:v�a fϘ�c�,�a��Q�vI,�|�x�OB(���5����q��k�F�T_��`/ʹf8��r�Ќ)��0���lܼY���1)�U��uP~���A*�������r�<b�<�*��}I\���k ���&�
�24�)��ؑ��pX�3��4�p̑q�_��������\�mh�D,]D����4tz�3(���
4MZ�����Gtey���D��Û��V!6V�L�uz&�T�,Ɂ��5ο��[���#����*!�i�`�����`V���<��6�:�)L;�D�}�s�����������[�]�s��W;�5�����a���=>Dj\I�Ld��'�����h?�,XUb�Ͱ�Uα/�r弐6H��*W����9�T W�g�W+񜦽#�#�E {>/�U�+3�
PX��^�����sJf���y���E$�=sIh��!4n��B�de����
W�j��s�A�t����j��8�<��\7*Q��HA�>mv�
��xyE���LzDCaa�
�J�Q;V��ږ�{À.���+0�Y�����V2�%�M� ��k��Z���F<E>�/7��V�TD,�Q�w�23}ϝ� F+�^�N`)���PB!�<�YAr����p�}?�eW\���}py�x�f�v�3��lu�d�H@�!&^��K�%�,Q�b.���<S*�d6��(��<"J�/�Fz>B24�c�t(.�`9n�����Ï�⍷��eW����n\��:�k`3z�Ζ����0�&�!�h�s���ގM��;��>�<�*Eb�Ҹ���P2Q�F�����i
��r����_s>~�q����{e��m� �{����`z��Č��G93�0�%ʼ�����Q��b�wo��6V�~[w�#W�!P;Ѭ�|	yέK(����`��uy�%�K+B,'S�8�t��p7�s0�
0��FC�����SE���'�>Z���#x��q��DQ�D�d����1Au� �Ӿ�+.9I8y���W��+V`��Kq�9�� ;?����2,xE��e ���q�q�_���̀�
�q�}r��8�"|��3�A�nt3ں����IS1q�T���/�ms��Nc������1y�}}A���G��OB}��`��#��#�*��B2S�{C/x�݀l,�K/��}�"�����[q��+p��0����ƅ�l�+P/Z \�D���Y�0��H�0������_ڀ�}�8�H}������Uu��NCgt!�WH�٨<'�KD�����@yYj�dGeDZ�i4�Ɔ����6�����.S�Y˟���N>���;�KC���n����O\�z�]&�i,q�(���*�de.���LqH/��LmJ`Z`�L�e�����wQd����ڭ�,`hU�����ӠR�=����g�y�*#=�P��r�@,$��r�9�}}ң��KK$���S���s��&{�pڶm;$�9\v�rY
���4�'���k�������C )�m6�9��YH�c6j���QeM�iW,܊�4KK�VTHryV7f�����&߫�T��5h>���&aUNF��D�3)	�r�bh���q��M���P�t���:Z��xjR���r�(�l%�d̚y�s%	���DM�h��T��C��(�!*_3������##���}�g�Wn����q�J:�jk��%׃�\�@ �hD���w��G��ꔖц@�Zm'�t
�}���F����`8,r|]s���B6#�B!���g��I�&໗}/��<>�������p�(�0iu O�jm�5abO?��i��}�B	;wlły���{����Mgq�7.@��D�ȑT5}�uJ�\"$d�sO;˾~*��=x�7�/_����q�M7c��Cq��.��k.��bF6[F*��^�ƂC�՗.ǲ3N�p/�?�x�ع����'~߾d�E3�e�5J��}��q�<����=����O��g�Ĺ�,�c�>����\�<����뫕�U�̙vj��a#�t2�Ä���{v��q�K/��g�(��ʫ�?��xM��X�E�UX�f����=+��>�׽bBK��*] w��Y���<�Dzp��G��ӿ*P�6H"z��y��Ko���oCu�XX�U���b���Ԅ��.8�:��/��Y�3s<3����8��Ð/�p���i,"ɬ$6:�Mf��!�mf$��5m"����8Ɗ��<��^Ay�gX��4DY譴P�J�~��_CwW�~�A�W���,Z�K/>�>`׎}��K�q��C���S�nBfct�t�N1������f,��0���3Z��g����	s�����]ӈH����É��4�N�sZ���Еqم�ā�'��څ?��&0��Q8���d��lHK'�*�jw+1+&Zn�Ĝ���4�P�0�N����m`Aebw]�I=�$ϸ"\.S٢�m�e���+V^�dv����_������2�\sͩ���6��6��J!q�����h�c��Ԕ�XQ��+YĬ���t%����HA�dv0�!&�*�S:RާR!i,tt+�xE^Rn���Xz�h���|�g���C���/Vz�T���Tմ��ܕ|����G-V�.'�Vտf���Q��h���摔9nV}:�]�N	<~�T�}��0���OL�Y��
k���l����l.�MX,�A�����NoHf2�n��n�x2�v�]z��s�E�|��y2�qM/�0Ǥ�(��-ωϡ2zC�Z���e��^��f�f�H�].�S���"6!FR�u`�O*k���;\K���z���E��,�f�.׎ֺђ0~��0��)��XK2H�B��1^���)Lt"JeC�Cz�W�<y4Iv>�$�"�"?�������`0 �IU�*���	T�5'��s��J��X��l<����6�l*�(�p�I_���g��ע ����J�)�	'�V�(�p�q�����{��3��6}�[n�!g�D{�H��rp:Ȍ����b���4w�u+v�ڋ��[����o��_��.\w�����W;Z���n�S���q�	,Yt8������MX|�A����7�r+F���Y�.��哱�tbCڷɨC)�@S���u6�]���xT	�pn��v��ۃ���]z�$;��QTᄂ���b�x?n��j����֛�ą!=w����;p罿�3/����F!:�\x9EVb�q.D}�~�3�O��֖1����={���P<�����=om�0�kj��s��̡��p��+h�*3%J�6m�D�p��g�2�]�&@#��F�3���O9M���z=�[߉�z;ww#��I��*o����PL��2
'�Z� �&6 ��Z�G�z:���.�%R���� ���gk>�|:�Cf���}Z���� h�w����W^E��&D�	a��N�����Ȟ�^�	��D�Y�,���Ɯ��A��}]�x�X�q��d�z�Syx�"�LK�Q�(�S���&�mF����I�-��',Ũ=���_>�k�ISǞ�P�C����p?xU>���J�F����#���O���5�䁧�&~����0N�W� L�Ϩp�=ʳ[�r�:*-K&^&lr���ؑ/s���EQ�3�R0���;��"�O�u�U�������]�uן��{��p8�x~Q����iU�H%S�D��DO��t��5"�?��@B���୑N� n`M�I�:�Y�
IaDI��ɬ&��,+8�a���~�r�wy�j�R���|@��\W2�
(BXQ
Ծ_EHȗ���+	K���6en s;T5�� ���9���vy2���^GP�Vҹ",V�Tw5�5�b!N�b]�rnocC�����Z5��5f2[�(����GW�@KoO��`4v��b��7�t�E�Q�l���<u�2V��R���̤��_W�?��o�3ᶴ� ���-Y�r����SI�(d���U�j��DJ����_�ؚ�]�9'jC:I�9�2C�_�����w���Ky&;L)T�Ng`��6��K2�-�fw�5g��M�a�Y�J��R!�L�_>rBoB�)ɸ�:���:��
����{�5O�|���L~r9���#��}��PV�V���}��t�K� %w�c��;���f�+/��X��!C��~4~|��X����~��iظ��q��F��><��эx�w������@JyJ��p�q���������_ށŭ$rE�?��]_�#�׍3�����f����z�a|�m{�!\��[E���e��-��2P������"X��`���RXLzt���칭ؾ3��n���<i��̂����j�j&�#�\6�E���K/B_w�'eSYv�\�l���W\��	���p(D���t&�T&�R9�C���o���v�܅��Z�5k��}��a�V�_7Z���RYR��J� Lw��y%�IKI�jG5 ͠��I0��Bp9�0�����cQXM:�U���G,�i˖�W�Ǿ�~p����Ƚ��A��|�.�m�W�Qp�a1�̳��ɧ-ī�w�WO=���~Ē���d0�i��E���0�4FI��w�at�/8��:
'�F2\��[�~�fx����8����z]b��۹�b�k1�Y8��`�Bx|:�]��=�z��bO�D��is"���Q�B��	.����'��䯝�i�C_��ʫ���B�B����f�d5#�L`��&��a��0e�,��وƁ�~p'�_�1��"W �J��ȴ�_�ʜ��c���էPY�$}��� Ǥ�.�j���4�J��/>�̕�:uQ����}��_�\.[����e|��F����~����|�Z���V�V��@��֣��NA2��բi�2������}�p2F��i=^~�
�*�r)u9V��rVllB�JӼ"ẟ����s-!�?�.p�WZF.���B�>��J�A�T5��r���kQ��8���̚W��~�T����vg%�Y��PP�ňh�a�8$ q<�n��S�do4:��#���g����C�3FE��}����^z������{;�3�m-:��OX��t��Yc�,I�RStEb��	�D��RA��e
��#�I��9���D���p!����Uz�����9��9�i��~�Y�;7g:#AZ�?V �
���~L�X�j3���������^-!m����w��.�B���>[
6��w�F�U�OB��Ȕ`�#}��e@�/��N���=t��d{�L�O����<^A�6��n�&R�����aDU�F*@����4�ע��KH�F�zt:�76�h�!�-���F�V�CCè���V&"z]	��^�3_��E���_�{���NI��~�A�ǅ�g�k�q��IF<�"儍e8�f�������F{k+�����V��_ׄtрp"��R�FA;hN��!I    IDAT�w��˟�̜�7���!�Y�6W �f%��X,��tz�I\slo�1c�D|��'ą&��Ilߺ���3��Q�2�7�� ��9�V�B=0�ʨ��������U����B�=�(��E��z���8ܞ
��S
qbo�-$���Ie��PF��H?�`	u�u|C)�I?��l�U�u�Ȩh��������x{���Άh2��"ς�:�̈́x�v�u�dM�"���ę�ᩪG�`�DF�ҩZN)��n�e5���t
��0�Nh�ζ��K8��q�9���s���?DM�(����P;�E�r���\*�xl����v�Y�=��gcL�x��7��m/��E��[�q��y�F�T�"D��C�߃R1�`p �B3��Á����5k1���dC%$�:�QͳJ[���yx�V�����gn�p �N�*#�m�;Ke�[����#����J�ɹY��y����{쪓4�3��B�o��e�9��i�=~�W>}�ѓz?�;*t��W�5k�]��xjņo���ĤWZ�����g�R�#cЊѣ�1{�!R��!U��T��Վ���W@��Q=�*=[9ԅy��LY*���>%�����oNX�֧�U����X��t�T��r$;�%��
��E�1
�(�X��5� �~~�T
O�
�� Ġ΀�jMcSכ�������צO6˼��P�Uu�&���B{F�nx��˗?y������&~����ڇ��'�n]��WO����zB��7����5��3�7��K�&���,l�y�A.�@kK�����ۃZBX&+�UU�N<V٪���#;*_[Da��.�ݼ��g"�!��B���ِ5�$����ϳf����l�t+�Ѩ0�m��w�Bȕ�(ȁ�J=�<��T��p�_7���b��V��>/z!N2Pp���H�{�"��?s��e�s�\�������%�I������M�uP[W-��E�?�ՂƆ��؛x%�9ᩮC*�V�&�f�_���6+RqX$ ���)�]�[�s���x��/��Չ4�B��T���A"��lF<8�t"�I�ƺ�G�2��j�Fww�#=�8�p��d�IȘy�.��CWH�a��D�<�/ 3�	����:|0�
����@�C �M ��TL"7ԏ���Gb�$�����W�Z_ӈx,#�k:I�v3��^�9�����H[.�M�x�O&Q�^���G5#�����ή\
�10R0�՚i�1��H`��s��X�ի�B9O�ܣ�sq|��8b�?���>P ([,`�������_�1�:ɶL�D�.4�\:*��et����^��6�KxuF������=�39���Y��P�"����ۆA��髐)�2eM�h�8��̠���dV83\'�U^� gb��s�Q�eODU�Ho��S%����dG&���8	e�<.d�?c��)��܋\&!�͵�MHJ�g��@��ˠ�Rix������E��Q�0u��.-�/J�R�-I�#����N��<�x�����_T
��[D�B�L�[(�R�a.�4�Ï��o�������3���-+V\s�����z�����B�yV�ɔ�wET��+�<�9SMX�PgT�n�8�p�s���HJzO�'�L���נL#!`�p%i���Û�r�R�n56'�����vԮ�N�s����fd^.jF�D�5G*��
<.$1USpD��+6�$0�S(�����Z�H���b�d���v����b��jv;�_ñ8��0q��Tg׾�ں��W����/?U��_�ׯ����G��λ7VW�Of��X
v�Ww�<05���V(�H��@�9�ED�Q�X��[�hp �Und�q4�nĔ&�F��\��T�L ���-�����X!4f�D8G���KA�T��=�A�δj�=yn6&���7ϓ{������
��hC��u�!�d˰9�x��a�����%X�q�/@}x�x��4�@yS�2�LJ�De�E"LE%�H"ݘcl�'�S��X���f@�"�j�����q˿�'�huإң�%�&�A�
Ya�S`g������ �N-����&J4_m�ˬz�C�r8]��:m�R���q���8b�i��Er��#bD��d���V����G4�	�\*	S�$�cޜ�2?�e?&�	x|na��uv�5���t��d���J�q�����_nZ�*ѣ������`ӎ=���-е��T&5r�s��5�!�	��P���}����E�.Z��a�����26��TI�Ľj�10؍I[Q[@���鴴Jx?�N�4K��;0��f��x� �Ib��RP1�uȊ��S�e�r!�$g�as�PW-�|�4�bp1�	���8Z��hQ!��`ң���|�D����{�f6TMm���^�C|�y�����kE����b`�>����Eo>�d��@r������j8��m�%Z��-�5�64"M M�^� K�w����@.��fFm�/	'Go��!<N=�ͩ��f:L��h��Lj�!!�\@SC-��a6�D`�������.������
1�1�-,
�D�`(�Em����D�t
�xR<�[Oge�8=>1��I^��s��D	W�}��]#���we;�㵌95/��`I_Ln�Z�O���+�>c�/�;��s�_��rپb�5�]��{^�����o��9���K�,V:�����r���Й,�X*�3l���﷙�:�H�#��D&«ڨ��dg�[�rO�ʃ��vɁ� C�E%��E�2�Sɘ��j�;�V,a�oR���E ������ő+%��*v飃$:�)mr-��F��$�/�C��8�f��h�`Ea���F�h\��~܄��H۾��xeR�.����-7]���f�?���yg����W���{���>�bvX���He��r��Z�+��#l�
ܮb|�L3gL��i��`֗�Xr��3{&vnێ�k֋�O<!�8~F>_�;�8�=����5$CX�F�	�hb8�o�Ǐ�@��1� ����F0$���p�Q�dC������0��y?i^{�ر�C�gI�9BxVA�(j��9��g���8Me<B��ʹF	�)��gOB{��j��!E775)��H����PM�@��P���Y9�g�݂o]x�}�u���_��0$���W]'���W}�Z��d�G�-����iSp����3�j;W�HX��φ	��O�s���>������l��%;�	���^�����nV2��H���z�2�]][���ނ~�(��#ba�p��F������p��1O���3(�3� ��J�����/�W����:1a���u������3�����Npe�?��Z*���1��wa���Mv^aQ`6�q��3q��G���B��?�/�{������a��N�����e,��a8.5��sCG~O&�&9_,V#��$�.'��1��NZ��g ���X˨�hjlFW{'|?�k�?8g���c�"��}_�nk���"��A�+��p�|�Ri��ݍٳg��$�Q��X�lٶ�]��Y�%$b�U0��%�����G,�"rw�M��L*���f�C��'W>��7nAss�\�~mUB�!�}.|�硐K������ol�/�rv���k��-�G��p��P���_>~)/Z�x���a��u�\Gc���j���݃'~�4zz{�HA�*��XPx�|�9pX��PDoo7�Z����?�/PC�u���)�{�E��e|(��Ũ�\5.&L�f��`�
�����!�A�VS9���m�l��w�s�7������n[�b��5k����xZ���]����"�0�B�P��t,[��r��+��V�!�?4�
�޺�B�lo(��e�?[̧�ϥ�2���� a5/��P��֚���3ǁ(�O!Vp���3-*f�n�:���������["K���ɨ��$V<x�CU�3*PAI�/���̝0:�چ�\�I�͈+�qq�m�������'��k����v�'�Rj�d2$���GKO<�ڕ�d�?̵�{��go���7K���]U[*E���L�RY�(��HW�+e,V�x�}	��NG$؋�-�8��y�:����@���N�
��.q��^�a6���vߴ�RI�B7D�I��Ҹ&��������>���$'*D�U��}�%x���a�M�:}�0l�^�!��<�")�m��3ټ�<+ҢNi�S�3�z�2mZ,I@c��B���~�Bg�NKN�g!Ȥ2�`���5+aa�d�bd��Xk+q���S��nWl�DB*/��f�������c�e�P�Ј��$A�7����Gֿ�풃���W^z	8`���1)5[��ޱI*?~v«o��!j���,������̯���OE>���n��P?��g��}'�aT�v����-܏��DP�$N���k0i|���)ek�䉁�6'�	U�,.?���J��+��,��<���&a�՗�\��5�|Q�.���d��\�Qq(�wlk���eW�6l���G?��s'�d-��B��C�fC$�DӘ&|����p��c�7�)
*A��T�3�fs!Oݑ�B"	�Rk!�bB�=_���@���<N� 7DL��a��8�nXMI����aX��V(I��Ő��}1��"U6�����hM�@�B!9GE��T�u���I$Q L^[%�D	ۇCC��IY��!��on�C��d*�X�g��b�"&�3";L(�&�0�9	¶�hAo�F��>��b����|^"�ׅD4��*?���0~L3�0Q�<��L�j��d�����S��� o�Z��`H�xT\ �y���s�D���[�ף��C�p�}�y��}]���'?E$�$��]�2�".��Lƻ�(tlu���T7�6=ؓ�Ll�ݐ����]���E����G@�]s͍S׭����=+�u�V��D�H'�|�����j-�r�r:�)����^�+����\.&�����7i��M�,=�kwO�k��Ϩ��惠8��3b�5�Cu�*��Y	���|wVA��e^a���k��1��y��s� ��_���Ӧ)"��yP�h<x��Y1P�nhxi��u:XE��$#Qu5U�������E�'D�̐�2	/�y!W�����WC�(�P�7o��L���Pv���;`��D���t�!�W���iӥ�y�}��M��ԍ�7�q��g�s���C�ۀΟ?�W,^�ẟD㙩����	���\i�T�T��|V�� �$"X��q�ڲ�#q������O6n��mm8��%X�v-v�ܩ�)�|%[���
��'̮�!0�&���#h�3�SQ(`�I�;Q�nB��Ν��0 Θ=U�u8�s�p��#�c�����-�tG;\�!91�s����H���2}�#a9���p��`�E'��u���P��i��l~�r�9?'?7L^/�]�_g"���%���J��sh�BQ�C�'M�5ŀ�ր/P-A��y���[���7Dʜh0��k�<n��	����.A�Xx�6�'���v`���x�ױz�:�\nD�1yVL�Hf�G�8p������h�+(z��u��h=
� ^|�%̗�J��`��H�c��+_9Z�i�G#���Ԋ6?���`��M�[O� VF
�#���,��K�����\�XB���&,�Q�ڻ��b2i����, ��/��N��w�~9r#�e�U�
_��)J�>��? �KBn0Y�]$��:�|^���=0)&�ˑG
BQ����M	am_�^�E�km6��-�H�k��`5ڑ����&��T�tFF.C�� �vD�qJ�:�	z�V�N&E\[|^l�����x%e�սـt2*/�d&}�|~DA��mj�G�Q�S�Y�D�D0a�ړ|V�Lt�mV�$D�D�@��(]�dg����3I�leJ"�#�Y�QF76�c�@�6[�_Ŀ�h��i�:�"0SWS��� 2�Ƶ4���D�--ryX�s-� )6�H
��u�D��;�w�s&"l��=>�b	$h�ku��4,��D���}2��������SM��s����:�������?�M�ӎt:M�gS�����NW*�J�r���j\�+���r�P,�r��J���������ydd�1���[o��{�y��v�h���{�g aϚ�֢�� �ROT��W��,��� :;���e�=w�����^��\F	<������+LHB�Rɹe3���72�බ��>���\�<_�׊'{\�;y �����V��aȃ��/�is���!F4Ö-[Ѿ�SfR��~�շж����_��008,	�1K�EsS�z�񛧟��6��U2���u�W/{���V�+�9_�Wޜp����h�?I�t��,�t^��I ��(�u�(ƹ�門��q��Xr�|t�ۅ���۶m��O7b�������S��Q�^��N&)�c8Mk'(��I�[�{�=4�7(豿_*�u	�3������,��������?����Hg�vWcTS��}��Hbw{����2�M���VW�I�t�^|8>��CDCCRmp�Nf�M�9��r�(���x��'���Z�8�n�������MǞ����ksܸq�����>���U0T��	���n6�d���}1I}D~x�L%��ۼ��:P2s�D<*�ntC#R����l����zԙ��F��� m$�m�ҩ���>�œ��F��'*^*�2��%9d�h�IXR1A78��q<N���& za1�bQ,V�in��9�ʽkl$���jՂ�`�wE�P�p@bY)�v�T��Y��`�������aU��tR�m=��x�E$��۫&8�"Z~�"z�;`��`�;��@���b����;(�ഛA{�d,(d�Mþ��dR���vz�UI˂�ހO�m.%���Ӈx����������2ii�����"!d��E��@�"�i0a�@Y�̝3��Wָ�2�
��5XWS�|� {I*j��:�	�]��I�TŖN�wV�L.��2!
����C�(��ҁ�~a"R�l�XP�E��,I'��.yn�p�M"����D'��1�����S.�[\UU &�J�9�J<�	�&"�� �����.	��)�K4j��vX��n�"C��.��H0��6'�=}�7�������<�K@���EY3EV��_l�w"Mo�l�������G��������yL��Q��)@W2I� ]�RN ��ٿF
�XE�/�KI?��E�cΌ�d!ǣ
����nf�ғ4(�vnr��za���4+g-����5�Ȍ��
�5׮���'��7�_r�g���r0k�=��:�a�^�Q'߷��S��_U+��=��r��Cq����c�������/�=�ӊB1�q��o�p�w����_��
��۽��=CñSBѴ�@kK�M�1�ѩ�R�R33�4�Y�W����,_v�=6�u�K.��?���WI���D:d�h���D:)����ISS���$���C�+����@'��C�)n>~��$�o��#�0����`�Øh��N���ø	S��Ï��;��	�Ӈ|��ꔋ�\��9�~�hP�G2Nw,2����xs��:�7t��T���B�ȝ�X���~��N�w~�#&9����ُ��ߠ�p����V<�٦"���$ٔ	cgO�T�����z"BAA �is��J���J�?_��=z^'�n"���F���Q��\&/�/��c�qȦSBc 䄄��V�V%1ϓ�F�6�y�ʊ�&OL�X)��F�K��ܫEa73����DQ�&Dr"�<�ʆ���YC�a�C�X�~x�tvt���V<*����_�݂�y�C�A�Ln���&��[OL��;;���. �A�S�n���(�I&_t�#�p¸f�m�[?b +[f�©1�e�&���B�5����Q���R��U6{�D,� 9�n�����0s`��Ą�������d&�$SQ0qb� ,4	�=��*?��D�iykC$�ӥރϗ��\th�$�z��9�@�@,��Z��,�`fT(�HC3Qͦ����A��    IDAT����t����0�MJ�ʜz��ߥMj��sV���3�7[0|��dF�-1N�8o������ry� W��N��s9��,M[v�IP��Â��&}X��&�.�������'-�G���_��¿�{�o����[��|�l�6�ql��\��9�$�e<E�aO[z���D��b��cF*�Ic�J H%�hooGpP�s��#@���E&=l��U�;����
��|kQfC����!��~� 8ߜ/�1<8�ݻ��G2u�cV,�YF&�Fw_�C�Q�ԮohB��]��s�#�E6_@8��7I�WE���O�a�y$����Oo8b���g��ϟu���z�ݏ��-�K:3L6�t!�A����$�pqs��Kp[͘6y"�0��U8����E"6�=����hƯ�kI�x�y�5X�2��;��mh((��I �ۤKW����tf�<��|1�R&���!�Ε��h�F똉2bt���W�s/������{�uW'l��mj�M� uj @翮v����`��q$�H3��J9OT�(,�8eؠ&�A���rQ���@(6D��\;��:�Ð=��F����+�^T?�ʛA9ǃK���Ȕbb�_���a�sz�1q֙��U�C�O���<Dy��g"�������J�љr6�C5�Oi#�r����c�#i��7�UFYa�v�^�d^5I�LT�kb�1
�)H2��KR]W+r��pD��!��'Jq��$�EZ�uau��Ei����K�ߛ��s�oA��U�D�Q%���)/�����/�*[�l�q�l��ۇh(����%��k�ط�
�u���p�qG��G2Bb�l<i%p����,F	\�!�5�m����D�H*�D>��� �+��X\M�����8a�ʐFd�iL��*�����Q��M�<U�L8���Urp��o�Z�m|Nrp���s��|�
\����۫T���W���j$
U������_��9�s{�]�{����\�=�s`��D3������`:��#�4�U�(lÿ3�Ϥ9m�{�v�"][wwbOG'F�k-茺Ho׺��F?|�i�߿��S���T@�/�7�����`�ق�J�O})��P��|*�r���2�Vts
�M�*�_�$E����B��C�d8~���V�i�)�n��l>��!��=�]�C����ϳ��ޓ�*����Cz�9̘9睷\z���y[���߈��aF��z�=���XLF�@�$�<��00�����F:����&'�	~Nf�0���Ȧc��:�+{�晓[�iv�%߽�~��K��m��d���U:'��Ƚ��O9��a��౛�����aޜ����+�Qd���jsү�f|�4< ����� є�P��(�QVRYU�X��pb ��U�FL&L�<Y�7�u�>��]#��!�*c<�Y��3�J0%r��a�S�-/��.��Ǎ�����T�z	��c��ͤ�K^�V��ט�D��`;E#�1)�:RbK�
�߅pI�d%!�:�=�8q��5*k�?�5F��0�ȟ	�/��c	��H��Ϯ���
J�����~���FY�m6��^S�� L�-��R�2PH�,�qU���ʔ���&q�P�~��2�T)���k�J��dR
{�M�g��ׂ����2�k:亰j�~Ir$�Ҝ՞�& ?�`��̨����4��2"٫�k���BZ,���w�����@J��$���2�c��$�y�3V�S��C�Ԍ���n5�b�fK�:'��+�|۷n��@�T���y���+�$���"�Q�HDa%>Z��$�i1F�b�gV�AM�p1��}$��э�n��Ѯ�_�,�`�g[�����C�26�{�����EÄ��-I��2�"�GEX�6�1����>�#�$K�����]�`�mۆu���as����y�u4�N!����$�U��r���HB��PK��}L@�Eā>�o�5.�d�F^5�=��j�y�vރ��[J���_q�+�-;9��U�Q}�\v~���oxo}ۥټ��k��0��	C��B�,���n'IBS�S7<�	*�����+��I �)59n2B,ɈP�6"4�Ϫ�j��׭�|i��)ՠ�P�S���ob5	���^z����uI�_`X�)Y�� !c~�ԩhhT��۷������u�ln 2W��cq��VKB%��<��H'#�����g����V���~�Q�Y��/�.��p"'�iT��1A���>�*��)/���7p�� Ǝk�E睃��=8���`t}֯�@���N_���/����c٠:=&M�$I,-���1P��0#7���[�sV���^�N`ynF
�L�2E6��v��$��uk�����/���2:��[3�!,J��*�M�lY���!XM����*�ʁOkS9 y��zU���I�]&�Z�a`�*t���Ow��GX�C�Ǐ���ە8��=��r_ Y�oM�����i[2��V�v֭��r�)����5hh	��!��x�%�m��=5�I	�yIP2i�Ak&�`l#��D▱\�>;�yV�21#{�^&y��3�*�bQ�ϦH_D�؆���c"M䆯!�1�g�Z�b�H<q��dE� �X���ƷJ�)�`��M�|^^OZ��d�'��0@y����0��/U<Q$޳�={%�;i
n�ѝ����ko���7�@�\�x��#b��s�ګ���c/B��r��"Q��K
�j8I��7ǌLyT��vw�b�2�"��F�2��eZ��M���98��G�	�������E��ȵ�XW/��*�Ӌ.�C׾n�-&�mA����z�޳���Ȃ:�D�d��X�)1��C=T$����ׯG}}�T�E�U*$@C��1K>S"{�+\S��A�~��(jA!Q|_������ƈy�
�R���q8|5��k��X��Hdo.�\y���{��sN�g�9�?*�r���gW|���{�����_��p_(�T��񩨈�ڶ	AF�6p<���*읓)s���+JlL ��/*q>@�sFUEt�b���@�.�_��
������Z`�d�r��MȦY]B�<��4Bg��)�j63���4f7_;���r�ò�x`39b����"�/$���憪�V�|⚙���
��[�Y��g^��l󎍦rR���:�z�]d�����#	E���^�b�f|�����|Д�8��Ӱy�&tt�,���o�����_�=Q�H���h�:ܼ���H8,=7?*L��>nXV�|}�;4�g�?�/�3g�LX�}��R���h3��<���ػo���.�!�hїP�w�m�c�����D����
�ʬF*^�	ټJ�����ƀ�)ש�F&{$�������L��d3u k�9�@Z���w�.U��bh#��x�Z�����7_�����J�{�S�L������a�k)�D"]��|	�H����H@)��u{��Ҋ�]{Dc��"�'�?�KQ�1-Q�c(�}$��,j�Uh=Z`Z^;��:EB�D�����d�$"'�+�qA����س�]֡�*A*C��L�1���z�[2��ѽ��&�e��=m2nF�k'�V�/(�b�D�6�pȣ���͜9S�I��!�U�"Q�)���{��)_�:b�4�tv���ϐ�Ʃ���N;�d6{^����DU�}_�-�!�������s�sOg���Z�?�{��y�{g�^���Ŋ��A�~�݂x"��qP�2�-��t�&�G$ƖcQ
s�/J9c�dДs�B�4�4T��(�J&欖��L¹_(H�qF�OXTѨF#`�߀����?��_YN-
ro�1"���Պ��V �^2k��OT�HT��9N�~r[�NX�Q��pO����#�GSS���zz��o@�z$��	������o�?���z{�l���.�h�r%�3��fNc��z�)%�0�U/Qg��M
Ŭ���*�����Ѡ���p��b]H��aW�i�*nn����j���ܭ�w$͐��*=MO^��*���{21Ȉc���yN�؄VT�T�PU�TA�BQA�Hf���V,II�c���5��JI�|��L���Y����?���N�?��fQ�����e��^{�k���F��՜Ε���M!�~�pB�t���x8��OR�-����]�hh �ݝ8��31al�}�]��yh�رo��\|-��^.7�6k� ΀� FaF����C� �/4n@<���G�)S���L?h� �ׯ�_^{U����⽏?Żk6�[�,�Z�.�C|�k��"��>@��(s�J4������$����*���;~��nk4�Dw6�"�3=��&	B���t	%��H�N��OF��z��\	bTt���E�]}��h!Z][#UNK�(|����X�$Ty��� "=�bN JB�R�� �Í�1�s�nA[4Q&&D�RIz=h����X�o��|>&���m�ā�̙,j��?����OZ`��0y=zv��-ϕ����3ߊ1�{-1��δB���'b��O�8�QP�m;Q_�(S-6�]>���� �M�$t�"��M��4\�ZgN?�>�.mx�����0��y��.>�����
�F5�B�x_=�d,8xV��)��%����5���|���jː�Ă��d^"��N0�ڽk�̡�,�/�:��gL����ɔ�C�k�a����J��u�R�^�t/Ͼh""�<�ĉ���t�>�o�**a'��'Q*�u�3Z�g�52�J��R[McZ����k�_@B�L��['����� R�J+�f;H��,j���_B����\;DFEӂ�Kճ��������9�:��8���vlڻ�u�l�gv���>�`���U�o-��w����[v����#4�f�}:�|2�b�$�(0RԄ�F�@[ܬj��?W�X6���h�-�y��Sd*>8�m�}f�d�vw���Jo^�|lj�Ue�)��r	N��ᐌ-q����u1��
�KQ`�U�$�)����z�|��!�%B�Zd���M&����B*,���5W_���\x�{����vk{�-����O��Zf4;�r%J�-g�ńb�T��I�q9�q�ҩHG.8�}9��`?�|,_~�f�L?p�~�-�z�mp9U���fe����ySf�Ա�x�$��Ơ�{�{M��k����O|�B��H�I�ј��~���ڽG� H�}�9l�k᭮��-m�tW�:V7��h�#�@S�.��;6���
� C31�J���0�#���JVX�oݺ3�ӊȦ�Z5�A�J�-�<!"G2
�Si��=J���s6�`��k)�7EZ��Hd�,�W]C��zy���i�'�lTΜ��A�WL�}h>^-1�L�Cр��V�ص[����$y�>Se�$}Q�Õ����k7�U��Fnd��AH����9j�T�T{�۔r]}���R<HtQ{S��7�wׂB0T��1��Qy��Tc���IV�u h�$����o5�Z�z=l���J��]2�B/��>Xmv�b0��������uk�e|�������x��٘;sV��I�k��[6�X���$I��qlMT;����L��r����TUKR�w�XMʉ�g'+��!	df+'7*J����H�����*@Ʉқ����bQ�f�<Hg8��%#���XPgem�w^/gƹ�8����?�>k��<�f�Y��I(嫵�N9���څ�7���f$���AN��FQ-�>g�~r��������V�S��&FLfd¦��v�ɤȇi�jݮx,-c�J"�y�6T5�!V�a(�7�y�}��~����?s�G����G�r��=÷E��z�����ۍr<�|,����@�Zn0ᾪ`^	,\�����Q�m���.�C�}:up
��d���>�J	T+s�v�J�+�x䆋3�*����-����y���l^�k���d�_���p������Qr���A�O��Q@.��I�����ݳ�Oz�?��ᚚ���Z��;�n���{��Ҽh"宮���40L�F�
<`X�����:	3�s������Ѓ�MEE�2I2w�l��1�~���ካ���գ����А��0�H.�y��)b�~�tB����#���	�'�|��|�;�?>^y�/�ܷO�ٻ�m�Ã�q��W����a����&F�*:̀�iF�ω�}U�2L% 3��ȼ8�D*.	����9:�k㡰w�n��Y�k�&�}�������a��!���D}m��X�{}%xc4
tMȞV��b�4O	S�Jdy�~�mWA���dO&����1��v=�edU��\M�಻1TP?ר:J�G�R�v&f�kj;D����ʤ������s>�{�3D�\�_V�'	NU�����$Ol�+�1�d2�V@em�^��%��!����9nذa�w��aEG�[y~i	��3�`�)o^k94cƠm���H;��p(C���	-���9�l���n&L~��8�83�bwI��JD�8�^aB�$Pc���{.������Ͻ����ĶͩdEG�P­T����2ɉ��!C2�d[�m?~��}�k��0�����*�Y_�q��W�\���ٵk�$�\C|_&�D/�٭ֆ��E��B/���g�p�B�5_�j���؎#׉���������+m�������t���95���k�9J���}tm�CCr��c�Jlp`��������>�k�஫��{{Əm���>����uj�����O>������5����QC�m(���Dhؠ��Q9H /�fX0�
�[��t�@a�z�d���Z �Ե1 �.{�2�Q6(�!Q�Rc8|'pS��zbe����Sa'��i�b���T�c�Rz*A�뒔�ɘr����;+T~]���y�
�R�z�gIe2J!�-կ^��s~��SO��O���c���u��ҫ�oA�25�/���EXB0:�hWI���*y!!Q���X( 90��g���E8D��,��,�(��b�AD(^}��Rq�K�,�,���n6�.R��+s�<��H��A4��"5��D�[�|�	�c����;�`ˮ꾯3���ƞ'�$$u7 `cىQ"%"�r���+!�q%�*���/���*�b�P��Se;W�8�&!FBb���jz��ݯ_���霳������I�R�I�Z������g�����ks{[�:h�Ko~A��?��G�����"0�I������$o������W�_�XxI]�9����t�z��t��|̢J[��?ܶh��z��2 /�k��+��ҟ���îr	(�d��r�`�f��v\�H��1����?�r��$.��q3>?�=.����O*
F���Յ�֒'�9�}(Tm��X{O�	��B~�����|"iP�]�Q8�-�J��j���ڀ�,Wã�2&2�Vib�Dt��X�'c��yx����q��X�o$W#A�����=��������%{�P� �c�����TP�G8���(�R��[r��1-�D���C2m+�G�q��%M#F��u�(/�W�pn%sY����r�`���1���liMy0�|�g���v�M^~�E��׾�ϓV�ȅy�cu�:k�y�+鳞��TM*T�\Tq1�u�l��Z�#�J�a.Œ�x�q�F��>4%U�ZE�3�6J�d��h�������b�8q��_x�[�!o~��Qk���&���}��K�N�:��}�G�����g���a!~����;��ۏ�_���e�8��}S�ܸ|A*�ӯmJ�A'R���K��S͟3��)��AI7ˌ��y!���@����NJ$b9�Z;o�ڐ�S�jd�	k�%���X�L��Pm�g1Ă��A��@���
"���d���jwv7Ny$U�S7a��5)��I�B����:s���������3g��҉8�~瓟�����|cy������g��v����:�Z��)NT"���{�Lh]���y���/�ßW-�M4�[��Mu�    IDATvSS�tB��|�y��~Rst�����bZe�C��(�q��l놔*$��H}�܆Zˉ�����X`��V��h��ܜ,�=,��܃���%��HJ�.N
�!�T�/LI'sr�[ߔ)J�#�����mR�4q�J@+ZS���yC�� Z���N�ǲ6�\zjjZ�UBdޒÇȵ/Iڱj��sB�E&���������k���Ո�1�,�HB�vX��75�5�����J�Օ�K׭:!0�q�����U��*=��j 3�8V88�K����l��q���`̹��(?n��a^[��8�xgLh����q ��bo���7�"���Z��ZǱ:�p-�Fb�Ơ��o�A��b�o�wS�����m��p�-{�{ޖ���ʕ"aKj��	
v*�o���\W��!M��a�������`�ێ�g��pj�H@�g�o< 33�*q��щ��:tô�$����Cmøbй����H����v�5漵�@ I���?��`nG�4n���v_K�ol��S��q$8w�9𔧭�S�=�N�8���]ɞ8��?�����<q+)�k�O�������y���������~��O]��7s
��v#7_�(����[}iJ�5{���P2ͩa̭m'��5�,�䴕�NS�i3����j(�j��I�d"s�a�Cv��PV@�!�WE��q)�kн��8W��9���b�9�!�2�s�*���|S��
K�!�B�R!!P5d4q��&7�����������{�{���N�?z��#������o>y�ݾ��ms�l9~Jn��k�fH�u4B�Wy���:N?�H���-�6���w�;����3]��3=c
U�� �7ƌ�����C,�l����q����
�0
��a�o&�bDD Kj��>Q���|��e�#H��ˈ��o�r�༴�Z�h[^���̷��j:��PIR�^�]�]���L�{D�/\y޴ǛZ|Mι��`D!8G�]#��H�9��@����4�!#�����{����
p�x#�|�Iٟj���5"5U=�j�'q��<m(��cnl�\�+�W�VEG�A�!a.������8��$X� ���R���"S&q��}���	��vD�DpZ�Lx���~i�=���l@zi��H3�-��qb*g�o�kfЍ�����s}lt��C_Q��QW�h-�!Iё��*:���U��9�J���$�X��r���i�rcI;�!�j�,�#�J��N�	d��tj��R:�JE[B-�J�����^�#��ǵ��08[8L\c�1��t&�;�x��K:�ٿ��d���ҧqAO@U0��<�r^Αc�s�_�롁���Yo����W�ȝἹ���i6��A�]�{�ʱ�(����&��k]��ޣ'��篽����/>z��s?X��5�{���/���=��6d�v����CY������T��4�!��L��Z_��dRQ�F�k��8m�����E�}ǋ�,xxf�Ԭc�a��hEtZl����U� ��+�*��U�<�-�`��	�'2��-�����;=%3�=��1��D��ڶRw�e�t�W{֚{A���Te��������ݻ��_�s�V'������?���?��/��Ǟ|ߨ*ι�3;.Y�wP^���+�Л��^�%���AG-�U��2�ZY���)Y_� �7�ц�3uX��5�0u7�Z��Ʊ��O��?FOJ��%.Rq�|'��&6����5�Ĝ�۽�:��䯛J�gZ�C���_囏<$S��D�a�i�kr9�ߣ������O�S�g9���p�� ���d,m<����r��yE"(���bd�s� ��ݢ����B;ۛѼ�����Ҡ��-�[�q\#L��8h �����S]j�ᓰ���Vu���.t=�ֶb�c!�)c��Q���t��P�B�eF#t撊x|�A�AtG^w�u��0F�FN�{�udC>�}!`�/�p1z8�Q������eeuS��6��wў���� �e<Eh4�P�X�\dm冼��U��'����+Խ���,lRs
��#>?�!��]����F����A�H�~��ʞ����B�c^�}`|xdƃ��O����~s�M�q��!�w�<~6Q/F��ii�E�	u�#D���X8����sC�������7�?��\�n�U=1�ёP$-�Z4N��<!g�8'�]��O9�)$��Z��1���o;}������}�}A��������7^�ট{c��E���/]�RS��2�'� �T����jCrS��&����6&q�MәZZ�ߦBe�{P��o� ��
���54�Ù���17�́�<�##s�s�J1��X�x�x��D����נ�
JH��L[U}zA{iʫs�O�v�ؗ��_��O��������������~���3O<~�3�ş�p��{��祥bnT�2��#����-�	�aI 5�a��b4N�h� �y�y7C6�[Z�Ң����5Gh%��"�
�I�J�
U�
��)H�Vk��ۜ����}����Y����Y(p�ZI�9`rՊ
�G�ޞ����E�	q�q��l�-��ɱ���������\��٬{���SX�5�%l�ݹ�D
,���\���9%��1��M���4��6Y`B�3�j�7�t�X��LS����l�u�`�Y\�ƕlJ��nKn�J��Y�̌�h� ܍���;��w~>x���d\�CF73��pR$#��h}�ؼ'-V�Pߧ��/_�h�1D�T�d��Y\�wG���/M�h����~V�;�@���`i2�g�{������W�x������p�F�	��!����>}Z��gΟ�Z���EY�ؔ��uI2�x%�1D�j�U
���f����q_���7��W���Xo{˛Tǜ��v���{��x�HU"8I4��Y�3V�����cc�wR1��Y�.?�\VJ@��}Y�~U�x盵�� �u�T&�M�J��΋fB8�
m�T��VW,*�	��lij�
�-��81��Y��_�M���}��E�ν�"qN`�!�F�="Tс�fL�6eX�EV�s�H4�㷟���_y�֓�~���կ��ɓ'���_���Q����O<�+�r����aS��G��|]
���4d!�BN�z��4cC���L��_�TV��%n��'��5ȩ��$t	��ӼKc������6�l�K�ǈ�V�Id��u�2��Pe�c�ŉȟ�&1���-�:Rl��޻g�+"=~#{d8ڒ�M�DѳW��S�'�������Աc��zݑk�����YVu[�t{�.�G[S矹x��Ͻ�ŗ_���͵;GUs�5yw\g�H[ȟ_[&%�t\]lՈ@�Ay��0Bd�a�+8RKo����LO�#%x����V��W��U�F��֦D��e����C�W���') �7�~8g����
��Em��f2��䝮��*r/�n.����\O����r�W���^�v�����w향
qsr�_��7dvq�6�Q�ܨ��?��E�981�!�e~����ϢC$�"�C�a����4,�Dd�]K�.]�sCKcuˑ[�����v�puhX���^	���$��q#b��q;o�P9�����yH�J�c��D�]�Z_��A�����]�v�Z~U(������lZ�L�f�"'��ͩ�u�%P~ī� 8�8�1O��	5zx��1��C9h6b�<�|�̙3:�WVV5Oޚ���`(+��K����?7muC�h|� V�8eο�Mwʳ�|K{ҟ{�����mhy�pZp��/�z���" �t k��lm3XY���̫9\�}�gN^3\�L�q腁\����t;S2.q̌/D���ı�ED����Ր2������O��Vy�f8:�9�cͼ���w-;F�f�^�v�����t������·<+8r�S��8�w�c��p���I ���)�Y�i�ӷb�/�>q�?�_?�{t}������3��Ǐ�y��?p}��ە����g�Ѐ�$b557���x:�y�9=�Ǻ�J`���Zc)���Z(*�H��+#g]���A<"."ܘ�-F�nQ�=0q��4Kn�]����1Ѣ�l��t�S�<b<cE�#�x���М�'�ۓ�ׯʩ[O����RSӚ��e�✌˾L����n���t�ҁ��K�3S/�I1ʓ,����������������pt����d8b�r�L��bt}M��E��15��+�h�Z|Q�HΘ �gI�S��V�2�^/cA���9��E4 h{�^9�>�h�݋}�W���2ob�X��ތ��էip筶��  ��#u��A 7&��0++7�Mw�^^�V����D�իҌ��ӏ9T�?����M����k<tp��1d
7�4�(d}sKk�EאO�Q¦��d@.螶t�@����c9v���/���������]!LD��������U�u{*��):��$Pm4S+�O�(�Ű���fR{'��J{�#7��uʓSe�kYT]��܂�o�����A���m���S��-�����?��)�jP�Pm��i��#t�C�5�c�Ղ厨���Pr^p�L[���ǈ1g8�hh��m|�h�y� �8���C�-�r*��r��9Y]_���%*]#[��P�A��9�L��gv�'뫫Z�wa^���7K5�#?$���A[��@��g�s@U ]� 5�V9丙��aߓ� i��&F���4b��2�14��5���y��m'����3*���G����gypK�X�����@�����9{V���+Wԑa��<�S���Yu&�����WQ�L�sjN�eRK�C�q��)��5I�M�׀�8Qt�Keq/�]jS!I8<(x���ZՓ7�	��MZ7�~��4:t��H��:yJ����S��8�K���'��{1���9���K�>�{����~�箯�Ni�]��Q��y���f)�N��,<�6�� R�L/ݑ��C?d�{��[��n��,B�@��Qݍ�ߣ1��N� �G����&Qy��q_J�����p�BnPv4d�����,jTy�5�HBA]s?U={��v+���y:L|3N���gE��v�\�9���ȶVp
@H9<���h�E�ݜ�R=P�A�'���8�-i�ɡ#��mߍ�k� CX�C�����a�zB�yƔ�ޫWu�����#̆8dj��Ñ��-��^SJ�M?����R��d喌�7U��H$��a ������4}��Ȱb�P�A�bd�ʔ/-Ggs�Q#!j�>��7dn��v�Z��T�.��(�%�@6�����G�Р���K/i�!�����H�muZJ��e�VJmR�`���k��Y��G�H�����LJ�D�qO�L#{_�4���F#f�NPQ�{*u�M��EL=����PYNW���JP0/�s!���"7�w�
�>�B c#�̙۵�'��} ����p�'@N�*K͡S5�D*�� ���R���w˗���,�\I�-�䶭���g����>�����V;�u��w����ȍ׵��MK9:��ˋ/�9`s�r��,�q����J�UP&
"D��<�on���ix�w�"@�Ք�u�����f[[���0?���u>�����8��C1��g]�HB�)gG
GG�{%\f���&W��,y��@�66� �
Ņ�=�N_�7��z9���\y�\x����ط�O��n�o��c�e��ե�� 1�*[��P-I�֊���b��W<��^\P5�Ǿ��v�\�̵,eρҙ��Wo\�����K��������F �����Ͼ�O|��=z�'WV����nM�y�/���V���Rٿ�^��+����j5�(�9�љ�,���z�H���K����ݧ�s>,:��¯n�kT!���D�]������@�A$!D�!���b��<%�P.ԩ�\���Y����[�(G%h-7O�"0�m>�H�O��Z�-��&+,�Gei[����;�~5���8~*�����Ϯ���Q���,�Ǔ���a�
F�y�r�1����Ӆ�2�MP����x\��^V��<Ӻ�.m_�Z�ҥaQ_�E��!��a�a�2r֌9b����l)�A4o�IM[��	����aX�9��7t!5�j�Ɔ���!'[S1@
 �8����� y�L����E��֛c+	eQMr�nA��E��������o !O�� �07�7D8~�f��'b�w޹^���ɱ��lD��A��d�e��lmm���!A!.�8v$�ahL�]k�+��8T�_��Ź��'�����p�i��S��޽�o����VǍ��}O�v)ּ��G��O?#�}m�A��]���!�2�88������u���Tjǭzƞ�L��&U n���F�[�~4U1��	�RU�Sj�Ky8F�D��;���;N����k�^`���<�~�y��P����I���cj��2���l�=ƙ���
�L�d$�s���y�<��y�"��Z�������7�e}uM�ǅ=��1Ϛ�ĀO���1P�c}[�\���E����f�����S��������b��"t���^���������ñ����{��!d�F8�°ӳB�݌4�Es"t^�8��>�AW�&.�U�o� ��x{b4&���\��پS��@5V>F�& �
88@:j�5��]_1����9�������}%��<��6N��\�u,�w��̐�CX�	kV� ��C"�^�ߊ�݉���e�܂��D�":&��Q'*8P�	c�� ;HF��8�vo�} �=d�R��P㬍{����p�L�pvn^�_x��bX����V�xԮ��S9s��@�~�x����W��|�k!����K2.%W�A=�@�qW9�$��1�X�5�l[���Ѥ$���߉�qF0�8�@��J#;��aZIB,���VU䆸�/��p�:yײ�<�ń�(�g!����"��,nSĐG(CN
�k�`�XD�P" ���g����n�����̧4��}$B�`���Zk�1����8���c�8ƾp�X�c.�����Q��A:Z�bԩ���t�.(�Q��3Cꆹ637��2ה�Hn�1��AS��ć�kG�Q!���ط2m8Ų���>��������j4��Hk1��8M�qC9mtfb�@ ������4Vb(�mՑ�<@�z��<�H������d����Ls�+��ǌ�Ӏ��~_� �G�; �����*"Q�Km܃��⾽2?3��}�t�,d~Ϣ:|8�ڄg0P����0�A�pPT\h<VGzϾE���< O���a�������?m�?��5i��/�������>��3?5�߰��1?�;UY���τ*K�}Q�7>q�rM=v��W�M�F)B-J�rU�(+�7��Υ��I��l�^�N=� ��J�Y��׮����4��4>�)��L��z��#>�AvE%R�������ȥeH2��G.=��o�?4�a!TE1�m�T�V}����U���f^kÓ�����vg'�S�_���$MӤ��P,cW�G�����x���H���;4��!�$�f��S���t�,Ip���v��4�b���o�������{����
r�E�јO��px�Ɛyf��6�Bf�d��`&��$M}���O��g~a��СC�[O>����}R�Y��[�G��u
�:I�������sϥ���4M�fYA*�W�l�)i��-aH�����I曄�����1�3i�i�]4���窦�k��n��L���d��d�c�X5�:Emhĝ��<��|�S$�JX罷�u��z=_�u�el��`���P�����	��=_���s~�]T ��Ѷ��3���X��de�Q�	�z]#�q\��={u?׮]k<�R�G]{���m]1D�p0ޱ[�����;F��+B��'��r�7&o:�V�ҥ�|(S%B�M[R"s��Q�&��ߡ-^w r|��A�4Kڨ�L+���s$}Zl�bwׅ�q����xu�]�u����US��S�  EIDAT��B��$U� ��i��(��9��x��!�j���Xؼ�	jX�&$V��t&��
ٞ��iz�8��0D-�H�%H��T�2pb5�*�@���e1��c��q*"jg0����{fN�ܤQ5�\��O��=�?|�C����ɦ�Y�����/?��oXn�����x�qU���%�ڒ�N�n���,Eu�ŕ��U;W�q����h��q,X̰J��Jj1��4.)��.ɜ��kI��L�&M \�Z�����w94�&�iU��NKH�D�t��ƻL-�-&޻$�I�z�1�b��5�`�\�ڎ��RI�
�5M�j�z��4�i��M��yZՍG]��F��Ƨ]�M+I��V�iS��I�4��`I�|դ���?�7�2�����rh���3n\A�&M�����.%�d� b򤌊���>�����0�D1_5M��#p]���[�s��C²��!��9�{������,���-pS=��o��x:6,K��4���I��]����]L�z����a�q6�
sG�4IH�����+�aѝ����y�����v�ݝ��<��p;/ZN��G����\�""�p�����)ǰb<FWeE���ոl
d=\�ҷ�|���z�W����&N���%k�p��$m�W����+����[U�j��I�gI�����ey^�-�� &veV�.�&�\�a��I���#�!��7z�Z��s-�t6˕;�a�S\�Oo�C�vU�j�Y�U�I��S��o�VZy��,m6��y*f}�E�m�*��|��o%Yޞ��Y!o;��h4?7;�R�UQU��j��ʧY��*�R�G^�-�\ݤiμM�<V��zM[ĒN���I�4�o�̆��'i���֨v>'�H�2�{�%�{xEZ���s&^^�ֆ�%����A��.���G��ZC���?gY���Q��CXWUYM�˝K���Q�"`��3"��)���6�c��
U�#o��	r|�Coz �EҊ|�4��׆F���L���岹�"R�t�:t��b�)%RK������s!�j#!�HHS@�D����@i��Z���)prBZG���ZD�O��,͟.Zş������{�?y��Ø�����������e~�����X����!������R�FҼ�V)e�>�/"�/H�����Rמ���J���2=v2��O���P�o�F�����"�oK~s��w�֜��oԼ���ܶ��h�����lldk+�daO9���Z��s���R>,���a�yʉ��z�瓥n790<ꗺ/Mփá��r{&�$��tZl��jn���әi����ܻ��n���i�}������qϾ�}i����h����B�k���W�>�X��"���7(��+��ߛ�H�J�w �Y�ߑ��d,2ri��I�hCu>rn�sߤ�V��n�ʠ;���lQ�V��ޥ���4񭼓du2�6���|c�5��;D��|��"O�$kr_ʨ�����e�W�ϋV!-I��p�$I��y6�&f�N�N�~E8\�%i�\�e�uP�-4j��Ns���d]d��M�J�,\���@ yu�,�u��aʽ�2��ʖ4�*]�v5����>˲�j�y]�m5�i�nH���HӜ�:�*��"��wS�&��,K����>:HJ���4�Uy��U�)��$^��EC�h�&I��ܦ��wV7�;�zy�Ӭ��zB�N���K��7��8	Q��s8n��d0� ��Ay�x���L��:��wp8��omod�N�y�`��w�s.�m%��v�$�CP��!}�4M㊢(�v[[[I����4�z��<oF��{�]^pپ"X��Q�^2�ۛ��6b{د�{�O�����o�q�/>�����՝�����G����\    IEND�B`�PK   Ŧ�XF|�X� �� /   images/608cf678-e816-4d17-98ae-736018483bd2.pngL{eT�����5�B�n�]�[ ��[��Cp���;�;�3�]������j��^���>]u��{WuG���b���  ,y�O  ��ߞ����b�v�����,�� `���å0c� ���$�����j�t<=�'`�k�A����tY���%JS��u3C�J;�ܠ�csL{!\��Z"��a��p�Mp/����6�%�زqyU�6�]���m��ש�;������R2�K���WB���	?k����o��_G�(+��� ����_�5R>�4�����:�1k��������9�X��e� t��,L/��tl%f�_s�E0�������gǜ=/X5�F%��Q�1ٺ�5h1h�^.��H�e�O��/h0�����=�\�M:_��jl���7Cj��|�����W|�@���f���{�ʑ�`�ROί��*Jcc�*�K�����!̯�k'����@,�%�kJ��P����Hbo2�2^�J�3iT8��ⵗ�]=Ay���<R�\��-�#��>c���J�e`�����YY^TMS&�kԁ�/��y��'R�.�.��`�8�55&�WKO��r�;?I�����d�2��eZj�|�7�o�ʥ�<���@��5m�x*�����j�C�2A1rm��u��L����fXc���zÎﯼ�"�e���Թza�Pű1�E� ��/e�0A�?4 �^l�5�Ԏ�����*�s��go�2�Fw� ȉ�GpٿA����K�-��i����E@��}���m�u��μx�֠�F;��w�{�}A�A��%S�嚥�P���fٖf޼�9��;���S�U5����Bj	߆�2�6���8�v���h[��@Sł1�
�`|��,+��C��v��H��q/�߬����	�����W~�����y}>�皊���_���<�_1C/�~��܄����_���۷�,��dp�F�d~���3ʹɛ��ey%8��S����SUGdD���,�Kbb:_M٭��<O�Ϧ/����	��@-�F��mm"QAJ��cLO��XU���f���ʡY�2�Dņ&6\;��7�BM����g��oNߊǂ57Ý�tQ�Шf�����c�f<�M�S�H55Pv�NL��v�.��n�m���fي�#F���~�"h��r��up;�)�s+�����S�$�KQ�p�h�QN1���Ǵ�y=룘�^X�]?8���:��	�����QTL4����@�K��p�3��Z�FQ*@�D�=|�����蹡���o�����ێy�����n��eIe�H�	���2�7�N�y�9ٳh��Bg��j�!z(�L����YYYg\�\����hp�c�r���H�N�qR�.��T��w�,�I��l�����ZV,䖅���	�[rę�_]=T��( g�s�a�����[,M��14��^�8!�[Ό޳8-�7i!˹�W��>kn�o������h"��h�q���^Tc���������SQ�w�8rv�9�=�+;`��O7��>���k�6A#�iW��r�c��yHU��;rѕ>����9��Y�5�X�4��&:vG`�b�F��?O��Fs��! �oR+�dKp��8�Ek���U���^o�Y��-��mӏg=&�w�x��n_�l}Xؙ�	��f�m��y�����߄ܮy��"3��<¢8�e'�8�Җ��E�y����M#��!��4)Eb���r����`���֤18�eV}�E(��5�R ��>���E����I�d҆�\\Q���m����s�@Q2��Z������;H@Ղ����z �lr�r�[�3�����������}�_M��NM��	����C���0��+�ш����ҵ�o����d�2姩M����#pm�!Q鿉�0�Q�^�s	a��wp��G��w�Q��XsgM�»vᕳJ8�o�C���ڢ[�y�����:�F�#s�ĵw�:����ږ���#�a=�>3�$�N�b6��bFY��p)�q��A4Fe���������{����j:�2�nkj��J�c��v� �RJ������?o��ŕ�NҢ�}G���D\Gu�tPv��/��y,0*��B�(��C&��:��t ����|"l�ap��{�w;	%�Q�V�S�|�~�:��������j���;���8Qm�'���<\1	�B��	6��T��b~+�a��f=A�É=?U]��x{)m����dq����zv@�>A�q%����"L�fY��F�"����h7���q�S�Y�|���*�T�����asή��Y	r����}~j �ӂzZ>��-�}+aI����ւ�3ν{e|�U�R�'8~�8bZi5�ԝ�oQ���qL'.�Q2b.�d�$��x!UQ����p.U��\5�>�s�2��E&�5*�ь:*v�[����S9B^aMssG9ղ��FZ���5pl�2�v����(pr��������J�5q�(���.Z6=�:՗�h��K n@W/��2�%j�]�������,ȸ������')��V[�q؄��z����^)@^X(�X��4�.�L�r@�!^��a߁>'�!,"55M�Y	[$��$�,��g׎X��!��^P6��z��Q����<q���L @�fI��[R��S���޽�w$���B�,��P �y�J�!tA��:�͙+�怎�$�&�ιwc��őcl��	���	{��S�z�#���A����3���^�h�~�nԫ��KW���������,<<>����X��x, |L(�Ʈ���sܦ�L�ߵ���{VM�d��t�oZTk`����c�7�)I�E��VF����;��������5z���9m���ܹ�9�x�횁����͑��?��,�ӸH�&����-�_y�c��b/�*��Ɋ�`����pQ���]��ş	R���dȐ�W�M�׎!�Iƹ>�$~L(D�=�~4���ѯ�W՞7��k������
�i�>�B��u���M������)������i�x�%~�FI��hE�E �:X�9Ͱ2�-5ei)����Wȳ��ab��vI���-�4�����J�����A�ڍ�4���>��Ԛ~�h^	��	�/���nޕgkS�ɼ�{��}a�z�~$#s4�<�3!�D&_�������_���t#~�x���	��쾤"O&V^���R3n�A����1������R���͎�Vu5��R�������XZ�ʩ9�R�R&v�*E����dId 6T})�(D�b�5���<5���&�7���PKØ���%��9������H�^�_'�x+�"ݕ��#�p(p�$�}5�y(1�G��qo�:Sl�|��3V��o��p�4C�p$�%��-�r�pȺ�L,�Ľ�[���������}a�:���g��̢dʺ�O?���4��}Y�3���M�W]@7LI��r��b�N)��F�D�ș*��y�n���Y�O�ؓ���{.��F׷a_3��u������2�n v-��[��k�\ֆma��#���3e�{ײB��,V�Xqσ��S)B�S��	���ҁ_�����m�G��*<��~	�V��	K?@5���e��� ޱv�1��n0/�ס����R�5�J�u����ְ2mu�
�Iq�����������u�	�w/ǋH���w'E�
�+;B�qR�w�\Xv�1���pI�4���IG#��^��R�t�r7������W�)�E�RB�ˍY�(��7�#,O]2t�"D�4�'R�F�M��g��6�ƯDUJ�n)ۊq���Za�4k�9����Ņ�dj�oc���������+\�_���x��P
���B���anJ
D!t��5���9N��Du�1��XT��ז�L��e{��rg�*��69���?�qS�Vq�<���}KCkQ&���󮡳,���LSȝ{"{o��A�R%$߉���Z�f;�����QH��� �=�#|DA6���|�
h%�*�>��1���j J���:<W���7)�9U/�!9�<�Ǻ$G�6y;q�=X<H�����W����+�)���E\��ʌ�/���bI���Q�܆} �ᏺm4vh{����2P�#}�ͪm4����G�̃�C���u�xx�SI%�aևrv� �|���i�k�	�%=�L��K��������e\�?�H�{��F�f��U:�
����oT,�G�U���(:pK���� ��a�N����$(���U���=������T<nbI����uR��0꼤_�$�?��k�d�ӕ\�P�ae)�:���n�A�5��V|�vd�)Ӛ�͘�#��]�T���Js�~�w�I�͖�Hˬ!^�r���_�:�����۔V�O�8�s�n�?|�o�0�7dKL�
K��g�*O7�� �Et{0&B�O���B;�}��H �v�3���XL�_��O�	ZYs���t֖?TM�g��]\n
<�56Xz|� �v��cG�f����1��.[�5�M���٫��L~�T���4��N\Mb���h���[i&(��G	�ms>|��n&�-�aH�1�KҺpT�ȁ���a�;��CBrs��N �58�<�>��)&P���555�{8�<�u��#}i�wj�z�8m����`���&ds��gWD�ܮ�Fܟ�d*���|+'d
?;q/u75���59m�&��Je�m��X�1��+c��FuG��}b |ܺrNn�X-xCvm��\ (��6��U����U�L��X����I�K���a��a	�;F�:.�����ZY�yKW��q���,-�J�Ͱ��=�yC ��T�XvI2��R�P.�I-�ӿ��t��w�t�4<�f9�\�8��2��r,��B�p�L�(�
Ƅ݄�F�^P#���~���3�S}�r$Ըpf_6��b&�7'Kz��{xz�x��t�&�u���߮�������Q
M�����ۓ���
1���2����u�~&�")+�R_�`s������0�ʶx�d���|�_�����Z������2���]�em�t�yɏ�h+Xm3��ch��� �`�<����fI0e��>�N���[�N�o��^�~��҂�(�X`}����C ='+��/��#G�6�\��~T�F�(�n�m�`F�9��T��c��<����E �ſ��<���}_�9w&�x�(T�bi�_���^a���5�{�Sg7��cz�3bs��_Z��ߏ��"MEe��g�k��L�y�M�O��{��4�'6,e\?�&!,�vlY�XQ�b��L�0�<��nCrOȳ8��)����5-Jn\��х�o�Y֘?M�!�o�R��~������Z����!H���xO�>����ݙ���C�UG#��}�����[^�X��!�(2R���Vq$���l�\
�"0�;]�J���E�|���؆��z5���i���Ĥ���q��;aR3��x�v<�6V9������"�.�l��ߚ�e��X8�4c�<&��Ž�	���m�G�8�_?I����S�|���x�"��[ˑ/DG3!K�P�.�1st7{�����d��:�������v_ �����_s����I#����j���:k31���?s��N�x�C{�&��w��t�?nll���MB�@�++���ܲ��:��2�x�ի��lƿlMSb>!�	b�k��$�d
/��W�÷���aP(n��t�m�˂� ���ͩ,�C{�A���A�oRJW�Ɍ#;�����͵����I���IF]v/�M$�Mݩ�>#>��آPU���Ƽ�^�;�V�;�\h��b!�dv�����j[�`hN�o'v�6
�X�G$�ۉ��R�������Ud���� ��{���H���~Wt�Z�����E�~�+�`�Fw�X�c�Ix��2��sϖ-v��R��}*�}��	D�8 �K��ᣈ
����M2��8j-ٸ35e㩞G�"���S����u�oi��l�P���jE�
�Y�'������6I_��z���#
���5��<��[��D@�u�]�'���#��j0;&Ŏ�~s�Uc�5�Y'Ip7�ʶ>&��^]@aM�<����<n�B)۞u��N�����~Bj53��vs��|��o��O[g�X��Lyx�-�sɋ���7u���٣C.���
'�|s�ٌڟ6j�7��:�q��bɵ��⹡ �	N�4���#%2l��mf]�{�Tĉ���b��Q	�ۙ`�s�ճW=�rgv/,�t͖-������6;�Ƨ�fX�
�[6Fc�v��f��X�{*���$u�@
ճ�5j���·j]�օ��N����e?n蚘�<.T�k�ԙ�:8yy�jfZ2[����.���E��W�m�+��1�����9O�7Q��IB�lù"��=����nJ���4~�ߥB#Cܓ�t��.w�cj�U8� >���$}�kbbb�X�Xэ2���䤰�m���V@O#�"�e�3@&�c�i��|&�9'����.N������W��@;W����Z#)f���9�7r5"�	A"w7��������9�h%��iZ��e��z�������Uw��/k��4�Fc�Ž�{$E祥&� �9�u�N���M��LS�v�C��\����5����N��#5� >��Z�I�6�-j^�R�:dJ:�|\�x��%y��^�U�hD+����Cs����Li���)����ή��&V)o��`���a2�tn��lXXY��t�|�M>>��-\�Mm�+�P_?>o�]lVeQ?if�׌���E9
SdE�$%R�6�n�'���;��k��7�İ��iO�9S�M�M���qo1�����$Q��mį�|}�������$�ƕ�C/�ܾN��&m{!(�0�b �X�˟$U����hGe�g؀������2&�<�i@��.Kv|`\�U���J�8ОlN`SsT��cq18첢�Y.�,E�N �
�_��_v+k>� ����Q63I�6���i揃�ԉ4$^ݹ,G���F�p"�b4vVݤ}E�����k����$D�"�X��Jv���d��-]��9�XWm����x�'����
c��u����̮�������3�Z�����]�"��f~0��r�&�ۊ���z�5�W��bf*+�X6�dT�d��� Wb��މ�L���2?�R,�mK�w��?'N}��f8$
g�%a��Vf�ғ6���|yx�* s��Q����!��K���Bw�2��y���zV�'���i�R[V�;;�Ꞇ���tg�C�@+��h���U}�ڳ0
�QX&|��+�؜��Cʊ�C�7$�ι�>�T�p�0g�t�_y?�ņ�ՙ3q5 ���I��<y��������k?�!�����h)J��+�'��������8��ɓ�zim�U�V��?��(�#yc��pӉ��T�
� ^k��u=�a쳓;=%��٥h�S��6V!����Pk1�t��PE��C�YŖ���P��ae�Z�K蘻��9V�? ϡeѠ@%�(�ĩ��T7�Ư�����|�!霱�1|��	8c�I)Z8�YYY��_S��0R����w1�tp�F־[p�U�D����o���;�<F��Pv5S� dn�G���R�S����vʙԚ�U�57�{]���D�k�C�9l���1��������S��߮]�y�iG��i��>zF��1M7�@`�Ől����w��e�ǃJ��B����_����T��p�A< ��A1�69�}l�+t�MQ�Ӌ���O�0�W��w��
�͍��\16T'�Y����s��eo�s�Hd�.ɞ��~s`�#p>v����2�cB���`�giMS������st�$��+��Amh3{i�F��u��4��p�Li����hM�����M������#�tUZ�+8r�?���&��օ��/�����:�1���^܊�!@P�@/�[jjN�W\;�-$��̽��������l���嗗"�i�o�w2hZ���=_�H�%�$�S�cSԌz����B�������7:�_6h����0�Y��O )bt߯��DV��,%���՚�('�|�(w�>D5���\ӎ%<B��<L���.���'�6�_���&�G�Я�G!k��}m\�]5t>�m�Ί��إ�^=k�<Y�`n���~VX��1�8\�u� &Tм�0e������AՉ������D���,a�*����\I����� i�a57�����c����7Ӡ��	R+-s���F�����\�uC����S:��)�;<!�������������>z�+O�l���iI+-� s	h^�@����h�%q��#���O]��9R������uf���!V��Ёׇ�]����5��B�0�(��HX�>/�ܾ�a�ʹ�]w�?GhjE5ۿ2%��dT���&�x���۩�r���|9�P��%&X3=h61����G7�h�9�000+�`iя�:�|��	,�T/b	nR�<��Y^8�<M�نoy@�J�N��n�t��7d�} ;�v��iy��-��Ⱦ]����j[@�ڰ�֎�+���S�P$\4�����-6i�3H2�0�ogGn��K'��zl�w�_A�G~+��L@/��^�N��$�mh�^כ8ɘo��L���:<��q�؏��K{%r��Z�_,�!�2�S�X�Wq=���W�1�`�r�L��2�U*9��~P�8��q_[�v�h�H5�B�iv�[:C�@x�֚�������-���I�E�Ύ�F���ŏ��PZ�`%�'���+���$:S���"\��Yn]���2�$
L	�c�?�/!!�Tn>�q�D��߮�����������b�n����<b�'/+=޷O;&�B͝��B��2��~J�v_���_]���S�˫5��;����S`��B��I���j��l�F�.�/�F	5Lj�-�}/֤ݗ�:��\o���~;&C��P)j}�Mtiқ}B�.���֧�1�mszq��5�������ą �q�c���ax��g��������z��ȸ(ɬU�_WG5��P�#Z����l��ߐZ��ǿt p�0��&�վ��՚�?]�0u6w�t]X�@��^ӽ4��SU�(F�AK6��55�֏�Ch�$2g.��E���T�`��ZdҎ�ur>�-4�eX�=;�j�5���}���~��͖�Gl�����>WrJ�ңVr�1�Ms'��`a��ӹ�����xZw��4�A�v��$w����(w�_>�����;�g�
sZ�Q~%�,��GI��t��Թ%��9J���9t���	i��T�����$^��&ht��$,t)�����ݣ�_]竿q��߈D��Й�a�o��6՟�th�'M�Xjt��h�`|�U�~k����舿.@���S�I����fc���Q������9��g)3�x}�t	�:�J��H6 ⮇5�J���_�G8���1�](���k���Ա@��u;Y=����<6��K3ag��I��~�,�p&�ӶGd&��,-P9Ӡ�1�"�xL�E�%:��;�[�S.^3�<$ݟ�h����;0ȝ�DT9�=	�ul\�:��8���u�R�Y9sj���P"`c�=�ڋ^�NBA/O]ƛv�b2�=L��-3g=����$c�����B�x�hvK$S�C|NU�?�5fp���W ����I�fjm&����d̢8�rԓI���?)[��
���]��G��p9�$f�����293#t3Ik9���'G���\�/��9�0�L��n�[ƇY���֗��?�"����,�OÁc��j'����t2��C(�	� ��?��ƶ���|�9w�4�|�`��kѺh�L�"6}�Ϲ�SM�3��68(���R_��_�紊�;�v�=��c3�_�?��U-Cu�+v�5�#j>-�+�`|�Ɖ%�+��<�'v��Q!S�Mk����'��+)�q�.:7�S��h��(��D��~��֘�(�]�>��|M^��jl��CPv����o?���A�A��&�X�[������EG2!��8����iTK ����̜������[�RU
G=���{e�:6�P>�5;�_��8�'���hwb���,�T�$$����Oz���s1��xѻq��L�<G�ڬV��'
���?*o�G��q�aW �ej�l�fA[�BY:/�~�W�3�@����v�����5���y1����Ꝝ&33���G
����Ɖg��f�5m�giVK�bʽY�G�dw����?��Oj�I����g}�[��(�X��Zs�g��f�n�S�.�f+��]�!�$���M"��W[�jIi&�ӻeIL��_r��A�_K�:Cþ1�����Nu-�so���a�e�n�}�c���u��̑5�2�#Ԣ�WZ=Y���JT�D��
�q��ư��#������ǊI*���{;���!G����q|@���}z�(��1gm�.3|Ũ�4i�<���\�8:�t��Y^��]S�N=���p[{�Y
ʵ�մQG�!Z��f��LX���א  ��	�ֳ�,u�pv_G-���R���Q�E?̄�C��6��z^_�@�=mm�0٬���M?N��&�F#c�$)����lƝ�E%�ٕ�	U�g훵:�,OJtG�,���"���~8�=
7�1�J�p�|GA�H �yLj$ Pf#�!���,�	�8v�+�r�����	���ɧV�u#"9��:�F���J�k΅�Y�Mm�j��x>P��z�'*�����xҢCo-F+��̏锥�����ң�so��DU4�<������u��NY\S����m'|�zV���;z�VO���p�.8��zYY]���>�m����#�����`�e*��)g��45b .o�3�L�d����SA��Wsk�{�O
Ż���)�A!��R�G��ĮoT�`���_G;J������9���^�7V||��(�x�<LӛLޔ �	g�^&�D����Q��\��03GĶA���3�Xx�3��єh�򮜁o�0 }�`y�9i&��{�COa_����<��G��,�
S&h��(�vEh�8�R��;�C4�����#,ȗ%	@N�_�6�3�Ž[t�1g����r�q��9�f��vݯ�ƙO^�M��aږ]���>(|��Kd���*�u,�\�aG:�.|�e*	�L~&b�[J�6-ǁw�T�%^�w�9`�
�f�>��ŕ��;����d*B�#t"�8�/YIlk���%�x����(� ��m��:g�+p��S|V��w����j�ms�}�n��,nͬ6#��7Fq��x��0���M�ߩ�646��TWOX�4�����>���+^���b�8P��K��C)C���R��jQ�f�p���RX�H�r&�]��'��vn�0]Hw�=�%)/҈{I���1��{�ؿ�l�£����w=��I�r������%�r5U��тq��7�oh��A����f	T���!v�Cp�:�lI�<��X5Wמ��������D3/,f�!��:q�aΥ��eJ�@b�M�#�5��18��ı%�����8��o��u��z�L��)Ɏ}^[��HF�#��Y:��|؉�d��9i/�����ӷE�\��i��,���D���i-&�f�?�/�	�j(w�q�U\��q?�:�t�~���tԃ`b���A�+'U��jM�\!_rĂ� �\|��\��^�`���Q��.��c�É��f��)�Q��D���V0����{�-��Uh�t�׍�j��H�ƺ��J���!�����!��d�;�t�h;���U�};�Aw�j��O�S�~�>V�u���a���^�9E���M��"��8p�NHqC把^,��,s��Q�1,�!�@t;���ٙ�2��2:�7g��� ���z#L����B��LV�� Ū>�t�E�h�4N!�C�>���Җ���1��y��MXw\����_�	1~Gڬ�@��T��S��[��9J��|Ч��nG�k�͆��#;��xz,q-Q? 7.���D���1���tj���^�D9ȰV|��`1_DQ%�p�!~g]�/��}^��ȯ2��K�nc+�Cg~S� v���,�v�D`zS��=� F~1�P���f���	�2�(���qY�݊�<��Tɽn��!��iR�b���hn��i��-2;��Dȍ�.�#� �>2�T@�vV:u6���m�t��!v?!���S'�7-s�o���+k���A �d�����K��_V��T��֬vj�4p�M�;#ޣ���
�;������e-�,ʅ#/�ߚ����������3Qh��LP��]z��Y|��6��D�������)	@<��W�	��V���ϤoH��~/+�K�_�: ����'��r#q���,I�yz����T�v^��<0�rj���[������ޗ�}�yyU4 m��X�q�vm"D�L���yng,M�nk��8��� ���Y��'��-Se���?+cN�����xq�/�	�۪��w%ձ��	O����O�����Q�M�����^���s*G�3㾼ߏ9���GA�f>Ɠ3�8dM|ԣ-�C�]�Dkb�@�/�a�.�,�Vl	n<��	�S=6|n��%�p]�_�i����B���҄t�@�t$;�_�m��]�jr2�כ��x�� *����IfB1<�"�t�yx�Z�Y�������as'�����9�>]�@��UW�����w/2�?&����i�c�la���.8˝	�X��Z�L���ꑁ��c��� ��B,E�8��&st�册v/gx���U:�݉�8�Qۏ�?X>��:9j�<?\�F�ꑃL�j����V@,"��#�J��3}��Yo����V��l���0��R���b�:�J��ڹ��ԡ�c�����j��(�G�"&�v|:��t`A�J�(b�C.6�mz�����ݻt����b�r����`����:]+�1��!��ap�,��W��/���]H�.����#�XZZu'W]���<����KP &RQ�k�u�A�QIU�ؖQ�)���qmI�E�M
<)�n�Qιͬ���&��,�
��Z7��S)V��U_������N|�	�B��G�1���<fA1�(y7b�"(
����N3rd���3�1�/OO�yA���[���Ze+�&����_9��N�߽r��n�7g�̓��!��Om�?�ۼ�I�-v#Zg��NZؼ�b�<=M�`���ca�g`������~���%����ۢ�TF�϶V!_f��w�I�GJO�i�މ EZB���7����k|"[T.��`M���\um��'ҟGf��sq�DQ�4L�F��I�*|���#�9��*4�;}���M�Y���L��U�k �<n�J��am�G�>fI�^/Ō��2�����3��7�MW�$�R��k"���2�i�8뻰=������Uh��4�6
��<&Kw�)�2�̮p[�:ps�@Xȑ>�})�;>�:�r�ƙY䂎W����G<����$�f�G��^�[6�����c5$5	����
��L�4��{�F�ݰM�9�y����u�X��6xa��;j���x���D3�BZE(�p��Kq��U�"�����g@�ݦM�p(�R���r���� �(��ў0Tp�͒�힅����E}~.���9/��yC�V�7:��WAHi��%�QU�Y��1n����k��>�FL9v�f�sJFA��?r��Эj�Q�����6�'g^��,+H��E�������7�^��Q�~�"�cG��6�u5)T4TVc�6���/N����c�*W��f���hSv{���PSg�����뛾���-b4�	���R��3s��eL�����f�=��#�c�s�ȘF>����7�H��^:B�W8w4�7?��ȯ�i�6�Wwdi�2
��#�l�<)dٞOb�|N�^���Y��G8"��,���t�/��@F��ۈ�/;`�Io�V���%kn��|zE�>�S\��c���z4�4�
~�^�K��;�{����✞����BfI������n6��j�y��jEݨ}���������-��h׮ZR��sߧ$o��~�4{�~�R�-�.�	�y��d���#�E���T�Б��^>�t�����ʉ��2��+'5�w�`��>!���#�W2e���P���}�t�R�G�R�X�2ɻI����[c�����!U�O��]��.��$�$�����8�1�G�{��/��:	�yˌ3F���]>��J�qm����w�I�mr��͸K,ґ�]�f_:�l��w�;��4b�}"�KՔ=�~#ۢZ8n�ʹ���mA=�8�[�-h8�3gm)�C��/�<d��_�����O_[B{_6QJ��#;�3���Y	�=�p!P�xcwx�A��]ˋ�O�3XSV�l��-�!ٚ~���˳�6ItG�fK����B=�8�Ԏ���� 5L	�h��7]���!��"~�I~�T�v��n��3�>�х�[��q��j{ �Ipڡ����D�L{*G�B��;>�����
�j�=�_����b$��6c&Q�l�;:}�?t^nV���� �R��s��Ӄ�V(?%V��p�ݾ	V����Q ����/��Cr'F���^;qh�,�<y	'�x�Ȓ,y�"G�%�H�T�/�_H��x�b����
ڠ�MXQ���} M����8������8��gE�E"'��u�=G������`�<�������0Ύ�ݣ�wlװ}���-�u�!�[�j�+*_�}X��ʳ��'N��zl8���>rɝI����4�
)|����ɣm2tq���Pˠ1�L�^��<����#+>���=A�&Hý:�ǳ���'p씋�>�]�z��M^��z݆���'�5N��h��h�O��b��� �f���xƊa>�iA�1n�����S���Y���L�X�4w9S<vu�މ|2~���w[O+�0��͉$|��Ra����Po����Z\����RȪ����!�%S�y�����=q�����d[	��©���1�^Q'I��.��ɇ5�`�,@��G�O*��2�G�U9Y��އ��'>�yN*ն=ЙlQ�Pg�[4@��6����O)�ZD�ه�����gwx���.׹P,�j������Ξ������7�db19������E�E*��m�ou q�����"��"W��>M�M2��C�G}a5�<�������t����v�œN��(��h�F$�J���=�\�cCYw�wO�y�Vq��^7Sr��V��F�m�gW��f�~:¥ v�+#�2�B�0�#���������ҏ���Y�EE�W����9F*Y�S�Gd�����C�>����X�X�w>]���.7Z��Gx�zܒ����q}�K��ޤ�XU�^�����~�&?(畚��^��c��A����wm�<�h��%�a�"���B2#�*Թ��?2ح$�D'�Uo�Sl�z�r����YG��v7�};4r?P��₅���n�%�L��J� �<����d�2s^���r��Q̿lՉ=��t�$�������u��I��W�����v��߾�����8bc�}��/���-���1y� 	�F���u���63�,��鰕��}���4�h�)Mj]�]��F*>�O��K/�r�b��WSm��=��s��7|����E=��,P��&(���S�D>R�gꕇ7�g����������ڷ��T ���h���� _p|��5���F<���jɱ�X��F�j���y.�lY���~4��*`�Im xB2x����e-�o�A��5K�/)L�<�⺝�`��/�(�\ ����*
<��*��K�dƵ+W�̝Y�S3�Ԧ�m[)Ս�ql�ֵ��:8Z�姫�9��fM�e�I>X�[�3,�b�%8�/M�/�Q�����VB�8�&N��K�wQ.'��_�e
=��m����=n��;z��������;87����v��*
a�#�-޸9�������uvH�E��L�p�4k��n�=�� /�`���4s��e����;d��S����?�Z�)]�l)'�m�>6b��I�'/u
�p��ف*�5��7~� �b ̠2������Ҭ]�)�˞��˷��0��:��qF��Re�j,�Pt+`��n	,������O��,#���d���]*|��A���i��>��.8�����p�n�����`a&8��1R��o@������_�U � q|b?���E�~�Ј`�À&/��8N�~��X!!@k�4}�ͭ�?��`�jiy�ZV':3GM{�{_�6����n���PQ��o�w,�0s.U��4+�������-&�xZ�uGG��*����w�F�^{��l�H�+t�kt����zjO��a�O�W隧�:ߠ�z��s���t�e¡ 2���$�?����<�[(��VE����[b�U	ˬ7)���n�ˎ��H���"�ö��������9璿m���֙�{��s�띕��"��F�Jv�s�<Fn�\î�`�'NL����$��klE}��;$�V&��>"�q���'��GOg�+4t|�}tN}|�<��{�ߦ�^e[�\|�S�zi��8����8I�S��~R�<y�L�}��F�s@�����H��D����y���=iķ����fv)��4}(j��/Ц��m�f��̗Y~
��� ��������î3�7��c2M����v��>�D7�@wg*~�LCbS|"鋊��������4Zi6�gړ�f����:/�j���~p���Å���ƕK.�k�i�-���8��~����<�.�'���R�7i�U��q���d��`�ںnɻ��aMIr��>�\a8�� ��),m�B�273�wt��]��joPr
��ebw�4�Dw��Jڣ9�T�K���%���?+�w-�S�qvm��5��\[�O.�l?K1F��4O)���
�2a@���~��5=�2K���J\�h@G"z��E�h�u�-��W��1�&-w8���1s$�(_��1G�>��C<���F9V��ʠ���6�6��V����$ ��>�����<�E�h֚̈�I3ǹ��T�����HOk��V�'ԩksw	#�]A�ڇft3T���oW�L��1����bћY�J�+�qGӛL0�Ӧ�8s�����
X�1�"����v�d�^{�������
	o����F��D��OZ�a:߃4FNӱ'��q+��}u�	N�i���p�h��� a,A(�X�X�tu�x�����X����d�i���<�d�;5̘����0�Ob�)Ӛˎ����c�����+������5�h����j鿻
;�~�qn[�l�??W<��J�$?���g �%EeJ�$��d\���t]7�y��g+�{E�?� D���|�11(�$�������[M�sž�/�������É��F
[��o)��Z�h�� X�|�a ���+@Z;L��������u�����c�\;�1W[3��lB{�E8{6V��ӄ`',���g�Ȳ�,��e6J?c*q�g΀�h�fɺ_ũ�5E��l��>ޤ1��Q2Ųl����^b-P�ZR	lQȥM�j#��{�~�n¸9�v�D�k�~����b��:�!�F���@[F�&W,�>�6!"��]�m2�ڷ��WP�t�@&d��w��}���I���G>������ޱ�� b��I��y��˃l~ߜA'ɺ
����o�9�~Zc�֋�_�U� ��r|��j6-mӭ�W&���ԌPcw�+=�V�9��ҀP��u��������e�4N��_W*<�}*@?�Ԣ�M�ё
bx0o�[���槥ŅT:a Kw50؍�E��ޫn���������%���l�0��[�\P��q�� N#�3�ڒ��,�<�p�>�RJs�)/N�Z2��ie�F×s�߻�r3�ZV�6c���S-�/�5Ӱ��J�����~�Mj���x��.5k�$�$���q�Yw�wM�8��D��8��]���kw�'D��}8B}4Nc-����ESm����Ѕ�3#�&ΧUe�m�o�_J����Y͎��,9�,1��Ŷ��&�"�;��ɛ�m�R�/|���RъPfM؏��pV��\.Ee��f~'3��4�M���2v\����u ��F�=��GZ�"1�6�~�<����
��5�5����SfƹN���a����%�b?s�.��7��8B]��=�0��^�O����|�5�V���&m7;�1Z�D���Sg5�2�ō���ͧa:3���)����Y&�5�H��{*F��^X�-�=w��S�hfz�߁�/������1���m��p0�u����>p�7�����߷ab4����u�IXr�|n�dHu ~����?�
RN'�9��9$�,�B�:���A��N,1G���G4xUҶ��DX���г5tkmn�X\+�|oC�U���X��.�����/gdcA�ӫO�E*��n��ǙR��M�e���\��B�:�0��a�h}�}�t�ȑ�G�]�LFu5ё�Y~3ZtJ.���� &��ٳ�P�y����w�  �onm��r�&x>��#⥑�����ô�K�Ҕ�z��sy�V��c�8X21����~H9�јG�[�,
瑁�|J^c3�yLY�"sdyl��jƧ�vk�X��F�{2&�B��*j������{j���u���0 NFS>/�0��=�:�-~k��"���^�O!~q�����X突���9�#�z��<�f'���'��3�N�0�eKqu�v�
�`D��=g��&\�~��?��k�E�ь����/C�b�|:g�L�w]�dQ����S�6�{��]e��k�fa����r�{����5\���Y�$OY}��+�Y8t�'z��S���tcg�?pu�A�0"�t:[���z#䠠�hLYW����2��f�Jmc�i�T�T76����.6�7h_0Q����;1Ao������Z2���.~�Ņe]Qn�ptq��d_|�If|�h��cDp>0�ĸ8�\�'���9��������ё̸.4�2�!�NN9��n��1	��O_p�5��L��l'�1e>G��Bi>t��(�D/%�8ez�I��n$qd�����ǁ!cl��tq�+�y\�ƚt��������v����U���/�OL� IG�M���u�P��yLg3����=	���2㡬�ӵ��X��(���3��MK�}Y!2���Ȯ����h���ұ#�j�s�)Hkq���C�t:v1������h7����1l�/w,k@�����4{�<�Ŷ�-e��$�kL =�7��2�HǱR��b�l��bi�"!�m������
��MU}&S�n�ϖĻaP�_���#8W�fc���v7\�WP����-�&C����l��`'�&�^�~��Z�����?�`ƍɸ���"1`�8ґ��`�>�� �i���57�ƅe�t^F�߰�ASBs��ǚy!����ݔ�7Ge~�y�4	p���$�`k�%�-���s����4��j��]kS<��|��%�$�|��2�-��4�N�@z��-�0N@�uK0�0����9�������)c�~�w���qɮ�y�'��?�>v��59[ ��Q�ě9�Z�צ�pM�
%��j� U\�ʝI2�:�ϑ�'!F7���o%�se��c0����djWp���C�A����pU�~�h<]���cK#
�`�И�x�߸�Z5|���w�57S��M�'��ӄX2���T�B���7 \���:��vV�]���{8k0�Z��D����=��'�����s�2*{ֲ���qJ�I��`�L��O^������i��QRQ4����VZ��A떖R�*�I0�P��4֥Xu��q���𖠥��`b*��m�}��R3��R�v�=��76?�x�{)��uf-S3s��r牬��%�r���;>�|I�Kj��;[ָ��U���q9(2�i�%�h����_��9�X�LP�H����ѕ+W*@���$��&ѤE�o�=��l�q��`�a��<tII��3��r4s'�\R����U�/�S�Vt�WI��x��A�N8�/-���.�D�l�4{��G(؋����]~�n����o3�y���Z�\R�G�ѥ� �aLH�@���7��t3��l+��se7c^��i�؍h$W\���F�'��Or������� �S�=��q[r��Z��f~.e��&�-?��瘽�9�p�����ݣ�}/��G�}��Gf����H�T��1<v]o�O����{��[�*@?`4���4:�;3�H�+�X�A
?8L��`��O����l��ڍ4��fV�M�!���i =�?K�F`((8��+���.W�������Y�X�Ջ��%=E;u�7�\��uߍ�|Z��GE�M_�u���y&F~��?��w�Zy���@I�@k"���Z^���uı��{�ךx��c��s��'�����۾���{���j�!�Ț��:���M9�.}�O����z��'�35�5�De ��Y�~L���Eͷ8V=�_wT>���b��n�I��Efrsϕs�a��^�w1������1�$7� :ϙ$Δ�2�(�u�@��A�0�E�K��������.�
0�f�j7�^�H%�����˥�4���:�9��Mse7���Vz�2)EۓuI��GE#[���)�(7KE�,۾�V2_!ɝw�=�׵��g�M�IJ�J�vs1-4$%/��8����鎮�~������O��o|�v��gj��AvE;��'���}����R���cKw�(3�y'e��y��ױ�][���ywP&��N��&�cma��|6寧;����~�\|}D� Ie�I�)}����P���#o:�4l@�~�f��Y9�2��b=th9MG�~ zh^��H5�-> �ɱ3觓 ����G�?�Uz��[����s#A�&�*e{��~��ȳu��V_��~̗���{�:�ʛ��~���͇f�������#w�q�ƈh���-�ˎ�Jgm��ӹ�INO��$�f��ѕ�8��0��d�[�����lkOٻ܍����������L�����ϵ�I;{O��{���o-`ǹ�f����I5n����t�KE;c��N��Y^�&g�Q������k-�u3k!W�t�Y���\��A�d� r�3Aj=�T�#b��d2�o"�q\����1�x��٪�����c; ]J�&�$ME���Q' n���o���`W&,���6�e�*߹��� Y�2i?�y�fM�e��Z�:n��M�݀c1>���7S#�c�\7����Q����sZ7��#�[��E��[���W������>���1�&q��x��jW�����|�/�nW�,<�l睃��y�t����>W�SK��/_��-7$iХ�UжB�s���>�L���NV�^�o���O���bJn����S������u�yI;��Dp|6�������m��em�2�1��Fźi4�m�T��"5B�'�l0�Y*{�3ae��Ke�ü�!~�����cK�a��T�]� +�62M.��3ۘncg��
$ Ϩ��(ņ0���wT�����k<.dL����ͼC���r��n�Ur�9@��0i���o���
i����UlA�|����5�]�oQ/��|�̴�+rm�H����2����	`��i�u���A^`ȿeU`�O:]X��H�I��P��I>�:
h%��o�&�w�$I����
�3v�����Ȁ���W�b�k�k��Z�N+�J_A=L?)��:�IL��(���P&W[��)gR�ݮ?O�+3�?���K�7���V�����ܤ����C��<�s��V�����F<��N�n���n���g�=�h\x?%P��P?�E`�q;o��/���9�,R"���f�9�u����Ϲ��;�3�HH@$�A��<*Z�s�$�AT�Ȕ5P��°ͺy�G[^"�<b�)�6��{�-L�$�̹"XX�y��3�q�]���̔��,'�������[l�A9zczl��/��N�Y�י��2�_������9൛�o�cmr��gd����zIQ㇟����AD����&w����<��$��a���}���(Z,D�+��y��}�'w��HvA6��|X-�f��>A��XP{�n¥}ûY�W�1����~&�_]�(��7�E��37v
2@��ƚ
j>�#�2�b���2��v�K��;X'�2'�&�Fc��-UzE�r�ȏ�؋c=#$Qʈb�V�f��p Xl�c@�$�69��O�[�1{��nR�mb���/�u���RY���L޶��x_|�$��6��R���_$ۄ,�?o�2mg�<s��Y�.����1���������o�����8�}�iT��{J_�'7��sǻ�����E�Ҍ��꾎/ݽ��y =�,*�W�ǽ��J�l��i�k���vٸ��P&�(v�y�+[F,�궩�PjgX�M��8u-JwH��0��{�4�~3����  �c �����.t%7?mj��#�Z���灮Ǯ�͎f�k�����F�	M�w�s�; �ǘ��u���ff���i�?�o�A��N�wZP�rH����O�<�O׺�.�U�~�E���,0ؽ@���-6��ڲ񿨳���wF�aOPo��~s���F����3�����\���fѨ�t(�>����/������Ai���:ݾ���h6��=�ˮ�s��~��Zӌ�Z4l�+���o}IS�Z��׬p��9|i��z��}i���޻��y9*�s}E�!���JC��7C(�JQ�iZ5����)"�R1pŴ.����l��5l[���d��}R�M�I�
 tT�ߊ~7�|�6.綵G}��Y�n��@ʟ��n/z���v�ws��>���<h1RS �2F�H����ZH�-1E:���a�q�~��7~7�x�<��d�����8ϊP�.c{�wR��'%�+^c�&�y�)n�Ͻ�7;HD��Z�f�+�^��{�Tn_�i����k[���AR�`��Fq��Q��׫ �����t��z҄��T$w�M*�:��6l�E��k�������noӦ�,�T�
��%2^�T�*���(�ҊG���K���Q�\�J�2�ty^{3�]DeFSK�w;sLQSJ�ɵ�5ݱ�c%�M�f>�Uo��8h�gϞ��h�#�8BX���}�*hzS��;g{[(����~��f��v7���͘��X���ݧD�kh�Z��ǅ�!�&7��"'[�y�ys\��$�,�#��u�8e�i�B�'t7;t�	�Su@��D4����_������4ƀF%�U�q�'�M�*�/�<�f�,���o˧^�l�8�ҹ :��)D�'�)s���tVs���NM��ӍŬ˛nP��q�$lץN5|�M���5�:#8�Gѧ�X�.��UYz{
�ڀP��,h�6S����O������fh�v�����a��ݸL�˺�o���93��s�e;���q��7��b&M4���HeB�*h��U���TzN�m�&��f�/��s�����x�`oo+�7s���Ӂ��X��-���۳����욱����\�sjA23�#EEe�iԣ�8 � ��ϟ~����^wy���fo��d�Y�M
<�s�h�z^d~ִ���J�G�h��5z q���Xx.!XU�Ä�- ڜ.���'Q� ���|%>�$J8�1��-e��q�ۭ�QQn�����c�r���%)����޴��L(QC�1��y�y�E����4��pL�F���b���˂�9�����M<����Mt�p�ܔ����� �@v%$Q��T�o5��V[Z�c�׿���裏X��1h�#Ld,�*�4� ��Q�ޙ���q�#�Gz�'�$y?|�wMߋМ
f��,���I�> �9��;/!�~I>�eɐ�;�s�6���t770��^j��@USCB�L(�^r���9��P��I?�wO�+�/�8�}��qm���oL���B�Z��A~y=`�"��H��I�3#h��HkS��E1� U=G�9�X8Q=sc{�$[gXoևo��V�}�t��a�6/|i���W���ô���R�<�
�c7��v�u�b&�h� 2���Xb4{i�!vi�@�k�1��k������}B`���$N��;6�2`OrE�-�3�[�g��g�9��L�1�M�����]'�H���eZżmn2k����Aڴ����<t���/_�Xsn�k�A��Ǐ��J�L�s��~Y(�}���|���*�n��mMУ��N�s^�i�:v��n�jO���t��X�zJ��ԅ�M,们]�\'&���@����v�G쇱�$�=�2�YG��ɟ�ɟT>�>�t�R@��4���t�� @G�kU%�t�2�Y����E��^�mO�����0}~s��OM�ऋ�(k��>�������F'�d�o�G�-�3��&�I]�����Nsl�SqZ��w5���T��a��\3EqfΚ%�A�p}�[`��/��/\4V�,fA�5�p���g��|��t�'I�u��
��ˬ�E����1\b��7^���8����ce��y'���L�����}���<��tlY�D��,ZF��n�n�c�#�%�$V)`�bMӹ�
��	�2��������vZU�~��4�pg�wdE��c0���4���$�e�3�[K� ٚjԌ� ��d:����x�}ަ��k��k{�k��9�O�2@/��kN��q.𖯎��,���7N��@�T�$�F�[��#�m�ܧŷ��m���>rϞ�^tt��� �YK�U�.֗��d��������>w3��N�X|��i���>����gn����{�o��^v/"�&ŕ�~6�#)���,He�5s�@l�����FK2��j�V������\3)G���Fq
�R���s�7�i-��USCu���D��F�ӆ�zi�gZĥ��d/*3��fw�(S��ڥ#ט�u�1Q��A4�Ӕ9 �])N3�K9qd�e�PԔ�~���E����XK%%���t
;��}�tA��|G�uٗ��߉sσ��n�9`� �2��y�q���Cʴ%��L�3��pMXr�2�ŋ�F���Xm%E�R�o^ʼ%/��N���/�����5��gN��y�i��
i `A /�U�_1`0�j�dc�:�D�g��}ʹxU��g7�������y �-+F��%��;��(�uM���&G�|���\����r�{��5t}_�������m�u�����x<��[TT���p쏧Q�&k��L�\��r�hQz�����dkkR�%e�Tb��I&������s��%�^_[�Ƙ10�2���ʘ����+c=q��"��뗕��K#)�^�~�ȼ�˶�|Y|��@�b�Ec��y����r�K��׷�E�w����S�|�ڃ�`�����I��f����to[Lʏ+
ni���S9�c��^P%ml`�o.fx�O�[P(�U��)��m[��(sKqZ�x��AO��P� � ��N���-VO�f[��% �ry�h�l�[xj6봦=L#�Y��r����$ҝ�t���Fw�u�׵'�}/ezQJ�%�#5��_�>T���S���_'���ȳO���䙬z�s�1�Q�����m�c�y�)b��d5�F5bv�q��B� }0���{G]�t�#���@z`��'H2&r%`5W����x�E�F�)7�\~�Ԛ����mr���K�)����4� �� �
&wy�sn���l)�KY�����{n������7۵$ǲi�9w�1�!�TU�[�'��OH?Ѐ~C�*�@
�74$�u�R�s����̈��2"��g2k.��ܤ�fv��q��l���k�F#��Ľŵԉ�`�h�i��טP�����?��1[����Ə��.��Y7�u�lv��z�}q ��"Z��F�Rk�%a5�'nY-_�Q�=�քc��ڨ˱�ݪ�*m�H�N�쇠W��]�7fՊ	ֺsQ⪭�D�[��Y��H���#21�n�l)m��v��=R�DJ@sA$��{����܇�*�~��H�H�cL$^�J%�����	*1��j7a�g��R�)�L�ؘc�\�>#}֘�f�n����D8��߹�7�)� 9�������z�S羚��ms|�; ��^i0Gԃe�z$m�;r� ��u�!Ψ��tNn��FN���3�0�0O��E�v�o�9H�6QBoT����2�u1�76�w=����"� �6�Ie�l)������&CJQ�\��u����𰦮u^%��Z�&�����WϮ���zѪ�ɱ�E��#��g�|�>��3��7�F�e�ͽ���۝I8�.��������zgީ�k�$�H�����#�+Q^��{T��g�?���}��ɿS�4=��V���|1^9���W7d%d�ªj�(�SÈ����۝�ŀ%�GG�_7cﻝ�[��uf�+�y̚�-����٬P��ۜYpS����.Y �Q]o'��Z��_"�<���dO@2�N�D٨n �	c���v+���-)�p?�� &���ZrС�.e,��~x������%�+yR!�.q��2�g͹&}��R�b�K��>�����7�1���V�Ҩ�T���޹,'������Sn�FT���ʋ�ٌ�O�y_'��Оc4��9��3%�rz��� X}��t�l~���aN\������̓��~�WC$��f��l���XK�h{O<@$G�s o#oe��#Y:��r�w�y��ju/��T�)kCN'z���Y�݄�ua�R�����a9��%|�J,�
�ȉ$��DI���^�HuF���D�����9V+�7g'-�l�ݲ1�U0h`ʞ<y���^��>�H�|�\��إ�*hq"iο�x��*�U�]����~������ic~L3�u��^�u��ۧ߱�]��仧���%���6�a�K��߽�B�.�0�빮g~��;�̲��5�Ȍ�Ԩ�� ��\�rV�l�zEtqq��|�vNB'�x�UFG���.�ܘ������� M˨P�W�[&A s`�"���폫�R	�e�:Tp�J���l��sCU��G\'�IU�~?y/U�{��y��4�d��it>�ӧO�7���O����r�X���Y�'���7�rϵu�1�n_���=�n�}\�!�]�cE^g�+��1Wof����:t�'u��gVZ���&��N������f���������N ����ő�w��	.T��ن�j[z���[��'�k��^�RI*�+��T���껭�"Ќ�����D鵩
�� ��Y�D��JLL�z�FIU\&&Q!�ӻs��Ș�9G�����;voZ�ν�q�s�6��F���{�LZ����͒52c� >�j\&��7�vn�mf�o�}R����H%���2�T\�9�稰�\�k�̔�Eٶ��`�Z��~����Iu��T74��2v�$-�e�5��U\p��Τ�,l��&�L�0:���3����k�gԹ�¶Kt{�}�iT��s콶� ��م��t�.�Ԩ�]xO	�T��;�8m� 2����֤�R���`��?F
zg$�8�l*��#å�&9k)���ݧ���X*�_
�U���L�e5:�ANo�k�@2DS^�x-M1O����pP�#��@�[&�r���y%�$�\{��^w4�vw��e�HS��-3������}�%rR}���4J�q���Js�^�����)jIq�${�sRc�<;}��,vgggw�c�I@�G�%��{�e �ƙ�D��x�w/�љ�`n9�&Z{�Iߧ�J.�l.̢�(i����^�~����N��R�8ݥ��J��u�p�sZ>[�%�
v�̻�*����3u��#���I��$h����o�I�v8���8��ܘ��	�F-a����qI�#$�������S^��P�J�n�\�zu�p��u���U�=����~~�X�'田b�y
0�Ś��$��'Nk��򻺮6�������vP����?�i�7���!K)��uN-Iޤ�&�������T�}m@�Q�X�h��%�ʫ����X�\LQ�ُ=�K�^�XE�a2��\rw�q���U�l�T�����|_�4�)'�vJ�c�9RD��W�R���3�M�}��ϟ?���f��S�l�����0��4��5Rظ����?��gӂ*�����@c}j�L�ޡ��������[]�����%f�rݔ�/�TpԨỈ���F����Nq�}���_���?���D�7�l�X�./9�Rt���s3i������k�f���z���ugS����pw���'g���q�Jĩ���ٝ�ײm����L/�&o]�d'�8W����m��j&��lQ/�bp'U��]2흂��Y��=���Y|�����hkP�q�5fx�q��c������%&o�ګ��&v��#��5Ad~�_�g��h ���Kurt��?����#�u�����<�Q��:�m*{NӮ��L �y�U��xb}��T����LrbS�����$��S�dJ��^_M>a�|)�|Ȓ羽
�P��e�wcB�_�3Qٸ�&}r�(��y˯{_��ncI��ѓ������%�\��$h���#�qᦍ)�mL�ʣ���`���X4�����0݃'=^���/�~��'-a7�?���J�73��W���^[S��)���H��a�
�C�X��g4�9�6p�~uO�ʞR�G���8iĿm~�U�	�o?��v�R��6��l2��p���7T�3x4���#:�'���ɮf�-[ÄS����pB�g*I��y��T��2��T�Z��ʒ�^2��n�����3���!è��;�+�׌�����d'{-�"'N���Zϋ۵f����}�(q;]nڨ�j� ���t�m��|�Ӏ�%gLS��
�9��	�8�	��QR��Ξ��i��l�<�QB��kQ���\SU���|=��S�J���I�=����}�=d]%����^�y@�6�%�)�e<�f���z�'<x�#�+�3�LI�\o b��<�!��~���������i�_	䫮�fUx���xIA�N z~�Z3 Wx�i4Nv�n��� tu�� ������v�۞�]�`G�D�8���\�%��A�%��v����\�ty^�*+J���s`'UwP핗�(�P����]�nJ��j)ƮL��I LSb
��ߌ����.uCXL�>���C����T��[�	a˶��7�Pp�u`�6C�۵�LD�n�c���&?��Qn|_��ffmjo�l��g��d.��	�]_G���܄{���� ��� �z5��wj�Y���֧N179�:�`� L�Usɑ�Jj��x�HI����{�v���V��y��u�y]%�XU7����s&$J��������4 �Mk�K��j �9����J���g~uC�qY�|U�Y�X�y���3�|x� �������b�ʀ�4�����[�F�����sڼĄ�7w�l^'�; }X';O d5����=@������V������j�jW���H.xLJ���	�(U��kj��$R^'U��VR�B{�u�����$�)*�%�4.�w��(���T�6�x���3DG�R���_�.L���);QСV���믿68�l�;b!7J$�Kf��.E�G"����3�5�g����4W2�dr����f^�l�0�+�}d?J���7���c��
R���t �{BZ�m/�ϟn����r�v��*�4�+�}LrJA�r���(9"Ӡ��c,���н���[5�p\1���k]����P�15}�Wt�,��e���/3C%�2_���:>brc��o��_>�~�_X@_�%��v5�w��5���a���| 8H�w�J�W��R�:�{��6}�r��rq�N�p7��jk~�|@� `��F�Bp�ֶ��s}�F�s: �=���]o��4H�o��
�rl�X��a=�Cl�T.���ħ&Ҝ�%��� &���^,$���:����Tǩ�%5����P�$ߟϡ���4�0J �V���O>QϿ�^����՘t�1�ԉ��*��%0iv(��� X�Z��8�ݡ��v��
�&��H��~H���wd`�^x�� �.ty	�@��v�E[7�!���;&��(r�9۹��v[��U�L^�r�HTx.���?<�������%s�'��o�k�#���x���k��r���8/#ե̈� H����jZ��%���:�s֯���&�Ū�����R%.7�U}��)V��:[��Ew,E{�ͷ�o������^����ڵ�gg��tn�a�l���F[�}�YQL.n�U'����o"�|����uO���'�������Fe�^5�1U��G������.vI����$U�=���}/�;ӿ\r��˕5)=y���2��pgm�ȹ>��C	����k`��&B�B����hZ#L8� &6�ܯ�s�� ����Ͽ_j	����&���ؔ�yI\��2,c%S�w)���`��W��9[> ���/��uJ�n��^MO@Rr�i
Ƥ�t�Kۥ��|�����R O�ܢ�!�����B%%�+T�0� v;���>�`��J9������Q��*�]��Y,���������)x[�%l=F6Z ��a_A@�'��˳����T�o�N�%�)�;��vJ��Τt�w =J������K֐��	��Ui�-����:�m����K��TzM�=���o����T�܏������H��Z9�B��d��'�nm�hs�l�w�?��������)wm�=8�u�o̀��(�}5 �/�4n�	��������������1�I;�QZ.�w4pvާ�3���Xy`5Pn��`�s�AB?Ы���/h�<�\X4����7U�� ��2"��4�� ��a�M�� H~�\��ً~�'$G��F�k�~�F�g����Z�;T奧�kߕj���;�����l	�ҤB{"�����g�ٳg�^��:�NЙֱ�<��z��=���|$l9�����o�nJ�s5�9�J�G��ý6a�w��{m&Ie����a�8�e��5̨{N@��_��]������(��7��\o.m�$	�Re,��#�Q�l9ʨ��+�$�v[��hb�SJS��jby��ڪU�> ��7�0xR��<F��t���/�4�1[�/+�˪��ٰϢ�o���8���f�@S��|�(Ge��:)�[I���.�K�C%@(M�S�\�q�����o�0�-ɀVv,vX�^uZPh5�/UX�ҋ��o�Q�.݃���'fqA�vP��q���{�t �{@�~�i�Z]�jI���H�/j^�R7��ƙ��R8@���3�u:�B|���������̻�����)p�ir6�e��U|��O���$�����19�N���;�c*�!:��pO�<1��n����%7!�RwjO���۟W��A��{��.�U:P ؖ�,+����u�ݜ�1�C�.?*��^�_�9���~�WB��"lݒ����J=�o9�������h��P�Dε�#��μR8��\�&=��L������$�{WIs%�!8���8��Q�z2>c`�2%M ��������9���>�k�ڜ�}� m�}�s&�e7��%F!w�Ա��t��%�mqV����A�:��-�n�TT�bN��3��WX��������5 O:�F�C��*�ؗ��d� �����#\j���<h7A�L;�群�]ݛv�q_���ͫ}i�R1�2�r�N��%��?/�^XY7�$�����~��u|G�<�e���q���e:ۃB{��%Ʋ|�wL��3�
�;J}"o�?��Џ�X�ѾH��>_�&��Q�0�:�n}�o��߫�ʞT1ձ����R�羝 ���� ��}ҝ����ݮ��Υ�t�С��3�� =��C������w�o��4�5\E�Nm�x��E�c�T��/��ܗ
1ڱ�*��v�$D����@���2e�1�U�U�{�ڽ�����kcy�W�_��*�ف)I�r���R��^��.ݴ�)� ��i� e.T�4����@����]o���Y�ԭ��z����n�S���}�����?��o���B���@�m�sݲ3�Ydj�ܻ�����S��D�ڈN����{a�f���mƿ 0A�n�f/wʌ�8s���b��I���ě�Ю�*w
l'����w�L Y_��*q�ܳ6)U}*]�=����+Ø^��&B\S�߇�`��"���[�m7^�hƣ��v�XSY������t]8����~���� �@�O��ݶ{�w���aB�l�%P^
scK�g��:ۋ/<pé����
׀d0��_W�d-��xn�:5�[��n����X����,���o��<,�cL�U����p\Vs	G��U�WѷX6m,��#���՘�������Ř�fj�]c�t��uusu��:����W���|���<����$���=MI{Q ��ӂ�m�Nq� ���Js�d�
b����B�q�Q�������m��3)c������V��/
Zg�8�>O:ߗ;�7��%�����S�$$Īs����i��}@�vl���Ki���ҠZ�l	[�s7ѧr��(�`~"�����[��"�ܫ���Ԩx���(��E
{OJ!i~��(Ml1fFyH�<����B-�R���Q>��b�\�4��M��Z�!��.�U����wCSM��L5��r�6��֒+r��Q��Or
C��iS&�W��n@ܬS3�x���oZA.��!C�Cm�e�ґPp� ���.k��{,��N:޴;�jP�m|�pQ�J���1(�Ğ�&�6��|O�V�Rw�L�|�!3�7+�7D߿��Y[��w$�3=��<�9�Wt�%p�~���ڢ�`�c�3��e�3�rì:}y��� .�/2��VR���6��-ʃy�h�_�F�Bs��݉ϫԎ����N�Z�!�k^���f�c����պ��z�;0��-,���倝V�C�(rh�{��P�6F�`>Y��TOn��M�����.�W��	Y}{y}BR?(��1t�9b$�����Kq��E�о�E�E���lN{*�F�U���}�T�x^�ӻ�c�>�^��?Bű���.}tb\�n?��"���y��R�)
�
Ԉ�
��^�}��!�d�T�f 1/�b#��Vl07��	t��s�s����ae�W��3�E>&cž������)<BJ��fө6�t`��c��$s{�q�9�a�Y��<9��갺"{@�.�ª�Ă�Ϙ�g��0��&���/y�ռ��m�{���.�AJR�ۯet�܎�x���.�w�O�Mt7���5�Uq�B/"�^y��EL=ؑ�П1}2�����Q���/����g��Y�:Oc(,TfRf�Mzi7��g�uh�ϖk�W���HD�v�D�<b�Tffl؇TҘiĪr&_l�!��n�7��,�o��Ŧm2=�rC*4MEL�4��U��q��j2=b�`��8��'�4$�9�Y^�VQ�'�[���(Mw"�6c�7s��a�m��L��ND����m���N+P��с���Dd3k�nߎ�T�d����V������C��D���
dc�;�(�� w�
�s���n�;��i�U���/�|�n6�Z!uc��r��L�VE�	=ܫ�Ff@E{��xMfIף��1'��G� e�Ŋg�^�رK�T���{�\�V����w���N��k�"�gIC��;���;E.���]�|wSSZ
�EΟ��|�t��=��� ��`)���������@����>;�g��E��-"��f���l����=ȎDo�߷-M�B �ڲ����U�(�MV���%���t_����ˈf�/�
��5�l�U��I{�GX��co�-m��{�Z��΂��&;iE��]&���Q@�	�n�̩����a���
�T.��0(Ŭ����iÔ�ș�m�ʚ^�wQԣ��h�� �	��5CqR-K��ˋ��s�Z��[nw�b��Ddn�ser�BI��ϱ��W�;jkN7�c�GD��*dB4G;ت���Jd�||��D�$,"<�3��R��+�(��_�~O����e>��:є�G@���IH��4�CHF��`�
��UJq0Xʓ_a[.�u�j�qߍx_VB�2ɼ�Њ��O��\[��0�=��F�Z�ž#>�- Xǈ��%� �I���g0�+S2W�I�8�ⴸ!}}w�K�n�j��Q�[�qv�p&!�7S�J(���f��*��,i�����0]��?.ɢv�N�4ݟ<�����i��`��.���0ώ�g&McC�~!>��^ކre������>�v�]�{]~r����?X%�.�:����P޽F������'���!.8R�`#K�yq=C�3���l�j����f��ﷷ5L|�&	.m�ܒ�;<bxA��dZj��n��Vh���ݢA]�c�N�m��!Bkj(V���|���9~s�����NH�t�@R$[��o�y��A���L�~�b�R�O&���wQL�_��)�`�9wO2�`^l��\(2����Э�d�*����l?�ia&e�kP��g�)��_&8�����~��,�y��{]YYK�q̆��ez-�,u��Rq9�DtS�Q��ey˚��E���bb%�B���	���k?ڠ+\V;�%�t�&f6,ŠV�)����Q��e7=���'�P��s�t��㻬�߀��~������� �d��Ra�+ȇ�Zl�X�ƾ��I泇��Y�+5��<��M���)�>v|[~����sb	l�'5��Ǣ���l�#U\��;��b�V��>�g���q !@���s,L�Zƒjn`*J���n<�W[IE��Q�h�O��{G�q�)��K��;���O��Q��SZ�&Q2A7�d{�����$6x���U@X,��	�>=?�'�j���0�d5G�1E8���q	�N��=Ly�h��pK{!m���o�������F�T���c�_/�ء=����)�r��y~@`I�O�L\�_�?=�����m�U61Gr�_ߟ�˂1�ALIhL�8Q݆e�ɪ:,Y'��Ǖ����Ӹ\��s*vg"��m`ۗ�E-G&%���A���ʜ>r!(�i�]pNewA��׋6�����S�X����˒��P^�Ûֳ�������l�!�V���i1L��/iÝ�p�6�:��j�[���㓙ot��/o3�`�߮o�ޱ\��X�#}?:��X,�q��%��C��Z���ά�x�#Q�h#�G�ry�w*�4��ձ�2�&�$H���H� F�BG8�(4��C���Y>^�2�S=~����%�v}�(c�	H�:�3u=�]���e���u$��茇@�l�:����������5j���������-y��<���b���*��-�����,<����O�t�!7�C�><��͡��Ү�̇��8Ѿ�3�֣�Θ���E֔�<V3(�x�'��J�>�K��c=G�~ގ��J5y�]�dC�>Q�FQ���&t�gj�kC�A\�Ď,y�$�e�?acU��|��^�u�e-e�V�L����"�Lf������ES�H��I}���D1ȗ��.y�w&�i���a`�Y����n.~k��+�flH&xU�n�h��h����W���Y��裑l�PI�!�;R0��~2�%��D�A�yR��:��Ɖ���Hٵ�����6F�"q"�)^��r����Kuʲ�g�-&7�owK��2X͕�\�*̯@A½����^�{Ż{o٣��W���Ud�K))��ov�O���(���v�WSƿ�_'�����q�S�BENn�~����.�ˎ$W;GU0J��6����#����4ܯ2�pRNi&RhqqԔ��㘶Wɍ��W����g{��l��4N�癰�]Ł PӇi�p7�KV�7��Ŵ���R�����g����V�,�������YF�}_�Ywn=�Cvl>���3�&il��ԆYa��_)O�|�$�q!4�l�i�X��gR0�/:3���l޹�L����%O���-� ��Z>ɋss��?vǡ�m�e��_��GV�����х�Q<V�	,���8�e,lꧣ�a�ݟ����K2����#�������v��ϻW�S�(3B[NE$��uP1V1��Vh���I�k�ԝY���X�u�ur��UB�j$�������O�TE"oRq"�+!�o�A��A�b����!�-��]ʩ�����o�Д���XH*��m���g�z�7;����'��D��"���u����37W&]��!��J��B�o^�܋Y�҅40�#���~��C�����_�j_@ɵr���j)�Z�ɪ��/�Ax?h��9Ҟ�+G���q��g�m�#��Z}�n�2��=0�U�g��Ln�+�K�l�S�]��ih�M���,]x�P�����̍B0��\�r�$YG�b9q�l-N�"7��⦣[���}mX$�>���1+����?�&�2�8��i�L���<�@HQD!��y�3�l8��l�.�t�+p��~���Ӝ�O��$���DW1��#d����h�FA��� %If���!ƮC���m�A��KZ�U�rw*O� �*�#o�סn�v�աGw��2�9�W�EDT�- �x1��Jݕ��Q�y���}3�S�z�t�(섅}��gɓ�Y5��� �zM�'����o���C�Z���lSF-6��5O�\�N��Z������|P Q!��ɳ��Bo�"~`t���'/�V�.����-�<�n�r_�����O���Gp���YD������.?��������Th�� *=͝���i0���[,ۅn��� RZh�6+l�t���5p������wx�R[��E���G�{��$k�k�\��M���V�M���D:_,gțY��fы�@nR���Z�G����C�z(9N�f��mO}��[��^0��8c=�	[�c��ދl�� ��՛�U�!'�$�4�j���K�]#_���0��3�"f�\&���v`3YK���}������F�Fn���{υ�n��ν���N�^Bɘ��s_t����x���QNI�:\�Y;{��#p��:ʊ��|n��U�;���R�h�T��b�	
�Rx<�B}�aN�k���Ks8_L^�5iZ�6��} ��"HC��;
�@~Pf�-k&M�jN���zzT󓖫j��Q�.�I���K	%R�u�RCc��T�*j����ҟ��f�T��5Ą�W�'@Tm�5Q>ʻ���>�տc��٦�0�b��y�4������8]ĝ.�O�p��j3����u��}p(qB/]��Z�Q�3s��G�6�qp��	�a@Qxxxm��z��}�]�h^�l�o^+�b� �Nۨh�Y��EUg�R�!��d������8��Ojպg�tݮ�%ʚA���oI���~u���g>QHdO��
�5���]�V2�!�y�o���[��?q40 �?�#��s-H[��}���2�0�����i�p{x�|`
���n9%:Q����0��n�˪�m�$�Ni���rD�!��5U�a���^Rr�4ND�;��s2&�ؙH��yr{�pє�ap��3���u��`�z��� ���E�F��\�Y�q�B���a�'��w�]�8���l�O��i{�N����F�8�*ۨ�_�����k��V G/�\�͒W��7�k�~	���Mb���8>߯�؎��E�,��W�f�\L�m���~���]�E1��pZ�V���2�:�/�����6j`�6�H)�&V���!��h��8�{z�5p�ȯ2��3A�U|�ZLֽ5��DUJ#hZ$~�h�\�z|�t� �*5ZS'�<�y�\�P��L�n��)��Ȧ��P� '�������7��l�����PA=Y��$i�*�5��<�2
��]������}ֱ?�1o1���j�tɷ�M�<d�!�� >��M�i�E0����L�K�fTQ/R�!L�|�*j:2<���E�}�(V���nE�D�(��%����߃�f+1A��F(8��2�t-h��bq�A�����{g���-����M�F�20��W.W����b�S�㢺��[�ƃ��Ud泼���Ш�;��Ч�I�vt�њ���#C�g�zTQ�[&޺'�q��*�F�-����`a!a���Gu�������]�V�,��s{<]��R�VHr+�EUF,�G;OD���q�!չ��F�QM���~�>�'
�ӫ+T��J�DK���MQ�N%��Un!j3������'��g�g[g=��^������y�+���YSR�ǲ���~L�CR�%���d87���=�zvܚ&�M���t���t���>�^ɛ���M"���y�T�{vY���ƫTO�Y!o+S��QknO�������YDN�1���Wi�.�s�����M�����`&长B/#���M���E�fF����c������=�:��
��-n��?v{a�y��\=^�������ׁ5y���!��O�%�C>�Wzcq����vl��W:asˊ���Q�%��9��|�
g���ӭ1(��+�t��p�T��7H#_�E,�z]�G�0��k�v�O�5�=ZM�~��?�~VUm�,0��oI��y/�s)����
��l�x7x��fsU��+���9"5-�\�rw�b}fI��L�NgS^�O��:��r�$;��H�?=�眻�qH���DJr I�GDm�NE��
�i\�S�uI������'��B�ܖ݌�gB��������좲��v�[=��89��7�F��RX��3�oI'<㉾jG���)YJ��G�hPNM/��������N�?�h�=���p�5$����2u��h �*v��rv����Z��T6��H�.���ȑ|��H���C��G��jZ���#��;\bBv���e��Y_ܤ�x2פ��R��ڔ2m5�o����^Ϲ��^x.+�Ո?���u}���>�t��n�V��㻛�ӎ!�?��S�mը�W��2o1tM[N1���Se�MME@P(4�m�@�!���{�=Lt����e�����ͺ<�]ۆ/��g��;��1{�cXBQ�HX�C��.�X~\�N����/(w�[�}m$����O]w�Pf�
�܎�B0M��ܚ�Rn˧x\��.��V��3�$ս��Օ֔�[�ۑ8EaATԋ-�4V\x:�9�-)��v�w~s=���0�D�N���\�2�*6us�AȬ�슘F)���'ꌚʗ#4tT�xz��F�e��6����k����9ڼbR?n�S�sh��e��	"���%��;p�
��Wq'�^�?����3F;�/����'Y�B���t
�D=vҝ�jdKБEts�KҸ��[�c�����l.��{���4~s�iV9H�<�K2	˶�ھI��Ʊ?�Z漅�.IL9�7"�Չ����K�͸o���QrԹ�Y9VǿN�m��c��K�w�1:�BË�����e��x�s9�m'	��vv!�%�:nao�tJE��UQ|;+B��⨵W�aR@�5I�L'�4��pը��|���t!�]��{"������v7�頩��;h5�mX�P�3^��h�!�a ��!,�/w~9	�_��[��yk��)a))��Z���Fz���+��e;�L�Jn����VD��������[����<�T�-�	>fO��{�0��iA���źU��	x��'5)Ր�'�?���LN�)Ƶ�۩k��q�G��u�Q��w ���3����q�5�y���/�ʌg�u��q�l3mi>���i��O�2�z)��c�ZzE��gZ��� 7Tn����k�M?�w��u�1:��"S�O*0lWlq�s�O~L���p���v�*}�/n�q��KʌںK�V�Jf&��y� �2��t+C�'���_��}�&�p,Ő��m��x�#QҤ��®�yC���7ywJ����SR���&����xz{$��k��s�Z�BV�n 4�'F�\{��)���,D�#:�Lgz>����⥫7�.o������-�c B��x������rv�~~�S</�x�G��/q�]B��������.�`���7$h��1�.-��t���0��ė�M�Ū&R��8������M&&
Չ�1��������J���y?��%$�53�:�[>ș��:]���/&l��_���9�)�|b��p��B3�f_9���$���.,ˢ"c���rK��n&A٭�������P�N��n���`��[+�7=����l��k�e:}W��2f|O�c��A���q/�"kCG�vo�'�������n�~�]uq�L�5%~�
1��i�^�W,T��w��m&�ם�4���&U0�Z�'�&G&/��e˻��l�����5�/�:�Je�n�Q\�}��c��$�����;e�5-	���`B7<����X��/p~��g%�h�Դ���⥽:����9�$�VBuAT��ne
�ܸ2w}9�y)w�4K��N����d���kj,DC5�\��@�Ɍ�Д�Df���eD��z�������z���[-e������N�	f�M��	�� ��+���^��~�Fٝ�x8O��v���ړ������.�99񛕥�2<�$qܹ�u�2=�+ғeCF=;�n�V��X�g�e���}��(~@>ե�jj���n
Cj�<5Q�q  +�C4j�#��۳m���Zpz%el/70�h\��� L6C٥VbNG�˻�3�ҿ`�@���N����I��T��?z���;_I�>Ҳ��,3Qlh��)��HO.⋏Rf���[e�#O�R{������� sݟغ�(A��9z�n�]4�1T@�oգ
y�mn�3,����)6��4����%x��v.����9���f\,�}����=J01\|x1>��"z���ӅZX`tl�<Y_��ˠ�[��4�����w����m !��[��}����̎���P�j�;l�䩜������]6�%�BAC�1�M�(\uW9ҿ�Y�MJ��4n{Z�0�������TX-�1	�d����O��8`]�=@�Ȗ�q[I�Pq=��1�N�#�,�L��F��g)$�$���4�h+�|��!�R8i(H�~��T��:5a�'�7����`�۝簦`j"��,�Z�c9ڦ����zK���D�Ћ�P	��G1x��u�%Q�Ul����%�r�X�@'і��A����z �H�MH����̄�C�Pz!%���k��ci�Y�^�nO ��-9�6������T������ �#�Ń��X Υ�+��p[kb���d���f8E�j
�h`.���{:�b�ʗ����[E�0�S��"
��oXW�2!7�c$��&1;�Dw���TkN2��FS�~���戾�9�d���	
�s��?��!����9�A��G��D-����<�|N�.U�K�T����4�3��	9_�#5�;	,~c�T�~1C�To襋���N���;�yϸ�j�3�v]��f�pP�m�Ѝe(�ͫn�uE�D_���!�~4.0/���(gn|q|��~����r�}Vhޥ��\Y�o��֣�)
�2�h����䘧���� $갺ye��`�qoƉP뼱��ݗ-JBM(Z$F�\)D�����f[P��D/����c��Δy��-�a�q��PXɂ����[�xW'�>u�U3�Ǽ�O{�7+N)'�v�W��Eϱfez�4����Q����J�E��e�L$k]�mA���Bu��C	�����A9]^�}�1�'W�:�y��Ho�?nS��~gٸ}� ���d5.x���q��Ni��'�����~Z�|�4k�8gB�/u����y�	؜S�sqY���Rŝ�3a��VhOѡ�����*�|+��Z��wOy�1v�E�;��=�d_��Y�w��x���>���Tq�'j@���Ѩ�>/�ѷ�1S�}�F&�>)��7O�1���a{~�W+�6*C�<����s~U���H�M4�w��"ݺ��b��aO�J���]ƶg�#`4��P��;���2D	��+�.�Ru�U�����P4���Lb���<8�D@�J<kx�&%	_�|�9��k�Y�&0>�j���l|�����4������T��� ǭ@a�x���^xڃ�Ɓs,]@}ڽ))�����C�F���s���$.i�cY0�~&L2\�-zE�}~�%��ԍ><��&�F,��mUxI4ү^��V��*���4�:]��y؊�(���=�.� �=B�W]�仂�S�����f���t��q��8���E<���_�ELh���F��HՐNv[˸D֯n/b1��E�V���7�G�u����DY33����G�0�-Ƞm̺����u'�뾼�/��ώ+>���'��P�W��6�8w��M8W}���Kw�:�_9���ewV�.ݹ^X���b,��{�<�6}^�O��ة�9���'i����L���6fK����4+��Pq�2�(�jO�i�q��^�R�XF��g�y��w����{H��ݛ���z���XR���Dg�5������ 'G�����L]G�eC'ΓAZ7�԰��j,޽,1�{0��r�O��;� ���E1�$���u�ם�
o #�L2��Ow/����"=�_�S��1�y��
\��iR98 �2��<�ܵ�.��?߆����G�>����t��Qq���P���b�ͼ��<��y/~H���?y�2/f�ta��1�����,�~vg�G��e�%Έ�L�����椆�m��v��ڸ��" ��^R��^Oef��̿⹗�¯P�S��Mj�p�V|�{�F�ƧF,\HӘ�H�R���$�몤�����Ǻn��7��䘡c�!����i~o���[c&ؓRq��'���W�A/.�v|�#��iޗ�(�����.(�y9���1Ǣ	�u�����]h��u�
8�#�z;���3��yà�=�~�!�����xj�����g��xp_ �[װ�,d��<Uiա��2��P�]��O,N��.~*/�*��8��
�9�]w8D���Ɇ�9��H��e�:���S$.(|L�C��;��\�K裸�5��ˋ�!�ynS]�(�+>�A�y�8�D���%���[�xin���%v��[�U�<"Rk��n�WR���х�<]�&v�l-z�y *#�u,cTDg�ϕ��&i4~���x+���%z�E�_����<�z���8�b~;W���Mȃ�J�x�5��WU�>2	�(=��_��ƍ���Mn�HA߅�vs<NJ���gE�J�׈Sh��x�{M�h���b���f������)tkrQ�5��;R'$����;U>���^���RxE1ᓭ	J�E+�;�5��>/;x�WW�����=r~ĳ^� '���ht������7SM�a�Pd���r.~]#Y�Y_�k�b)ٍ���I|�V�NHI>+�J����Ahx;�ƚ��NR����$�ןZ��>i(T�kX���¢��'6A��*0G+���Y����&��P��~SP�ɱY�����z���A�ya!'��ѯh�gQ��������]��o��[������DV��w#�+fK�/'���\�rL����x2�BҦ��z�i�Ȑ�IZW�hX�<�F��^��P%��N@,���B/t�+uW7yUv�>��x������J�Ue�(&H��gSu$c�-M�}&c'Y��6����X�T6G�D�o�P�;_�x}�fP2Eit��vU%�����ǧ� Va㙎��IS�Υt/ɾD�mt�Ö��H�u���</�0�h��Wɺ�Gt�'c�q <ʮ)�'�
�˙U�U�1��AzãF
�!�u%��n� ��8��(��Ew5�<;A8`2>�J�Č!���˴��>�T�:骩B's4�mz:��'\Wo�M�x?�����?����?��S0�"�O����ޙ��Nׄ����A����.�2�����,����*��/G�+�D�E��=��MIi%dt.Uǽ`��An`D�����y�|D ���*�M����S:��m�pV�)G��A�F�N&���PO�ˀ�I�c��Ԇ�9<����������RǦ���T6`�Xu��{s� ���h����S� ���}���˴/��Ic��L P�N-(�X���&owc�2����5�y�!��(��Ǎb�d��f��qT�ܽ���C�.��o۶�{.�&��j��ʻBw1���� ����SD�Z,���u�)��Qm��{�`d�b��J��V ͼE>At�j@t�^�����"�W���-�V��d���9,��aJ��6�m��"�I2#�7���44��P����8ĎhK x�	^��3�~g�ֆ<m�����(\�/9+�c�uj"'D����|.;�^c�vX΢6u(�~���􊽄:���� ��\�gG�5�l�}Z�ʧ� i��Vr$���Q8>+�xO��O�7��|�f�]�:�����&�]���h�4x���/������e|�#{t���4����^+#a ����b/��=�-��c����}nٚ'���y�,�ɐ
�����n@���h��/�iO�"g��S��Z�P��"CECt�<�:6��Jx\5�=��uOڷ�F^�Lzmh(j_cR&��O���0�Ԫ��c�{�D�hx����$|��i�k��u[Re�5�Te��3_��1���_¹Gy�(��.����H٨s���|6��zD��Bd��rO4`f9sz���k�=^��Y�����z�'�LLLR��b�b0����]?����x�6`��|"�_���O��U������K@1n\&�z��e�F^���Tk��-�6�^$��[�+�Ff-*��ϧ�y;b+�?
����Zd٤Il��\!P.��IVT���Oo^��˟�Y����6^��.�3a�}��e�		�Ŭ��2�䄻L2�-��t`�(S��A�˾�ls��ۖ����h�R�8Fu��wG��a���/�!�ΑQv����/���r�N�ă�iuhH�+:�-W>w�Ҟ�+��!��x�����	�f�CS���*ޙ\��btҧo�[����'�ߪ�Z�L兕bc�w�B�J���
���""-7EP'�4SJ�v�n%��fhis0A۶��;`�j9)�#���2`Ԙ7���3�n˞��.\�<?j���7DL��F�z�xF�[D�o�K�
�x�m���5J͢�:b��2�?Xw��c
�s�y���񢑙*������X/���*��q���J*��Y��Z�?Kך��I�N�EP�x�=+r�s���;1�:PyOLf���ϾZy��e��D��z�Ϊ�x>b�V�1�{ݐU�eC���咳��q�q�vy�A@>00V��_���-f܇,�b��j�qs������ղ�{�y�څ���?R(c��6�$:3e;_���܇K��>�Yr�_�Z<���(��n|L5I�p�#۩�݂$�����T�U���D�oqJk��aq��u�������ڈnQm�-���D��W3�9���e%�ڷ�>6֢�S%�7�c�Io�$���"U��Ƈ�2O��[��z�]E�#�b�[����aփ�N�4���Sat��j�eu�1���̈́�6V������Ī�u�[ #�8�����lA+Y 'W�ڔ��m)���d$}8�,�0�fi��q/3�d4�p@�������d�am(IQ|v�7BL0ݢW�)��H�]��U�������=��)��sݗn�q6�~���؋��i�&��5e�� ]Hw���J:=�"ZZ�*��X�p��@p�4aD�Ӻ*�aR�H�ÛZ�S������k���\�`:�$Mc�b��yh��;��f8���n�i֦�	��?���.a<T`�>nΧ�+�c,���d��� �R5"7_�]��jǧ�|Ø�l?"w� {=�g������{��&c�G{�=mLI�7��2��<&�e�>����p��k��<�ļE�
A�w���W�Ǚ��ޞ��c�/�T��19mV���h�B������ʓ7��
��3����CH�����W��=6s�$tM(�ޞ�[ ��i�J�Ҭ{,\`�	��>�7:�7S�\��E�q+�)�d|�t\Ǻ��`�V�
f7}��P�����k/ ���%>�;�KC�ۆ9����F�x=��v��;�{4Q�A�^B���;i���߸8nndrD�]:���θ���ǨZ������A�Ω��>� ���m�s��W���%c��<��Znî5Ŕ,fA��Cww�dl'��y�y�����\�g���YS�"�D������Jp�C:ǳe�Ӏr��0d�m�1U��|�*Q��慊q������?��(;���b��f��!��<WNޖ��s�|��;��c.%��q���~�c�F�L��O����&�vS�;= }�q��犇q�3\��Nߗ h��O��p����Y0��+N�4e�|��d��,s�Y,�>9��Gw�W�����m�G�q@��;iW4�[$�X�E��!�l�P2����΋���D������ز�Q�R��6�yoenNɾ�r;7�oܾK����d���	�ei���V�����߻tj���j�U�o�I���Tt1=O��??C�Q�X����_k�)eu��{�@;��o��A�_o:�;oj����YTsS��1��Y&2�״ 	����:��or�ݡ��Ԧ}���WU'J�I	p������n�Q��R��0�#���vQ'	��.�LZ���g<A���&c�Hlꕏ`�b�ܶ5�f��+�9N��*)�c*}g"j�7������=�k��?�b�l��5%]s��|�5��5*�(��0�<�]��(�%����n5F+o�V��\j�)�3�����_�Sg[����r��>�Y
A�݇)Ϳ"�[TP��.R�EEY����.��u�.�;כYŞm�� ח�*�w��E�P�Jy׋�w�����G�i�>9�3N�Β�e\�|������7�p�;J�k�K���*QA����Oj������ݢ+S���[o���QԂP����h�yܴ9f�NRr�j:[jT0�@0���4��$p�77ǆ+�I��`^�4�l�����ti�k�5��'�7qw� � ����=C�꺯M������5�>Z�m�J��z���B%lA��p��iM}��c�c�Ty*�IQ�s�1+u�
n�v �Z�&#��?s^�w
v�w�Wj6��$�x "�-�.�x��S�m$|�f���\�����r.X�FӦ-�	D��?;���Rq�!�8� 
��/3e���\/i�u�OZdxV�b:����,)�ȫ�	�1!2����n��eԎ�n��bJ$�{��᫋��^:m�}r�4l-�ׯ<~w8+&R4�	m@�R��{D,k����z���ۣgи���x���}
�2��#X���'�0y$)��!���6D��,����;�׭��:UA���Gͱ򥸽H�,6=��w'�iA��F(V�k/w�~�A��G�������<P�5ȁy���Xꬿ��m���Z���}G�F(~7m�<6>
����rڸP+�兠9�e���o�;�Jc�#im|�]f{s�L`!7�o�hNN�{����/�����lHTAGb���$ݖ�EW�LM+.Up����5_����R��Ԑ����Ce*�e�1D�3xX{��<���G��N��U�贏q9]g_��CVh������IՖ��fƷy����/s�;x.�< {W����Lg�Gℕ�<j�����tDۤe�ξ翐��g�����<Wq���\"q��0t_ャA�����&NM*�T��1�K��9c��R�l��k��?'#j���w�?.1�x��|���zjd8}������539Z����������=Ho�3��H ��r�3Q��6|���i�!�L9h1�2��X-33}w4[阣�5hA��`�,{H�b��k�=�<�����O�"f�N�{nX��F�B���tYRoN}2��쁨�[�1�ky`�g�Z֡'LFF����=&�U������؏�����J�)�&E��it�	��C7�.Hj�1�1S�>Q(r��'l4|0�^3Y�����S��\�C5XD������d������������.'R ��i'ө�D\T���\w0��I�*s|	�PO��x](�c{U��.%G�f��L�ќ�_~G���7^������;x:�<���֊�г���Mm�D�&1�� 1�7����	���X���3,����(���&�
(�t�=�p�Qs0fE
��Cq]�ƣ��UO�K�*,6l�⏜���%ϗ9e�k>�����G�UsV����5�D�ȍ�L�w����T� [拾��v�zs��v2��o����zo'�W�W��?;����{^��Ž��#� F:s���F)kQ|�����-�*Wa����� ���z��Wr�67�QW�S�j ���rg�*FhO�*�� �EM���>J�8(�agub���&��4�/��dF�=�=\1�t��,�48��U�-?X\��F2���������{,b@\��.+ �ChM�Q�/����4�+��3#�˔t0��S�g�a��-]*�Ŀ����p�_��5��(����Kqww+�������/n����Hq�������\ə�ə9��u�4j��׉���0�ko|ƌ��n�Ϭ�l$|�r%�dJ$�^,M-�!G�x�。� )��q�g�Z&Z͌_�$C.6�Z���uf�qP���38���g}�]���y���_e&:t+6��v{��u��n�����32�O]J��D�\����愈���"�w4�u�W!��b�c� 0k��L*07��K�qfB��J�X�beC�8R6���͠��p��ѧ��1jꓓ�0tV=��=U�v'�V	e9Q�LN�%�4�o_���q�]�֫GS��l��a�|b;�W�6��k[7�1ޮ�jx�y>�}�K�u�Ӻ�f�k�Jc)7�7ǹ-t�+��)�pݟ���Ǿ���̢�B_�2�h���Opk
"b_����Ѱ���gN����iO{Z�U�(�$�mzmk��*�Ik��h}����Ժh�m��5��^� ,=ؾ#�c�?�ɲ:��A�1-Uȏ��{��	�˟ȌH?���(��{�����0	��De��LVZw�����l�1t���7���:R��d��������<33/�5}��6�g۞���-��ϾH�}%jR���s����@Ch�L�g�g�T�$*�>m=~���1���3!�Q�V��0�N��˨5��Ĭ0���$4���Z9S�puu�Z+/���譃x���S=�Z"��O�n�G�yi���[}C\2�B߉�%�na����観SNsy~;%|���`��jhw/��#�\"�}��(��2��\���;#�}v�N�#x �v�E����Ah�-��C�g����/�ل�u��Dh�m�l)�y;�]tD@7:Y�U�yDU�W���E�.sT4/�~5$������e�[Q�?�ո�Б/�j�>�o������K� ]\�4��ݦ�o0�d[B�����M����Ƈ=L�a�(�̲� ?d����W@��s8)җT4(�K/-��_z!�A8�%>aq�/?[�X%�%�%26#��ʷ��MC��{���7�g��*��H���:վ6s�L�X��ߙ�_S��o��5��=:�ρ�I��޽�F�P������s��'Fh�ґ��{�����P=��{�W)zNE^�4�\�����S��LVq���{��ws|s�cg�#>�v4B�FN*��ۨ�����)�B݇�6���ϟ�ʆu��@���o��re�;�H���4y+GP��<�VcE�*M��ɴ��u���ײ9q/Ē[�i�܀첤�O-�
KP��z��	3�4��p;�d�n~���҈��*:󾊟x�2U.e/�D�n���N���T�!�(t<��Ͻ�V�qЅt�]�m��Fq4� ���ζ��s���;��DxN�Q�k��.�}1�؎��
'	�I�5�a���:!�;8>�>�i��j�:/��m���s?�R��+Ub.�^���+}�&ۨ�� �X��,r7���^X?ꔼ2|A�r�A��,&��&o&Zߨ�I@ٿ-)m8����h�5��I���[ݘ�Ⱥ��R� _�Lv��ۖ-t������U��a��j�Q��DT�5eL۹c�A�
jb�h����zͅ�6;[�w�).s��y�2���ߏ���1��j{�����Q\���nk�q�!�.wo�g+��d���Q��e]*L�߆�n��D�/ʣ�a���D��$�#u�g�� �j��
�XiG@P����uv�⡥3��+HN�<e�m�IYo���G8�w�px�7-����jWG�eV�*��)_]+s}^CZ�P�N�OQ�U��fl^���7	���b�|��'�[�2�HE�W�g�.DSc���%��lj,XQ	��{���!/�i~VI��y}$­G���8��?��;(�El�A�ýO���p!ܔ~sD~IƄ]WC^�H�a�Inـ��+18��+�~�eR���k�7��\DD�T2N�f�?���YV���&V�� �����nJ�|#�1�������4����F��{�~���L��o��5��5�Ǽ,�����t�ɕ[[�{�-'B�u�a�b�Թ/��45k�C�hCtya�L}Y�5ʘQ&�=�nf���B��o�%*N��߯�����S�ީ_��V�e� ���Qi�5V�[���)SF����y�����S�l���fk4nܞ}� ����BVO��\�����yC6� ����_�Z	������B��}��L��;�\��#$V�e����j'|܎�w�{�[���5��I4n�kD��2�Gi�൯lG#'��恫��k�H)"�B���:Cz�脔y��؞�%�4��w����r�����*vkf����i���ϧ�c�Gh�
�Ӏ㺝^kQ2��L,ۋ��
��v��o���&'�/HPDǌ�s�I���g��Qh"YV|3]����2�ݸ;�����@��MO�L��M��9���7	M-[9�����r��P���W��[Zkʘ�K�G�+���Mlo�AhN|�����_��ś�_���l��i��a�)Mhs8��~�/@J�X���;vv�5될�0y����16A9*��m�����ʌ�B�![��'�І��S?Ⱦ�߳�����{5������^]�@h�WE�c"9D�W%���ۜ�d�6��Ʌnʉj�"���Jږ�YDD�x_=���73��&# �=0O�?�ԁq3̯��]�|��.ｂ���^�t0|(B��b>7��2�<���������4ݚ����F��L%��q<|�i_貓���k�C2寄��AQ��U��>�����T{��nRu�Ž��v���3u�������n>Dw�b�C?�Tb���<�~�^L~�e%�?Vi}��?���^�;�\Y˅J^���f@�˙.�Ȝ#����+.���R#֕�6�0��f�(Xo��QB[m!�ED���v�-��m{SBU�!��0|�7�hKG) ���zWx��*'��ju1�;@<I�8�=�)��WD+I�X;��uv�dJ�c?y��XN1pWL�+��ҩ�1�F�"\3��*r5���m��{y���n�'��cպ�2��ĥ=��٩�Ƨw���A�
��׈�;H��F݈�Z�E ���!�I.�Y�V�(;Py�>sQv1s�󔰉��W����t�#��s*����������'����N>��*'����� �ʙ����t�x	��)`�ԯś�^�_;��ͬ��u�a>�}a!%ω��2S�kQ��~�d���ͱ$XwDkt�I�Q
�<r٥A62NIF�+��U㨘�N4��Z�	��˻}�` +�r�4$�d�Y�s��6'�\S�hq�p�4��$r5���X,�|n~������x��m��7x�J��ݺ�}H�ω��o۰Y��RZy4�!���������|��^sJ�x�6�eoQj���:�i�ҥ4��~�����B2̺����)�\b]ky����Ճ���T������aV}PAT)�7�R	I�<e5�4
1�,����v.�9�!O��'��ktIU0c��^�S����&���ӕ"���Ը��hi�ҙ���
G�_J��`�f=R�s.I�E�}���g����=�)��泣2'�7㯬R�c��Y�I_�◷������z�"ȸ$�#�&+�lݾ���2�h���E\�^��z5��w�@5�̟�zd?�Ez���FމnU(�z|/�0z'D��������p�	�tڒ��24�ľu]R��U�s�9輯���a��@~�>vZ�O/��&ߞ�����-uǅ:�����#��'�z*���f�:�3�w���������Ղ�^��a���W���6�Q/���fg���	�2��T��%策�ǔ �����\ c*4��d#ݾ ���F3�(_�")��V9�Ձ=�g�u���Z�k�? �N�i�ZD]i���sǰ�p���J��%	�E(��p�������b%�%�H�\xΊYIOh_n��`ͷ�L��i�ުLyX;2p{�k�zJ��˜�
���n���
�1���{WH.6�D�"�+U��W���t5��/ �!*�bup�>�8�]�7v�m�z2�H�v�iG1/��RfZ�xk���qO�)��b��p������������7巓I�%�m�M�*:̂���{�=�g��[���zT;�,H��Ƽ@��!��O��y2廗�N�ϵ��o������h)�CE� �5/�`u��q=���N?���s��`�~C�iB�%�'V}����S��?��9]g�GdwϿ��,ğ���(�)sj�&�d�����~/7ѓΚTl=j�(�V�D�ci�[J��Ziq�����oA� 8	b�mLI�>Y^��<hQ貯!�T�w���5�R�鵧�-2a��A�rI�ƹ����9�qr��O�ace�����_�(b�#ӹh���*�|h�=ֹ���˾@�� q�x~��t�2$IԔ�X�c�蛑� 9�r��������(��JxrԉS���P�]�D��5���[$8# �|	Z_HN���D$��l��z�M���`�����&�Vvzc��s��=&G��,�p�(w^�����jtz��@�Uz�f�A�}"=����,Q�y��!���`x?C��&�3��j�@���*��kC��Y�^�%sT�R�\u����2#����,�r�2�"�p���l����'���� ����X?:C�"�'�F�e(v���I��&э�d����!�&W���]�����")�?�����3�����r<���C��);Ga ��o�_]��>��vN�J=;�C��%��?O�%��݌���هRW1��"_f��2%�@�8vQ0~@�8�jۈ+df]��8�)��5�X>-�v�q�g���_��٣��� Օ}���C��;Ѿ���l�|u.J�����o���Ο˺�'�1ۍ^���M6l�	T�'�bm�g�Ag���V4z���Q�zŜ쥻���8ͼڳ���$��awSQ�)�0]̘�`�z�Jh�݊�/�b��m"��x�>���P��>U�� �o��B��>�y{Q�>0 �zYҰo��G�W�����,>�D�"v7��,U�\f��"��}��\��q��հ��]X�3�4�hh�����jq��]�|�tDHKrpd�G4�A��J��|#��	e�Nl�P@�z�$�+V�c�(_6Ndu��w��":v����Q@Qr����zz'Z��y�����g;�yOl�-2�KB�M��e��e�D���,���_��
t�k���8V��Q����^����c�گ���J#�%O)w�G��SmC�(]/Yf�65xF�����n��I��7[W����w=��g2�!D+;s�}��tKݸ|	����(�o��xqa��{ġR�6�_ N&0{WY�q�@ؼmɠ՛���8����qex���J'��0MϘ��'������rqYg��䴎Չn��4^';�����>�w�����w�1ӫ)�0iU�bDZՌ�#���i[LT���n4{X�˭r��YМiE���|�èYkͱ��b�����f��F��ZW����@�D���[d��xX���������)�q
�(�k����םR�Z�b�{�wx��N~o�n����'YwK3iq�
��獒�͑�5J��H�α}b"�!�beʼب��g��!�ބZ�~�Z�o�@���_�~ow�1�!�N�\��u%���*�xy&3�l�r3΢S�i��+����H��v�iU���oї�ڿx;�K��*F�l��0O��
^b�C��p�b�=�S;�[�nT'�G�_��r"".ŷ��ᢴy(�a���=Ą����sT��QP�/�ܞ����u��Yx�J�ɼ����?\�	~���F��ƭ��ϔ4��d;"�ހn����$8��)��ö.���.~9�7�\W��w�ۀE�ʂ�s����e�"2s�������Px!�)	��:FO��C[v����8���)�C�h3��g�H�J�%4i��`�܄�-�s*�j���=��_r��6՝m��D���z��\9ks2�e�6H���42i�"i�L�p��-��jF�u^�e
l͌�E���U��z5���m@�+M��eM�������>���ݖ����viC>�����U|	���'}���_f���_!{Ŷ���3dބ۹�>!O%�?�9G� �H�ɯ0���Y��ť1[-��M�����Y���X����2�<�{g�k})āG9�ل�=i�d��������i�V�ߔ�܁�i�;n^�];�0�OyJ���R����_�|�..`����v0eV�Ѻ����ێb;�l�,�%�{�k��Lպ*�U�qn�"<$�o�Χ�!���r�o����L3m�>�n�u���{�V��*�6��O��5wO�by�~s|@)�����r����d6-��ъvө�8�J�xn�u��6m#�4�Y�P��(9�O��w���E�m`Vڀ� �$�(!Jl�Z����?3���t���� 	
�>�"��[��(D��g7[^ID_��w�/��V��zw����1V[��5G/qb����=�T�0aQ�FV00Ci��""�[�g,���ہ�y��ʗ��Q��� #�
e/u �ڐ������@�Ѣ�W(���E܌���nٻJ��.7��@�܋�}+ۣ>M�se�s�-m��IN\�D��`��+a˘��/���,�FJ$�A�HZ��/��Y �����A~���+tf~l���N�R��I�����y�o�q/�:���OsZ����Iw��پh��\��ɲʅ��!��֐W�N7��WN�O?�w󥞿�؍�+�/�s��)�*�Ӱ?Np�L��&��Hk�_E�V��1��PF�C�0ܳjD1��a�p�;��)3�+�I|���;'3����X��-�ȱ��]ٜ���~�8�pM��z�V�'�;��z�]���[����H��w�Q�B)+�i?���䓳��������ǖ�� �B�^�o�9��rr?0�9�<a?�ud������4�y���p�m}Ny�o<��б��N��&'{U�1:Tf׶�hѮQ�
��iH�w�AQ����=��KP�2�i-8�>�	v
J0���_n�߉�	V�o.���֞6~�o�'�H�xWȽ�Ս^0��ӏ��_��*'�3�lZ��9'�����?�B��c�6b�<��ǹ:�@�ח!�+2���.�[@,%�-U�Z�1;y���M�f=ǿa��S$�yPx�q���_�����M���(��Vd���4�ڵ:���r}qT%=/�d���.�耷�����t/._<�=?��G�Z~R��L�8��\��#�y'
�MF��o/j�<��N5����/����s�8D�-gR��e�ק����(Qo���Ft	@� R� ��3��vلB��#�gů�.��w}�&�6�O2E�
��@��v�e߀\� ���׵�"�ː�az Ĵ`?2!9�@o�)�~[�F��S��ډb�7pL���.$��}��ӫX�!Vp-���C$�&���-��8�)a]ͩ��w�e��|�M`� �Bq`Q������D#�����R��*����"ś#���\�y��7�������;#��diҼ*x���a�i����
�z�'�+��c�̡�'�-�.뛱�X�E=�4�gW�#'�"��xZ��q��?AK���1���"hWJ�bi�Ǐ��s�Zu��ٱ~׃y�g����;q_�Ka���2@:�����
[�i#	�^��p+�m��bT6B�G@����>�E��.�ͯ2���W^�T[�[M��_m���|A�����'7������~�px���7����⋊/�LSj�Ek��b"�ʥԿqq����^�>s��f�LC��U"t*��v�r��B���l	�[b��<չE�J��eA��z�?=��޿p��*k�Co<�?����ƺ����n�E��ff�:Y�:}O~�:"��xK4�ͽg�����y��	�!ځ�ݴ}6hw�¬ �/^FO�}7��lk��I��mjxy�ç> 3WW"�E�[/ɦP[��$ ���mu�ô_j�*a;�����y�7 vj38��+�Ӌe�;�RJ_4t����;���a^B�n�5�d���Ei�Y)y�W����bz{���)�鱮O����Q��F�'�6��G9't��IW�����%em����p��X��8+{���{�e�HA�gɰ=Z�@ѳ{!eǲS��8L��B(aBъ ���V���H{;c)a��BdRA�z̺�	�x��Ǡq�1N��o���g�l���(��7�S?�$���r^�<'����pI��j��m�,oPQ���y�ۗ"E���{
Lx�Ls��8���2��p�>���������Z���/��.�K����섗��.DY��>��͋-[�Y܌��OHrb|������ L�I�o�t���d�ߘŝ�pr���_M#�Lkv��C��hs� �]�G�O�L�&�hr��=�B1&����}?����P�_-�1E�OExPz�Ł��a)n�;M��賶���N5�?⳺T<惷�e�"�[�6�N8s�����o��$�H|<̢�?���g��*�N�ȿk�L
�i�B���xQ��jAe�zd�8��Ze�{�ո+lϱ~ ���<�Wf�S��]᧵\�b䅊��wJx�Tzͷ���J)F�"9"�gM9ʼG
�W+s�VL9�+R�<鏒٤P��,R������������2%{� �[�����r�'��}A�ɽX���gbVx�%u����NW�tA������ng؎f��9g�ntL�a{�����f�H�K^m$���0��G�^*w�S$�V���Y͒�w�%Ő�Ӏ�!>����v�B@t�Ԩ	/`�J��a%5���$�7�ˢm�KP�gw���ĞּO  #�A#�νHM��W�Q��3�@l��y���v�;+���թA	iRQ�����b)�#�0�n���/U�km�_��{�s�6�( -A��=��%J�J/��7*f��_j 'p��㯗tX@�䪼A�P�F�o�/��Dh�Qb���H/�wfݠ끮M�M��V˳���G�J	���hv�u�%���H�&:*�±���E���lxb^(�?<͉�x�:�:Lݞ,FT�*0����z�S�t�q���r�@4ӽ�t��ƒ�_���,8����1~�[ZՅ��k���6�u�r���Y��@'��c!g�cD��V�����.Z�#������ac-��w���$�Y�l"�� Ah������H�����f�W���w`v�-X]9J�/R��>����0��T���5�4ͧ�rTq聃�i�_��C��[C}���y�>��5~�&����C�{�'E��՝:+�=�pu�TӇ�!j6����P���[`)^��{}m�%����v<KAS��Q<8N����2j>����E�e�6jd�^NF���)����J��P�ɇr�وbr`x��3�EA�S�H��4��/����NU�-P��8gU�ok5F1����E:��ۣ��1אW��Y��V&g���8��:���;Է��B���{.Bڜ9���K3�s����b������mJ�V�̤��~#���w*�C'F>'��[t=u��c���B0�b�QZ9H��(�}n�~,��AFK�$'�7 +T���t?4`�V~oy7ܐ���&Y%[���Α��L���״K	ψX��A�ߙ_V"{L��мu��h����3�^������;Xy8���!�����P5c�79�L���J�����&�����Mc��Y������K��e�;Pi���G���(,S�_��v"wj�x=��}�*�>H���\G���
I�/�3�!A,4 �$u�>��*9�/�sE7�H┞�KO�n"w����uA���	~ZP�9�``0 �o�\�~&;��;�[��\��K�۪P����`�[6�G���c�aΙ�j��ت�P�}�]|�h�*oi�j�����Hk[6U~ŭRr�/�o��
S����Q@�lluz�$�r�ߞM�:��WԼ&�b͆�f�Q·{���B�f��vs�y������^�0��� � n���d���P�9��p͹t��|��S�f"�����j��Rԫ�
��>�����v�O�D�U
����r��F2���0'm�XHQ�@�|km�O{՜���e-�HӇu
_��71*��)���a�����}�2���e6Ԣ�س�9�s�;=1,��n�>VG�˦xy	8���8%�7k��T.?��b���Cdw���,���uq1�l����&H��Ά�g�P#� Qth!u��5 ����Ac����T�x��0�KX�����Д`q�`�$,�vɺ�٩\�1� ���Dѿ��"�R@��;1'̯�����Ke"������1l��>=$5��bT�i�Q�C-�.P��i��6�����2_��< $����o�\�uj�7��v�q۝������o}�j�g6��\!珅�3z/�xH~���V��!��0ҫiZjt��o��UM�P��f?j*Vl�`���qj_E��f�L#��6���RH.Ad��_�
{;��,�ӆ�� �x�Z��U�Y�n�Ƈ�@����w���_<AfI��4ƭ��ύ���8���׵ӥ`�	#����r���Rر'W��
#>a�;�4�S��r̋3&�UG����8{Z���_��xӝ����q1��O�K
x�<���c�L��!��N �O��N�I2��S �{�ة�!FȎ����9lWI��S�m���܌E�W�Z��F���*��R�͆��B�� ��U�X�x�{@[�\�Oو�S��N%� ��B)k�kG��Ie�e�?�g� +�.d�9e���3�hu�Q/W(�ݠ����S�f��+��x<t=�T��I��8~j��|�I6��|��Ɔ�0�-I���2O)�ߺ���ۮ��]7Kg�v�#EN� a_�?��4�Plh�Ũ���ߦ	ӓT'�ҧE_'ɹ�<������_*.e�DW��쐮aZ:zyy�ɐ�P?v��2Ԙ�P6Y���a�y-�6�<	�k~�����NShR�L��K�D��>P�����Sk7X�������j[2��wx�w-���p�ډj����0߾Kl���F�Ӟ��,�j�;e8�}ڽ�4�; �&��V���̓���{=�箔���L��yM�S%���^�%c��]����̮%���ȷ�=N��k�t������y�{����nr���>=5��[�����n�{��z��c�w���*�W{�O�����2�Ĺ���������<2�n��6,_�C�f,������툁�U� �-L�@� =σ���`�뭷��C��к8��ķ2�����WD��%1#=��׵���������T)	R
��P'�?����l޹C������t�<헚�/b|	�������i�lI��>��x�6HB��EG_c,Y�>׿��M���$�.�>�����Qf��IΓ�,֛��1�
I� ��YU�jC� z.�O�m�	�0�Aܺ�<��Ed�ź���� �u��}l_�c?Ѝل����jD�v�-�(�E������c'��Hº��RlP���_�X�4��O�*�;�.j#~㔝u­`���ۤ`*�myc�P�����}kҎ���~r�v���+�S�
���k�hq�s���;jY�r�x������2q�/;�ה����y�^BPks3�?v{�M5˺%����F�=^��8�"i��ғ�0�y��˓8f,�{�گ�����R#���-V#��W�ouu�Z��`� �W3�����K�exq�"���q#�,zZm	�j�����ώx�p��rr�%Dἵ���Mt��p�~1a#�V��0�X{�����3�G���ˡ�����9W=���IO��;=s�p����~���L��8�SAC�^}2��@�+d�bf�'��Q����>�6�V��Iy�V�=���<�����-� W�9�ԯ�}�,C�Rp)s�I)�<�v���vS�/sF94�/����4i
�<��S{�!^{dy�`ޅ�܂$��i���(1��wq���ܿ��4J�^��ZN*'
�$�f���_kʅ"{R2���$���p�5To�SY�=�w®��q:*UN^��bbH�k�߳��y�p\�CqP����U�@w֎CP&-K/���L���A�PY�N�<a%�X�j@3��`>��k�"`>���E��y��룘�}��wX�����0m)=kX�"E��.���\�]�B�@�h69lI�05�̹g�����ڔ ��U[HK��,E%��"��ЕQh�:)�NS���,6j_�șp�↣��TRW (�)ݐ4u���l�m�sd a V1��6�.�*L����f��u�rC�i����s.�g�Zn���r���)@Ƣ�D����)cz�`�wZU�k�D���v�%`�"��_�:F ~65����_Aޓ�΍���ݹ����:5�/�)����N���jƆ�.�8񿠐][]=�j��f�&��n�q�n���.�	�9zHû��h�<t�k5w�x߲>уҞ����_��*�{��y�j��u��&>�2�&��Y�o���u�:�[� =\�Sʲ�U �։|��2p��O뽴���A}��	b�<Q���bF����d �H��?2�]��pi����n�p��.����qXpY(��%1x�kO��}��>�(�0���qƦ�?�w>خ�����zn�ao���Ly�����!�q�I.y	�S�!T�d���C�yپ�y"/�|=bu���.�X^_r�<���=Ca�'Q����M�e��6�e(x�&����d-���z=`dx�	����Pj�8�o�o����{��s����%KY����+�-��	0�3���׃=vj8���$�Y� 8/��A���s��^j�"��ӽ�X@����c�^g���A�c��{"e&�*O�M�����CA�D ��S$\�(�*���L��9 ֫.���- ��tK����x�e�>!.�8��z�>����_��V�������He+S��Z���3�d~S|ij���K�����I�o�@���ј�h�y��k%��z�����l�iC�/��G�$��À�p�k�X�;#&���5p��b��ۂ���y4lln&��>��y|J���W�z�������8<���j֍���c�lF��,Y������A� �`Q�A?lk�:�He��23��U>t��?rt|>Uy��tXg�
/EAR�H@������О���<N�+xq��w�A��)_��O����_��H��s6Ü���̹�x��)Z�"1ϣ�
|�IW_�
�Ȫ
�w\G�i���k���0��a�q�p�|�B�PG�����a��?'�c��P�/o�1%v���f��d=��.���z>��1��Z-6��"O_S�0g�Z�N]�&��t��v�}�h�/���|e��	��W��B�E�%�8-�ab���//&]�4�~2O��U&h��l����_:G���1y����� 8¿p~�����c��w��kK9XW�p
"�\'��<�
_��v���2թ�c���I!x����:��Ԏ.+;�
G=:��evx�d2c%�j<,@u�5�C �ˏf��t���S�"�K��$��:�q����fs���98)���d�F�ȩ�E�i%�[}@����#u�q+g��/�?�V5�r�D�����V�)�9�X;�����(��B��Fu���)ul�d�������L����.;�5ʉe�혊��l���q!T����[�V8թ�W���iqQ�B���ϥ�a24���`w@[�Qv�rF�v3�O����B�yͺ�B��%�酝�ݧS�2���,��H@"�F�G�'b[����S���E\�}�@edߩ�io���n���:34���Q��?�������&��)�k酞�Y7��G���)�/�+�z?�1��ek��R�m�լ	s��2��r֬\���V��e���m�F�Yn#-ki����f?����}��8P$���2>b#�hX�D�4��{|d3)�~����9�1
&��G�$,�O9���~9�P�cU5�͖���g)�����։�f|I6
���V�t�,X ��{�����x~����ٗ��P��*/���CZ/���:��_��%A._�'J�k�c�r�-['�aY���b�c{q���>�q�Z��Q}q�m[�3*�b�+ڮ�UvH¾v��u$x���6����C�v$4��Vv��L�L'��oY�����np~�Z��r;������ێ*&c�|�_�ML�e�G�K�yϮH�W��~D���gn�jفŚw����r�p���%�buO���/�=m @l����P��(�V��	Ud��*���/�Zn��}�޽G��p��H} ���s�ֆE^��sYr��ſ�.�B�HWM�����@� ����v����F�@��l`ζ�����m�3`�v������U��9dѩ���������Pq��a�L]CUg!��t$�U̓s
�������E;У��<�D�]R�s�M�_��M�sB!y���������o���baM�*����o �;�[|qC�Ӟ�u
���/�z�az��<B��,Q�P���&g�UL���r	�R�[Ϫ�|�f����G�8�����P����1�L?��I3��"�buEO���L�y]���j3��NNO����R�m��0?v?Q���p
��q/�����-���2%U��(�_�X��F�/����8���?N�ǈ�tj����]ov��n!4ͽ��w���#]�t����1O>7�6Rh������ϭ��fIA�ދO�z[%*��M/6 k�Gt�i[�<y�_���v	@S�8�ы0U���Hh|����9����h�NBGފ�-�vq0|��K��S�}a�!���E��'�ܦ�dVL5z�u� 11��	3��2��J!�evUZ�]�A*���+9�x�u�c7�Pđ�d������^à��Ӈ���Z�r�j�H�D=9�h������3m�����s�貢J�
��B�E�DW=��<�O�s}ϦӞ`ECT}P$�W��@�e���'!@	����d�&7&��-��DX)fG�0�0�|֩��K;�6[V��\�y�?;�#��)�uq�qP�7EC������
����z~�B]�y�_�u����h1
���g[�(�����
��l>Yl��>�3��46�j~3#��g��/��"�����P�6~K9q0?�
GBYY��[{JH���|XZ�kd���a� Z�;Nk4�)�����9p��߬9:)�ȯa#��e[jXV��+;�5PG|�F�ls��sc^��� �S'4eӈT���� =Ŋm�l��L%�U�1��N/�MB3��Fa�N�u���GBPF�K2D�����(=�3�ށ�2_e�T���`�h
?�҆\>(_sm�f$����[�7�(>{�"����^���I��y�9o���<�ʛ�끗�Bl�-D0	e�C��ビ�6�� ��X�{k�J&�qX��5:J��k<Lt�~�m�V��.�G��fR�uB�5�hX�)u�7�	�����o��T�D?vo�9�qq2�=�@�;��z4<4�h��C�=�|����qo��|SRB�V�#�a@P��u2������G̛?���רJ+�.�5b\��ߦl��i��;�Q\pŖJo������5Mܳ:[�]���R5?.Ę=yL{{�M��V� ݀ڌ��K}����j�����&��u��kp���_�9�YΙ�p5�8���6x���T0X�y@<x���P��Oqi۝�$�H��hkRc��@,�y��bl��`�}�U;4_;�'9kw/Hs{�{�%.�A�lC���|2]���h���@@:復�f�S������_��O�챴���]yY��фh����P�C6.�Sh�y�I�%�'� � s�P#؅��Җm��N��ޙ�B��Ʋw�;moۻ��S�)�z��l��`�솆���:�0w�����R�5E9�\z���8Y��e�$vt���-��, �L�R^4N�@&��s �/*h�n���*�_���[���lR%f��,��$$�Y��z��E��?�c룼n�u,��!���ָ!1��^��,x��S���G�U0D�5]QJ@z���n�S:P�T��%�k��fai�%����|����gΜ33�	�]��ס*#�\�	jé��NF�_���L4bدOQ� mm�'�����"��u��/�^�<`����j��D9�����0�H�_:������Ϻ��*��t��"?2�e��q��7�:^�W������'d�k��;-MON_C���ŒN�����s��8��zhq��+�m��K$�|��/M~{��"� �+I>aX���!�(G
�i���ؤ8�[G�wB���I7��e���Ժ+h07�z��@`�(]��(�kD���HEU.l�b
?��Z	�]�X�*_kS�m�tg����]�q��<�6��J����j��&'e����睺�|�߻�^3�^���+����U0X����۟������{���6%���Ϗ�S7���R��Ca?}�J�޻������_��%���NN��~C61����)/�=7���,\��&i�����P�"�uӒ����==�����ĆXBz_�w�(3X��=O�FNΰg�:��׏v?ˑ�V���֓���=��v�;��:8}�_��De���Z��VQ��t�e�E��GZ������wT���o=ДN�d!5�Ƀ�{z\$�[��x�$�7��<��,�}F�Ki-vǛ׻�7����@0ߞe�opc��+1��o�mqԃx���˟�}����W�n7G7����ؔ@Dz�a��E(�� �� ��6D�@�ۃ����$b�0sRl8	[�#^�R?�������|�N��Eۆ^���s�å(�MM͋�L� _ڃ�V6Hg�r�u����Wy���}*�����嚭��.!�r��*��s�GpF�'/��NL�~��ǋ�L�u�j��f�B�`�&�����нL|����_ɥ�uw���B�fz���y�YK�PN���l�ٜ�t>^��5���W�������ؑ�i�ʩuퟔ.�H���k�{%5P_T"���Q�V��4|��cn*�Pm�rW����<0�	g���&]�H?ҽ��K ���9�U{�u�}ƍ��������g�������bA��%w���&Vm��"ԏ"���6��K��m�.m����W�����������qm<f���r0o>��߮����@7�?T�l��W��b��������B*A��Y։A��K1�'T2/OϿ&KKzN�׽��]3<AAQh.5^�_���k!�x���]I܁�X�0�4��"�*"�@j�F�Co7��%���9�(��,
V��TSW�|��;�T�/R��.eO����'(����]��8=�s��Np�Z__�#�yY?�片�fB��D��W���\�"37']ݷh?l M��Ҋ+k�9	����&Tl�B��� 
�X��tζI��i��ڻn�|M�֯5�O��=s�|����s�mQ�q�f|J>7�����3�L#����A���=����au��D�ACk���P(%Ш���U{t��nT�H�O��-�^��L�82R�_��Yu���h���S���v�="ٜ��XѰm0�?�R������s	��H��JʚV0��!�)Z� ��U�������Kpysg.s}�� ��Rw��$=$�l!�oD�(�k��}��d�>��> ��|{�D�?�W�Fv�����[R�[zx�m0��1u6nk�' ��CgU�e�C.F�Z(#֒��VK+qy��٬&�Rb^7s;��E�<[�4�v��Y��-�x]�Dr��f0I�˯�|�Ԕ����3w]F�����oY�OMn���Ԥ�#c������3�w�Ď2���R>@�D	!��er���M��4@���=�Q�$8^���F=��֐����z��j׊H�x��t�!9�uH �CD�Pefd��Qa��Ȣjg�x#�1�?7�%\�e�f���Wܫo1�tj�F��D$�ut�I��_�lyu���
��E\�DI�%a�f�
�X�,
�v}H�OІȵ��3�v�~�zg?1�&a�2����kO�$қk���Ҿ�Y��pª���h��T��a�A������5�goV�hiR=Q���E��w��������[�����sҾ9�c�t��Z�{<���X[!.²���F�'��YB
A��ذup> �?��2�N��1��s��)����ų����m
c�Y��&��%�f�3f�L��2 �� ��z¥�&V��ZV
�9���0	*��Zc&��kگ�Gi���T�-7� �t �N�s4��(-R��r�5���<v5FD�)g�Uݰ���p�	;%vx�6Cܺ�� ����敖�3K� �떶QSfo,��=w��?D���i==}L{\�?��R��|f���Z9@�S��������:������r؃��.�\ɼ�����G5�#2�� ���$
�֦���vPo<���Wt���..�L\ R��o��z<1�0.t�w�y�JµD��"��'��qK�� S(��e�u�i��~���닋�'FP�2�Hb	��7e.�
�
X�W퉸�7��d�9y
��s���~�]8���RB���N>���S3b�g�KV��l�AH?����*cH�Dr��m��{��$y�[�cC��O� e� �o�����������.,�h$Y ��s5�/ 3�$+��$���pcn�arJ�^Z=�AM_�d��٥K���(� v5�8%1KZR3�}i�c
�g8��u<��z��)U��LS"N��wI���v������(�(e���RAᡆfpXm	�Ɣ��d�U������	����%��V��%@ێ����~v￣f\���w7�N��9�� U �_?�-`�7��:<a�����j��
6=�Q����!��W��bȄ���Dc@���ş�(
�!k.Wt7O>��f�4ao��p�%>㽩Ü�^M�T�J<�/�ߦ�Ɩ#��S���:��`��f96����4��f7���]^�\-����[�Z`p��������XE�T>���[���*�F�;i���1Gz�M��OL��7������dĀ�S��$T��+�Lq?�7"��(��l���<|`��c���xU�4B����U���f�I��0rZ% ^�-��d8d�94`�k�NA_w@e���8^��)�o� Q<��:�8���]23$��� ,N�Ȇٸ�"~gr�GB�:�n����\p=�q��o����(�*��ڏ~���qM-۸3_�J�+R�E�6��
�퍖X�í���#!��+�L�7ݥ�ˁ��)���o�鿢W���u���-UJI$�瓈+�����L��	�,d<�����1�������L�UÖ]h�oH���~�j"i&9�WVU���T����[����<�s�SѪ^�@}t�������_{w�nJ|���w�2̿�z
�ÅXw�ki 8!� ���O*I,�)lC�%��l]ΣcP�٢��#8 ����ˈ���2J ���Խ���,�*��}�A���Q�H�8�/�|0��S@4ǧ����ې�@W���Ќm*��V�įr��kR�}UV	ܢ�
�s���>V8�Tܓ�4#?�0��3��Z��r�#������)G��s['J�):&��:eG�4��~�*� ��w�tE���j�|����� К;k�x��#!J�k'-��WQB!�A��P�R�7�C�G(�d��R�(7����}�Q)�O;��ڴ�gU*�0, �)���}��5� n7�R��_.��T����!qLWϵ��j�>w�	=�q�(v峸ء8*�M_�>߷Ի V������Μ ��B��$�@��
��c���`�@�R��Z�^�5��5fxWy�b�,tk.����fm@��?R�pO �<P���MV|�"��J��T��H�/i�(h�{�Zr�ӵ�j��O͊�2���$!���v��\��TR���1��m�6>[�o�[���@t�0l��yi����=�X�O��"n�$k�����A/���;���
M�z�*�(��ay.���Xz�u��������"�?��4��\���B�-98��B��s�?''q(����|1ϓ[8�:W{U�p}�)�Rm�*�AW2YM&�C��]��Ij��\��8R��e����ʤ���^Poxo�S�#)Iוϯm<Կ-��������m��k9xV9b ����;1�v�_��+�������A������	��:8m�6�������AH�^�j��WVE$�mbU-������-_�Z�Fa5� H�b���s���y+��|�|��Oʥ�x���7����%��E�L�\1��V��jz��5'�ø�5�p L�ƙ����A��ȟ|e�泓v����",6.��>��� �������ox��#n�N��tT,�cy�1��T���<��{W��0�Y���#>gk���κqP׮Ns�TlNNÛH9�᪭�γ��� ߴ�W�(_��ܙ��yz=�!���#A�A�b��fh�:�����$b>�nv�<n-�b�5�iջ|P��
��s���Ϸ���C��-qqrj��w�bh�`$g���_����;w����;ҁO�~q�7�ig�v��U2���	�����O�� @�Z��B���3��z^鐹)�v�X�#��٥%����%���v���:��Qϣ��33��Ϯ�$4Z�|U~,�;��nK���H���:��o6@2�����e�:^Da÷�`K�""9a�|�����C�ѹ��Q�� �{/Y�gh~�$��Կ�>	�X��\l�k[����bk���LC�OB����!&�&��zFFȇR݆����3��pⱪ.��J�h�mHLd��fd�&��	V�a.�>"MHk�q#���~�l������C+CnK�`�Tx���j���Y�Ϣ�9��I�/`7Q2^(�߾����Z�H`]�\ #��5�a]��π����vO����1;��t+Z�S�^��4���U�Z�r��������Y���Q/����jb��"�y"�,�
�������~|Rҁ%�o��?Fc��_R�ù���1&�ۢ����7-6���l�0�W�cZ�/q@��0����m�j�I��k|�nCU�Vqa"�g����uU*Y*��}�N��y�G�kA�B�[�pn�l�(*��"�U�K&���m�YR3$�L�j�}7�F�S�A����\	��zԿl�=V��+���7�X����ƥ�"͔|� jO��f�R�<C�h�8��I�N�w��R�ٺ��̓K ~s��nc���6��"͂�dL�WH�ߖTn�y�&��o�7�#6�L�dɝ�_�+�a�W�$��������br�����x�����X<����\v��)^��H�$��pb�H8�|�ܢ�pF��.;��x�ӫ��R����	y��`w����3m�+P��# j�&��ɉ���*�)����Xk?��;�E�֟l8[��[x�)7M�u�v~̄��%�vZp �k��L6�Q�8s�����|�h̀��*��]Jdͷ�R{m�Y�k��'�ڐ�ܩ���8�Q�N_n6y6���\���K�.l�7�ӷC�xxVOh�4�$�>D#���˕��sw65��V�&�����͆�v��j)�� �Ο?�6�D�d����$^t�t�	X��#�#yHh4�|432r��V�|����y7$���2Ab���p6����PD�=�R��E6n��E{��q��\}P?��[���nr������H�ᕛ�/�aZ��<�����A�Frw4�6�T��O@���*#`�R²:[tΩ�'�.ծ � � *PC�:�k���x���ёY�)<��4�B�r�*�.R
 �P�/GoQ.���o쌐�9S9B?��un��mQ�<NlÉp3����,{E0��%R��H�l0�:ױC\:���A:�ƫ��m�,徊����o���^�2���'�����4SȤ��kGs�k>o~�ncy�+X�FZ`�w���1xuVJ��+�5y���I>��*��őT�ka�=v�]ߴٰC|9{ؘ�ݖ9w��|�:;�����N��:s(a��z=�>d�+%aŝ#�J���KQ�d�ܿ|��Z�DRX��	o	�OM��G�?ۧS�Ԡegg_f�B|)��=�J���K������Q�<���嶇C=`w��_e����ɢ�F��ff�bgs�P�~'�Օ���Ҁ���� �/�O����W6�]]0����߼M����Kn�h�Q�u��,�߯_���(2�tC�*�n���rt�m�4!+�D���r�D��R�;�7�L���"x�-7�ֳ�����x�kk=_��sA������=��W�d���r7H�=lz5#�!?����0�Qf+p�PgL;<U����y��_�`\�?��M������y�G��G��A�� ��S��\"���2�⺺�S�c$Z���X��V�<��Ֆ4��#�|G]�����Ԕ4��b���r�Gv $zw��C1�&A�Ej[����#��d�|"�-i��!@L�J�8B3���Jw/�¾i}:|x`�)�sҕţ:!�Bv@A�ͽ�[���5cUPK�z4�t����|#���"���9���S�q{$�MdE�iL�0^ǧ��ߵ6�Э���o�V~(�d�sV�����8�30f�t�uАu�����;n�>�j�#�(�X���H97⍎$�r�oK��<B�M��Rʧ�g��^���>�b���v+�vb���8b!p�Y"�I�L���^�7
D��j����'���H��B˝���'��h߽Z�ў�Y&�����e�zV�ج�gd�zM�E��/��]#L�u�,�<���5�\fi�;b���t���|�[eAea�y>L���Z��wZ����[!�FƊ�r�i����t�@�&Lop ��\�C�=�|!؄�p����ߢ�h�'�Kp<���+wyc@�4�NN�0�_J��$_JN.���;��?���� ���58צ�ٓ�}����U��Z���+Zq���5���F������'���0���3/���C�v����c��D%�p��ŷ�9�Ώ=tzqA}�K�I�yk]*iy�Agվr�9(�m��2.m@d�i��|�`������0�=�f*�,z�6� d�y�O����"�g��)�����j�Ii����͈l>�ahP|Q���3�'���g�b� (3ڠ���]�^�+%�M�U����1���T.)Rah��./K�b�t3��J����)�tM8���f�!c��%H�Ꮛ�e4·�'�|����4��p�%�Usӷ4�l�cUou����>|
�r��:�D~�?HOL+���U��-�~��S
!$��/?���L@v��ǙCɑ�fd 1(,H��YfH_��4�#���b�{ˣ}Ү�Tl�����?{�b`,C����G�Lk����w]�H��^<82�RD��+��sV�^p
�s�����v�qH"��Oד?�V�{#��cBP��[m|yyG�a�ޜ�i#��d�DLȆ(��;���}�y���)ԃ�[� ����5D�Q��PeH�m{o�F�S<co�&���w��*&A���)�b9(:s���=��j��)�MlUSe�al����0"yr�zW��ԣ��ũ�x��1�e���"��6=~-b��7����k�s�,ƫw�lA�N���@�'��g�2�?���`�����M�K �o�K�k�1W�+�zO{x�WinY������K@�SB��̹���0O� �]����p�%Z������7<Ԏ�sU���I(6�j�(p��P@ ��}�O�a���#��x𔜪hP�Y֭�Z�0x
0m�S��!�O�5�3n;m{�y�ޡo����W|g"&y����mD��c��0�X��<{�_��Ͷ�����FM��)7��	Be�U$X�(��h�Ñ���]c�v�Bud��!{˘���8׵���X�0g&��JV	g^�����q�7x�I�~�,���A��k��u�`rXlB^L,�����͂9j�@�<vVw�9�Oc_q�S
�����ڀ3wo��`b�J���ۻ^<��^����k\�z�Gj B�A�|�nr}�u����-l��¥sV���z,e->^���ו4ӷzv���gnm�/�<`Y���c��%�|�dEFx\\��Es����ﱱ9F�L�zP�J��t�B�i��╝c�R�"a7�"�$(�L��ܔw�����H�����$���H������*l�MwY�$�Ƚ�a� Ͷ�y�yZ�2�N*Ȏ��71�h����FꙌb��;���D���d��L����2B��Znڹ��Юz9�f�2
��mM��/�T�}��!+QSnM{�����Qr��0�
�m����ib�K1(a9%�G����ՔDf��fΩ�T�2c�2����ux�@)��nT�� a៘�-0�gI���e���kB���|�n�
�.�n�d���ӛp X�q�u��꛸�~Ǵ�1�eG���O�³) �-��E��8M�?E9���)��˷�]8�@͘%����E*EF�Ĝ�s��3^'rK�uG�r�.�mHUa��B<�Y=!WXC�J�8�mn���Wm��5}�X&�<l� `[O��d?�n'Q	����_U�za�^��3�K�3�~�T'���/����e��Qx�Z����f���Q|�,��"e��-�.%fPҬ�I=�F�c������X>IL���Vcʔ�R�Q�Wߥ�)��"�*��V\�Ӷj�������X�3�;���OM�X8ݳ�ܬ��ʝr���J����H����<<�Y�����P���H�����~`��������P��{��AnM6M3��r��ǉ*.��?�V\|SfK�a�B�ݓ_sM5���[U�aW�aW�o:�k =׹:�ɘ>��	���&�����!�Q�tE�}� M�o�xו���J*����?y����Շ�/mk!H8vj%8X�(h�<��YG���_���Gn9�|#�v��^}8��H��Ԣ����v�K%�ҧ8S;�b+f��	�Q�ah)��etub>#ۃƄ�t����������}Kд��V��7�nl���̟�(={S�g�(���=�`r�&??�<t)��ڨ��Tb~�$��ڪ*��������D3и��!�k���H��|���Ù�G�Q��2Dkx[��=q�Z�C
�A�dy�x5����t�%�����_+R��������U�����d\���G(Ց
	[L1�$K#k�u�;�K�KfJ^b�9��?��`���ٕ�M�1ӕ��m�����ԇ;#yI���`ڲO�	�D�˃�a�8�6P�ͅ��vM�L{2��_�˥�kZ@\�ůV�'�sS���x���n��_��~b�1���b����$�蕳?��EYSk��&$���s鹅4�7T,Pn�m�S����	{�U�S�
/��O��$Y�⒮nNO~0�e<18bpb��R?���GN��n/I��w�y�7�T��>�(��^k��?9���������RQSYY��	Ɗ|]��Ta�Β/ �WR��o]O�7?7 l��y�y�956�_9����K���'y�gn�i����b���E��<#2N���;w
�0f�F�i�6��'ŰQ�H�|�)������W�3�҇�9�f�[�t!���vV�lLQr���?b�
�33�a��	W�U�0n%�L"���rM�H�am�~��º�C�xO@�W{�(���R9Ƕ�rW�~h\��y^�-�}p. K�S].5�!�1#�0J�|�y泈	�N��b^�g��D}��G�!ݻd����>.�O���������(ɦ��>��W������.�1O9$B�(���G���h�d0���^Օ*���m6���CT��2~�f+��(~(+�t)��_<�JjUTg���@�lS���ř��k��@��JB{�}����U��մ�0o�b�����3�;1��2�1F�<���'@=?x?�O-�ũ�e�W0�
pEu�T��z�9��y����GMs�Yv�4;۩�S�s���)�k��d��%l��G�}P��BI����9T�7F���*��h���P�c�\��XYvwΈur�򺪪�_��|�"�55���&���Q��%�2;{�N��Xeq���P$PR�}�S��$���]c�䚰���x����N(H�Rf���ې�<0K�����f+��^5���Ύ����f�^��i�	�����{{$��)gB�0K}��|9���-��Gliφ/���"Y����,�[��^b�ů�k\���>��M�?q�'D�q�!��|(�T&�����fG�tQ�!�}�HS��8�#v�y-C���8f����Cq	W�ŝ��X��=��g5OވQ�Փ�m�h�@���n�3v�`w��bN�]\�W����e"TX���E*��X��N�V1J�˼�cl�*$2��4��x����j�^�c.�Z�S���c�vF���~n�� P��c���)|sE��gR���?���\`�ߞ�5è`"b6M㻥%��ʼJqly���[U��W�h\��Nj19_H��� g��׈�c�
M"p�f!_�?�ɒ~��QXʔ���R�]���Jz�۝*���b�FO�h��<N�Ch۵v��<�jT�fF`�.�~T����y˰��Ψ#L��qQtxj ��Bx	��M�]�^D��I*���`F㸯wiۑP��'�X z\n��|8�⤑�K^rV.J=��w< ��f�لW�]���77��N�"b��s�,YW�S��?�:PZn���3\ܼH�d��}�,zP�Kk-�~v��ْ�Yʒ�v�)E�ٸM�<a����H���F}K��nmǝІ�s���2�w>���(=�ٷʅ�4�;����e��1�2��+V�_�g��>�N|���|S����w|�!�������sۅ���^�u���~��h���ψ{g�I�㨚ٴm�~���p*�+�W++Xq��w^�^�����-��������G��x�v�w����. :�F��>��������<��r=��n<ܗ��%GY�#��@�Ƃ4_K�5���eŇ�jW�g\�x�߆B����3��N�	 V�U.�T$�|qR����i7����lG��#4�9��7���X�E �F���=-i2�s�Ỻ�I)�?P��T�ēm<@F��O[F+��O�Ŗ��I�|����O~m�Q�H��[����������ģ*�;)�^D5���!��$���9��0�ؚe�xC_�W~�6�U}��M�dV�"ם}���T�@&��)�(���ʖjoA;�Kg@�S	A�����n�F�,���"-��mh�s1�o�g��\�������Y_�9@��ҽN�n���pt�W�ȏA�L��
���޼�$O����R������[3�y�z����E�&�T(b��33�V)�;L�>�
�I�PO�u!��'��w&����KA��U�jNs�����N����K�������_}�%�{�,�
��Y�4��΍����/j���մRGw�9%w��RO�~��)�����n{X�1��-64��)�w���O�ĝ`rX�]����FK��r8:��4&8ϗ�j��#��7N�*��n���Nߥ�·חw:  ĨHƗU g��AV�7$��'���j�pO%��$�Z�����/�fG?(Y�ְq�`��;��ˑfІ�ӡ׆Ͼ�����=��F����V�A��M}������:�Q6����Jv���N$w�����<$�����ק�gj���.����&��wtX� m��D��O
毶V�1;����O�/��= �.ї#��U����\ݎ������]iv,��|�,�/2S����e�PF�mr7)Kw	B�b)�<����7wudBR���}��sZI�`[_@խ�P�az5��kN��J�U>��T�A�e�W
٠R��Z���[\�*x���.��vr�ܢ&<dXE
�DV�����퀦�Y��G��.VJA�~̧���4�laBk1�"�P�WS�k7��״:��_̓��l�d2Y�X��W�h�	l�8�	<��K��j��>�0�༷��e!����'�y-�~�6�����>r߲��ֵ����$T�M��Y"gt|�+���耦Q7Y���h3pL��4�:�~�+�У������t�v ��p��?��k�V�wtd��}��t]�u���{�O�P)w�W�&�BQ���*_'ī��)�mcdX��Sc>��!G����@��_�G��6����~�W�3�^��`�w���˯]6Z9TNo� >�����N���(���>Ib���[�!��f#�v ��C�F}��]L=�>�̭���jR�y���	���c���ـ�'xё���Ć���;�AJV���S�s~Wg�}�X�f���)���ZG[�p�c������=�5W�at�#�e���	�������x-f�a#�ꒋ~�e�J|[n�c���[�a{����{�貢.4����k�7_��a�ϻ�X�}�����7����H;�}�5�s�Dy��W~~���2�/q�|��GX<6��P�K>� ����U�m���(�v]s���L��.���/[��n�q�����$v@��r��^2B/�w���CR(M�N����x\�7�`�DL�n+��'�:��]s+��|s2-鏻�)�tO�1d���w����~�
��+�l&�Ot!lfE>�/A��e�4u�KU�بZ��0��=�P���#��|tF!t~t������uE�Ga[��K�p-C��;�`5G�6�X�O�Ɵ��������7v�޵�H�h��6�N�c8�Aʳp����4�υ�AT�h~�Je�ѝ�8�]�c�Z�~�Ң��7;��C~�:��k��$%\2�r1�������r W>�1p$����fm�sL�ܨ)�Cc��W���9B!>�S �ܧ�oN��pWo� ˒�����cA$A�!^��w����hT9B��xA�H�]�m*L������tw'�����Iv��¼������La`���#��o�HTڔ��%�_g��w_���P Аs��>�� J���0`� ��\q�v�0���"����B�6��7�,��q��`(.ɿUXF�E"_UFv��Z�9x+@-SU�(I-�}�������
�����V�kky�������&*��t����#(���7�])M5>�;�����^�.�w�W��B���W���gχ�χq��F*OUI��#�|���7/���rKj������o��!��c��m�a[~�Q�o�?Q�d�X�I4L^ �d���ϷL�
I��P���1���\�����s��=������p(�K�ē�,�Jo%���+r��L&Y��v�cZ�hcTo�s��$��?�f{6����|z�~��K^��K��	����>�E�N$�;`tb�b��
��M]�>�All�O�߼����B��Kw%ԋ>̧����r�#��N�}�q�L׍~~��
��O�i���@=�$�w5\�����g�}�[����"T�<aª�oa败??�U�I���]����l3���ؤ�ڸ��D�vP�2�l5�}ŷ}<�����	}w��N���\[�U��Q�.6@|��k�в�>�x+�
���ք��Mq(#�@2��Չ�)�\L��$kKꬠ����D4/g�`N�_������h��������BV�:����ee��\2P��>;f�ɷ�b�*��)/���Y`ԝ
Q�o�B;����7�J�n��IB�
�߽�^���Y<��
5=��Q`5Q���Z�ؐ�I�%�x�w��_�_uX��U��^�}w��] ����O��"���{{{;�#V)挄������?/R&��J�w͑��+^HV4��t3��nL!���J�_
)F�d*�6(u"rz;�C��)���j6
o�A������ǧ��q�,s�h�q<?@�wr�_?�P"��@|�����nf� ��~~^����;.* �#xx�9�'g�K�f!��b�QŨ��-"��!'ɺ�<�Jzs=n�.�x�p��R�����=���<���n,�e�[W�A�M�%]����2ö��8�ܜ��<�\��H[F�L��n��Qjx�Y�4��x�8�B���t�`��=O��]�t�<^q���=�N16�
q�cc�no���.�_���W�g�%<E?6tr(r�L�}Z�{�
�<A���Ь��H9ynvln�߄�My��ͼ]EX�a��U�_x,ĸo���%���:��j�t(E����o-}n���`�
��� �1�f�9w�
�fv��b��U�	��&ҌӮN�
��2ʧ�f:ϗ���c���
��8��*�X��#�
�z��[v�S���`�,��:��S���j%��4T�M��@�x�L�Zn�fs�X��f�܃Rgr�O)AB��((s@�� �����m�FC�tQV6w����Tl�f� �e�4����p��g��={����\���XP�0u���s*��� qc� ����	�b�p��u��zֳ��������π.�|4�M�OĎ ��~���i��%K�[�6��}}K
��r��<�.E�R����5Zk#"����Fx����� O;�\�٧k�N���'��}�SO��X��3� �*3�ft�+��2�c���9��qpB�%�%�˷��̲_�r=Š>�^H�uL7Y둾>�@g;v�T��{�X��A)�%���	i�i�����xi��~��T#-�S���;G���ڔR-��p�&T�+>�ou����Y�ņ��MYt�����CXz�Aܯt�\�tsw}4R����؏��Z�i�l�4��	,H�xg!L�Z)K�)��	�H���-�QO8Z��+�c�>o9���j@K���ͦ�ɱW<���q�[n�YY�v�u�9�f���W>Zɋ�������S�Y�6���s~��[~���6�b����O5�W��W�|�R�K^�&�l��zM\�𣏕SY���T�t�[X#�z>�+� �&V�%Ts��Ú)��L7��*bA�ELʤ�>�j(��2�8 �"^ġ�֒�k��#�+C�"T�L�n
� �'�?�mD&�-�a���o��B�a�w�S?-�F���i���º-��ʺ-�ޏ�`9�8R�>_͒6 ��T1Bv��L��z��N%������8��&H�ܺ���UD֖���Q��������{�����S|~�3��xZ�| ��
aOO͌�V�u���OL��$y�"��������Ÿ�5sY3)�J+���*׃	��pB��@����o�Q#e�x�IQ����J�8�=��UO�ruk���zo>��ɬeD���T��[�%Pod���M�vCØ�����cǙ͇��
�!�I?we�EH�>_Lõ���� Q��I�y�� 'q�����4g镬ޙ�]������;1�·��h��^^nw�#j���u�!�=q��>%���]��E�Æ��c��ù��Eq]N�����9�x[W;�?a�mvy�w<��غ�$�?���քA~��4��Cmu1_�!c�i�_O�$w&&�yn�k�I��^�cFX��pdC[�A%���v!M��%Җ�dQ:Www�a�ot�ԆQe�~�x�Dδ����qo�L�X�]B͵���E�"Hñek��6�רU��J�Ի��l���=3Ds�cT>b-����5�c�+5yp��%µ��N� �DTeOl��Grv
$*7�`��*d�,��%�T��%b�֛��+�m�*��-��@F�W]�[�3$g���N�5L5^8.�'���	�&~�k7���_G�!�+N����s���)*I���4A�@#C��\�+gO�ϣ���;w"6�r+b)�>���_c�.�&��}�V=���+uͲ2L(�Ȑ��3���;4����U�V���� ���RG�}Ic�5��_sf�n��&UHf�8�aVq'q����8��'L��>-�����gUFb)��N�������c��AYI	��17�}8��J���`��E�ɲn�X�x��Z���R��7C�_2߶�9�]aǇ��_@9&!�n45ci7�����b����M��O2�z\*��<<�I������Sv��DL�Bh,n�������qHPZd��b�?.X'��-G�ى>M<j�9At��������ڍ��@u�ū��e �����#�F1������H� a�猀�5@ʿ�*�/o����]DF^ֱ�r?�Rll�	)u�y�]a"�{��	m��;V�r]5;�����kfN=:۟����j��A��90ϻ7��&�7�y�����^3�Ɲ�&E�H�͝7�gwO>e���]Y~�L�+:n���΁��]@�dmYLi��P;��A\Q/&��Ee�t�}��4�8oe��1�L��tGH��ó��yfb^-݈]s�JyH�����K�i��(�R��'��?~����󇇻��7~�7��ꫯ~�S��Ԟ�_��_���_������~soo�f�y���PǴq8�F[e^l]�v��H������ã��Th�tR=��Ęq�z�C���k��=nQ�p ,^�%�KT�q�,�����3ĉ��J��H��j���q�(|CS@�5����Z�1}2�ۚ1����ٵS���C:�& ׃X1���6F��׎9ZL`��y3�"�{I�m�����#��jmD�i���O���D"ӉA�y��B���g�\6���hpf�N-}Qk�ک�+	�f3�U ��Q�#ZY��f�"�Q�N'4�>�ik���K���Rh�c�<�1�5���`�-]J�k:@�̕�a�5LԬ$Qǽ?�7�ެ?x��H�T���.��5�60�C��y�n��ct�q��G���uD��>ڎu�|h�h�E'>�#��Z�NC����$p���k%J)�H�s劋���N��| �ڌ������)qCc��f��Z(��aD��GhjS�Ӥ;\�~��u"���/w��&-�'al�@R���<��Ŵy����ӶW�~/���e�ᣏ>�_����9���G�o�����o�~��p�+F��y���ڮ�
%A.d��"���AD�U-��:_An3l���F'G,m���f��� t.��Z}iNcYb���[�$؉�Xq��_g�yxb��nr.%'ij<9��7o޺v�����կ���|�g~�_�����_x᩷�g�%%��_���u�ߦ}������}�M]�5a��g���;�^��=�ϏG��,���޽��ppҎ\��Z�V���JT��$Y)�����J�3/}R1Qy=��1'q�#�Z���;�^��c9F�҇s�S�T��K�K�jYX��d��	+����\L�9��._�T��\���5R�vܼ$��PSU���.�J�"���Ѷ�~�>Y]sL��m���d$x]����mPs,�*?AP;�iS%Zd�#C�*̺Z�$���]���u{!���%U�o�����	��~"���<��K�C1�{���"k�����[��SWN�M��:aZ5��xJ�d�(ajg;�q�F��#���0��A�@W}�qI�BFI'�Ab�"je�p��Ӊ�ﺵy�1~��O��aDAh8���w��=Y� t�%�q�h?Vc�Lj�>Ʊ͵u�AC�e�!��0q��n��N�v�bc�S��Ϩ	���������g��S�(�$�ͦS�ñΚo+����g�?p�{�m�,g5�S���76/U}Y1�fYS#z���X�ɢ&�,kf�f��	+
+A+����v��2�z�̏5�f�������� �����{��?�}���=�����[�Vg�hp���d��A���^��,IHIhH�����NE t&"@c�#}�a��WR��Õ�/���B�9�3d#j�0d3�R �J�QqsT'A҅G�Yِ&��y=K��۷�>~���g���������͗��ͯ�����>�ʤ��#�3���_���!c^:�<�ލw�z�;ߍo޾#�ņx7�&��$�ZR�#���XP�M�jvJd� '��o�rl�9�9bAi�q�y�HM	5���$
�6:0&n��
T8�(}PӢ�Ո(:��_P�ςf�\�!Q�>�hg+#�O�\��8�VDʒ����f�8FE�~��Y�q�!T�żf���v�4���O�m5h�>ln������ 8>X����,ǀ�ک�:o�@��
�q�=�K���RKCI��A���餥ߛ�D`��Aޘ#"�v�xB� pd���G��489<r!���L�'�u���K��H�+!��v�5�����u&�:ڀ&-�Ǽ�c�#��!�B��5�14Ƌ�~�ܦT������}�b��V�p�1��0�& 6rF,aY�����o�nܼ�4"d����|ἤ�I�k�6��ep���F� R�Z���$7�ٺ��o��0�>�Z��Z���]�w��L hNg��w����;X�9u# �h�6�Y�^3��V��s�C��t��hf�3��g���Ѐ��o}k���������oƓ��"�B�IH��F����*_�(j�&�'�}�LI�b�Y��wdA�	>K-`a�L�j3���k��f�Y�e,�;��������)dt�=#�N%��Ɔb� u`��!����5�0�th&% _�%�Ss�CR�����'�������7�{�;���o}�_��_��_|�����O?���b��O�m�4��.&��˗$F[�\�d8��m˙H!�*�U;�N{��:q �6þU��D2�J�p&���v�W�B�s����#w�����c4;����΃�冮�G�܂�ׯT�A06�wp��r�ةa_�6}�?4���
m�=h(�|/��.
�m<:vDjF�������<V����V{����������&J�Đ6����2��㱁0��H��	c�b�p�p��p8�����ǲg"����Ďd�-qߚ����׫W��=��s���n6i�,�_�X����~����@����d��7���;�m���8I�21
z$��������=�'DB"0�e�&&���0/���K�NJ|�vN�`��s�#L� ���g��7�����n�0x��|���P��um�������|1X �	��8����� ��*ႈ��	���z��]p-�})��N#b�^�dD�S�h�I[�IZKEw����ul�����k��(�5�@� �s�sҾ��h��%!�|Nzcʝ��xR���w���N���R���+aQ	�>Fc��+���t� K��w^�%IA�<,���C_�K���Q �G=����Us�:5��u ��u��ƅtНQ�7���\7\y�󱼞!Ի�1?��[���K���T�7�q��a��.rS�~�2����5r���딧�0��U�j�Rs_?w^�����l�^P8�X�_.�}��v��|��[@~`� ��a*��[`;�7�| �L�/vk����/,6Z���O?|}���m�T��?��C�n�S���2?p�3�s[�z	G�dBg��AJR�{�܈�����bwkM뷶ni��d��Q� 8��A�Ҁ&��B=�C����#�F�<Kb\&�Ҭ9Є9wFJW�����D̓|����믽^�q���[�7W����?��?�ҝ��N������vvG?��u��v�����l��(P����ԤH�'��$��GCР����_�.�>a���F�:���_���� $���&W�n�1��f�!�kS�q��?-D(S7|Ǔ��#*�KG��PK�|��2cڦ�y ��:y/���P�b� ��!���K8���S�2ЖXȆk AeYfJ��M˸�,w��:�k���r@��(�$��i_�2�����:zy�L܇�����ɾ����W���ۍ�3�P�{�{��k������y�RO��v��cL\0���$�� <�j�m��Ę��dO�=�������vQC!R�Z�BI�zM����p��ޠ����QkZ�����RI�'�� �a�P����]Npo���l�g�����SN6�\��r�\F�S���c-���1�ED�}�@��=�-Yܟ��_'`��g��g��0�y�{(���3���x����	�R�.# �W�.4�y����}K�)��V�#�I��5a��m�k ���{��l���k)m�
��ǘb8��:���p&�T
lL����{춁qo�п��������G����Fk4ᚢ�+�M%t-�Ulr8�r�4��+R������A�\����.]����]����]ȡ����Sl=Ru�(�jT�J���^��9Į�f���@���!S֙5�@	M5?�I,0�J0@kK�r$o�9y<���~��{���_��W�~��88�\��ws�����v�v>%/�#R[Xe�F�_*?k0t:�5\~(���t�v��۾?�с�D Uk��E�Ĥ�&[4��:���>F�]>�;Nd��4��V�,\q!&t�ȓw]!i�P�D�=��)��
c���z@�0��@
&O���&����Ea!B�<H�<F@�I��]���sx���\��(E�f�e�2�a_�i�<��`�@��xD9��ׂ�?�nȵ?e̎@�땶�Ց�2����.�c�4�J���"���	r��5Ip�.���U_waH���Dc����o<is���R�\
�-���S_�<�܆JuL����q/%���s��(�XF�Q�#��R�1��Ԋ.�
5�a"�B���B#!�[(x0���%I��s� ��"�����+���cb-��<B�%�_�ĉ| ����_U��j��Ӱ} g�~��V��Ǚ�?cB�u����j����ln�z$@��#,P��"�a�pܜ�WIL�=Ԧg���z�.
�+C�\.h���@F4���.���o���T��kB�ַ�5��/}�`�aﴉ�5��9���(L�<�u�Ǡ����&t��_{�5�A�r_�d��B_0J7��6A}�1���8L]C3H��Y� �\�',|�X�����w\ʔ½�)�.ĉ�P7K�}����F>�FCnnm����M��\q���>���K�[7_Xn�':;��|��ϋ��R'�Z�%MΘw8f������JALj����њmAKM�B:/��r7�9(����Ёj%�%���3>�|�A�}��f��bG�X��[1*����a"@��&V�k� ��
u4Qs�PH����4H� �e!�!�i����q,ý��|z0�1�3�k��u�la�>O�3�r߉ہ-�2�{h0SN���fz\�ھ}M�"w�����z�8�*!�Ӱl;�vн��蹉'OS�. �b#%sT:��w6��،5��1���Z3 ˁf�Z3[�0P��}��;��f�%b� P������ۄ�Ѓ H������'�]��:�>m'h�\���sl����9�B�:��x�rv���Ò�*P�5s����������=��,lWǹԫ8��9sF���9���\c�C]�(���%t!��o��0�q /������*S)�#=O�%�S�%�ߕg��.Tҹ���}�k��Wy����1K�d������>8&
{�)�7<�Q�|�:�p�	Ձ,<Q��)8�>h!�dyb���q��5G�p����GRa��_5s$u�����f]�&#�U���(�ʜ�T��CI\6צ*���7���ZҔ��R��sr���"�x���[�/�}9��a�0���Y^�]��s:��3�R�tèk0��:�2��I��PdNU�H��q=;0; 1��b�@a.�pL��k��#�!ˀ6T�^�iu�A��^�3\��Ag��?Y6��b<Ae�� ��e����W����âE��k��7����V������5T"��>W�1����ZZ��ʾ��.�P�l,8@���
�LpL�ǧι��3ۅU��M�6��ϡ}M��Ư�����֦i�l;����_����D���B�����	&tР] ���א5T�����!4���?=	HC�9�Mq����Q�ܓ�`TQώ59����V��	7$�+�I�T�`	"5$�d���*u�%��9nI�s~���+8["��}X	s�m�a�b^��8���PPP�k8ЕK�B����i72וn����ٖ9������r�p]�~�&�`PT��=e1�1��`�{Ƕ ��a@s��s���[����5�l�YY �z2��W��X��]sm�`cz؂���An<:b�M��@AS7�uFKI��u�(���$Q�3���]������'���A��<�E S@ٴ�<��d�)"4�g��,����+���{O.��'�I�!���iD��:��	2�1��}j�jx�c�D�;B ����FD���DHV��� �
�T������Aw����|�_��W�O�:��je�˗_y��h���z?&~�Ȃe9� JTҘ��)���iC�������Ϥ3��}8V]��{8UB��8�8�i��&�@
�w�uM�L�@ҐH[�!oK0��i6��W_6+�X+��=A ؀����I(��?��]4�|����l���g�
�����ji����,����P��ָ����狏��5�����/��m2?��2�o>��w��l����}RТ�ɭ�^��cp~����4ٱ+<8�\���xq�w*,�=��6��>qBqq�- �Қ��Bl��S�L��\#`��O�J�
L'C>_D^5m���%h�Ѕ`��=�'w�}c�^���꾪�sA��I崭8�Fb��I��1���8깄�  d���j_[n-
l��΂|k,4����|-�Y�bW�*сO���Ɩ������]����{v�@�5P"WW����< �C�
�o����u7IpOp>:4��sP��矡Us�+1�|�g��X ��w:k+k�Փ���\g9��"ty��r�?,`S�bӬ���04��=��w���5r����	��^x	�s6�F�~�@���Ep��A�Z��[axF�G���\��7
��@����KD�hL����$�I�L0p�,�	��Mݫ�~�I%����+����f�W��h5j��Sp���(rU���8�G̀ )N�b�N+*�ea��4�%r)USe��c ��?��"�~`n�	�(��M9W<3��m�s6ΌI�B�<PsT&���?�{�>�
�K��$HaW�4Q6��g�(�	n�����/
��u�&VyF��Z�
��t�b.�ϠkE����S�b��'w�~��@E6�2)ۦ9xV�af�!��|��֧v^9��b���篠;:DI�ѴiLVa������1�u�5-^�U�����~�3��$�e���@\�>�儶��1�3�g�*1r��TY֦&�Ti�/��ǩ4HA�vy�����s=�;*q�	&e3��V��- ��ÊE���aBV>��
�c��y�.�Q���e
:�:����P����:�P� r�s��ߋ�I$F@X��GP�|�qMv�3�	թ���ɥ`��>!*���s�q-<&v�r�;�+����j��QPf���뀅�E�n͉7o���#��U����Δ��J���`A��{N�P�8���884�b̍���w���������Xi�(�����
��e��Ǜ�����=}m����<���qW�.OtA�M(a��b�������T��BmҶ�f��å��*7�~�Aa&$[��K�Un�pǔ���~P��Sʄz�IK�=ǧ)�9�B���yI�aO��*Da�K�-À����HJzE�~�R�����s'��da��/�96��x0*?��	����;J�vR�F}E�B���a�̄lm�v����H�,����A�E�r�R��^6����kx�zE�3���kD�y��.�4TL^N�]�>Q�B6g�y��E�7�׎U��>/���5k����6m�i ��$�fNjt��o��N�O�<���d�,�^�t;������~R>N��ʤ��Eh �:�gk��/��h�O��a_?�-���y&�/@��;ӱy�+��wո�wj�~�:&>��#k��>��u6��LM�<>?L�l�������D�]Dj=�l(b"�dӷ�C�ƶ�H/�������~Xy��Z&G�sJ�r֩��R95^\f ��_�/�n�1���\@��Aᘀ��s���0�0�5�����/�Ǖ7��s¹�4/�,*�=�	�4o8G@�p���0�HU�-\�	�����-纓�,`f�{�,���c!�
*�A�)b���V܀J���Z������wz�}q��+B�t�R��W_M���z�nMZ���Lt%�p��=_~ 1�ܒ��DA���Ͽ�Z:�ԫ5�qs�Q ��=ᤅ:_�3>hw��f9z�)�8(�W��BB���u�\�(�q|���
�b3i��ĕ3���m���*�r�a2�nc���?������G�ܱ��x{{;���@�-�$�� �4�d>($�[�9kn5��?�8eL��&v�E�9�)Wm�o�҂q��<~���KRu1�sOݸʓ?5�ok(H�ɇv^L��_cf��s�@Zj��t#& �F�m�]��>6��p{�6�d������7��&�����	|���Nb���M��9]m��6�����1)�zR���x?[��}�ι܀Uc�����Aq|��5�, ��f�_toX�q�^`{����1�YKd�)[�X+�sŚ9m��F� L$�0QZyM�ڹ*"�	 �a:���+�$�s��������ɼ�B޾Լ�������j���(��Ƹ"n�>�:�|�T����1]����,>�l���}��gQ��dw[�������1,��Y4�K�>���1��7�T�
,�p
mU�wmH)]>�����q��-��*���$ol#��D��ň�,!�
���e����+j�X#Su�y������^W���Җ*�K/�QT���k���ر{�X;��_�re��K/m��9��	려��M�*Bi�2w�T�y�,y����0�Z�4-�L#,E�Ii�Z1�y3,d fh� ��8ǹ�rJa�yɄ���8�D{��di�c�nf�F����u�裏V~��*�kU���G�M3��P{q}�Z0
M�	m�TB�x�BQ�i��.MJg��xPh�$�F�I/4�W�H�pC�܌�F$��q�m$�
<&[��&I�NZAȷzt4v�~�Ϗڒ��;�w�|�9��qH��/��M�f,�۵I�l��E9eOߛ���m�<�X��>G�d���|_L���X��]�	���eE0=�>�]��;���8�&��"̱���s�����/�۵�m�ǽ�.����>(\��+�w�GUX�4ۚ�Ǡc[ϣ|�T��!��c���Yh2�xQ�U�XK�:pw@56��CYH�X��s� ��4kR�F����q���fz�q3��E�ಯ,�,H���3F�+k�6[Y#�Yz���7��G}�"����|��0�S��2P�G��,��q� ��fA��o�o�q��u��|^��CS���}}}��Ԣ�����#)�������AM��C$ �\x�-5Ѱ�rUA����N�(��rX/�T�2X/�'���[�xuu��g����فz�,�
 �8��qT��8�a,r��W>N�Y�RE	��ͪo�gR�����,+���g��R����.��!W�b�a"�@	 NH���8���Wϟ����?>�����\Nx`X⇛�"^s5�XdQ�IO8�qIR�����Gj[P���%��fR�)�`4
5Q�!�H ��.Q�����{�<@T�=%_4G���Awn^(͠P߹�M���%4a+�KA�,�%�G����)�|jk��جj&1����~w�m &��ǖ	��ӧ#L�,c���a_��'��r��0�M#"�[��b˄`�^�Ԟ�y�e�	v���%����p�~�V��p-%�wP�A���ާ���	��d��eO���,{l� ���d3?�ۊ6���j��"O�$$�U�P.�р�o������D�@3����x����E��2"⮢�����ȱ�b-����q��bc���GP-R�����}������G��{����ن4i��h�>���o��:�Qv���Zs�v��)���C"�9�7�'w�D�;斫������D+-��ͨ�")x9���*s*�Q��
E~vw�H���[���J*S�!������>}��x��+B��_�ŭ_��_�ʷ������=���s���}r8���3�$7�DE,%L�w����d���ls��Hk�lp�Ze�9��1O/+�����@g��'Xr��E�����e��X�$�_&O�0㡼{��:�`���"�c��%�]��"�V*QB�����zr��z�"D�B
%r�ÈryS`< <r�RN��g�B��BI����q�:����R
���޻z���*����̅E�����*H`k`B�3k
8�Z8߸�E(��أk/���E��򛧡�>73�g1"���d��r3ٚ:�;̵�mk��4�`����Q��TM�0M�ױ���˚Jy�;p�s�%��:���5]�ƿ��ښ2���-����8{_I:ߕ�ɕ�xv6,�ںe~�9���2�ʚzni��Ε>���[˄�9��}� �C]1�-'��4f��Q���Th4dϴ���n?��r���[2uLu���A���(q��r)���$��+:؋s�I��k���=�c������1�a��I�.>�z`��t/�H����y�ɳu�M�(;��I��U�,��"�s�N5cWW�TPFc]m��t��y	Ρ}u�CM*ٜa��}�R����9P�;��u��N�Ap�ި��cǞy��9^/q����>"��}���Uy���aʇ(�����,Hz���qf�r����rмU ��q��[q��\�U����񨨌�B4A�L��S��]zR��xIn���6��j�9�'��'Ƒ��qyy��]�0M����˛6��Ԫ��z�R���A=����?��K/��J�$OQ�țR��k� �B��x�F�!-�Y̙P�d!:
�7qN>�$���Ŕ�
�8O�h�K�����2{��|�d�璹E!���䔪gk�ln#ilim�;/Mh����f*"�*�zem۝�©�v�!l*;W���\�w|Y�gW@���wָxs�6�t�������t�P�{C4�`�5+-����c�ƾ���y���)/'Tvf��U\�KO��(\�$���q���ǋ�.��0�잇�S��ܾ���j�2��iΜ�v|�aCjΤǺ�g��JE�فfM�^���b�2�	�]�v:Ƣ:��N���w�����sj�Y���[*V�^@��zU������"<(fQ�1`�A�"5q,���,�vw� M��u��w�Q�*6���8#�(��CS��Ԫ��k7o��]���q���u�<'7d�k�t�l�B�e)�U���HK� G�h�w\F�DeB���x�V{^�]��͎�}em�1�V�Z�-*�I�ӈ���R�fT�|}an���߷�6�H��'�� 9rw�'�}���Z��k������� /��<[�l���7&�mA���V�_�#�p1"K�p�Z��x9���49�'Qf�L��0�=ڏD~�Tk�߽�ӛ���-�P����j���M� ��L4���v4�)Z�c��C��ξ��4��p���v�a�����4�&�I냽���_#{�屦����akv��S"���y6aOx쿹�z������^��E��Ok�y�S���
�(tQ�E���	��t��9���B�4}��6�k27�l������&���8U4W��{�Q1s�)-�ϤA��VY�b���=/H���˙���v�� bL�P��s��Gv��r��%���9
���F˾�j�.��6�5���*�M\�T�=���������~r�;W]��*��L�5�G�
�Љ�9s|�C4�SIh�RYp�%(}u������>	}��\YH��r�?k7ۿ�l.�|'�ϧ���q�7�pck�`��:�z�Zn`�)�����!D�T���z�E%t}�B�Q^�͎�� sNӐ��(��|eB�A��盝��Ч��DݘF�y���\�ne�1j���e��$�uܠ)�Qҹ��k��ai��ʸ O�eR-[*����t�'`������u�e�up�?WI�&���|6�>Z[+�����?�<��T����`��yR&��bU���"v��D�3�|�=�M2��Mm0�J0���$A���Z�k�*M��nu�D�\�,&ʜcI��h���y#k�����J��p���Hi�c����:��rj|4!l���\a�:�B��HYB��&4	�甹������l	BBTE^`<' ��U������kC�s�,�}�U5=$�.կ�=2�y�U�b/\��NLq.�\3y��&��$��5VA��]Kc��!����!v��+<
�����;�V ̻����VV���'�5y�����?sf�?��w��V�'�w��nggg�~�����,���d9ʰS��ƋJ���2g�M[��������&R7��(A�	0��]�kI��.`B�?j��	c�x��EfL^������|P����dZ���4�8�va�J�t�h�)�5պ��Q���UTԔ������O�d���lIC՟��
�����fTW������,A^\T��G9�n�q�6퀸�v�Z��H!�%��`�Z����.ǜ�`��tJ%p�Yv1	��ԲI8=V"�V.U�"�=�ҥ*Y����/vt;��7`����C�"4Y��*t�dʄ�!����)�����۰�c�
)ARP<�9�j�����(�;�	�΀`B�t=���y��g8���@�Z���E���~�J�sn;�S��|��ہ����8�(޵M���oh�P�y$�����0�z�T��9���q`~xA�B �]	!j�-�Rױ�>���@�X�@�$��
.ԃa$�+���_�����2�����;*�z<���w����?���}���/��C766�9}�s���G����Y�Ul�K�� x��^�ls��重���I��z��uP��B$�D ms����L�dVSڹi�5���#oґGU����QB!��x
�X�@Pl�ƺ*G�C
�.�SdN�t@I�uih��k�ߋ�
�d��=�09�A��CKfy�Чy�'�i�D�y�te_��uXI�H7�u�oj�E3o�U��q���9'ڮZX��C=<�*4R@��u�ЋI7����5�S�	��er܆���ǂ�ȋ#��fi}NÐ�t�"�X��K9E���C�G�e�>���LY�V�SD3�޶Դ�T(r��:OA[��NX�4���(k<w�e����O>tܖE��.M|����`�'�Ʊ㣠��#]�g�l�
C]�1�6�x��nfc
��X��z'�r��KF[P�!W�k֛h�H�c�Q��'��v%nm��.��-����u�Sk�5�p$�q��bҟ1��Q�y/Q�h�m�a,c�0��X�eljر	��*�g#-���EU�;���h!�S���D{�� �*Zk��AN;A(�VW��$N^�V*�^���Ν|����iW�MxB��{����Ϳ���x�/�����{/_�z�࠿G�镵c���j�J]�(�f�^mTk:�"�#|�i"�`}����a%< L�'�G��&J��3�厣j��L��^���`"�!�R��T�ۑ�>��=j4����'�qޭ�`+�3>��"�����!tM�t�ȭJs���ۦUaq�e��<����z^8��\�Ư;��fk�e_8��hU�4QNk���3r�o/'�
����~��c!�k���]�î)`�� n��PN%�m����XB���ɜ`k���#�Z���>��t��](�V�J�Ɣň�?!Yɂ\���[x�,������,���0����Q	B�fh�4l�-����+!�U W.��گ*QfmH�`ff���]-�=X�v`��J&P7X��M�)�2H#�� p7@n9�ʅ�=X-Ѐ%�d��>\����ɡ��F�R�n�Q��V��WgO�_����-G�O�'�w��_�
T���/|ᯞ�����srg�s�`�?�qs��8��i7�����Z��j���\�%��j�$ ��T�sr�aE:H'
�O]����BA&=Ԅ��ݠj��C�c_p�JUN�P���A�,T((V���T�h��RI��b�����.�˧\s&6��쑠0浗}�<�N�bs�T��R�V�X�F\�5p�K�T�&���)�� ���e.��'�\)���O`��5fA	��m��妛��*H�籗|�Ꟶ��u��,�i����(�}'�7����Q+Ρ�ԑ��)�1
v�
��{�۽ ���h��T(::��u�G@=T-��1�&��l�(r4!�ߛ��s[֎�8�%T�</%�4��T�bUYj��&~x
5������s
re���1X0��iז��dU��o�Fe����
UAM�I��q��p7s-�Pu[����~E��׵f��=�z�[/�t��'���wL�����g?�YH�����z깃���׺�����Jg�{�?�m��Z���Iy�Kr?٬��I-����U�Ҁon�@�EÂ���ᆄ�FvM�Skr4�Ey$8X�&��Lr09�ʇ-Ld;��U�qJ��!ʝ}]t�K�8��n�D���D�8���qј��T9��gi��vs�S+�ږ�Mڛ]HF��9�0
�|o����I�������y�����X�%aR{#�à���JNz�C���w�m�^�0�a���m�O�~C��㻍���a�O��Q*��v�L��m��Y)L�v����>�h����B�L0�;��wp{�! �Z��eQ�u@>� ���D}qcs����ך(k��6�38қj�+�\�9�x�e��-��̱ueh2	�n���6s	C���µ���sЅ��m)8l)�ʖC�y-��x$���O�ʂ��c��Ƭ�J;���sM۳�n��q��ʫ����vG=��
<�����OB���_�җ�$	��q�j���umaw������|@ޘg�\�~2����ı��Z�ծW�(�V+X_IƃL>|��>F_Wፈ��7	"T�7kf:�]������|��;Ǻ��'I0R�o(-��Z�@�c|��������1��9:�D�?:�Я�<,�=���D��e��ڎ�V`kB�c�fm��L�$^X�Y�u'�ΐ���V�&^�f�sԻr���l�d�-�VX~q�vgkՎ���\��ۻ��(`z�Ի��	,e��(����Fo;&;d�@R�]�6P�0�B5.��Ca�:?��7ɔ�f����͹��'h�)��6Je�Iaw{G����:��Z���~���vPa��(}��C:��p]刳���Ҹ�@�F�zSp�]�N=G��������|�Q|�~��A�Nf��`Z�z�xj�-gch���Ou6��V<5Aq�T�su,cy|���x��T�lii�kg�<t�'~�'6� ��Mq����O<�*����k_���_��x�y��n���������v�߿v��͛7�Uk������|kq~�.	��kxǁ�Qe*�M�P�/L�"ŋf}��y^J� -'p3ǩ�c��c���P%���zQi3F���P���S�<7|q{��e+����n.L'8��]����L�OƜgZ8�-��`|��w{R�ߔ�B�7�%�j)ʻ����&Ӧ��b�u4h%���mB�fRw��w2/}�0��.T�oe�y�A��8��駧��M;�҆�f�'@1 ����!�/HG�
t��tD�Q$�!�/�c�{x���w�"���p��[Ș��M��R�p�"Қ�[�8TV���l#��up4��H�Q����Q�7��=��S2�CvPXe��\9���c�-�\p�,�{�"��u��r�ݒ��rݿZ�o�����������?yW��w
O��3|��;Ҟz]����H�W�^mnn^_������ytkw��$��'Zs����bmn�]��͔n|�N1���%F�fp24A��&:$vE��*E�Bp\�I�b"q�Ƈ�|OY��n"xS���]d����ԡ.�-��Z#b��{hgBk��c�{䦻��`��	��:��O:��oM�������{�yF��Њ|^�|��k��L�� ʄ_Z��V4m3�U[\M׭q��!8A��ww'��6B��4�ҸK���i<�C�ѝ���ૣy�V�Q���uU�/�,��b�ֈ��3c*���D�!������K��y��c�`w����$��+#2q?���$w��Qj����\�����5���$vv� 3_��
�re��Q� 1�S�� ɠ��բ�qɏ���?/��h�÷�����E��g�n��%e�;�b��0+,q��e s��X�2
�T�q�a��7��$_�?��h9ܺ�Ǌ��ܭ�nuŮ�U{>H���3Q��� ���>����P����4=�����Y�0�s��k4����utu�����.�QQ��S&�3�	D�{?+I��L��AD'�q��	��"Mb��hh����~L���v�.�'=k�>�~�k��	�A�.�Դ��{�lٹPC���	�M�!��X����V�{A�ٲ��#�� g����vF��V��P��J:%���Ɠx��ģ�����1�2�?�2��U��G��訖��D��E�����V���̫g�{�`�^�"��P�4Hq{�<�ZaO�y6�9�|]���-������L�:����c�a��Pώiػq����T��	�dS��Ch��~������P}���e��eu��ص�����\4���`Y��%w���	J����C$gW ���ɢnO���	�;�GX��F��|(��4��6|W�k�8�xn���Y"�\�)�KM�3�W*�V���ʵ�/����<c�w�6L�n�J:��5L�YNp����'|w��3ƙH^ϸ��1��_aa0�mpR��$��;���Z�j����K9ϓ�2�j
Jr�#�
s�Y��b��nu."��[[�>|��K��8"��0��dt�b]���[P
ӥ
������Nt���Y��.t�{T��fZ���uPg�Z��_n�IO�K���������K�^[�&VZ����O\�nyH v�k*��l�j��/15ޏ�#�+����Km>Q���ޱ�Y��ã��-
������:a]=�CD�7N-�+�}��{�����v�J�7e�r?�Q�DGV�\�Ñ��-�������l�	��EۂO��O�%��;�.��Q��3���%3nU��b[���%�չ��{6�������-i�gѡ��ꪝ�y.����bcu5�j��VT/:�3����y
��@܋L*ZQ�Ye:�������*c��N~�}e������W����$����7@Tj��$'ԉ�M�^�u�k+��4)N�^�/Z��<�����	��_�bGE��{(.ʸ����VKX��0S�\��N�r!أ���|(NRK-�Jq��zࡣ�?ɚ�#=�m�~����x?ϳ�`�m���׉�Z�}�������7H�瀟2eh<2�CI�����ʞ���d�=u�a��[�����i�G�?������ïv�؝1�gh4�ı�`�*���=h��n�V���m�(�� �+~���S��g`v$�;�q�Mh�'�8��,�Ǟf�I_�:�*����3J�����M �#'Mt���J������������ļv��`6.�k�L/	ʏ��v����>�9�ɹ�ZX��>�+�R�G.�vu5��>9��aR�fo2����u��i�xa�":Hh�4�+I�C�&R��;�n�ڼ�C��VեD�,��!�hk��i)�F�^��AjI(R��m�+�D̢��Æ�2v"����9��ʙ�^EZ$��v�����P��2�>;e��
--aQ~�L��:X�B�3���}O��R����[�q�����mv�]�m�u�Rbk���-����5�{���3�mr'�)!������#hMRV�U4�!�9�y�?�ZyŊ�?�I�}Ѡb��'0��n����2�vEa�`"mf�>��Nz�w}-�x�b�����> Q�1�O�M�3���!ɵ � w��"ۼ3Zef>��WΊI2%)����n���1�:��;^����;$6�L?�$3���R���k�RH}�m�>�����;�l.]��bNN�m�'��8�mn�`X;��V�l9�޲6i]�^%�>C�4��f-6R?q#j?x�Vǂ����R:��fV8q��k����+��Ax���K����GJeR;��9=~�hZ_i鍵dtt��lmg�Lb̘&نX=��pk�t�����մ�U�q��|A�9|
RYTȗ��`@S���c�+�-�E�����ֺ̯W-I�?�Ўy���®Ws����Fxw�gv��Z497�?�]k��8<1Ȩ�Y	Y-�,c�`� ��/����H��b�HD\]�R���^�����W�<ԥmA�M�1�U7{���?/V�����Z���{�,�b��|��;�����p�آ���Mʹ��G�rzXx�g����(P�������t�=,[=�ގ��8������G/�.�~L�"���boM�^o���"�\gT[m�n �C���"�/���`��D�I�T�!>��"��s��vn��+�qV%����K?x�nle����%W~W$0��y����'�(�,㴆�4�0bWNz�,�.>;_�n��o���3TУ�^Z-o�l��͔Ω��"\)��݃�_�=j�c��eֶ鿭�ȦT�"i�V�K��=z¼確2?����s�>y��h2�����D&���<6̵�q�c���	}h����Y� �:�£É������"��)G6@d7��ן��˩��@�m�p8g��@��0��Yq����as`F��Lz���}����#hڄb�����X�\)��39��Fܴ�s#�HqN�FHg�a�)�5�� �:���%.p��觖�	�͆K5՗��nQw�p����N��6���������Þ�eN#J~!�𻥋�� (���hֽ��{�I{���\�\��+�������/.���>W�\��7�o���
�N�/|���9m�tس�Ņ'u�:5����6ª*u=����ß
�"?�B"Tj��:���Ɣ/=����m��%�D�j��?|9r��E��H@[ ɏ�B��=���B���^?F�_�g��#�x�/�{�;O�1�-�$Ȝ9�iw82/f-e�b#O������~H��`����I�7�n�^A� ��%�]��d�K�#��)���&��%EVKIb�x&�~��Xן���V<|�sT��Ҷ������&9 ���&��*8*�j���Ŕ�x���L^�b~p'Eٲ�d^��r���]�{Z��jX���zD�g^,
@��4�|��X��q�\�V���O�~vm����S�4����4LY��j��sfvd�u@��[�P�'�C���ft���G��J��~Dc�c�r�Ju� D&�f.8�3/�b^���6D���e��﹍=&v''��*ymB�S�gmh�#�1A�!1e#LԜT`MML	�WV���VI�`b�J1�����%"�gE����6��r�4����|����얫�ݖ-E�/=���%^V����,����*��N��?i+cJ���3�&���:�$�>?:�/�D�7��c��n}[�!ތz�lB$M=jTV�Qz�5!B=i=�x�����00.>��z C
�X��c5S(`]��뚼$��� �>:ci��4�x;vlM1^נ����6�:q/�퇋���0���f�d5��_�[�$��>Mi�o?35'g�|m����������*(�^�C��1�n\��������{�E�\1�\N��L�FX�%��U����	F�?%�嘜�@����0#��qI�1�EI.f����A�f�L�����U&�L=���3td�Ctr�!Ԇqqț|ƍ�Tx�xÖ�OK�Uj_�$� R����f�!��ǯ�fG��[p�2 e�X�I�0���γ�Ջ�����w��	>k��q�Î�/�L,�̀�<ɋd���z��Z�(6�*���F�\9kN�	H}�P���^����jb>�˲�eˈUg�����rc��;��`�A���U7Ҵb�'a���pr���DKЧ���Bt����^`>�<<Y�ML�!���� ޠ�I����\�aYm��Mk9���n�T�Y.[�w�o���[���|���]8>~<3js�W�yY���a���oc[Q��zݶ?��u^���]��O=��:�]�U��; �A�ЎV��j^��vk�f��ä��|�1�VX;%�8��h^�DDi����c3�cr6����6l�Me݀?��'I;)������΅������c�e�`�!�G�0�&��a�13i�x �.T���p�+��V\����H�/kУ%���.-�إ��mD�a��ܬ�s�F�ߗ4����S�L�a俕��I���\���	�DB/�*�M�#���?\m���1&,{���K��y��~�U+dM-��0i�p�\vY��c�O�2�c�F��AO:6��M,�����=4@u�q"�!�+-"R&|[0W(��&�[�(G����;�0���9(�ófUܔ�����b��%���O1�w����G�YtW��
O��"x�r��?v�@9���B�w�C��
���EC8��@H�X���d]�s�N�y{�.��cqx��ƫx��ǵ]�>ћ�	�;ʹLa�����>=��>u+�g g�s ���f���u���Y[�t=C��X�u�A��H��_sE�(4c:����Kl�ax�U��r,[���<"��'SfZ�i�K3<d�c��bxv�ׄC��?S�-�����J"j\���TK�f)�SH�-.�_��y��Iث����jՊ�D�4��V
xvڰ�mgq�rG&��vy�L���P�����-���ǣ(Q�9u���}���"V�y>E"lpe�'0�w��M}!N�H�8��A1�JG})4_=���X4����4&��p�=������8	��o�����N'���i=D�ez�͖qbh�Z�#@�qm�I����7�f��:�;��M��=��F�
����כ���԰�l�S�o!�5Z�Ȧ����������7XYV:�{s��А��e���o����]�qQ`ٱ%N�J^��z������(y� K(��4�=� 5G�?���Q��<�7���|��`<|	�5뢏m~���9~�XT@��{W��;�7�)/o|�A�v� ��(��,�U�.u���}�
� ~.��,�\nt�Vz�,�]��>&+����B֭��L�`��ԍ��8ۏۙ��E�â93,"~{Px� B�}��se�BvV��,�����v�a�c�oq�����'K�p��ĕ������&�(��h�q���U�'�	+������mȧ��1�K%cK���2:��bX�O�Pt���ctm����-�C�p��}���[u���~=P���u�$s��_S�I5 ���%�&!�����nm�d�Vj�5ri5<�����66�w��k�Hq�����u�Q	��(��D��K��b�|�\3"R�Pc������&��gK�����t�ٞ��\��9�H)�D����$%��� :;(C5�����#�o��W�9v�&�pTQ�2gpx���9�8�v���j�O��N���>J�s��"@yZ�tEv	��̏������A���K^lcҔ�J��%��	�M�97 }�� 
�o�o7а�L:���EQ��Se<�H�|�H?�� ���@���_ 7��I����iv�H�:+K�r16&Һw�.]a�f2���y�����i������Mn.�<A�@%�9��-������)�Y/���Im4R5�0EV�"m��� <��"�3[,���m6V�l����<�0�K��2?��}������2�/U>�s1��j�-֞�'���j��D��K'����x'!���2�)7�R|�?���F$�N���@��y2+�,��.�~��n�B��/B�1��;@�p�ȝǍ-ٍ6�H{�gM��o�ADTs���p
��tfIH���a�˻`�`&q��)�0j"Y�g���L��E64
��u��1{;�l����ή�z�l��9�~��lt��4�H�\(}��\u���ބ;��@�ٻ�H;���T�Ǣj�� ��|݋x��pu�_B���#���N*��<?w-lg����W�V�V..r��׿�E�e�1����wYP����8mU`P�G�l�lP��P񝱛I��]F�4z�V0�
����,=����|.�r�嘨r�pʀ��X>cJC��@�{��U�D<�9�[V����o�'|��B%�Qv���������*��0��sW���̮3���Fe�O��m��:�T���1�c�]NO�C�B�˽�Tmġ�d��{a_��Tvt
=6�"�;$�l;��~D�_E���2cx���K�-�4�#���@�I�4�s��l{�/_66KϖPb�� ���L����V�Pa��Y������9R}��O��q�g+W_��o�&SMu�X�-f�楂e�=�?�w�-m�"�(K�NNN�5���sНL8ljjQ�ָ&�J/Ģ�Ml���?�����¡G��#Jd���X:c�>s�ph�v��k���1�*���6{ǌ�}�N6��^ *�0ԕH6�Gce6!h�:K0���}�h�/�20Ak-�@4g�<�HA���AK)��#�Ą���<�i���I��ɼ��1��*#�qG%�wX'��^�Iё��/�nN�@=�����3^7x*9�nw�t{^Ҝb��-N6����`��ѽ�@4�{@�v4�tMa=pc�ү�9��V<ջb��i�jyv��Lk7��8I�=[ ��PՐZ9���Nn�]ծ����έo##a=FFF�;���k���9Lyϯn��1�$!����	s�i�B���s�l�<d}]�ĳc8`��H�����v���:"h��3ɺ��H.�׉{�3�>guĨ�/r��@ ���^͐
İ�C��P�M�[q���������� �NF��'�{�&z�\��
������e1e���2R�-�+US�)��`'�Xfҧ�w�w�&��Z�ʛ�؆jc�*�-ߕ��g^V��	i!VF�#wE����ׯܺ���$z�a����:T�)�z�Z��U<�hۗ�iz��.����:iQ
��[~��s�mp,�V�BNcbv'�����)�o]QN�]US�z�kt�=<<��A����e~���k��4�uog}��9&�Rض����.h��wT����c�L����]�����q���+�`Tu�pQ�Aw߲�^R��i,���E�y;Y���i�}���	?Ic������w�wzDX���M&�0:�d;�Px��J�!lY@��/4�k�q,�nHI���yB�g���<n���r&H��Tgɯ$�/���s��S���V�*�n�n��^BE%m�.�t�417j�����@!�?|������뼛m��**�+<m[�Io��F+�<9�n���>SGh��j�����H����J�I[�T��[��m�{=�0]�$G';��߇�CB����"30z���X6HWc���Z1O�K��Im�m2��p��!%����|��E���X�2ۜ���[&&�	�;;�칿�Zy-{#�e�G��zD��QOA��0�ZI�|��4;L�@ ?����>iݯ/�b��}�9S��K~gǦ�C�R$��tN�I�J�Rtx�CkS#��㙹�WM��y��
���-^�_Jx�CR���H���v��q��p���zV��{���o�&����P���#o�E��7���� �d��I���BAp���1e�Ug��`���Oqf��,��~?eo�AA"d|A�K���͖�����vQWS�D#�wLJ��oe�GX<���������h���Mj�!�z�x�ْ�V�D!��e���}d����+�N.�W����Ƣ�*�@����n0o8s�� ����a/Q*b�Y9�(�$�����������Tq��2D��5�=�h�R۪G����w�l����KY	�'1��sl�I�Nֲ�R`��^��Jآ}���x)e��o�ft����������pP;�� t`�-�fd�i��ͭAˑ?'8S�C^�ڜEs~8Z���~-S�S:�܍���y����c��Oy�u��l�m�mP�N�vk�B�!� "�4LzWձ�%���4�TX��6�_,W��u$��w�χFB("�V�˼�Ƚ�h���W鱝iZ�� $(�q^x���=���k�����'ݳ���pI�"����'z��IjU�,B^����|���h�߷���U��[h���ml�.b��?�rO	8m`�Q�������P����4o	-��K��y���5h,�ؗ������jџ2{��E�Vׁf��1[��%g��Ʒ��5���dE�#�RIwhA�����k���vjſ��Ќ��>d�?i���d��b,J씥=h��^�ʽ�*�Bs��Q�4R��W�d��y��94�QXGO��#cb�j��|�eao@�U_������]"�K6�ւ���#�Z�B
�D��.�����JkL|kJ���vg���^���u��iy�A�[G�`��<�n��\'6~`Ny@�ly�Ϸo���e����L�x��T�GY�3���ݿ�? e�d����p��i^��`l�8�4 ''�Ѩ�����+xcc# �� |ҥg��s2��U�]��GB�D�8����z�ӡ �L\`E�r|,ɝo��CVÓ�̰�#�vmx��V��V�`+��eo���aV�ʏ��G�n��WTK���R��܃p1c��U�05	?�����rWM"��x
y�t�WT'fR���q�����q���z�m��W�"	���3�&�@i:�
���B{O�G�טʺ��S�.�!�Т��cE:T?�K��n����)\3�y��P����n����-))!!&!ykQ��g/��9�|T�nWGE�wo�b 0	�B,��7'��'^*�m�BR%�����op��vy0�=����М`]�ew;^"�|�8�UG��b2��(�2vΌq/�v�?SЈ���S��u�w�'K�$�-1>�� �>�D��Y���Pne|�*�Q����G���e���9nm�Xʨ`��¶j��h�~�>&���DuM(i��%�`���Nz*���4�r���,�PF𑋅6��~�2p�����y�7Z�u��������.5�T�&a�:�du������_��#}9�r]5��+�وa����8�M�X{����Q�nu�:���+�=�{��j>�Xzy57��x�����Ba��_kH�/�[��
ՠJ&����-dH�U���u�,�JVqc�/�.�`*�*i�ԝ�(m�Kϩ�`�� �L���4`��CY'$�.�^�A�����C�\9=sZ�4����-ldk+�|��*=��ħ(<f�ޫd=^^Q��8�-YV�>�#�#*v��F�q�o�N鲲����)˄L��[,�͝�Z�N��)!q>���!��@�ᗙUl��wjEe���1��H�e�q"F�}x<6 m������� ��p\��&�ӈI�� ���)�S����%=�o8���o<]���ޔ�������y��8��v��.C67k�:oM\fΰq E���ƀ��p��wRd�E�D��B 0�([��=���XV���ȇ�L@���V-�QX\�ŗ��}�Σ���	</o�۬�hBB���V �/ aYS�[lb����>�lY��(���7dC�X(x���̞���0����%��@�r9���A�{d��")V�{����*F��~�[�,l��E]��a���8J���z��w����
��[����o�ip��H+�E���$�
��]��'�|�JpV�#|�;5,�zz�;���Q�[� �� DwǨ���ǲ`�g��V2�oP@pg�_����j��RD�(Ga�:	�>����|fU��roP)>�UD�f��?fRz(nǩ�4.���&����85���2���-uQ1�co�a<�B\�����PA@�{q�G)t��/~�$�*>��)�;c���U�A�c�Y�0��e������u��G�9�@
ŝ��C�7{�D�t�Y��l�闙�^
�#�=�ݿZI�Q�Q�����5��/���n%��?[�Q�����$��x�/y��P����{� ]�~{��¥�d���ү�{`ٚ��$F���C�͆�΋{_�!A�˧9#;���e�c[�i(��7�A7-�xM�/��	H�����!��t�6ʬ��L��,o�q�<�f�Opfc�d��߾��2�1�4�d���������_�Z�)ZZj�;���D�%3'�(;Eۧ��B��G����j+m�x*���U����*�ӷ��zA��d�����+/�e�jBt�Ȑ�H��s��Vll컴4�`U����>�U�Gmb��?B�qeb�n�l54�jcC���Ī=��T� �����nթI���f�KA��p>� �r j�I�T�3|Rzv�Ն[�(�9]���������
ؑ����2�s���a��A��ŉ�`��l�_!(i�:�tY������oc�˙3�\���ٺ����&�m�I�K��ӑ?�W;����K��mQ�.2���X�̿���欩�{����rOM��v59��t�v9�D�/o2՝��n+�>j��;��*�F��G��J���[h������)J�5��?|�h�U��w͜>K�t���R��\!~�������o&��4�4�g���b�"�5�JT����?���]��H8�4:AHd�-�%��Z9�1R���_�8-	Z�{��^���s��_�r���vp���%�8-��Cf�*t�w\;���@�.9�W�o��/G�=P����+�/�_����ʐR:@f|��3V�\�0F�#�����s�sO�iB;�@`)SI���I(CC�X}΂L�u�Qmm�'��[�u"=���vO�9�`ce�ۧ��&L<U܎�jr?�UKἆw��2�>������a��3��IF����FMI����Y�Odz�b��輺,��+��#�Q�i������ ��3���i�~�����Y�]��<�EQ=0��F�N6�3��[�n���=������ ����E��E��S�/��e������ʍ�f5遟���~SL����lR�)�Q�f��+|�9�-e�Ie���%9��xT�q=$5:-�u��uK�6J���N�9�3{&g��͊��s>[��L��<^4G��^z��v]�"$4{k�Ic��3��x�|��l�q�%�ߌ|�7��i܂�l�Q5"�K�T[�c1� �IѴ,o��"���s���O 'a�rG�S}>��ai��� ŧ��C�v.G$)��(�$Vx�,i�R��OēJ�x����_�ҏWI�p��\��*���
���ː���l't�R�y��7�&�7k�%�k����K�Z�i�6g3/��p����C��<���$:��h��l�}�-�L��A�&���3�'���������b酭����0v$�gƳl�>�������Ϗ������'�}�Ҭ'ne�����;Wpa7�Q�4^��Ij�����G.�U_Pn���bp�F�`�0Ր���7	DmE������(a4S&����1�À�S�](@�NyQ�쪸h ���_a�q����qD�`�Q��I�9h��@�����y�K��+�v���W�Ǔ-L�w��_�.v9ɨ��0� ��Fn'A��/rΛ]���e��y_l���(�vCMEW����pP/B��	y$�-�)�-{>��#�{y�C��Z��l~�^���J�vY����]�K�(�������ǽؠȿ�;h��I��e�OGP�z�� �{xǁ�7U17�+�xO<B�VڇM	���P
ݟ�_*(,Y��K�VV'BQƑpv�f����iz��d�A��]x�Al���� ��|�I�,����N��k=�S}n�L�����@ 
D��2�B�=K~�������E6i]�F��:*i��a�
)�Yޝn��~��.�j�7	�#mBm%�ʏ=T�`�&`.*q������cE�H��3�8�pu@z_��44f>�cR$�#3I4�%	���j��1#l���X�ř�ʅ�5���>�n�������5Րc�Κ<����g,yw�;���S_d,+����Ğ�H�'��ƺ��_T����r�q ��Ҽu� ���w�/��S4�L�H	�x�了jX<�YYpo�(��7�I(&�=��F(�:���W��?�n��N�k-��ʌ.��ǥ������x�WW;;�/��a�h"��{�����������Ċ�R���O��yi��5�fa�PK   %�X5�3$ �$ /   images/8251b1b7-c97c-4929-9682-a545aa133660.png<�cp%\�5|b۶&vrbL�dbs��mcb۶m�Ěض�=�~u�]]�?��w�սzG()H"���  $i)q  l�?ゅ�/���#�?g/��  ���%�#  ����"j�Y�҉6:��MO�ݑOGݩ�*Zf�pf��pb�Q/BH�Q��Ef�8�q��8�9:�̶9�����Gk;�^f*�Wx����y�=Ow'��W�������\N��������/�������rb,P}�_�O8�B�wG�#�6�����e8K�Ż2)4������] ���( S� �\�ޯ�s������?�����o*w]�z����s�Mv:񛮼�B�Xn�Fe_����B[�	f�W����f�I�����Z��2w�is���9��F;��Z>!��xS\ْ�s�ݏ�M����3����7)�U'O4˽Ħ>�Ka1��ҕ�G�"����P����QK��?_g��n5_�x���I{ڡ�﷣G=g��?)�]Kۑ��� P�����E#����f( �r{�j֯e�wjY�QȘ�:���`�]��RFԊ��&&�y�M�8��<��s�z�9R��[O�ȡ���*�	^OP�oR7�H~�Zo�ڌ�.�L��1���&c�2�4�C�8�����[9iӔ��rܝ3'
G:��~����|~�Ef�H� x����F�gs?&����Y�yhK?��Y�x����s�v�m]ߕz�Y�>i$��oX�:k���^���\__������}B�����'��_��T<�ɽ���`�u�J,���֪�Q9;�W���Pp?�v&#���t�b��)����=�����y��p�v��BSȵ���Y��|�V8'����UE�����U!�%/�X�#��*?�6X�\ͶnԴ�G"s�����Z�Oj2����g�j��Ƈ%�vmk�犹av��0'� 䘙V�
�s�|�=:�gK6�rB!�z���{�#eؘ�z��#�ǐ?"�uJA�(#�t��+���!�]��7\�W��g���_Ћ��)1�V��ʭ{����@��H���S�����Ͽ%�ǰtP�����1��w��c�w�X��i�B gvy�e���e�u?؞�宪P(�i�.wK1rK�՗G)��3�	J�	%S*3��th��C�5\��or�L:G_@��/m+�Mh�Ry[V�0|��������|<�4�ZZ�q�`��!8s��H����W"��m�Z�SD���4�Q�/?�a����t�OiVS��[� �_�걝-�� ������`<�[#���������Fe��F��6���Q��6uc��ޒc��L���ς��& ����_J��;5��8����^��5~�7�\U���+>5��O"B�k͔���[I�������q~�Q��s�����=/{��(��3���rfT�@A�W�%�Va��N�v�h�_<54l w�����kQ��.Z�h5U/5iB|�jV���b��'���y�*B$��dGf���us�R�HE��2����B*��,�����O���X��Y%�!.����b��S�kw=H�O�n��-�h�Vw�8�����_	�t��Xm`�]�!\��R�q,1���^�h���<6 s�o�E;��7�`�ٲ����0���W�ݚ����=�p7�m�CZ���BNk��~+ܢ1��TY�쀦�[u|4�W�76Ma��إ�i���Ke�bԝn��MH��	��֨���:��'��Y�о\��X]�L^�#s=���v���>�U� "�����&�K�@����G��i��C�j[[�V����}�U.M]BN+�b=�޿C ��g�t���`�y�^U�+�jG����X�e��j�2�f9�%���XJ˛��v�~����l�`*2K��t�S�]��L~-^;%����7�����v����%��}���.�U��5���ԣ�y�n\���z�=�?�ǡ��W�$����O�9���a8�^Y:ð:T�2��n�?o>���@�����v�=fϦ�'LF\|,(������G��S�}�-0�Vytk6v���W$�O��r44�|���1;����L�����j`j��_|�G�<kN9��{�{�` ȓ�����0����ua�/"�aە1Q"��U���ld�dI�Z���q�&�Ja�:�$y'l�N�DݿS��QF�XGڧF�o�si�H=�D�d��$��!��{|f���7�knWK5��%��(Z�?w��b�mq��$��t{��&9�m9f�;�]��%�BbF��V��m�6�=-t\�dk�������(�[���o�=L��h��-sb7hg�~e?�W>�h��g�_6�`U(�_�~l��(,�fo$�6юv��j��\�X���r\$����$��\U�:N����P��$��Pڕ��'f�T�dN�希;��fb������mj��4��KI�?��W�K��WB��e�(�OA��O٣��ϫ��:�p�^�՞�]�>���`���	E�&bpeb�x�1&���&aA�}�mX�E!=�J^B���?�׬��ݣ�\0/J*�c�q�?^%��{B����J�x�
�ď6+��U)���I���П�5jO��PҊY]С:���%,�ϣ���?�����V^{�GY#۷^z^>o;�P�vbw������#ο���0�`B�tFT�R�+�p�93�8�K%G��B�x�}k��Usp�l�C�\�o1�o�˃t�z0�!��H�jf�];�2�Q����B�<w���X� �
%��MI=���CAo&��PRg���*{Oҧh�	����� �ϗ:�J�ϝ5������rDE�<UT�%<f7��� )N�s���&k��s���H!���-����S��n�C*�Հk�{�8��\���:7���_S%�5z��C�D��1l:磹��KKM�w�~����tI���c�n�Ol�f���`�e�
���=?��9�+6U��Mj�z������q����xY���<� :�0$>M�i�����MO*z3{�e�W������_ϝ�]:��i'DxX�PW�%V�"}�C�^b�3\�ۗ����߶���uoWU��~[ز#H��/�ϲ�D͌�+�ëhC9($U�A�o$Q���"�ʻrr�+O#�ҩ� V����֤A]�@D쉥�9��]NN}
�~��Ax���@q�@�!Q�kc�csÀ������P���tQ��)d2_�di��mZ���cr	ljlC7�4�t�p�Ѥ��^7�����9��H�Dds��ƱC�	Q:ǿ�AS��1����Q$n�����y�|�X
��LK��w�!Q�hbmhY8��*f��H�D�d��2���I��s:z؟Y<"�y����~ͷ�Q��K`��@����_��x�S�7>N��Q��UG�ֹ_je��y'�F��l� �0X�L�p��sv�9�?�r;�ED��#�!?��E2�Ne�~������J}G�}�2�N|�;	�c������ϙjaι�[��>�X"����.89�m�z/��9}G���3�ْsf���$�@%��2]�'SZ��
D=ݨ�~NZO�2��~� �3���.�ٗ.�o\��w�=������W}l�Һt�ڜF�����U�m���0@F��	ߝ���d%k�P};�J�<-A���
�x_Mn��j�d*V�Gd�Mr���[��+�_-�/z�^�A{̔7K����fR5�UX�J�H�W�%Ջ���R��h�F�b`?�����(�8��z��J���e�'޹��;;"
8��ቢs����=7����;r-c�OЃE	�����iA.������x4 \�:����p��v]�~�I���]=������b̭>H�T^��x|�`=�1�#{m�ód�+X�	CO{�eE���
�dgR�'{!�+���!r�'<�����l ��HJ�p���6�X´z�t�!V�CD�������� ��hm��햑-�:�=�U�0Y|�t���I4�v�v���;!��+}&7�ݖ��^�.��Oc�3 �uĻ�r)���]1�,0p��I�P[`e����G���bU�/����|`w'ڳr�8�-k��5Dihe0^����9��V;Y6�����p����]�+LX��E�:�ܞ��U*�;��֘Y&��±�!=����.F�w�T�Lcc1����>�����,�[��y��(n�R�^��M�������k�UG|k�)�s��}�����C�ag���|�j���4��ۨ�ѿݭ͊�<
ѹ-g����'v��v�.�r���|9Eގ�a�����iW�7��Y\���㛞�L�_�?��$�t�mҴ��!U��P� @����Y�����o[�DO8Ԝ}����*�|�U�:r���G� Y��>E�*�&�4lxլh�_�wy�I�se��['n���Jw�:W�ޥ1-9����Ks��X8`�D=dܑ�ڋ�b�U\����9�POʍؓ�d\,��o�ʦ춸`M�7��ۉ�֟�Ce���ry��V�x��X��-�aa/� 4 0?I� ,��R�k�6��?�q�?q.���]%8e]��@�@���O��c����֝�tBjT���,�_��IN,�� >  w�ÂY�qb��=r�j_�^�vn9��:{+*�`y��=�вgc��7��@@�`���ᄘ�c��
�ƌ\t��v<�k2y����hpd�ѫ�l|�|]�M7Q@��\R�u�1;
��K��YW������;&e����֦6Z�����`N�r&�Ŭ�ǭ�|��Z�<F�ʣzV +�ܰ�D��[~��y�ə��ũ�J��׻~�M�*hnc���8�ARN����L)�~�h����һ�sD��^?c6�������8��z�Գ!E*���gv}�z��A+��D��G-��ϣR	z=:w��|q�h��ú0P<�͇-����?쓁2j(�� (��	%O�7���tX�r,V5�,��߾)����:
nU��R:�r���͍�p[T��kE5�}��'�� ��z V�A���#YJPB�Ya���n�ow��!RS�T0a�������q���?���3�b��M��b�><=w�a9;P��O�Ff�0��l�.���4+w���h�39#紶Pg�cSB��Q��я����a�v�Gܹ�g�u�]�� 2Z�/j鳓��"ݐQ.&����*?+������A���-vf�[ߞ\$��Yr�GGe"Tio�6�E�3�x�J������{�܉@j2��cj
�3�{��lu��VlіT�F��{�L�,��Y��]6�q3���Ύe�'��櫑�%�UFa��q���[�B���x���6�g�b8ϕ�y��"� �i�EJ�s�˷���q��F��q{���B�
(�;#���$���p�I��'\��W֑B4�^rV�=���+��U���tn,G9 <�TT�o�D� =JB��3v���(��������$$��B�!��\��2܌l��)`���`k&�j��H�X�Y��z4Og݁\iDe�#�d�^m�0f�PNn�!�^���[�l0���Ć��h��nFٶ������1�D��2��G*��/�e6(4�"�����?f�]�K=��=��=�� �<+�(`��Tg��B:~Oڇ��?˧�M!�e��e�۫]�_怋�ԡ�g��Zk�+�8�4�'T��8�������}}LG����U�R�/�)X%`z S?̓��$��J�v.�Z�{.����� ��j�M{��g4"��y��l_j��������"�>�v�@�������7���[]ί�Y�vT�zo09�9P��^1+�[Qf���?��+�7��|�y�o}�������>�2B,Mw�-���Ay͏n�=U��^B��wo�(_�7�� o��+!n^������'�%����#����q��*�K؁�>����k.a�1L���O��~.��F ƞ\?v�ÔF.5buí?!AN�^� n�����F�j��y��ʾ�Ͽ���=�sjT0����<Q����B��_kW��'n�o�D�8{c�b�p&��\��d9�&���pǾ��ظ6���;����9�]�ӫ�4�,����ԑ�f�p�)���(�D���-WD�եD�C];���ܵp�s�s93�-ˤ]�2�ii&��,O�����r���c�GU2���ՅD:���e�r��P@�Q����<���՛tm�� L~�@3\MU��������eW���6_.3�  
�B0Ze�ʙ�튝��о<"^F7ٱW��V���%�V��m�,����׾��=%bA���f�֪�幔��74ha_�̰�&H ���vEb��ս����chjV��z�xp�Y�w%B�ޱsuO�E��<��}����[���X(u}�����`",���Z�J��Cs��qR���q`Lt��ؚH�������+���~�B`��3f��?֎�m��x:K�_��z}K��!�����T>Wnx[q�nݩD����g<���h�j"�c��i/��h~ �8*$�Ku�b;���x���	��X-�k��g��"P���ɕFrϹ�u/L#Upn�q:���M����F1�C?�wZ�!Q�(^�g/��K �M�8

qb�.�{�5� {C��e��f���̈́M�2��zp�o�Q+�Y�5 ����<�a�P��7 W[���A���0�jn�YJl6�bԃv��4*%e8cVGVg���4�OO͎�a��*7o�	m/�}[���B53�b6p�L��\�@؈[�n�O#Zd��C�;��0J�o�����!�T�П��W�}Іuh-�,ďۋu" {���P��='f$<��}c��a�9��߉��Ym���2ϒ���ɨ�~�>wcX�/��W!v�]m�]�E)|��}N��n_�(o����2_.�	��t���5�KkO�|6�˰\~.�ǻ�/^2K�7��_�31r}�Ю�ړL,n���jhA�}���C�럟��<&�x�ŷ�2$�Adⱐ6��U(sR�<��|"�~ަ�݉
��������'(�`�*<�D����n{T��D��8u���v,6l(.lY��Q.R�xs�-�~w~���=��ǡ=���1'2�\Ҁ���]�ts�+$��T*� ���=v���Ddܽ�g/M�\Lb�Uŷ������JB&�nvIi�`�}�2�yr�/�Դq%6��%��q�v�>^r��ڹ�/fy�{R����O�Od�.�˗�+���zWbz�h�8֞�{3=��'�v�yh�|^��[�G��-�.!,4/Q���/V��ٵP�]��\��_Hܽ�P��?S���>���>��ri?���#k�N��J�j3]�t���^:�~� 4���ٶ��9�U�Bĺ���y,9�D����,��N�i�0(K�>8�"
��\�Wg\L�H�F��MD�[LK~7�%�o��3�� I���Y�r�z,f��?ڰ�/ϿQ���A��@k:�&�:�D_v����?�3��Tc�t�@��g5��62�������#�ĩBXIפF���K@4����3"�D�pg�a��P�H���<�Pd d���ª�Kf;c��P8�օ����]I&r-�e�ů�7�Q/�Ԑq�2�t��Xl'N�]� ��G�/�9�kN�����S��H|�:�/ܣ�^�����Dg���_�Y��N\cD�D����NJ�)z�|�a���d�Z��X��'0��Z��NoZ�@"έu�k�F͉�Cc���I�I��_�>$:a��mtWA`X�kވ����ʘ�L�S�f�D�=���N�"*�P
a�vt&��(HR�|���+����o��M�4m��-���m���N�r!�$`��$�t�I��-2[�{9�����S�A_�v��̠�~��1��(4G�S�v�k��t��+�fN���gObK%7'���X�{h9L�&����c@`.�T�6Y-�zP���g��r�'_%���y�c2��k�v�ҵ3
P]('���Z,͹����4��lQ���uľ���C�٬z?�Z�AM2s�1I�����dQ_��Q��(>�*f��C�J�:�$�\��JP��<���J)k�y���H���1*dE�:����,�sDmGW5b�����)��'�r��,m��&�vM���moy�%�VeI9I����$���X䤣�&����Zgm���k�������@Rw�Z'g0�R����� ���Cz�#%�*��ÿ�|�5%cl��	<n��=׷�"/���ߧ�&���$�~VB[Ew����&�u��B��k��G�Q������*;z@��.+
��A~��	����(���2P���6 ���9Y������Y�?O���9ߞ��6�X��z.�D���T�k��t �x �Is���2tf�R�Uf�wâ,$��!^�7��js��s�\j�	'S7$�n�Hj
m��Ϥ���a�H�d���n�)g�X��]���S��Bʜ�q�
Ѹ'Gq?�f+��Ʃ	f#ax6vbS?���*Z��Fm���w�xVhO����7�8v���l�E6�Pg�w���-���h+�����!73/5:�0D+�m�5��s�k#�֟��4Ģ�#eR
7�II���~�-�]�(bNffg�������!$��,�R�0�a�%�R���À��g	Hyf�,��� _|��\�!������-F�݁�@���c�-$M2��M�۹I�M����gn��f�x*��!�v��&,&0-l)ѻ�sҠ�o̊L�zL���I^|��Rv�6fҍ/Α=v+�j�	�]A���{��?Q��C��]�俴`�|p�y��7�0 !ΩYڨ6�m�f�� Å)%�s���U�"�W/�O*����LU
��{N^H���ϼ�C��L���Hx쩈@��4P�v�g�1�3!��J\όut󒅁o�����v�}&�w\�\�7<�RcʑN7�V��z����!��y�w��� M�%��5Å�Z�E q��Ἒ�rd���0;�O{ _�̙X�+<�h�N+W���)��4]�e��_��gz`�(h��6[V�Q;�/�g�+wroo�#�Z4�ύ�媺-`�a�����F�K͚Z��+��ңvl���4���: 5�A*?��x
� y�#qTN�'�����p#���k"{@��F�Lꔑ��+��ϙr`�����dϔG��zd������B7�J���,�7)r���Fl�f��^�sC\~6�h:�K��߶w�t���E���m�Ϥr�r�g�I�l1_kH�1;y&��zZ�ë�����޲˽�'����Y�������{��,���.��7�޺F2�<�7����qǧ�F�dɁ�k���1�ą�%ޒT<�M@�ҋd%�p����5�O����Oo�����w����F�JQ�=�JH?dK#�������lY�� ����Qu�"k�Fi���>P/x�l�h�1�;LG7�������Ҩ�8q��@��dU?�� >�	<���P5��1bh�5�N;Y��=���ԣ��t���`v�������4��% ��x�5n�x;���B2lٴ�x, ��z"պ�Zi=D�E����D�{�ʡ�<�a ��:�[!��Fp��	�aX.�:�|1��NB�U�,�K�)=c��Y�4�	�]�,��ß�S�L~�����t�P��z��ϻA[�GbćfO�l��2�D�(�ׇGG\���d���kv1�}^��NĦ���7��Ƌ�+�OѦ�U����7.?���!�]�]����Nn�W#Gچg�5z�7�>O:��r�$�硼����i��&��R�D6������1U�K-�N@Ln�{�6p/B�*m9!9�>ìx9
���c�� :A��C�k�08x=�r�=�����kS��>P���^A��>��B�k���޴�N�T,iP���8�ә3��8+lK�rه�,���㮨�������QA�ZO�k���dt�^r��:�}�h*b�����]��j�f�\)>D<t|�E(�z��k��80�gS]s�
��J�.�FD�&����1p�����j�v5�)������f�g%P�:@b�I����|��Ղ,��z�,%>�\1�H���NvV���iz
���A�iс�� �@�d����EF����13vE������圇=��A� �}q��B��_�����Z�m�p.�v�JS��a�Nc�\_P���E��Y�iz�	�!�\V�"�9+�~��Թ�Y���*������?p���@
Q�0�LB(]�+s�1���1��%G���Ȅ�R�(ui�X��G>��/��'�*��S
J��f"Y�P�b��O�p�x�Rjo�1���%�t-+{��8��T%�0s�I[��Ǜ�3&�ǩ~�˨��Y��>��a�7�|��q̅i]����Ғ���@�y���W��3<{[><����79��]��+zdSPp�MG֖`fl@#���-�ْ5%���I]�X'��u1"���W=f�VٜQ�k���GØi�����솶��,�cQ	aᳱ��}aBdщ����Q�����9.d~|5�p#]�����¸�%�=�}DY�:&�.�Hn��6���&�@l����x����Ǡt��c����6������0<�A��r����������B+�!	����U�o	1�oPҗ��߻/[�U�-����)�_^�8?3]���W�R�c�m��iqƓ�(KŻ�q��#Q�-�!h�f�#
���L���ʆ��գ������@��ŃnhW�܉���2�Uy�G�W[�,m��K��Ir,�8fJA�@N�ӽ`����ɤH��g�C,��X:�&P�v�<Q�=��� =B�JH���1��&��N\��'\Ҭ�5ȳ
�ñԊ����쉗7�Yix��	]�M���XC�f+D
�Q�6���	�d�r)
D��F1�޻�I{�d6�q�!���_��G���N{��l��nY8F����&��'��B�-�jxv�� ��ص�t3�`�2*���B�x���9F�߫�V>3����),z,�y�P�i�����Iq�7�5O���Ÿ��d����s�iR·��J���귪��ү�&�@h*���qa��.�c�� ���ݷ�u�5�A�	�!!����d��\�|�Ecx�W+��Ӯ�1Q��Z?���+L��i�����.J����c���G�6-�`sj2��7c�4�ʒc-V8�x>C}�pN�ߠ|�[��-֞8C-���M�e͍�c�"9��V��}t��U|�?i;H���V[ѫtu��U��]�cծ�侻i�WA�9��J���I~�3"��צ:&_r��	,jr6�)�:�(��m��� G�}�%l����0Е�nb��y݊^��5w�ڻ%	�$��DW��Oœ/��L�U�k�O;�T�s#�qZ�G���\e���*��*��A"eE�-h*#��ⴰF�e���}w��bA�h�Je���F��"v;�/<r�r1�!<������I��S��y�B��6�t�cĵ1��z�yQ��0�Ay��	V��v����n�8���?X�ʮe:[�����E�ɮ����d$ھ�Di���������[$������!n�~*�@���ˬi�n���h&�]b[cI�� �^0��hץo���T#7����ovN����k0��y�ݟ��bL�!Gx v��������7�-����1%�R�c��?6@ \����k��e�u4�wC��A`/q׉�S��dȈ�URѵ��"�A��y�ّ��ߤj�5��Yb	T^\�!KXׯ�X|RF4�9��n�{�Ɓ�V�ʁ�(W<���[/��:
�++�x��x�0oB��t\�(212�����X�_&��ղ@*�Yټ*)����^��sJ�m9�
��v��G��N���aC:آLMBY��Y j6O|�-tke����(y��60�����r����Y~saRX�׋�!�h�j���y�Z�<��lQ��.�
0�s�է���6
]Z4Edu6�MzsZ����☪H��d��7� �m������k�Pg����.�I�@Íez-a���e�h�9���k�����&���O��uz��Yt����'�@���\��u�H�r��P9Ù���=ƮҪ:��"}!�4�!�Ta�(�������1��P_�>�ˊ����h��9b�����>�WR�2!�M!��ϔd7BaőV�/���7q3�mc�L��I����)F	!p�%��s�KBx'��d�iv0>�s�"���������f��_N�A���e=�����蝬ӷ,.�?�\�h\�t
Cw ��q�hj�&|�놪׷���S����[�����_C�i���i�r�[#���"TȋR������T�Q3H����P�!V��u3H6���cD0�SBa��Cp��n�:N�2�7]W��z���R�pA���c�����\��r���x�G�Ʞ��nI>L4u�YY���ތyd����0r�x�0�R�a���S%�Na)̒W���7ȝu���+㉁7(܈z-��W�_��"���E��U��ZE���ú�mLp��j���츍Ȱ�3k:/�$2%Ư��0k� _����D����!��s`�#G2k[cl^��V�g�Gύ 8�F$�8��l���a%Y0I�4Ȱ!��!�I��nJ'�&���ķ �5=��y��x��Ӆ4#��L�<kK��9m�rީ�uK�ҮŔϣ�Ӭ�B�����-[`l�-����q\�h��`"�6�1	�Z���E]�DŎ<-�����W}ܜ�Y�[�z�4���E��5�Ph�� ��_��^YD�g ���8���y��~��n �$f���R6��UֹV���y��:t,��!{M�`>��\q��q�6�:��z���ڲӭ��s�;X.���%j�:�&�0�����BC��� 97#�.��r��0�E�cN�\~��{��	�&#G�� b�z�%�Lb�ے�v6,z�^BQ)f��HN27��H.1N:
-~l���mu��+Y��|'�/:\'"������&��V����WƸ��`)b���H��]�3���D�Ǎ�6ч�F\����˹�<�2NrVT	iB���8.�$Ƚ��nKa[�'���b�!�W<�r������hr����~��$
7�Wmi����W1vn�a]&6��3����H�d,V2k�^���&7�X������XzG/._C`V,wm-�;��i�F`�`�PEo]V�!fB�'��Y��߼	x���n
���@�h��X�Q����r~�m*�����&tr�a��)!�/j�9YTR(��(� Ơ�FEw��LK��*���֯邨�S�"cC���β&�>�U�
��MԒ�C���.d�R�٢�&���c+gc,$�g;�����H]�.�Vt-:��*V�XczFǆ�̽ʸ��]���0�&d8���֧��`(<M+�6�yx���HnH8��������R䩐��H�,%eM!�����k+����B��ޫz���;V��6��5�C��l�$��PM�gB�����'�w5<.u2��%��5������	�M�	��`Jҫ����`����j ��;fȢ0�:Nry3����)� �EȨ^�Dn&�sV�h�#�3���`�E���W$�] ��,���`XiRl��Q����s���p?}<!�)*�����}�3�G�%H�D��[�0q�?@�.��Z�Ktڜ&5D��6f�='O#4pβ��Jf����z�IKF���u 9�=��Iv+H�D'Z};�4��;�%�bL1퐷�b�,枹�M��|�9��2���Uգ��W�'�Q�%������/��0j�^k�9����?+���:��b$�\�^�썶!$/��s�_�ޯ�4�J@R��������k%��2�����RP�>VCi#+s�5UU���A���y�Eü�٨x~���t���N[�hT����_�}x:~HD_�E�᮫G Be"�� ̇�GϝNOx*����-�5`���QY��?!�歐8C��K�%����<K���I��tg�CkQU�wI���o���('����#��|@��[��qu�|U�����r�XFgS�MO��3D���JS��v7@?rؑQ}�Rz[��yY{>?��f곀��՛e`!���h�D4m��Γ?�~ы�����~��@1�{�0�r��X�_w����B���!�$�o�k��m+�Ǯ"W@�!��KU�#t��0�2,m�e�nRZN���>,�Lo�D���C>9Zv1�=0֣Izj��k$V ����S�ԃʢ�.����tX����`�i�����^�RZ=bMbD�$�L��W�7v��b�</�7W�0�kp�HDќ%m�]��e;:Y��e����uM�����v���u�U�}��k���wDH���~;�I=���WլKcEm<�s�*���P�S��hԃx��?�懋�D��5 �C�Tmc�kI���1A	4��]����^,;oު)&)�H����T�u���G�m���AEs��nd�M������-�����ɧM��e'�^���.��"7���؋,�߁9ٳtA�p�mY�[�;_�(��p��%Rb�)'�7�GF�������DĮH��κuOF2P0< �$��͠iZ�K�P��lG^�z�m�ռU<B�R.rW�����VOC����v��bI5�iW;0�p���G6fs��t�]s�$5�/�[8�h�v�!N�4���&Qh$�(�����`с�8�%=�b�!����!�ʬ��pa(��i�?<Dc�3Ex��O�M��'�ɍi�ӱt���|D��E�p�=�֠{��b��ܓ��ll7�g��ʕ$B�r5����0�M��©ߞ�Z�Υ���ΐ��MZŸ�/")ȧ��F�j�ֆ�t�\W�	����~r
��ڑ+{lx<Jh7��y�;0@S��Cc�6Lx2��@�7{5�J1���:��ݓ�ն��W>@����G|�W�d�;�{�	��	�M R���k�8����c��-~�qG�=%?�\���[J��{�Q�y踲X�G[i|����r/U��z�U~��ލ��}��@�Eg�GRĘ@G�5��ɕ�"���]���[���^�KF>�e%+�䣰��"�q�p`���9�R��ʟ�'}��`�`�G*�3�|U�;�\�P<o�$z@"x�5ͱ�|���X��z���;�Xދ7��nw�eʫ�m}���^�~����UD`S�{��Sz�E�[�.ß�%r�p:�A=�F
bp�v�+@Mj�E�F��X6�����ZTO�k	;����y5�$�h�A5`�s7j��%��]����3�}���ȡ+#�nƤ6�_t?�Ё��W�_�H:�AjaU�z}���Ϥ})�!)��C2�?b���^N��bƑ�h�c�L�����n���+���I����J̸Z�}Xx��Rݘ���OL���2Vb	�Ui��)�c�V�&��*;���΁ư/JD�e�W�?�6P�v�O2R��(��G:�z�h�7�{g�,�O������G��~Y世ʒ��a�>�;0-<��k�'��m�] �T�>�U�Ёs�w�Kd��e���-oG�E_�3�ȫ?�OCͥ�����v�(��NG}�������!��y��ٵ���X�G�:.����u=��HK�����1Kޔ�s���Tk��姁�}_�{"�Cq�@
�E
�`��'�#�&1J�����n{�n�L		�c#nYn�V��cﹱ��4����:����<p!A!(Y�O�j���L)h�nAK_H����4��r�f&�Yg�B��£xI��N%fu�k`�'��i(��V0él�V��>JL3 h�����D�U89%��T���U�a�|F�򅯲˙��1t�ƺ���$�Ά�|$��g�ܭ'�Ǽ��lo&���/�!@th�盙�a���A�s��W�d���^{pu��Yb����l�5�^
ŀ
X���~W�%�����1-�U��O$3��� �I|ozjVHBO��Y��"�0<E�g��46�	����uV��}l�+�j�cOp�һ6{ݚ�7�{z��~D�:�.2�����K��yq�@vV����p�k���@�@��taLm>u4r��xSvj�=cAbqA��P���W'cc[Uȧ�AZ(H��~n6-�(�yS3(�ձD��X��H���D"����#
����L�]��n��H趞������n>J��������4��n�Q�;�va�Ka�D`� L|�n���b!O�hdd�5������J,J�����A混�^�P��"-ʌ@��G�G"-���v��Ʋ,�u^_���_��E��@F�	��� p;U����J.�����t��������A����G�i�9�hɈ{T�6�)B���T^_��WW�4ܸ�`RY �>4�p=0�_}�<:�W�[��l0/��+�cܶ+�I���-�;��۶�`�I%6�@�/�/�\�pgUD�pÙ�9��joOSNӲ�a8���y�U�R�]8�(��>mEV�˧5��[ ��� ���:抝��OG;#j��@�@�p���:�\�A��Z�~��j@���{]ОO�5Wj3'Xg���������@�1�Pv�B��µ��i�e�:��5���$����v��>�7�����P-~`aX���;��@�:��q�a?yS�ȉ2ۓٙzϕ�r��tƨ�u���[�r�F�+e��N�Є��WЛUkF�A�5�wȉ�WֱY0���cTU�|5��U����3�\3Z�1V6����^JV����<�ab=D\L�������,�gc8)�L�s���{�j��w�˗_�Z���� �jX���M����syyq"g�؜�1� �瀒�F����� A�n[�%�g���R��,f�,g��8l���f	C�����!9P+O�{�kg�Őo|��f,�YW����>ԛ�
j3)Ǐ�0������u�4rw{#��/�\���e���p��y��c��y9;?a�!Y�2h�s̦�{�׾}�V�zۗ/�b��'�gs���A�1w�q?ڄl�-1wM��8^�����# ��w��#��g_��,kC�h���>z�u+��K��>�󾾸T�l��;gB�����!8��,�oC�ʊa��(���0'� q�BՂ���6\�"�`�ZJ���vw���b:�S�� �R�h����ŵ\_��]��9�w��ӹ���Gk+���x!?��Od�v��G�³�
�
^��rŭ���7���c��$v��iF
eS纆>{�R~���x�	���|9Pkր{�Pۅ�G�}��Ƒ��
,��X��l�PF�(���(s�>	l�Y$�MKR�R��n��g�E@�Emc���&�2(Xj;�Z�������w��֤��X-"���w���9r���j���8.y���O���G�	m�|�!b��B�]��Lc���A����tg���#Y#����hZ��K5���v��5dJ�ܺ���M/.���;2��8��<2��@�����s}��.n����D��7��g�}��)C��C)�2��u�5 T�}3u�tani���ۡ[�zK&�dz�V
�
����@p��EΪ޴w�_���[=���$0�>��£V�3X5dg��}^"2<���Cޏ=K+e>
�\���&Nu!��߯^��@~����b��/����%�u
����|؎��uD��7���n%��G�AeI�$����ޮf���7�˟�\A�b�K3L8->[�{�0���؎8�aS� ơV��E�0<y�P���Z���0T53�$�ٲT��C��0t�${!�����+z��i��!�dSJ
��c��^�m�V�C�V�lfrhA�\.���F�LJ���̬����A�0�&T�%(+�Ѕ���q:���r5ГQ)�'����zs9�,׋>��>����K�p�f��Yx�m];��a�B�&�[l�����V��:�u�l�c�����.S9���	����Y��Grrz"ejM�c�p�RrGfvD1qo(#�C�����Pk��*S<`0��S2}~�-�^k����;J#�=X���+����� |���H����b�_���m}c�Xat̐:��4���@��iԈf��\&�)#Poաe	R����ghB��Td�'�<֟sn�"�=e�9���x-�f��,�
�-�zEq[��
*�Q��z��=��40z�N�3��FJ,C���P��p?�#�{7���;u�d��9Z]����.��.x�b-p�%�M�OK��ɧ�>$��9�"S>C"ւ�����!�E����ñ��x��^��~-痧trp��d��vA����c���[*��������z��ѧd��@Gq!t��Et�*��Aj�A 0zy����E�����γ=C���L)i�'�u���r���P���X���Bk1�D�,W;٬?r�(����9��Ȅw
�s��Qf4�Q�D:�
tB�2��D��#H(e�X��v[�a�:<�M`�J>>=��~.ˇ��kn7{x��$�A��1�g����F����&̠�X��M��{�J�Ņ��IJ����-�+���,��:��f���J^( _�\ȏ��^��(�AM	4���5���cNF��ݦfȿs�H�qؗ%�ZS�u:�żv����}hb�"������&/�
A�
�J�-��Z���Ҍ0�;��5��S2eJ�]y��z&�;X  �������)�M���K��l�y�B~�/�\_�P*�S�L�跺жd1Xlӑ-�qn�E����Y�5ƣ)���b%�w�:�7tP���gz:����p`?(����=k� B�A�b���K�0���5�������#̖�5C� 52�����W�����KS����_���5�p��Q.F����s��md��NY�
n�=h0�ʀ��F#�T��p_>�+��S��L�L=��21��7��ulw�+��-��J���@�!���[��X�^�˺ޱ�ߜ!�,���:յs��� ׯ^�� 8l6�DUHG�-��2�[��BDӞWo�`c��A��0��l����Ϩ���͋�@�=hk�ґc��ةDX4	��
y�� �CGB�r���Ш�!�V�~�������g���IH�Bҁ����ղۿ���q�S���?4L:f�" ��j:��u bi(D8{SkYK]�����ěp:���/�Ky��;��Ws:ܸ������C��c�{,l�49�q=��d�,�[H(��B�֩$ϙm^b�y/u�1'Ԇ�]V"?���L�*�Vt0�n)M�����p����u�l�X'I9!�d8Ԯ�@�z�޾�(��'Y?����)|����Cn��<���p��9�4tX2�%�Vm��栤��u<W쀄��6� /��N2_�~����Jp]�5*?~�9+���!*��Ll�iq�:����P�Nf(��Dd쐕��ˊ�,$����Pg��?�����?�3�:*��e�,��̉[�56X`^%t�)ʰM"r)ȵ����i�?_�3����^W�K��� �Hj9.����zܐ���v/iC����gS�DIy`G�vI�Zq6u��,���J]g�3�W'
�������ׯ�͛W� ʁ���|�L�Q#��/_�O�5`" rp:5ȩ��;� <�}��&��@�����V��[ș���YfWr�)C���
�9Ǵ���~P@}R�s+�e D�Uj��!���`�^�:լ�Np�-��GP��9mu������G���  h]!�^7X�":��zo3������K��
!�[�H�
���L�!΄C�%>D��&{cƘ?<](���x7�Tכ}Dɓ�����:�*�M��.n��x/�����K��qM�� �X6���{KpE�![Ȑ�������LǬ�0N�v��#���F�!��T{Կ`� ��>�E����uM�������Z�@�������F��S����ø'H-���ي׹ �6)@t@�M: 0B#WV��M�^5j_|�#qo~B��_��_�J	�m��Oe�cB�����8ο&I�	�����㽅�$�f���M����F��=�xE"��F��[W�o�́mEt��Z�˿��/��/^��}��W`T� *�:pc��2{����%+V�K��޿c�sߥMP�[�ǣ�X�b�:�c�c\��]�@�+?���u��GF;�c� y��y���4:�F�z��n�"��8���>����!>�s�H�Ij���X�e��gS�v�>(����6<`�Ibpj>�I`Z�O��4�hϒJfj���B�*�AI/J��Js4�ʫןq������7�N�ʓ5��T��P��ȅ�����r�(xSc[8�o�=Y�!O��F&��m�:�%M��^�1?��}�}��E��b�Õ:��0�a(
�'�m�:�ء�6�p���$�X�*���ϡ�#� 5�%�5�uWB*7[�}ǲ��8_$D�����"�[���oC	G`�u�J�����X� Ǚ�%�f�s.���齝�seR��"5É��!
j0ȑ���?Q�$�̆N���lt��m{��F]%a����5���}n6=��L�~E�N�7?��,u0��@�:?A��!Z*����{���>����4kۺ�i���
1��ķ"-���>��T�`�gj�`����M:�<���\{밻��i�\x/c�n���ӑb?a��ͮU�K�0�.�r��3��O�탽Ŧ&�����Eqj_n���5%�0�N`=�`Ajl���[��|ʶ�'�l��:T��1V<����%��W��D�6r���� (t�vv�V,K!$�\>Do�h�:�g�
�:Ok�u���w�N��v�������ڙÉ���&�a��̕��k6 ��{kF�0�32�F�c���_����������ޟ7m �_���+�|
6���#�F�_��Sd�a����G��w^񳏙u�덟��=��yІf��?jH|��
s
���Ib�8FP��D��`}���:b�
������ l|T����/e��H'�7��3~J�!�=�f-I�|����0��ݷ�5�ɚ��L��+}�N��/)k�1������V&�5lwKy��r�����H~r�O��ҷ4j���Z���z04tz���P���\A���M���������t�C5I�h�Y��	IBR�3�zst�Ø@��il���t�.h����eO;�	C�R ���ۏ�R�7��;s�+T��e~{����D��PY�A�YZ� �%�Sc����!���g�Z�z�1�&0���K�SC����پ���?>Ƚ^��C)|����D�~w,��l�-�� �Y�0UEP�(eڱm^b�����[�n56�zɼ�X�W���6�:^�mބ�X��CKϞ�-q����;)�����<�-�X��e�[��[�:j��w�����`�7��.��B=D��F�O[���B�leZ�^��s�ٶh��?(K4ʜ��B*WQ�0���dzv)Y9����|x� WWjfgJ�mW�]�N��I^�w�A��݋���%)E���|��8U���0$�*����D��_^�ۛ��_�U��c���o����	�)��iݱc�6��Kq���s��/��8�1E�eヘ�"#��|:�Ym1v�2�齮�wO�$���T�^���I���y2Q6�5f��w��F�a�!sk�b������m�����7�H�@��_��D�B��lu�>�#�� ��ܺ���Wz�P��9DW,SbG��B(�m^�w,�v����}�qΟ]������z͊
�*��ȶ������k�m`����������������6,�ĺ�|@9!�T�����\ǆը�:ĦK�!"'Q�������j �m=�����q���P�x\��cp=�S��@�-#w�ׁ�l0��db�G�&%	�T��}!��1����V�vB6[����S���d�?����X?�#w�V�~����7߾��x��P\(��k3Y�k�+��c�~_��:�Y6lG�������C�<�����A�O���0W�3�p���(�7oe��e�&l�v<+��}-�e-�>��˫+���`w��ţz%j4�������ԡ'��EM�J���j@0�I���3�d�>��T�;���/h@�`���Ã��[q%kX����X�v�{�'/&(�����@���1|ۆ:h��Z����c�{%�&ƀ�SA�MFF''l��;�/�B��1E�0�6"�AmC?l��֥)a.9	N]��%4�Ol����6�G9��cr7����`?��
�������/T�!SdZlc�$�������S�~��ދ5q�5�7(l�j�X���
���C����{K�A���iDv(g��;�
������t<GaЙa7���&,·��\8_9(��ЇeGp�Ɉ��N��[]�\ț7o��յ,�-Î�OM��� {,�����5�en�0�P 7/�J8���c��߼�����^�Z(�v6w��L�;@!��t<G���9��611Kl�	��^Z����+3U-�jXl�Z*��s�[��F�:��T�*s{�z���`/�hT����R qG�F��Qf!b�;���b�t�w�r�`m3}�s�i�	Zd�DN�	8'κT�z#ద;da
(h��iBG�����D�w9�%W#���~��v�T���ק&|��w����?<�V�p���q@�%�韞�������ku�f��&t&p��q�e��~bTV������g��齚LӰa��+�)pJ,R��oǹ۸n�z��v�����1�m��������c�G���Ci�
��ވJ��)�\]�����;�w�&�+�٢�7�)�u�������쪸j
`�� ���s�����NN�c\���d*#�78�DyN�3J�w_�t~�y�cr��� �zS��*��oe��7 ����-�Xw�p.Z᥶~�(]�q����E��yb@t��7h`�ۭe=)�{�� �*a� \2����B���~���Y���w\8X0�d��P%�:
����'t��Vz�.��7/�SN�>�z��S��.g�RP���~���X�F�^lr��Ęx�P޼Etm:n��zGg��b��'��, 
0?���\l�^��8�ӱ�}��ono����6���
��Pl�t���e@�!'Ǟ�YP�b�����a&&�kp���i0:2���J�4�n���/��a8�-�߷��&�r�mgM٭�ZLBۆj���`��D�!�N��<bg�|eq�X$�j����1�w�[Rh�H� ��)��(���.<Y٭P����W�z�=�s����O��g>�W~��׬7������ٿ+��S#�����z�l���% 4At �i8P��:w!�C���ým����
�6�5�����ؼ"��tSSK�aE.��؃2��1�N3��l0�6r�XCȧa�ݰ-�5p4a!C���$�M(j�z>O+��QO�p~g�`�<��ש:��&��E&��:su�D���o���r�(�Co�f�3�.&�,B��6�v�����Ou(0\�H��#�~&�}14�B��a����z"��l,\�Vm���YA���_q����O���}��'��|�ϗ�p�$��L6��n��h[��R�%�~�߸��-KmͶ!�L�M�=�M�OEW>�5�|�͡s���{�6���>~fz�ݱ��uM����wAc���Hk~�y>>3G���ɔyv����d�����,Wҿ�F����/t��B?ь��$�U;	!%��F���/���BN..��ťEu��g'����9�>��L��Ax�\9e9){sK��̴VC�R�pq�Z&I���Qf
z_��3�ԉ͜M�Cc���Xą�\nh�N����I������m+w�(�f�K�5@*K����9�<[o�Q�'(Sf{�
J��H���%<U�ZV߾�T�*���vz!Ԝ���d-6����k�;��]!j0�F� �b3:g�T�2c�}�X�wQ��J������}~���|�d�������� �]��6%��x{��F��Z�#3p�r8SU�Rս}�z���/ү���?�ͤn��ΐ#��I�CD���v�Yj3�2���<$<����Z�F��f�������{˾���9| ����f���r3S�כ�����?ې�k,��NB��� �u�`��[�&	��{�=k{���@I:��{$\zSɍ8�8�j_"wM���S�aD�~٢;=!(����1^�wRyM`��Ӌ*�{�Z��10�F�)�Twx��g���J#K�F�O�TI��g�������R�e���1@S�zg!���u��9��Y��n-� o3�1-�M��ݛaO
�O8�{ws+$U# H�Iz��Q�h-� �{�����>�
N?Ju:������B��ܞ���u�z��*ߙ tUV4�Fm��?� \x3�M��i����>'�n��L#%��r�瑐A�3�$�f���	ƨ�#�U#���T(���{����P�|��u�P	�B���	��pѠ����*���mO���A�����cX�kj<{���R�OP�zF�<n�gh*�v�>��y˯�tg����v�ono��ew��.+�lW6h��$�UQ�f�`(��F� �������lV�Z��[j�N����Ktt�ٗ=�����<���Z�X�N#t��D��M;/-���?�[x��g���T�h��>ƅM$ SE��q���S���}X�||�`� �}���>�9��]��٢�W%A���ڽ���U?<��O�:��o�}�b�����X�����>�T����� EIR5��]or7\�c]%�8�z>Z�h�dzo���c*K�A
�L��$��W��w�,5�5Z���e;��R���96s:Lʉ G'�� �0��;�=�m���/l#/](ڲ墳_U����K@�h�8�sT!A�}�Dc�*T����Psb�I�XQ)*�dRв����:���xSi����J�4y�~
�|7vЯ��C	Č@r{�g�"a��>qB�E��٥S�I2�0eQ�DҔ��N��(��ë�~ @q������� ����JNb�?�y���B@0F9X�TrD���e�v���3z�<0J|&�=׈���4��~����T_>����|��ѤU�i��d+T5��J�q�QHdA|���m=��P���9��'�A:���	j��
В�i�3g��ə�:����c3P0�-]&T��"�=�I	�D���dͩ|N�+�;�;�r�dʦ;��2>M,��;�}t=\G��^��lG�44;�����\\�m�h�fj�����[�SӲ��d�cɞ� )�	�s$��[�3����$�K��;�nhjK� ��W�R�:U��(	#�{U���9W����"8)H�t�"T/���D�41�)�X1�02�ݞ�h��
����u&������{
�3#f2�P�2�b��®��������X8���Gsʣ03ak0@�
U�u-6/��ݣe QV���A�f�=p�pqo�<��U^�����۠*w���S~�N����K2�����������p���⩢X@�������/j�|"�,���u��>���\ڮ������L؄�W��^�c�m�2ݎ������5�����AB�z:fci����鮇�9�/;�掆vW�cf��Z��
�=P���!|���p�����6����	�ꉣ��S��f��<؇$2���~%�^�)���d <���,� �a�V���X��R^;���\3�z�jn��(
�V�r4����O-��~�PYc��'"�R��Γ��GRwQ�K�خD"1�=]�����o�žb-#_���,���  �h$⨐9�Y�<��0�|xt;��/,Ki;_�ЮՋ"�t�1χѧ�ѝ�
@���� �dv��M�P�58�,3�5��Z���y��@��F$���ݣę, I���I�!��E:���+8�����Xe���e8��A>8I@o2Ɩ#�AB��A8yy���N�(������~0�Ms^��V�W��\�a��̳���d�j�1��o�����T�d%���{��Ə����t$Os9�>fD���'�,5�Wqaey�q��ӣ0/��"��}��x��i�0�A��	p�BqKj��x�w��ï��>����"m"��_L���d֔~d�3��5�jY@c�7��=���$��*Vx�k���������9�ޮ�,��Y�x�}Q}�%�$��PP�`�?ص=N"4�x쎪�#OA)��R��7����^'dA��gHt�E��Ŷ�=<dX�Ah��g��[�������� ��_�. L�
�!����^�z�vŏL e�i/h�!\�߇��G{�;�AM�q7�tb:���h�v��}��{�j΂k�ظ��Ƭ�e�kmیV8�����Xʄ��'Sf�%g�v��]�~�C��Ke��H�X���~�4h�q�����	I�	�����p��M�;S]�9>���lcܧo��h��������f��)���k	�>m�}*X�
U�h��(�[��w»��u+/�e=��#�z���S����"Lw����}m�Ug%�(�8�U�p(g88F̡�+�`)�eљ�9zq�$�+�0�^���7��.	�κ�����vA���	*Ȧ��);TM _�ٙ��"����Ύ,���tS�p�����l������{���m�ٌ��W��á���Z��9�UR��J��|�FhX��AKE��x�����_}�m��=����=�fj�'m�:e'��'��4��XQ��������2�f�u��H�Ԯ�!�X�m�6kN�C�R=�x�xQ�����s��q:����'Zz�J݃�9s=���+J��ζ%k{�u�,���A�n�X=�w7�ֲ���[�w��/��"�V���>��q6 �[�*��+�G
��Հ*�e&��� �Eל�J��|mYv5���H�^�և2w��W��uZ&��KA'jID��ؓ��t�K�.	�� �!�/�!�ȅ�],������o�������GH�(�5��,�h�����Z+���Xr����\���uP������2:s���Z�7��-%�q�ӵz	��F3 �L��t���텽ݣ����2�=�|�'���Q��e�2`C��XT�҂��`G��*Z2��I�4�^d����f�?P@#]���LSr<��R�0��8aJ�cF��A0N�*7YvR_�з�{���G���ʲVJ�RV[�d���9�������peA����-�y��TN��q���z�sU6�Ւ� ��@��+�)b>��4b�G"�y��������~��};�V�s�9M=l�(��|���G�Nt��F��vBc'�j�Oo�(6iL�)Di�����5uqm�SCX�,�1+�Y�Em
�7�VCx��˥+mUT~��څm�9P��^�T�D秬꿃�u��<�&�$������l2�������o�03C��p}x^�2/�A�TC9GG�>�� �0'�g{�e!# �bib���ޓ���b���f��;XZ�׻�£�<��
5��E�͝q��^�Mxt4�P�A$/�_���S� ���K�N$CTy=�QE�@yZ$�G	��b�)���eh��D��~����� y���0����cs�{B�Hٴ�P�|s�04��Zx���76 7@l�N���ZI.t̀[���Vd�G��?��n�o��Vs���e�yܦ:��,��gI��vD�f�kEݕ�X2_E�9C�Z�V>�ۙ���{� {Q����\�����<�̱Y�a{n`�W���(��+�F�ío�- k*�ڽo��g�ܢ]^SABQ��J��J��.�eSFqa�&�e�r��Hvx!�(@�[��{vvN�4����nB�}��ޅ�Ҳ�L>CM�'��0mu�sQ�t��'ar��hiF9)@w�h�9�ؾ�}�������Č�BU��������`�;D ���(�����ɞ�Q�|����DԖu�U ��`��,�ݨ�vs���)ޗ:ɑ���X����IX���6�~T�	���pg�2ɵ�A�G��k��k���u�Q���s�.�
g[��@0��{��ٿe�c��0�I�|�3��`-H[*]KB�p�d͍A!���6{��޽�2U���qE4�pG������>����ewbp�~vaj{�ͩ>��@�rgӊ�+�6C)Q%�j3NԌ��^!�6�g���B��o;�/��I_�����_:�m��I<���	�V�8��,��ڙ6��|�GI0*Q	�����b�Ι �W&B�D�HN�
k����R V�X�o�Q�"��D[���V��>��N��������9iŚ~I#qZօÉL���-%�cƣm%=��Mv`wzmV���O�J�/���pR	���%�t�Q�Hʟ{o�B���7��e6�)�Ǌ�����[�fhj�������٫�9W�c���ڮ-�̝�dv�C�;f9�^S�����L"v3�U��@���]vaj�����T�L�Μs^e���Q���l��*J��g �j�����*Ef� f"�g�����q۱�ke�����
�P�l'9bJ���E|4G�
Nͧ������� ���@��@7V�N�H{i�Ɓ`CS^":�\ѐԫx(��#��	g-�Z��A��:��j�o+�A�"�4	��Xٸe�׌�������lF�<�,t��C��0ǘ�k3^����D8��"��u!0��=�L��&z����TaT�ʪg0孬���	Mŋz�2���R�	%��h�_�����A�>��]�!�� hn�*��q͛�e왱�`�-�[6��T�,{���W���E�m!֓i���H��Y��U`�߷��Iۡ��?�Q����U����~3������`k�5E���-'�OT������!+g�y�)�8E؀0��;;=8s��,h��}\[�����,�{C��3�E�fE)A����qo޾G{�a�3�;;a���'�&;'�Z��!^g����V��|VeöO���}���zaA/�Q�O�>�gx���/U]��u?��=�X�7���vMd[T!Ԯ�HU��l��}.�y���Ѝ�J�IMil��ɇ�vSh���a,h͖�<'2��� 
��2��9�L>1����m#M&����2��DI�F�ܰ��1�U���8(�m�c��\�N�ї���6�%4���z^������١o��U������n@�*~����	�	(�آ���A:��.b8"�o�G^��������݁|C���R���L8�BYt��=�������e������,����W��9\b�	�P�ǈ�	��>�仯�SI�r3��˪��/V,��W�ی�t:���x�M��*�$}�G �68�w�g$��1�ą���3��x�����#̓�7��_P���_��ӓ�]]���@C��Ő"�ilY�(T�)�bdCIo��������~�駰��#��	-[9A�h3WJ�PE�:#����=I��c����w�i��YɄ톢���T��d�C��ss@�rPEX�0��2C�k��Dq�0����f���f�1�:4�gj�
N۞�>.ë�_`��{��������<���]�^�ZЌ!�����bD�(��A��C�rvS�s�@��vm�������[f4��KG��F㐙C�!���d"�Z�D���XG#��t
�0�]7Ų6�.D A	�n��R�K˘f8��l�u�%����vw�����ك8�K�Oߩ�bc�xJɎY�8��mա����˰��G��.ȸFc1U&���p�ƾ�� �]/���C)�/�=������ؕ9�c�=%	�F2�%�0��!=OHl�P8K�Ϭ.�<ٙ�����|vo���ݍ�D{ʪk�������dg2�^�/O_�- 	.
���������ugd��3j�#�}���W�#�߿W�Ү��_���/¾}ֵ(	����æ�Y��n.���%#|�Hf��Q��φ1*w^u�N{gӫǦ��q�tU���L|�#�	!�$�'�]F|�x�	�vjo-�ߺ��.��oKv�Y.}�S��������A�2U/S?;F}����ʄ7Է��f�C��5�Y��ؒ���	f�(��F]k��gQծp<K#�{k�H��a�U��&դ��{����ᖲ3,I�针U�W���d��C"e׻n�_4����yXv2�8��0u�z5hִPfG������>��ڽ�������P��ե9���A��*j����5�`4�P���^9�nfH�d���e�"F[8a}_JF|�m�qb<uY9�YK�NK�@�G�LpAײ��9:4U,�X����m��Y����^��W��pa7�,s��8BGY���ʲq�UD�
Ӝ��oxe�eY��EX�܆�FG,2�ol�f�K�d@EO��.�|\��o���!I���2���g�.o�G;�fNGz-���yJ���7����|7��!�̰؃�V���=�Ge��*�g���5��uP#��f�#�ej��Z�u{B��(I3o;��z��裙s�0�� 	�8<�A���-��C˼>bh�E�\p��Eaf�����#ڳv�&��D���Է\Ę3�!�.��N3�7Ͼ�e�r�:�^Vt��.�9�4wlǾaD�Svcz�\��*3�Yp[��P���#�`��0������2P�����QԻ��͸���c�K�������j:���|�k`T� ���>��j~߲J�:�)'O9dj�Nd�c;�Sw>~�D�89x�BP;�Ӗ4hU��8�-����*x��}��	����'��{{���똙�pB��[;.�L�L�*�������Y�֮g�]a|i����A�4{���l���w�D9KB��+������)�ڱ_&r�h��U�9 ��q��|���џ�1Fq��shK�� h��.PjJ�Z��"�[��2:g�h^~�m~��Ϝ�v���i�,[�rfX6}�9�g3�_:�d��!{֚Gށu$W���x��OVh<M��g�Y�κ'1Ӧ�q-�_gA$�cP�
���ch�ۢ���k��
'T�YU��/G��yfIG��<B�b*O|#B�%� �_(��2��m.�S�&�=g/�UU�ޏ�(���Ko�c�;g�������3�y.5>S��������~{t���b�ΰ=e5И�2>B�W����؎<���um5F�Ъ"�pg�X�����:������ݻ7af��]CRvv���e1�0�8-nv10��46�	�G�lx`�3D2�Q�8Bt֎%�¥���G�R �QE F:(�qfI6��K�cFqjH�C<O�#���7jG-/�kjـ}�N��@	���Ht��8������̛T&�͐o�������T�[:;Z:�i[�9�DT=�+4��0_t�lf�ԛ������24�k�q�-� q7� �Yx��Isx�:�2�jy,�=o�҅l��Z(���9�����5^/#������Q	!�-��Ubt�
�;v i���C~u��o��R�3SX��&QQ��p���f,�һF�-	����&!���0�<��#`�K~�q������ٵFӰ�§�H���=<��E�ĐQ��=�s������z�S��po?�-hI�EB��p_V��q�݅9�Oח������w��f���Rk�,(SS+΢�s 
g�DA+����֫%���^�
���&�f��W�fR�"��a���#��ڳ&)^�Jt�ij`�oԵ(w*��0[]T�O�")�P�r��<~�y��K٪�NE��U��;];��{{[�2:���I/r��Ά�~��e�[��%F�Ϝ붓��#O�eC����~_>��%���icW���pf+��ת������%a���-�s U�@�B
�Q3���&Z��*~$m��x�R��Z�d���%�m�G������Q��>N8����b�tQ�!�<!���
`���B]z��v)}�](�Ț*�fu�P�ax��2�԰�1XO��n �B��%&�\V1j�n^싨��YTi	����u��� @�� >�_B0y�%�&n+EF/1��'9J����I�ֵÌT"%,�2 �{��e�w��J��sQ�S1� �=���s�6��$z�Ͱ��6���g*�8W�?���1׋qiwʍ@?#��k9���u0ՌMgC�����(/¿�1gm���9N�/ކi�*%2: sSy*D>�h����N�?�#�kQ���k�eN���PH��\�uR�NՏL�;i�`�-�!0�sx���8J�)[Ks5���5
p�l���^Y��j�Y��p ]<�I0�LE�Ӎ�E�+�+0z;��e�tw ����Q�پv �f�A����c��8d���M��,�-���o���Ψ��./8�U�`�N�O��;�]9�YIYӂ�o�Y\��A�ZW�Y���g������y8>��9��QF�o��3��r~�9�)�T,�v ]`���I?=���װsK�xV�(�[/#N�%x6hp�����T�F�o��4-�3d�I���]�+=qMY�y�رτ�`S)i�Q#�v��y�����A�Ƕ�{�3��<cj %�jF����}��y����M=���H�J���h��:b{�5�|��I����5�3\ǲ7�άAB]z ��h@G���y� �7E�R�V�x���7�ή��y6��=��PcUMt�1�L�+�"J��8��;QH]?WlՊ��h¦��&B�Q�(�q]��� �[N�	�̒��;�2��A�E3��<{�`?�O��T��7�3����ރ �v�~������,�����}ݽr��u�9��/|�"'\���j�g�(Z���h�X$�g&=�t3|3���Jo�)���V-��Y�@f��� �_{?$�j2��fi��e�4���8�v�_����=҆֯R/�^��E B�N��!�;}JҖ��{��A�����cv�!��O[:X��=�4�YD(۷k���`��*�PR��Y_!�BjQ?�l���cw����k~�6i��AE�Qd�%�*���9��s��W:1��ǜ �A�����J�d��A{�,'�UZG�ʼ���zD��b3����K��s�"�h 7� 8�Z |Ԉ�Q�U��:�ّ�e��r�v���N��	���,��,�wo��Օ��P>ho_�֭��4��Gfp���`��}�ғG�d�r$�;:9�G�B�Bw�gQ4R��Ž���]!��'���e����\�^�ǖ��L���z��]��-��no����F�iw?tv��	u���iq��=cg~]E��"���%�vtpN��.
�j����`�^��g3&K�՗�̹�l_�m����?��}nz���|�z�G�0����n�A]��k ��N0�5��<G�Si0W����U�6�E2����[R�����ꨣַ}n@g��[@fs����jG�b0�S����	��$���}F@�'L�ǿV�؉:�򹢳��ׄ3���I�YԻ�к�:��w"�����2�lVE2�����]F�]F~�:|�p��lSV��-�ѕ���nn��SF���&'��~[�a��#��}9S����>�J�� ��e�5�}�i4K�:�̞��w����ԊT�O`�BD/�T��b�;O�	�`:Z�}� w�f8/�dZ��T�-W�Z�h�ש����2�(m!+π�ﰮ}��Ч��>���X��T��s��P�����К(�r�WA���/͊1~�� ��y,C+M4�I���y�[�#Q�nu7�z)��>�
��E���#�A�j�n�hRsʉ��^Rό�=ϲ�tvv��O��\˞�	�/އ����oB��)���~o��YIn*%8a��4�g��$��T" ��ȑ`$�Æ$��	#B�+@�ܐSG?��z����xnx2O7���f|(�u4��P���y�?�/^)+:3%�>sR����0���HS� L���0�׊�a��밙�X�w���@�5�|#��!HQrxV��S^W�<��(1w�,���eص�udAV�E��̣x�1�����!<~��!�@��G\����kehdnD�
*�k�\��U��NSH������a8{���ʮ@d���v� �Qҳp���!���!$��Ss��l'�%��J�Q��v��r��p�o�U?֞b�5hRa9�����Y8xq��V�[ ��d�,Cl(�r#D��ϙ����������V��J��'rΡ�%3����ZE���W��l'�o V�~�~|�N篿R  ��1��g�����yؿ��`�k���7߄����C�����pfg��=v��O?� ��>*�l���B�Y���D7�>"H�x�&^��չ���;ـ6����=���������6����Q֨@��ډ9�O�(	���
�d�|�ϳT�A�v$�'xtN�Q����}�L>�(-���	�t��Me��b'��#����������6e������ʖZm�<��3�Cq�G�������u�۽���Y��45�0{�il��z�G�^G�ù*v��Q�8�{�x�PLs�k�ԭZ$1��CQ��so�dè*��۰OÚ9m�9*v������������''�vڣb�^[�2�+�T�l��^�!�'�G�1g2s*�3�wu%�J���r����E"nF�Xl�g.Q��,n���8P���(�H�1E��4���γs���Kg�0��Nx�a�9�*4,���{��W�e6�.l�d<�QZ�>�7��#�g�*1fyU����:��#q&x�J���TŲ���k�{r�(�g �N"�﫼(������)=��'���d2�r�̈����zz1'l�Lh5�F�@�R��]>@�*�?@$�>���q8D�Mx�#1F���[�v��52�"٧2L|��'+����ұ������b�g.F"J|koFK� ��i�)<�A�-�==��w8pI=h	��d�.�'�tw��_hi��Ã�p0ܕA��Md�r��<����(\3�h,K���g�k��	��R�K!����@ڧ�{� 2흝�m ��f0��'B������e�Ex�ؐ�d�3��J��l�ý&[�w��/[]�d���C��	'��8pJ ���^���8�>>�}rz"���Թ��`�'�VQ���H�&�kWt�ʮ1�h$���o�Kx�fl����+`�OBd�K2�4B��D\���"�x�Z��v���<��bVF�  �Ү�������U^���`x@��9�o�IJg"��|�,����N�0�;�<��%��	>7�������k^�Sv�`k�1ld��`^��F�Ҁ�˃���6+}��1{f+�с��zUB/���5��S�#�]Y�F�J�&a��~s���S�������� C����(<��R8�f����V�����ml8JT��m�8�a9� ���O�Q��5vڋi��q�e�IO��ES1�M6\��jC�Mq��a�Q��
?_�߄��Q��;L1*i��#���YXH�X��E ����U�Ā��H�)I�L
CO0�o�K�����XT3���6���e�u!�n�B�2Ľ\�TB��_~�_���w���C��J�4��P9��|���)#2y+a�*�p*�㨋��uT�Q�P�Po���hƍ��w�w�Zr��AK�$�8F����wO�\i�H��"FO��҅'r�e�����y�i��Z\\]jV� FT��'�]�̵y��P�B��&/�<���3ͳ�Z@�0SfK�(*�5e�rg�P)/�|@�Ӱ��[���*����FtZN;`;�P��96����Y�z�X)[���s$f�׶����B�v���J���@(gu(b�*D�SG��14�'! W�AOӭ���?q�y�T�/k�"(��+X��B(��98����99p�a�+*@��+��|!ǀ��cCL����e�)1�¾�5�� �lJ�]<�$�=���I� ���S���̿~�]����ێ����cx{�>��s�WfЖ���p�0<yT@z��ܮ������g��������ʾ��>1�S-sr��Q���	��0htÕe�3{���~߂%�뛷?�D��9n1v�e+#iG�7e�%����)d�L�&���>���1y�
`3�Zz{��mfm��0��/��b6�
F%�j�~����~��Φ�[�@���G��Z��]�Rf��猯��v�=9h����@�rh� #�$!E����P��i |e�؋��Q>b��pg�����H�+[ѡn�<��ڮ�y�<9ֈ��������@�QTU���?Dv��۶�������fo�Uu�/�q��eEu�H����#�	��o��y�U#P��N�l�$�cK�3�oA6�q�����E4��["	��١E�h������EN�i�:pG��gm٦���x&\I4���6�۟�~~�s.+�΃� �N�rL�Qd8>&���xQ�M�D&Ls��ߘ/]�9N�q��p���iwv����o^�C3��?��ǁ��y�se�V��Z� ,ﯮ�[�4�,Rz�6��=܉���������T�֫�R����K����T�&��Ne���Ml�p:�dp�g�d\�?���P٘��G���2�����:gjRVI8A�U�'0�p��N�+�c�uh1q�V�eZ{Z"������ ��/�ۑ��g��^w>�|f�C�t�����Tk9r�0W=5׊�k����Ux����� a�������Fdh
۾�ۤ:s��,}NY���ف�dl���j-cH���j�?P�� YD��m h'�G�G�ҲE�C'��,bo�Q�9E�Ct�����ks ��a�Z2���>\�*�#����վa����u[XVԨ<��$����ah�kU���zk�����!�;�?^������G��gZC��c�Tdw�d�w��!�/3g*�|sw����v��Ë��4�Էk��t��2�A/�-� Cм�}I����T����V�3����D��49㚝f�)c~��/a�8�x���p���狏����UY��XXۂ�Y�Ld4�F�q&؝��k'ʱ�p߼�ßµ}6���ٙWdZ]U�R�^A�����8�a�b⢕�Tҏ|��܂�����8����m�[�
��I;g�O��<|��^���Ǐ.=9�v���Y�I����q��3=�5�)�f�dS^��$��
x��r���X���2�8���a_"����d�$Nm�m0�&��T?�+y�﹢�S$�'���*&��ul�����M��?�6t���{��w��o�������`�~��)4iA�h�P����E�:�8u-�ױJ�p,"{AP����7����eNx-���2�$��:�vĹ�T�,]�`�,��T~��D����=m�"�p<,���}er [� $8n�`d+7��l�qRO`�r���՚�4����S;������W!�aS#�n;�ȴ��Ņ�덒�^"awZNsvy�)��x.�׫�d�fd��h6�>^BE<L��ܬ�j�S�c��uYľ/��vG(�>�����ڝ�Gp��UNK��q�Dh�橳�b㠼ǃ�f����K�8a��gu=ZG:ɤ5+I�TƊ��d		]���R�c�4�5��� �pe9���L�_��,c���������Y(ON4k���F�b�;�j����Q�d�D�iNk�1�]���|{.���,C�z�-���!*�[��߿{'��#y���z��8�����Y�qn]�S��ڋ�ً�|-��KIKvNN����ʜ0��R�Y�5�K� ZQ����r����PA��j��l�u9�?�T ����]�Y07m���i� }j`=���ޛ�F#��S��;�l�/?��_����/�� �>����P�����>��H���������%���S�1�3�۳!��aR�P|ek�o�G��[�g��	����ޞ8�����;f\u��e_�&OR%�d:��YF?����mt"Ǻ}aR��HO�Fu$�X���g��H���^�s[?o�9(�L.��K�X��s�d��c�h`����=>�`?Ae��8��M�@V#sT#�ʫ�\��#�#
#�-�2$���<L��4�J�L�����$(Sf��'�/d�V9�3'm �%,�~��*�25�pUbs�3�-��P�mBO�p�S)�����q�(�ގJ�6���T΄�M��޿�J��[@��z���鐩��Z_�ȼB��.i��f�N�pn1IU��=04e�W��
z���ĞJsD*�f(ʛ/"(k-��+����E������O���P��3�Y�n�D�11�0z|
�_�6���2���m��-꩎�H�	n�"�H�	i	ٺm�1�v�Asɢc�aHB��Y���͛��凰lfg�� e�:����PYtg]�z���KkY�7NR}����"�EwGΖ95]C��^�&~c��-����@K�A�|�7K��"߬�6 b{����o,�ˬ G���	�lR�Ɣ�I��ې���#&C�9Q�84��gA�=���T�a���� s"��F����y]?N�����ѣ^��a����޼{�����)�129�~S���_����s'���:�y�r��݃Pͧ�\���C�f�ub{�1���M���������s8�33�"\	����2��ͽOZ2�X�6��x҂�g���XZ"U�pd4e伎=[�"��|�5�[T��ĕ];,eIf�8���n�w�a�0'�(TPo��M��.z�+˴LN���������xmY�P}�`IZ�Fɜ��n�h(mm�w{C�s�	e,�r�JOB��^�9��GX�9O��{���q��t�z�ڗ
j��+]�>W�%�_�maz�6^F�6횣#Ϝ��s���^9��BYi%&1z��� �v�?�^/��c �Mҋ:k���h�)D�4{v
a�'�)�'����\���JN� ��JM��-��)s��9!���p~�������d��-�6�ѩ7���<S�����@�3B����Ly�k���w�j��+�8Δ�:m�$����NG>GX;Q�97$��"�&#�h�bhu����s�ģ�Z������yh���ٶ���"��Z�bљ!�脿��p���u�r��a�HE=�ύ��!(��De/��K�h�Ɉ���Oë�W�l_���\���{������/᫯���B�(����EĽ�����V�ф�� fh^���OvA��d6�9۝~�ن��7�{
��2��2��B��`n1Xf�7��)O>���Q8؄�� �B
��~]��f�nԞi9� y�ͩh0T��{A3_X�L�����k�S�3e򷟮�xY���0���ܨ�$�5�����2";��U���ی,2d��F;@-�Z1�~J�\F����vnV���2�C3l��������^�އ��.�ǫO�T]$rv��F��w����>�#\s_{@bR��{?����۷�?�{���P�D0yǠ݉��B�V�\���x�e���{wsn-#�����?�=_��R�4�}uo����'3�v_�oO0׉�]]���������K2��]?N���+��޶C���]���D*l4{���X�v�{a%�,�ؤr�2A�~+��h"��r�
s Z*[�4�_m���7��F��糥擵'bh����XS���0���?��C�?����"xd��to�fE�K��R����]��� ���\����αʱO�3�,FvɄpFi�FB�ƈ�J�R�@��c"��j��3z�n:W����uߏT�������L���2b֖�������q� T	��-�{���t?�x���zf�ml�$�뻯�Qٝsy��c(��� ^<��=�î���#���g;S+��.����FB����ٖjn3f��p'�}�զ{���9��q$���g{�����Ib�,����w��\��9j� �<�+�*K��>�3��`
	^x�r��݇�㻟��ƌ����;_A�l�Ek�}�@e/�6�p�cV�r���f�R�����e�8!\��}3{e�a�%�-�O�9���S���PjlE�>F3(��ܒ�.�Q��g~#N�4:�{�[�ZFE�J���u|ʷ	
�Km"n��՜��յ]�DB�D����Ww�!w@f]JӅO���#�Φ,�S�(���ӱ���xd�k#�:H&�-���~gIwmf�zj�o�	�i��SG og݄pUo��̝�D�lؔohBJ��`���G��ġhl2\����s۠z���9�^��z�x[����W_}��o~�y�"#�g�{�p~��
��-\ܵ�T(ڃ(�ĺ����T(Z���h���p�p�K� x�y<��h@�|��y`]�8(�Y�LS���Ҝ�	���~3�%<s>�%2<H`D�NƂ O�	R�F3�v�����T�U`�� ��Z�/`py�/t��)@SLG@˞�������S����)����('AKf����t"�
��W�c��f�5�r�|eG;�R!T-��s���3��M�@U���ԍ�����P�Ȉ��, >��=���}�S��0� D�..��o����򵸔E�R%����KK#K���d@���Jǿ){�G��v.
�+^�(��VU���j.%�����:E�Lŋ����R�2n�/P��� �}�="SfĈ���i쟭Z*C��Fu���Ȟ�-�8�ut��Y�Di�A�'�N!٣2����q���(�m֪�HCx�}z�m{���E���忿DYo��dY�̐�߯�vP��+��N��z��ᦂӳ3�HH��ғ)�Zr�ә�녝����{������&0���ަB������I�������`�͑�M�F+OLWE��D[٪3��iф�˽�_ƨ��63�R��e�,��,%���s������a���~7�^v��ή"{ĳ)ǰ�v��	��/�`�w�`�� �1���F2i�����A��4�Da������f �ro�ݴ+;8�0�P�;?�({6L^58#� �j� iF��Q�������F� � �4�7z�R��@�D|�MG3��e�7?`Z��s�T��*�Sy̤͠Վ ��ZQ��0}/��j�?��%����՞ظ���@��K⡞t��\Yy)�|v��ٵ�h�ʜ���v/|wt������A8�u��}��C*0Wf;��3�s�Nk��=�ʫ��ʴK���o��*Ý�����o;�)bfm���P̙k��́?h�6�����b�s$+O�3X�F���Ƙ�� �Qo�=#�څ.%G:mn�pRT��rv�(�>�Z�*@�W҅�n�{�*�),��}���S�ͣ�}��G���|,��#;#G��$6bS�R���axqz&�:�n�%eV27Fr4�����Y��X��0
]���8�^q���h����a|gN��%�`��0!ȃ�j���HR8E�r�恾{cZm��ڹ��~�JPhk�u�vOZ�؞|F�͵�궅�e� ����Vr�-F�������κُ�5���!(1�$%$��ImCը��;����'��Y�e��F�l�a ��0�}��q��?���l�өg{�0:v=��f"������
����S�
�3��U��rz��B�Z�<�#�!�H\_8�"J���A���z�\��v�:Ù���F�<zNL�eX{P���,RS:���奝	;���,gZ'��
��̶ߡv�ID
PQZcLn.~���Sg��1#p/�}v�I�vJ�}(i-a�M\#�3����X�׫q��pȋ֪h��;Ԃeޛ�܆�P�V�C��m���@�h�y���Cx�>�~������I8�?пYh�+><�lǍs������[6�w� !_|�P��h������k���xb��&r�3,�#it~��zg�ԌƽE�h���-8�]	1�qjx��o�<�}Ec�;��b� ���vb��J��骨�3�r����gI�F����i���W�:D��?�����J��2�@����8��C���m��3����p�z�g��1�]���]z���{�5��	�,�����f8l��.4���2zk�Z;��[��^ڽG�G�D2w2|��d��e�����lcY�6�'��R�j���`���u�(uM���/���B�Z	1�C���]����_�?�$����d�����B�4�L��7`*F�P��1�r0�� G�����Rf. f 5�	/Y��#E*B��*�",�b	�B�a��G Ek�.=3��D����d��D�>@N���B���������*�g��ue;Qo��f[\�+0B��o�~G���V��b��Д*h�d��ik��z�d��E�Fѷ{���w��M�'k�V|��Wv�%l ��S@5d��V�}�d�K�nn�AD��ZA\���_kl�-`4c���+���OOe����(A8�4r���u���ݯU�ӛ��{�㈥��ʾ�+�*������:7G<~xT[�}���� �̨��S��ͩ@:�%�Ja0��`_d ?�ưtMЧ��)���&��ck�ȋ�@���.�G����Y��G��*K���lS�H<63±2���✨��̅�[��V	������������71��a�*V��lM�H�j1&�h���i�W��-5nvc�So�\j�NJsPݎ���/�����}��y���	�ڽ"ೠf]������	[Ըj5�sEI�tcɅL��mրC�ʜ�29 q�ԎzQ���%k�.��	�NO3���l�a�,V:<�ww!�����)�%r���}�t���o}�)��p��j'���=YT$��-� |��8CF祈(�,JW�$f�[q�B ��r�+~X�8$;$8i�nz#�XkW�H �<f��sM�ţӥ��p�=��r�(ɛ��1��t,�5c0�t���A�[?��Xף$������?��L���\���H;�8C\�i�:b��;\�2���l3��-��̉@�ݎg��{}9��� �>��N�L�Y���2jc��ok��{�4D	�o��<�kEA�H�"�<�Md�*��[�@�,���=N�Ƚ��rr||�C�,҅�s�������?�7�7���bn������1#�(�dP��� �Y�&�{��P��x?��J��ӛ��$��	Ls3ƔѦ���QMl �f��ͫ�0��� 1�ߟ�ވ8l�Y`��u���֎�l�$ǃ�d�Gˇ����XT����1A�Y���Ἕ��{�(Q�<��>31ӥ�����1V�+%);{���G�V��Ͼd}���Co���LU#�k�蛲�OO�	-�1G�R��7`>�{����U)G�X@�p��<|��o��W��.�ۘ�NT�go_�Gadgl�muxV7�m����{��}����0��WO{e���ec��' �h��������Hs�ث��]�,*��Z�,�v�ߋ��²�Q���B�-0�uE��U�<VG�X�����*��N��ǗNvS:��9��T��7���jd�kʄ�3�Y�#� K3N�)�	�ǩ
拳|Ü�Le��&T�~���йj�����V36�
�pb_p}P���'(xkg��_�h�V�f�Àb�i���G�Y;����"��c�|�}��/����7?~YO�,�,�K-|p�g؏�b�ֹNd$�Gt��7��؛��m�2��� ��hrl�(X��XF�r�9<� ����
����Ĕf��~$��{�ȗj�8��4R�"�vˁ;��)ݸz	���L̹����J&��^���S:k���B%��_�ǔjw|	�E�7H帆)��]y�v�zS�f!��r�'��:<�?��=�MVI���H��������C�.]�>ɨi$�ֳ#U�M���aia~ya � \ǡkWIowmι���P
�2�526��}@|�Fxa�ksX��V�#^>��)rS
�w�E��)k|41����MrU M,�}|�o߽?��1���]x0#ɜ��.�46%�H�rq��`�c�Q�w�Fe<�!�3��c'����2�����D�|����>f"��B��@=�<>�������s������1�u�v�!�	��/-�IF�s��\$e��2�>$pW�w�?cTd��?�g�4
��Щ������^�m�~��B ��會����̃]Tl�0∢�cϒ�gQNe��}��|&�V�N�y�+$La4�xL}.^|�0F��[Π�d�\��,+���S�#j��9g����x�s�)&뤗;6�Ț�s	 �')T�г�z�	�7w�#�0(�
`x/�W�Ӫ���ES]�Ŝ�)�|.,8E�܉�hwd��!9 �:�e�D�����Kض��ۏ�hӾ��S�{�W��mLz�6�:ԟ��#5�2�M��4-����KU��������R}��2�>ˮ��T%��w�eNŁ�7�����n�k�'��N#Q�3���ݮa�J��L���-$�c�����4����iN&���<"��T�E���D[�����&�D���X�)���͋��9S�����N�2Yr�`�UD��w����W��)*� $�=���W�'�gv��D�Yȑ�� ̡���E�+��Pu3X���#���EV������5����E�ń���Hp$e(��a�X�I��>,7S;`׷w�i�mj�J3=);3�X0���1��2x����LpyI�`�n�|W"Q6m������C��s"���j{_�}�}�����_��e&o�h�B+��������̂�^M�xN,C�VO����:Bf)�&�a]�447Z����A�<2�-*BkGL6��A�Fe�w��>}��l]�Ңo�7�Y���yƑ;�S'3jM[bw�p@�����++���K�6F��m>Y��
/��)C���!s��a�������� ˙�������yr�jLmo�wʂCD�GGiY��L�s`K�QKT��Z�FvC�/ }=��%I5
�$�m	�m!�v��UYP 1@��޳�
�
^	$�*�倛"쏆�����#��{/)Ͻ�<իN'�b�G�H�*��yx��&$�'Y'�v��i�7�X��A���,�a�ݏ��r�T!X-&���X��+����	t�ٍ��ImnN��2VH7P��s1�ts�I�kdNw��Й>��^z����A_�M���(�
f��eN��2z�6"�w����o�.j������:r9d�Tc�U\�t��:	')~�����L�01�H�6��Qv��%\Q�7L@�,�V����ݞ/ָ_!��X�Ȉ!��W򁒳0;��Sȃ>Y�;.	yٖ�6�)��~/f�~�-�,Bڣ�[p '`�nS@Jt����U�|���	�u��,jʒ#��(�R?Q7Zs�>a��A��˶�eN��/�gYP�(d��X,=RR��
�k�OO�C~߲�}=�v�������20ܖU?<���;������$08�A7����@+��\*���末v{[=��K&�͵�W�J�����w�Q������2R����_^��z
[T�U�H��2ʷW���l"&��U	����8w���	�#�z+�H����H���mEƉ�*��8������I�ݷ߆�e�d��a��KvyzpV'UF�+��8�����{!g�n���JZ�+sX �V�q���IPHJM���ƫ����Ȏ�����~��P����Cx0�8^LT,m_���XVMs��?��i��它��p��^���S0	��
��=��1ԙ ��Ge��[�Z��Q�7k���΃e�D�d�����ؖ4��Z��ul����F�{ܛ�l�8t��\�oAeI~����Ո����%oA3�� L?~� �U�~nS����;��/@p��b4�$�<'5�C�zt^����e�$M�-{�?�S^�
X^2�-�ׂ�.�лFw�i��,���������u�ԋ0������B���۹w�؎#��i'�eS�;�m]F%o�5�>S���J�
g��v���g��V��Sצn��M��N,���BR�+-�gZ]� xu ßUmٴ
��ƱN��%1h66�x6��@�	A�ܧ�"k��SDL\[����Β�^nl���6�����:�6A�#^E�Q�H�'�,�{נ��L��@�F��O[��8O���3WD��n�n��_n�_0#�)sJ01 ��.#K��ҽ]s��Ph�\e���<~wtX6��j%�M%�Xnu۰�I��f7��J=(��|b1��l�E��%_�:�][�ٰ7-��o�mb�(1�c�M�&އ��hy����9+^�ޢQ��>%�񻼹��ͽ�~<�<�M��,ʆ)��)ў��=��]oIt=� ���%یqU.C6�y���<o��깤�S! d4��*��Ĵ��R�%B#��v�� "��*
dp�����j�}����48�z���T��._�Y�^��Jd��c�m�z�P~��e����&��peN��>� T@
�L9� ��6�1���:=ǖIA�����ûO�4��4�-V�.�zR&B��ʑ���u�S	��Sͦ[�yEVy?����o ��zꩽ�uC�T��������u�yײ/xɿ������ �#G�V�8���И��ӓ�������ɹӆ�nlYW2����ж�f��H��ݡ�Qp
�]���ƒ!�RQj��> $U����W5�RtD#�pa�J%��iB�(&��C��(x��	s[�;s2:�z�{N�(�9�.�}	#E����~ �y�3����M,H�M�*V#F��B�`�����A�S��}Q�#Y��v0�+�)��8r�p�;'�	
�E^��6�@e�,�#2����Jck9[{@�J�
����g��s�ߺR;��J�ɠ7��@�����ګ3TX$t�Od29	e���W���]*7R���DFP�R1r�67ם��y�%e�ۀ�M�x�ʷ���3[��DR��j���1�B���ͣ�~�*S��aS��kJ�!�l\D7�2\����)�mBHR���v�F\T�j�R��t��m���;�^�[>�V(��}5�O���`Z�^'�5�=_YX��f�����RI��U�'��Z�D���x'�3Bm�?��c�~��2s�A��˗����.�f?\̜S� {#���no��� �_2a���b�A	�Y}�r	|`�d�?���8�)K\^�Y�5g''�����vV���+8��F�3�=k2]l�+�CXG��g��th3�hζ��{5��ن:�ˡ��n<�"�����¹֬JB��|�Ol���R��� (�(I7=���m�JPQ�,�;��b��K<���hȉ< ���rS�K�x�������{sH�z�:\��6,�hN�*�A!�8��e�1O�_���F*���;ݝ�:.�jY��Ճ9�g̚��`��G�v�BdW���	
����}����6��W��p'�x
�֮9���=���|�A��..ã���R׈R�L�ʽ����+�n�}���0�������)���-�q�3�q�Q/���ю+75�����%����������;����p��� ��n�G���
G��unn(e�\�|�4��_Z�9�8z5�u�Ɍ���^�o*�cbB����{��|y'rU�$C�������/�'���U�G���;����G����9��f����	�֢��Ϋ�����3-H��9 �A���l�N+I�y[�%�T<Su���y{�rd+�A��^4��ð7�52���Q�a<Kc��U5ڎ�������K��^O	D�.���R+!��#��� ���l����,]LA���2���
�X���핁���ܵ~ɐ��N����ec��3aMhl%_��$����V9O}�d���\������3۶�zcP��k�3�y�AGl���(����BV�U�S���@u��b� ���n3���c�|���*-�.T����J�"�
I�U�:���i��ʆgE��[,���������a�H���m^���8� ��lVo���D�40��'˂�`ᄶ(pg���0�9�hDs��+�?X��T6�������f�;��*��
[�%s�+P��гC���{:
W�WbM2��9>J�;s����~+�=�e͉f. "@ݿeG!n�*)�M��*�W٦�Q�nKrn<��=Ē�X�I��*� "Yh
I�{p��n�?�S9�ü C����jD*�z��Le��Q=c�b����ؿ�6�'	��G3�����]Ϸ/_�����d� ���E��(��� �f�U�Bs�d5)0�-;j��4ON�E���G!�ga %���%i�`�_.u���_�|^��2gy0I��K} [�U�>o>������Q���N���%D����,�(#*'H���B�r�:=����@80�N�\ʊ��ܵ��s�(��� �8�oB�_��8fÖE=����M���+����1(y#���[aسH�2���}/�]�γ�Vt�!�Mp��ƛ��z��L�����j������{������7cf�3�Й��'(w`�"�����_"ۇ�u�� K��en ��@ �i���_#ή훏o>��ŵF�i����F$��|�/�Gh?��|f�n����_m�]�����c��=:��r))��L���r��k�%b)�5\���,�A:cfyrN�&'
�[6�s���>J��5s\iܲ ϥڠ��K��Ƴ�L��w��[��&!����*y���������3Χ�,kN�w�L#���.��L��_K�2j����;�䀫�ޥa>|f��+}R��#�5�vB>	��{\V1��9�V�9��ng�Q�$�t5;x����q/8��T8��kk3;t�YGe�> �����F��R-.�J�48::����;�oQ9s�s"�ŕ�� �Z�؁C�Cw؜�
Ҁ�X��拷��էOr1��tP)�P��P;�6��{14����:b05����|�!g���2�ŵ�`*��ic�x=SX�8W��Kt�6˯'xT��l8	����&���G����&kĤ�f�{���������ɩ�{����{���RF�I�����R�_��/��𑾋�*��6�[�utΠ�Wq�G9�ed���CE:Z�S�Ǜ+e�ޡ�:��۵�U�4Ԧ��2��U���YG��mƤi��?I��9`��^R�&H�b����1�����㴦���<J�I�Ȯkh{�����<���%Ty+��h�Įe����Q�)�����O��cCօ �@����@9����p��7�2��N�$&눌�Ϻ�7�?��ѽd�\J�񐅤�G{a��$ώC{��kᖔF�b�R����z5'��|�
=/� �����=�N��ݖ��y�d�WWW�ݻw�~��޿��>|��xG3a!�<�l��7|���G�'6�	wt�|��֎-�p��~Cקk��S��O�8=�;R��}��r�gN��y�@s;g�B�đ�P��?�z�&�wfԝ���no�3k^
��[,l��`�#���.�Y�8�Μ�o�.l5Vl�Z
Y[��3ٖȼ�4�^�O��γ8~�z���Jh�M�t�	�ϙ�h�/���0�[���f��#����3 ��*?''�D?�xΥ� Na�qǂ�~�EkS�˲�x��4�
,��&��L �,�\k'Q�]��W��]�=0`��*�{�?&цX��^�B���kU7�\���^mU������/#�4^��Z�I�M���_0�T >̱��R�4;|gF���N��G'���\s���}(;�q����?���,�L����<d1�^���5���f�R�>[�Q��
����H��	����E�Wz����$���e,�83 m{�6�a0�HX��]����z2d��
�G��s֧4��H��V��&���3q������e�w2��Ly��O4^���q��<���_�Ɠ0@��m�_9`HJe~�6�[(!J�V!@W)F��2;������F\�6 }0_G��&��/FSe�߿z�����2��Ry�b�
�9Y��&"�B��W��x��w���Q��ޮ���4t./B{�U�Qb�N��4+ae�ײi�:[+0&b٢��t�͝� ��Fۅ��A}e�²8)���1ː���C�2��M�ȵR=�j������H��˂;��S9�����Cx�u���cW��UGs���x��8��о}FvR��N��3�,�Q���L��,闊�۵^�kz���^LS ��R�]*�*$f�d����γ�V�/��q��W{�����J����qy$h��s��~mg'���!���Ƣަ߷��]���CI��af�y޾���K�x��v�{���\*[|*�&��Ⱦ�W��=��a����7��u8�����0k�n�ٛ�$���>��щe�����<�I�Ƃ�ڂ������t������
K��&1NӪ+ ��Z��4�-�]��l%��F��vv�����L��8X29fRlb������]WY����Tʠ�r�^pMY��r �38*��$G�'�3Ͻ�1 �yK-�R7덣L�������#ɲ+����Rg��.���3�;C3�ښ���1�p�-�U]*5�v��w�{��-4��J"ܟ�w��D��Ν	Z��'�4�C�N���c�ߏ�c�K~U�t[�̂ ��s,�e
���YP���N͎P-�Z.�5F$�	*]��eǖT��fcS�~��[gً�q�ʖ��ӻ[�����퇍�/쿋�?���ݲ5.Ƭ^���{�vޒf&_�"��i�_��A��yG΀����A�����u#���ڻ�h�B'��:�C+
�E��2� ���k��=q���ҝ�4�>�m���<e���=���.f��9G�#{��7k��d�o*drx[!eF�"�2�}�r��5WB�����!����c�a<"�[:��F&r!�ɒ��D�1��۶i����f� H������pl�/m�,�Ew�і�|D�I���a�~�.Ա̚g=��Db_�'җ��H��E�s�Y,
t$���=�<�,ۄNo�7�+i㚳�XWν9:����Pd>�ô �ʲ��=7V����Ee,�XP�l�=�z�LAE���_T>u���W��@urs-��0?ϯ�(`��y���;T�0���l�*���;׿���*v-��l`B��d4?��	dXf\qXK�f:�Bo����p�ټF��,bi�0��
/��7aX��t��5�3c�6���
�5v��><<ۇ�a`�oNٍ����-��Q��,��SQo��c��3`eY�/<�����[,(�:��-��r|�!�ɥ�K�k�����'���F%m��%yI�aF���*m���?�liG� S�zFo�v����n�y������Q��}�%&��*NK���m������n��ޱLx�c����~	n�-fO�ӳ�3��'Ol/��K�ް�F5��jTך�R���Z�=�$3���5��Y%�h$0��Uo�$�l�hWN�3��U@[s�i�f?�+��&&!�d���!�9���2�(u���{��ٌ��$Sּz��K���'Qi����g�E�׋-?o
Ft��_�U-*T�4G�m�B�8�
I��vصgu�s GI�&: r"�
9���l;U,Ͻ��Z'j�̃��'W�.on-� �<~O}����9�n�7��vFx\���L}���n�j��Cep
 ��7�
{�j��4P��c������Z$ۃ���Qs[�[�F��[E���ZyQF���r �r
�����B�6>'G����
�l1�9]��RUߓRd^҂��c!��L��z�-��Ĉ��o��}�4pB�㼛�i�b���[��R3E�%!|Ŗ	PVő}��?�Ȝ&�ʓ�$t��BN��.�D����gDE�W��A3�m��;@�TP�*�*J-����P @  蘻R�4N�X�3xrt=R�DlYf�jS`��iC��J!fD�q���_xl��|z�������kEI�uO��ت��o{��o���%`^�{Q=#�b�"��>�it]�U���d�����^Y�nU�j�CjGb�:9/��F�+�F�Ԝ#Җ3˒�_;ا��r���]����a�#�j:�#%#�mw�P���^�Vs��o�%j^}aٜ���FLIbs��]qvom	,"|����v�!u�j�LF&̆�J���<�������Sźo'�Qe:����`]���Rl�E߷}3|8��eW#h��\Mb�ՒA'�MJ\�(R9��� gg��eY��!�n�;b���U� Ԍ틧�Z�L�>,sd��.� �Z�HQ��KUg`v������M4����B�pڔ�A��3B�b�����8�?{n��C��s��y�'��zk��e�]�&Wu+f����VJ^6�#����!4J,���@���*0ɴ��G��ѵ��i	 B��'-?R��L��U<�'J��v�DO%h��"%�^	����eW���O�2[�|4�Ը�G��w��_��J�O�Y'����K��Ad.񚅍��{x��$�Mbڭ�y&�٩����6%_q|��R� .	�CjC�{���1`��8��X�Y��� �LK",o�'\d�E�SeO<o{ S�� S�(fD+U�l5Drn�S�s���/?�"S�/��>�/�l}�\ڔ{q	}����!��o�-j���}�2���_��}ѥU��s���1�"���YF��y�� ���ō��K�tz.���2�!�ly �U�*�M[��E���ce��?�!/p[@�:�71`��l\�<�}d\\���^�,��2ܱ�?���8��w66B57a�I�V�I�� �4�ɂ�h�C��R��_rX�����l��p�����hcS����gmk{su��p��Q���~�Q!����E����0Ǯ���|r�2&�����l=?)����L}�n�Z�8D�F�9`������P��r�2#J�#�X6���措ǹ����g�����iͰ <:y�6�l�t۟�/>{��a�~� �����-8y��}xl��}��:����5�X����T��m�;�:?���^�y7�A�v,�ꘑ������M���Ie�L�%T':�?��cgǢ�Py����GX	�ⲓ�r��pr�*���3s��R/���^rm"����-�[У1�θ�7���-e"��\�#��+1a:�=r?�M@i���r��[T<>V`�z|�~���0�Ϟ�g�B���e?-s��~z�?�jTs�fp�K�){G�٫Wvv�a����F��d6�R�?��<�{~�8<�g����_�,����U�����gD�.*w�n_�˻[6�b�=����9�����v��p�k�3���LG����vO��\�rj���M���Y������ӢX�a�ww���ߏ�6}>�A ��^�A'>l]�����K����y
�X�kd6v� 69�[P$'���z�	��t��>پ���Ʉ���s*��*g�i������[}�`��Ix|�(���� Iߖ����)4�/i����G� g.��R0FT%��g�H��/f���S�n����nՔ�HZ@���jp��GdN:S�@c$�Qۤ�{�aی3�	=�*�=VN܁�e ���b���\Q?����f�W�dx�Y(/.*�l�s+�sf)v��v��0?�m�M�^s� �"
�Y~re��n�X"�a0ʤͣW���yrq�Y�Ү�ekWXBƯn������X�*�-0f!Z63�g��Y��O���~�J��(��݅8����Jq��ٽ���	�5+��e�DPǽ\�:rV��E$=nD��x��s����C��Y��y��G�-0nV�4�4M���s�2�vu��Q��?��t�m1a9á�Lc5Q�}��	������ E騿7O?G{�>Z�o[��g�l���gI�^T�]��FZ�4+��(�4-��	�b������ot�B	[G�GfEo���F� �Z��^ח���ݑ;�V&2�溜O���?�l{��蒠sل���e`@硜.�Q`Ш\Y�ʜ	=`*��P�P�V�\��d3Xgd�L�O���j=��a/
��Ȍ���~;���ƙ�s!U�LL���ef|s|�u߽��限����[Y#�ݲ�YI���q,����F-�����uڿOf�f��Tfe�bhv�7ꇻ��'��s.�n��`�û{�������-U������f�tlg�O�F�������8p�.�P�8(���£�Ga��U�Zc~�ք�N�1˸�f�3'o�DF�XN�5��;���L���,��DU%?+�,ff��m)�J#B�걊�m�p����?4�\�0�,��>�z�=�W�L`T��:=��q��`�?mm�PP!�+Є{�g�Ng�ɪ�Nc���/>�<�����#�&��������mo��\�e:O�sә�t��}��T3�^'qlyaC�@�-�/ ����a��Y�`�Z��7�j���6��Ff��S�.�80Fc�g����f��V�q�C˘����j��/F<0�<���Z���6:Ɯ��2Z.����� D8��K�f�{1jw�me��.O���~H:�;8p'*U%�@Ap�n[�v`���ᑐrU���e$�>K'�|�O����pD��v�J�����At>~r�rݧ��U�A�P �a���0f��ZO��=q �P=.c&���q�=$!my@2��?�'3�������z�Q�����q�2���POunF��T�"� ��[cs7�Ѓ�e�%Yʂ�^q��^w��!�.&3֭�t���b�d b�����1cI?Q�ϟ�y{���޲���E�p����#�ڴ}���IJ��f�5�Fӓ&��7���%Ƚ��вlil6�����ɫ�9�.�9�ϴN?��>��JX���`02��y�ʶq�.l�3;Cx�m�������gfh��ڇr`z�RZi|�KS��C�]��9��#� 4>BEk=��t�r������tV)��[��	��3s�p���	N�Vc�f+�3��)�����8B�� 	�';[˻i���m�G�gV.��]z����F��,yik}gϕ�������Ȍw_wA%�������^�S�86	£�ii�26�7"�Az��eA��g`?{||�ZչOP@)�C����a�s���W�_�/^~f���j��pɪtQB���ڂB�]/,h��-#�*	�9l�܌I!��������׿|���I��%��
�����n��O���~�+q|2���@wU�'B������v�	%�m$�C�H^�x!���n�V�̼��h��a��\Y)�#���o+��?~/�46������}MelmnH~��?{�=[�s��/��)�HI"���p5Q�L��j5�,�������ww��~��/,G�I̭D���>:��KЋD��~�<��/�����f*y�$��[���4z��a`8��9�m���`��<�"f��9��`�	�J\�+�}�7��M�Big!��eby��}�;�����i�8���)mon�/^���,P��������k�,||�d��@3NYˁM�3̼�����m3�G�N��h��Ӈ �^�5��2$tm���H44�nG��G(��xNd���xt�"�Y�:�TXKU=`2g>�@BP��� ��J���C͞��w�,nG����\삞���..�6��ʫ1�MLK��t����VI��c:T�U���y��O�[cG�R@=���%1��3�?�m���o7���[�{����o����L�I��h���i�7?�� d>qJB���*�ީ\�a���k	?�>bU��}&�M�'0�-���k3�=o Y �ږIQ[�h��q�u�2���=y"�]{.�مR���ef0�*�y���N�p$���8�3)Q���(w@�hT	 �o1�����F�6���8f��G��k���T7�8���c]Iǁ/ʾ��u�YC���+�<�7׷꣒�n�:Q2�T��7��f�����3��vË�G�pw�Y������w�W�X���<�nn	D��5��	���H;,�adN䳗��S[���1�In�RP*�l>}�<�����O���|1�����]/|��!\|��o.�|�B� �}�����ٛ�\�q���&%>�����O̹U�̢��P}4J#Hƛ�X�|H��ճ�>��6�jT��*��v��UN�6D�Ud����gZw���oD�;�ZgMY)�C��q���0"�C�\���Mя�����c�_���o�t*R����-�X�S���E$��5�ٱ ��}�˫{9MyS%��+V!rD�|�N�~��~�2'�Ȃn����b���o���m;0e�m��;�!HY��0�E�%�N�J[e�6�ٚmȞ2Q��7�dV�	k�b؅T����|+(�Ւ��+΂#�xndIk���[�6��˕�M����?��G�@�甎*��@�hD��r�R����/��ac�>W�2�i��,DfDp�߿�)���~|�&\M��)4rHl2_o�C��Ç���d�YIy
�L�[U�U*���!"�8D��9�� �#�P�@�D(=�FY/����L��9F��@����mIB��0G�P�-E�l�m��`���?~"�ʲ8+��|��5=[�]�v�&��]_��O�'h3��*�ޓ�-8���ǟk~�Pf���{����[�qr��ՀI�y�Ҵ��2�Q�����B�L-#s����u�]_��M��5�F��~��{�����[77�2�
T, �<#ϴ��̘ �	Ҙ`���.Aj>d��v_s�:Gf�_�QC2����f+�$��R~a_�!p~�m�Za�>w�H�i^N�j�am�������ֳ���0��?�:�c���eB�1��ږz�qse�-� C6o��H~M;@;�B!ci����q�o���N.���������P
�@pQ�Q[��?���d�d��;{a����:v���X}��}�uX �AV݅p�V�$����o����Ҝ�W³0O_����&�ƪ�q�M��v����pEp�\�µ��/w8?��}��"C���O�7�`tGǫ�!`Dz�0������7>��U���^�����ϪG)k��s�?Sk��4[�Z�3�XQ��G�	���� �~��lkG&*�wp��p&��D��ʉ��� 9k	�P�`V.����t���T�j�++��ؤ���������TN��rn�<}"g�=LH�B S*~����s�Āԃ�u2a��̴n�lwv7-�<���~�,c̀����C`1�z̬I�W���}QJr��j�YbDq���٩�"�p(�$��à,���,%�.B"��\Ƕ�T*������/xR/$o�h-� �l�6k�U�L��%a����P(�?;<�}������sJ���NTq^�#��9;�~�I�/Gy����3�ia�b�cyZ���0� ��9٦��;�y�.��Ԑ����	m��s`���9O��l-��Q>F%`��$d�E��!�XZF�q%���5l�Z�kAV��5oݎ��c��?ن~���4�!��=77(�SN>99���I����FJ'5���1�s�g�Y�z!a�Vâ$�f+
�C+Dj�r�0�M$��Q��6|6�Nx�Hk����3�x�)�%��T��|�u��GhO���<)��}^�t�}p$�����lؚ��_`��TzT���N��K����v������W5�k �O)��5������9/��ʬQ�b�%�d����Ap ʙ}ތ��I�ǜz���=�Ȑ;��m=/���������Wt��2l�؏@��@��U͂OV����[Q���M`;ן-^�~0�'9�L�gk�� �g�=Иd�lVДb;z�n⨋Or�1�������0�ӄ;�$��<��H��@�!M���h����c��q~6����,>� ��dr���N�D�j������c��߼{k��:�;y�+�����g��w���ek���}J���<3�l�)�l�h��Q���6�R�ZpC�$pV�Ԏ\��IP�ȷ��k	��EE��g�\�L��v�@ >�`����!%b��YM�
.��|[�-$9��?�j*����HR�f�U����a����*�~�V��w�>��x����pf�58z�H��f��{��eXڳ�M��v�;���/s�u٫�-�e�kC����f+�Wu�\+�R�-�9��.M�c�P�G�bT���s����-t�a'j���`��z��n�^W�w!�ԥ���(�H��?��ۃ/�g!��y*�9�O�Rd��u_�Ј�O]��R&�b�-']B��,Lm���T�ڴ��Z׵�;$ٹ�
 m�Y��]FD� �`i���YF�LwP� ���a�=��(�!sF��x�-ZN�8$��:RH�ZA�c����8w����m���6�mP�:��1s���У���p8��GT����m߂�c�7@]���a hA����w4�/TA@9�l6	w7.GX!�E-���4��Eӎ`�{����=�fɰ0�	e�w�k��-�O���p�8L�]��@��g�b2����ƥ�����4cO��^���E�[��w��I{��y��_��:����{t��H���mK/k{����ր�PS����@�<9p��]ŽG�I�������q�OJ��Nг�3�2-<ݒ�Ђ��R��=ǅ��܂�!�����w��BT�!+<VG�h���Z{66��:��|ӱ�]N�SK��Q���0��3���&X��tV����<�����၂̀�
�a����&x���( g�\�i�R/8P4�n��J�ќٿQ������w�k� AUR�L��\t�t;����B�*Gт� B"��ʧ	��g�^]�Û�{Q�(�{�!�ތ%���9�%�#�)g_c��-u\�K��9 ��
_��Ԃ���`���9[q%�n�R��u�I��Gz�}��T�كru�-&Tt)��*[.��;�5U��G�
�AU�pO㫹���G�l*;����>o�"�h�,���ӭOˀ� -�F�A���Ŏ�Z0�m�Y����&�T��pr{��ϼ�m�v�� R�{t�v�93Ϡ�-
l%j����9�(��jS&;�4'�w�� vq��garw��tJp��d(�,jGD����u^�z]�����!3tn�d�H��:�XQRT���	P��DX_����|n��*];V����*	x!��Ȥ�,��5V8RŤU�{$�~�7�T�0$�C�azK�X��:1?�C`�Lx@��/=�"�[z	�^�|fN��PP����f5�`[;�1[�:J�%t��!"�������u�3C�p���C圾S'�Eߊ^��G^GP��������R��Vw('��d�)3S'%+�>�-}.U���݂F���hUI@��4����2G>J���E��h	`�sx��+����O��a��16%a�v�I��e=FPa��m@B��1����_���?���7_�}8�t���A%��³���~(�"b�2<�{��������5<�0J��&oF���e$�'B?0���P�è��:?�ÿY�~�(+� e�>H�М�6Z���e�����8c%��*��1�����X4��h~�
����;�P �D�#k���4�.�a���h�I���5���������T�) �l98x���M��h-浐�To@�/�W���3w��'e�,sU��J9����L
?�^�y��M�1ڞL��|�+g�"�P��L]�����" A��������&�F�(+��!L3�K����}���$8%XA���*���
�����,*�H�v��^���)Aa- ܩ�<1���2 d(�L߿�y��sa{��9�=��*����\�4io�3Kr����U�l��&�K֡��'�V��U��MIC>9a�����'�7��J8��l\
��idqq/�C�oHn�h��j� wv���:� �P'�Xro�7�ˁ�+1���)[O�Y�-�������߆���p���M�u_4a<7��q�b�
o�݊�ns{W�u�gWr�,�ٯ䄕}����"#�((�n��￱������r��v�VՊCC�����[��9ڒX�Nu֚Y$�ZDf�M�MA��ͨ��m{d�9ec�	4��,sXΖQ�a����LR�ԅ"
0��ԛ�s�W�a��H�5�jܠؠD �N���MG�%{�������F��e��k�z��lor|x�i��H�ҢcJЖe�!�`- '���Yt��p3e����)t@�̐?9:�U[e�U�{��1�oCW�������w����f������d��� �7kwy7�ى��}��{��*ϧ�ۀ�+A�^\c�d&=a+p�s�V�b�|=�*0H��^�1�J���;d-��9;ֆ���%��E�8��˱��f��E5���V�V+�]���Q� v􍘁�:�`4��@��3=��3��	������NT&
BVK�׾ߢ f��V��j��:]�V�$��n�~:<86'��,(l��	s/�|iM�h�*K�XC�����Ջ�� Ns���hEJ�ё�/�N� ����e/�ᾃ��V'"����N�P�{�����\ k쳷F�7_|)gμ+��
{��o
{��N�h�μ��hT�H�}e$r.�gܪ��Gș�Tޯ}�"g�ȶ��MyB�r!h]��5�z3���w������Y *�2��{�nz�Lڱ��!�et����l$�ì�P���ً�@�znb&�zo�\|�y��;s U*}�`#�Q
��}>X ��tZ�{����
qj T��V��d҈QZ�ĸ<�p*O�٬n֙��,8}n���bt�
�:�cQ8K���ňp�8�*��S~&!)ʎ��Oo^���lS�j@&��(!@Bb������E蟼�����w��6J��*�� g�1�A�]w7�#S-w3KΜЈg����]��_iD)�PڜQM��|%�_��뫫��7߄��ONpO�FHG�4�(0�0���=��pWH?2����2���Dk4�D��Đ���^�;J�<JT�k�N,�:��)q,��5g4�yXu\��Q�JY�/�RFP"j�6Y��s��d؝|�q%'��e�&�m1����"<9~d��Fxn�mU�X#�X[:N�1p����<�3e�j��C�Cm��F{�Ik��b�ك����A�h�U4y8yd��;��h(�"��� 4C�o�Վ����m�sv�I)�\�mQ$�y�_�I��6��:�W����=��"��0��iY`���<C���ϙ�µ����pv�|��&@)mW��Q�P���ЩD�z �����c{�4�xwu���k��Ζf@�.u8��V�L*H��PQI�=W�X��,�Y"f�W�9@��Ϩ���+3ʗ��/��
�6�g[��߅7?���`�&'R	B4OkO|8h��|t�X�*����9�A�~�q����\�^�Ha���\��vm�U��{AC�؇�,XT����c5Qƒ��|Pʸ3�F5�o��h�ݸ2SUy ܊%`!Y���9H�����o��bf��8�gEi���uc��2�C��B���Dכҁ9+�����J�� W��S5�2ۗF�(��E*Y�(��΄2�p'��y��{ﶄg��� k���w��b�м��� �Oi����%�lZ7Ty.��7�P����pP�^Z���}��؟�N�l�%e�l,�;�8$/؏����}L�{�t���7x����D~"'Z��;�IO99aٹ,��&I��g��4��j�Kة͗J�1+N���).�7_�X�J��髬S����q�Q��󮩎�3%h�G�j�i�Ǿ��S-���
��]GR/-�����٣��]u,#����n��ys�=�k;���@Hxc��Zs��<r�6^��~��.@�oz7Q�W ��|�΢���gO��?|����W��Ɍ�J�|P�K�W�M�Ulc^_���Ƅ�r=`������J˝q�w	V;�p�Y�}p�0_AG�R1FjE��O,�8E�/�Ω/��ݗ"�Br��5��*��W�od�N`
1�ֆ�ٸr66���v���ak{W�f����\�x��jW�a�kw �|dMەm
��u���MuM]�Qz�E'�$�f�>�?|��q�*��v1BdB�#����ml����4�@�Y�Җ�1ݝ_��3�0��a�.)�]K��l��/�f��X�
�x*6�|�{���BP��`�"(���vM^Nk�E,�E��g���+	���?{&cĳ��2Ck��Y���=��k�	����JR��'*@��V!�k72��~:��á=˾�iy�s�@?���9(9�8�̣Ofw"���CBo �������0fw��c�� �۠�a���tl�ON70"����1
R|bܬ���:'R���N��dU(|NY%��eL���4d�Ih�^с�������̃�%��ʃ;pF Xt�o��hQ߼~N�N�M��xq��*�޴�8�������p\M�h�Js��]�mjq~Ȃ��i���_��p��7ډv��uJ8�1��~�v�ˢk���Z^�i�>oK[袶@�Z(�&����>�k�����oOO��ݲ{��;~��K��'��*��˱.�'�&H�2���!��[�G�t�)^�W�,���_����zzʷ��}?'1;e���R~��^;aNr��~غDơ�`�o)�-�����#��
���&�l&�K]m���_�Ĺ�Ut��x&�j.[�(^I��	��aZ�=����Bt��:��e�j n*�hY>���N���8����ӕ�3{���X~E��vؔVϲn���U�WQ�I Ⱥq�e`�2aP�����"�����l��:� �0�;vÿ��U���Ke"#�� "XP.*�����(�H��p�\o[��g���2Rao:5��	�y����X�1d��M�#���%�W���R��qʔ�Ч��7^���
N��l�r1c��FUk���/ʃ8g@�%�IBd��ix���E�R�_iOrg-�h*%�"ғ�Ws��X�e��6�h�&:]w��(՗��
�x�)B����-�lEŦ�yb"��z�>��!���2���.��7/�V�Xâwz�.��\+����HsJ����f嵕Cln�(��S��@��e7x��qx{y���u�^���؉/����n4��N8ʻ;�5�Ƞ�Q�y)���_�s3��m
���	��H|��gN�����qas�������@ws�8[�L��Vш��6څ�5���
Ǟo��.(.�1G���`g[�6�H$A�ۀ�L�"}e���F��bEk��������4��ԋ�J�x�q����d����z����;�̸��V�����d�N�f0��kGߑ�E-9��m*?ϟG��:܌�"��q�Z�zO�y����m'�~���K-�����s�	!��J�7�����4-a��w\*8�}�:�ť�N�1be�<k{�O�OP������$�����V�Wbf�[x/������n����#cvt�3 /1�Q{m��G�D
\�e�I8�`���_pL��p�����Y�ź�&�B�I��{�Nc���?PFzȈ�v�@��	Х�eQ�5���Y*���k�5�ߎz�I"I���4�$#X�,�NU�Z�s\a��W#p����ni'Q�A�-%C�v�G���Boo+d�o���KXP�-ll���G}��l�
�w��7abY���,�-������p��>y�;>��34�T�M�а<�Z_~�Exn�ik�)�+F(�=z���Ȝ.� ��Yj�F)��VS��g�/ڳǏդ �1�:�6\Ӄ������ח�=��MD�lTлW]��%qo�H�qЩ�7�C��R���e���p�5Yd���N����_��F�+�<U�B���簽|�E��o�.|��KGc��h	⮎;RO:>�L	O��+��;��x�3
A�P�"D(��I�X���c�8�&DRMGҋax���r9�U��T���b��h�{e����$#�� ��|�3��-Zo��ڃnµ9��}��0�3�@6��ށ��
��E($+zƛ�{��<�o  ��IDAT�(v#`�ӧ�f������CY����Ks�R�M��Ђ�����l�m��U��S���婮���s�6��Ȝ"�S��߼7��� @����������'�~��=�x�/T4u�ц�F=�<64�a�#`�v��ɽ�����FɈ,�)�<��{��H� 8dl���2�s���`;1�o������ܿ�0���i��eg��`k(v���J�<�9eƆ��-U��@Z[�OT]�M5��R#e���Щ/�K�-_�@�����ǪUǞ}%���ǌt���E�=�Ri�Fn
WJ��p�+Q���j
�Ӱ�	DS;jZㆪ�^�b�rE2�� _!�2Z7�N?	��T��r�,܎�Q.�P]��5�1K�� �ru��$5���Iʪ�*?��}��^�W��v��!��#��g��������}8����b��a�f-y�L7����^t�a�,�v��F�E�mX�`H(s��e�8���s	@��U��]AM��s���a����N-�gcw��Q��h���̸��m��z�tE��e�������+������ך�f�2��҈J��^jU4�B��"��S;4���|�g�{�-�]ޘ�=��W�!�[��b]���" 77�q�X���5���1Gy`��\�Y?J��W/^�ϗ�{q�>��|�,��a�)|��1{�ӏa����=˾�'�.!@ m��w��z��P�����`M�]��=8�<�p�T�<3����[�|g�q�5��v���:ux�m���Sӏkҡ+�T�q�n�@(�g����cը�[��o�(�(�!3��}/��bP��6,�Y:S*&�M���X$>U��`5荆�^�|�?�-���@I��^Hh�Y��2h`W�y�Ne�H�'�-[?`i�m[�AK}��Ζ=�+E����Q���کo8/][��M)��@�ೊ�YXdS�$�t�<{�@��ZV���o���[�֒uxb����WrT3��E�J�B�������ߩ_ة�DfB�B���4����q�7 �,j'�`_V������d��aW}�C��F;a�����e��/G�� U�}VM�����%;g⹚s���0_�����
�p	�8_���n����Sg��Y�c��s_�YA0��7c��0��Cm��^�4u��k�DI<7NP�.о;���?��)|��f�K�GgEG����N���7��ܱl�e�+X�86	p��I��x��k��`J|�gR}k�I�r����C 4�l�s姖�+�K�	8�Rkm�I9�%����Z��l��#�B�;]�	%�PP��ߑ�c@8��2�{*��NUv�S�
�b�n���?}:���5�mϒ]�C\�,�j&���=�۪4ҙ���,��׌Y��]��>I���6�[�r�Vo�=Uq��6ռ<�CG'�f�����%�_�����x	V�N�2:o�����ɀ�UݸvF)wF����;j!��5���;���(� �x�F������/���m3������F����*3�������1�����2_*�&k�gQ�8s�-��M�5)�Lٌ���`5!�K�D���OO��>�o���2I�aw��B���Ň����[r��f����۷za�P}�Ϟ���N��\�q'����F��ϔE����o�����5�*~�#�4�CL��y��A�5�L*�z�=�|�D� �o�D���� ��.3x�c�lrg]�c��ch�^o-���E�D�P���N6�9.,Ym6��ү�8�kd�l�(�D�(�7@&�wmc���D���û01g@agW-�k�.fk�A���sAo�c��8>�];%B�j��Ԙ\���^]]�Z@�`@""��n�-�Vk��Zyd�rcw�.�@í���-�[!Թ�
"�F��d���W����6{[}��G�j˒0� x�`$����ţ'�l�=q�w�}/o�$DrԦ]'�'׶ޢC�<��͉`�g��ak�7�9�=�5@�#��r-^����\kL�9h�W�������:�l��)����]��a����%c�`O��Z� �#�7��B�ӻJ���]߾��]\�[Jh�)�hĳćg]gWҨ
���D9ҽ���ٵ��Gf?7���
UI�|�,Ļ.�����K���i��TfΣcDJd~�XC��Ț�!Of���8���m1/_�k�e��8C�]ab@��Z�rx�o깦��,w�]G�S~����T������PW�ZF (��i�g~F�r�9���\텏���X��ɒFN�--����pY���Vp��i���,��@�d\�3^%Nк��q��V���#~�S�~����N��ƥ��[_�"9���ƞ�g6���4ʊq��s�yU� ��χ���ܰ�����J$-�ZZ�� �o9@�%\	���d*���~�����i��0�Y3�DE�������g����efn�Pg���a���f�CӦ̚�����<���䏽ai�����Xv��B{���� �<��ž%�E3C������	�=Ԃh�]\<����2�?�����R+y�,��?)#����}{������+�i�Ҧ�}��I
*8zM�36N&�e)2?��8O�������o������9	����d�,���1.���� �,���U�N���,j�E�z�ZC֝L/���(�Q��{V�����i	d� �w������+!��=W6��eޔ*{Q.��u�{��jp��k����#Rvmo��q}}kF?
�gIZ�A)��M�/� ����W"z����������"��Y���d���1�8�3��k�ﮮ���NƓ�$%��R$Hz���R�{V� ��8=ۇ�.����|��q}�����?���@���}쨺��ڞ���-{o�ڷ�"Z�C_T>w�����{ug�`?��I������.�;�.�(�ۿ�s4���J��>��d�H�wI�]D��}���b�<܀����3+u,��{l����Z���Y���y��斪�HP�	�؂@���.d/�D�S���ʇ��d�����"������b1�H���ek���s:_��ܥ�V+x������!�`�k�ݖ+�)���6���y�Mp�{Ԛ����˯�9�3�B�[q��}ć=\�S]%�Ѧ^W�Tyućh�{F�_8j��L�ĽL �R�拳Xr���> `i3��\F	安?�]ơ.�np�W�g!�pe��0��'�LrҺϪZ�~r�8�N#��+��,]���m09z���S��Jrİ�Q��$�s�~o��~vley���x�H�}WD�Mˢ���D�����Xݤ�hM�U4\$!��D������'�\��*2Y�}vyN�iA����'5��^;1���2�T��![F�]fao�c�1��ŕ�נ��R���"׹#�7\������y��C�>�[����c�J�]�k@y6$+3H3���=T5�Xl���"n�1���>�^K��>3G5�������W)��|�#w�f�w��������,*�M�l��6�<�������=��s�*��xV�U�>+M�L)�qȘ��-��v�s��(/��\ň��cc�9~�@-3�gr�zh����GSpP��ڣim�{�J�	��/T��hٖ�v�r��%�XҞN��P�0e��hE�|����2R�J�PF�����s���+��d�2]k8u�K� ՠ��tu!'�9����2����ެ�����eؤ$
�a �D��\������	���}���;ͅ����27gy�l����G�a߲TD
z�2{��A�Df{6���a�Jں����E��� h�Ar���;{>�����l��;�)��;g}��������G�]��Ϛ"����p�D�9d*-es;;�=�鵽��LB��hm/q�=r6�.͉�B/��X�g��}8���~]�������7�!�c/3�YD�&�����3������4"����ѡ�H!p�8)���I��2������S	Jb`�r�r�f�(	�OY\��"�ɬ�����+�U(FU�dm�� �Mgpn�%�A�"$/�1ֆgAK����e���o �w	�{L%�&f��ݤvV��*�'����l[r�����Չ��i�W��j= ��u�:9�����=H��2��>�^<3�Q�,���Fwij��E���Zڋy�WubQ|0�@��d�Ί,~u�\RU%�5����_�-R�ʲ��'<���iv�ʇ�A�Kt��[���jS�!�\NE@~c�NO�%��+Fð��\�|ah�f��X�p�v{r����mZĽM�����!j����[��<hi��u\�1��7:t���h������(;I>��i��aN�"�)\��15�`>ܸ�ÞS�\QT���o*��
0i�O,�8⻛�:��E��J�A�+���.}����/2�[Gz���8@:��lpy�0��s��^��hP9rX�nx(j����;�œ��o�p�]w<|���^ht��GS���ۄv��=��D�+ߕ���}91wv�&�0	A�[��Ï�������d0!Lɛ���2z��(.�~���Xn	E�^B!�2k9�ח"I�f���v�G�lJ��;�1�Dd���I��_-�����j=RG@PZ�U�۳x}�Q�=�'L���0��?m��n�?�-f�]'����3�$�8��~����W��2��m/�,�c�*@yc��=שj��@$)R�"[%#n��gYW�ۄ�hC�2{f[�Q���f�W7���q/m��@�k�۾8:ۨ�l,����
l��_EL�g�zۮ�Ft w5����x�m&/Ȋ�+�O�E��0�2C��Ι�?D�Fs��m��do�����W���'^��b��d;[y�S�^?N��#&5zq6�c�g�\��0*�[L�_��QO��pߗ>>����,`	�5� ��{��Ը�	��˿���O0O%,���j#Vj��+�둡��'"�`R#�1;���ԉM�N��y_~o���W� (?%��	I�����H}�(?�4��h�|����<VS���@��r����P.]K�g�#�*R�ӒZ���	�{�B���W>���v���l5��:�,�+�C��v��T*n�·�T����؁�N��c�p��
���|6��^F��1��aq����WB9X��e'z��p�{=��Q�2��T4�Id�7��q�|ߎ'�?)�s$}���?���f�{�WJ���p*��|Du%j��Ћ��;c9g��pbƭ���O+F�lT��HB�6b\;�A�hӲ[�(Ďtx���m'�z��gt���µe܊��ZՑ>.�C���\�f�&
���§�'�M~�� Hw&���E�@<ϥk��8v2nT��>zr_z�Mzqs.m��捸��oc����y	���wd��gq�87KKd�P^�' �����FI�Q�R��T����u�
����C��˿(S��G�o�kسg�G�dk��CT{n����d>�P������`{���k�\^2$߹���!{��>6'
��� 1Fn�m����5Ϙ��c{��6�����d�)3�#V�e̡�IS�L�d@B���c��^�2�L�f���pz.�9ա��=v]s�p��FE	2�ʜ+m����������csTm�/-���΅N�1�Ǚ�Ʃ%o�+af7�a>*آw��S}�o�F�RE`d{�xg�iL����w~bk6[�r��'"�zΜk���~�b�QAb�=��X�7����w�Yg���>�ci<U�(��b��B�x7q�@=^7�����+��ÿ������S�h��rX$縡U��<h�"��%�G9a�N,���qw:	I3"�yU���n�$[J)���@�!�U�����6�.���Ri��'�����V�GAw1I�,%T��J��JY�c%�K���˭ց��5>!V:��<�5
4���x/	Vx�S/|l�%���BK���a��V*K��-,*��7���2'�~y�`��>\I�5��-b�����g����e��ή�����'�
�K_dFU`o:z�D��<"�Xt�sfN�l��/���Y���j ^D��/q,�Y���J=(�L��vS�A�/�˗����]��GGf��Yr���)_ W6�O9|���ui��}v�������u4.�����2R�qH��u�	6�ٶ�#����P���(9��,E�I�(����ۚ�ؚ��|6��,]c'3H�l���AH��v�d�ȁ��{R���������|R0����ǆ��|��w���e�P�����&�����!`�"��*�j)!�TQ�U��c�h�_�^Je�ׯ߆���{�G�D�pO���_��gn����]���T�� %���)h��)�*�!�)-΀O!@���ii�]gt"2�	
N(��Uz?��q:UovgAX�.�-\��H�MƗ,jo/��o#e�ʁXS:Z����c�5�a)1η9a�c��$��L�%\��۔�ww$ Y����UTr���	#j=��oޅ����Gǚo��}���v|&Nxn�E���jO2M=\���� �8�������|�%�1��H���� ���=�3�-����z�E,������0��ɆHy�y��3�]kGT�G���/��G[�a@�B��#�s+�U����8&�D:1s��X�4�*����>@��ףp��0]������6�$�dG:IA�а���Ŷ��Ź��~��Aꗦ>,U9��V�׮{�1�m's�l��X�̦o��=k�8Q:o��	�l]"�{G�u~&���cŖ+��|-�?����1 HR���4ݐy���O�TD[ ���uӛ�g�>8wgӱD� �(tR^�Ҕ��s.H]�=�ħ��+��f���z�v��ob�� ��z���|%��]�0G�؀��yx6���V*�,�z}�����a4'W���	���܅זq�f���O�E�������w���BC�0�W0VI1�l��[d�0*�O§<���W�^*�x�|���G22����o0\Q��O� ��)�3͖ڐ����|���p�d�E�I��+�����^��P��x�J���mS&���,��̽?���	8x�="¯ȟ^R�,��`����}���%�ƷB,S"��f�®���L<��)�u2r� ]�(����#�����kE���m���اi|d��� @�!���p�d#\�0�u���C��Y��֒�QfP-e�0Z�v_7Z��YA�� p(Ia@)��3v��Z��m�thA%D��dm��aRc���-����N��NeW�@�ܞ��"��ߴk�2#haƁ1x�۬�T� �)1J��	4�F�0�+���9����s�XP�Ѿ���/>�<"�T�$�����c�Z@�т����V�-͹V��-�����p||�j���5�4�o�{�ioAk��JU����)e�U��	Fn�%�z ��C�,�C��L��!�R�H�0�!���4J8�:P9v�av#N9s#�� 1��lA�L}�I���D%�T�b?`�^WA�Z��y0�VM�c�.�w쁖U�D.�aW�@D	P
��{,b�r���4�G?�N2_����^
�@�lbEV��lz�q�{M�`�a�q��;8I�(u_�-	����u����2�_���ys��o��*2�i|��ɒ8{|-9�hk�)	p ��S�g��&���3�4�Zڽ������K͚�e��t�^���������mV���h��4������9�&d"��EbBvƟ�Q�.F8�户�����w�z==H�>WeWd
�OCnNU|�D{���@��20��r�wʩ'N���o��h��1��k�vɩ��|]3���L�V� 9e$�0N�|�o�1�/�l�7"�6�!	�7�^�sg�b|)2�ןޅ�(��[��lmi��*g֓ٺ�A�	����<�4)�7����O-p�_aM��,����O��O���b���k��z�s�*pN�q�,c��5x��Y8<z���^J��gO�
�va����T��ܣn=㾓�t �hwEG�zNlsCF�(=T�B�hM��v�du���F��\1eQ٥v�k��ӈ��������X�y��Č�`M�G�6�-#M��{��9A����������-�ߌU7i#��9�J�JzKw�U�[��PQ7}�[x�7������X��������:4��Js��H�}����S�0-xB7�[2,�j1�z��H�;s��JD���f��I^bq���2d(���uDE��gbh{��i8~���F��7��}89��������u�n�5�K;���BT��}��2\$���ե��Ee�!Է�}̬kњ������}���T�鳳�v��F�#G#\�ev,����K	+�pz&�oH
����MT@�+e��$�L���{�Y`Gb)s��ﻊ3Lh�����tmW��5N'�yc����v�������.4�a� v�}��~��䄖���S�UҔMKA͜63̙g��d�-�V�] A �XE1����C��O�h�9[�5�N��N����	(VĲ8�;v���զ����_�ѻ�eӧq�#�Z���X��^�z�FB�@!.�I�-��QA!X��iU%'L���hpR^�}�ڱ�y-��4��
��M�A�C@���;y���	W���x�^\kT��#�R}_�N���'S���m�_���z2�塓v�RE"�vd�L=�q>#�1��\n0��|�c�lBnn��d��X��QcO3B�!>1ci�D��ƳjT{(�}�����D"?ڰ<��g�����L��h���9��2��|6����>�"'�>��������Q%+I����Y�<"43�<%8a~a󎲶eg7��һ�gf���Q@�|��`�u�ahYwF��v8�I%Z"���Q��+��gq�ϕ}{oӳJ�W_}����޳L��؁9��Z�=��L?H��؂/��*sԥ4�#�/i1������I�E� �kVx����س�D���[�z����P��������Of���eF��"
����`����e��_~��0,�/�h�55}��cV��h~�t�R�H�ٛWEZFy5�wƌ�3F��p��{/3BEO��]>�6��(m'�߷��I#���|aʂeiᆞLd9�(0�Y�E�:����WfA�j�=�z����ty��6���p� P"��Ui̽��	n��U��	a�������	������Jͫ3G̗(`�s�;���7uC�c��y��@u/����BGv�ע�pe����6U�!ڳu� 2���qbO6Ӟ�r�!Y��g���R�E�
M�\W���X��>e�71��������l�<�1UM@1�3�(Gx%�����(b�N��y, ���c� �U����	X]��f��]}W;�8�'/�[�i�����@$m�4�(�	�b�_��B�!μ�ىҧаOFQ�[v,�`��\��;�3|>�����W0q|<7�;���u$A��>8V��({%`n�/�b���l�c���l�;T�����TD�I���%'���C3�߱}�;�, ��hB�'N��uG$b��oM����Ty+����K��/SQ��z�b�(D7N�}��aA/��txa_����)���N61���qH�At�)"�O�]z�6��� ��3���?>V�}�t��2�`�,��q�)ѳ�&Y89;-�}��T�e�T�I��=�#���e�C˔(����)/]��nA�����$�f����e������k�>YH�M�8c\lA��&DpV�F5���r�S"g���e����R��%�N;t8d֗�R�m;H���� В�KKu���0W�T�[k�c�7�b�]��dA�^ڣ62�ڎ���^����8�=��p��$�u�s�?�v��<�(�Hi*�l�f�	dw���.�Sn��^�zA�C,�����'��B D�9��՚h����.�����g�g�E��ǛI��q���:W�Js��p�"��tڵ;�5q�q� ���T�aӲC��-��N�hW<��H�EjPq�R}�����d�I�����#�[����ۧ{��xe�_Z��k�P_�����O��\���Cx#j�I��D�kYi�{'�-"�H���e�m��.�L���=U�^>{!^wph�~��p��c�j.�z� �S��N6���ke� ��],5�v����l�f��kZL8�i�|��^붉e�7X	�T�9�az��%�g��7�u
ԕ�8�߆�Yʀ��$��7��0�ߧ=CŌ��B��>_]d�1�|ȯ�����E$�q��ή]Ȁ�J/֖��M�XCZ �"������3'����a3՞!(Ej��a-	e�#U0=pF�6̆i#�)�'��H �3�ݐ=��0Δw��U���D5��C���Py  �,ͣ=�k��-k��;�ɩD����`{�k!�`Y�9�#�u�T&	@���TᔵSζD��n1�?�y��X5He�4-FB�������o��EN�6�틼�JI\��"�H;	���E!@4t��7��k����;�PyP�prS6�ť� �ې��D5oߪG�� ��=�"Hx��Ge��j}��[fz�L����6#�A�^�h؝�
�<s��oz�֌�R%�3J'v�..,�U����J8�� u������Q���
'���6-C +<�@�Bߚ��%�VQ#pnS��-{%~��I�%l?���=��޳���~.0����8�B=8�ڗ���v��"F?X�,�"0�L_WN���>��A y���e���<����2�b�S��r��D�4f�3/�(-)�BP_���u;��ּ�Yt̅��V��<��̪W�	#�����Ǫ�F�(�Y屽nv}���޶"x�T�gsd�u�@ᘐl�Чϋ�|��ɢMY����:{����t�*�1�����@m)�ˀ��U�D�- V��3Ҋ���,�[���zGu:�sJg��^j�d��G����#��Q�܂�gǇR;B���& ~|�����p�R���	�z{>��NFf�a�+Š�)�nC�`k܁���L�.�����=<��l���X�0�r�B��������Sę�B����#H]�b�v�1��7��2��G��y��E��W2��wc����y�f��8�|٨�R����Ftd`Sۥ�҄�(�+������|�8����O�䛰����H�Y�Ey�>�
cP�*b�R$ۭ�Ȅ������s�9Ӆ3��v�7��QME��S��)?�~-��|�J�q^����Y��S����#ܥ��5�f�]�-�`N΂eL�W��Ӊ&q�|,��c��m��%���=�PVk6�"�%��G�ԥ�d�hONX����$]>��h�4qaP�5�gS�N @�Nx�������s�i:E|A�,kx�A����H_?g=Tp�jw;��/rnV����5�Ԙ�&���՘z��6�n�������G�'D�d�|r��II��f�ᮜ$��!��G�*3��0�p�8D+�\������U8=9xB�;��'Ї���uZ2�.{�墅e�C��_���&����4��8�d�ݖʳ���f(Q���
�4����0(��.J�W�=�fDp�t1����,܊�v�(����I+ �3z�[�m��'�ݏ�K�L���BA��n8��g~l��p d48�2���d9`�N/n����X��\ƞ?	�v�7���E�
κ��g����]�(w,����J�^�mW������=���3����L�9? ���5D��(���f}��� �$h'm�z2˫��PZ����G��Dv���������B��v/S��+�gNl�ߚ�����O͘��jdIP��;�j!鷳q��2�jC݊Z���5R[�ke�EY�l�>�dDY�1��!2u�aL���5CslQ��Ã���Ga����٩9{�g����Yt�r~�64&4�Ϸs".b�*Ę���|�@����]�f߲�.���(�]�s��gM&��."! �
 `���!��O�{P��O��I@h�Hx#�H���?��]kK���[�f�@k�[ 8��1����u1i��t|����w�2�Q��vrr�*JV]f��ʚ�_��=U��\�åo���ھ�攣��KVD=�L�z>Q�8	Q�{�k/mZ�l6�����|��1�����٩kض��@Sۃ��ۻ��ע��*�������-�B@BɃ��3��@4$��Nt�4�Q�k��`w ��Of�?�K,~1;UI�{��":R��o֣�Ǉ���P���D䈘Ded��%3ǎ �j�Y�H9I鹎�W`+[�+UrN|�+�u�th���̾�ٳ����s9O��h�^3]�2ظN���U>.j�p(8X��.�G���g�����?9a&��g&od�q��A)y���@��c��G��D4�����3y� ��޾'��R��< Y5{��N�)-����'2�VX�0-{�����*�
ܘ�_�3�x	/��o��r^�K�YZ�>S�z��ќ5v�&D����T:q8�E�K��7��~g��2!�*h�B�R�W��GG�*�K>M �J�ȇ�>u��ٸx5� ��-:�/
Y�V����V)�k��^���,x`f��T%@�͜������o�a��e�zۮ��ّ9s��g���q����9��֞�9k��h���>��H��-��Vk���E����p2�L�O�I� 6/�Q�4~��cwe�l,}v@��L����0�X������\){��$Ș�ؠ�af�*�*R��n���C�ߞ+AϹ_g'����.t����7ڋhmH`��h{�`b�����;\��3��Ým>�0c<�hI�T%��|�B�h�2#)���&\TN��(E.��F}0�3�oS�m�ed{���vxn��сD��E8��^cFg�eZp�,�,F�1�M���l��ǘt���}�v�E-�������qdY��	�	�Ul3=v�ht��,���HWwz��,@�����a��w�H�Z�R�����,�@fd�9g��@�F�swЕ�9��ڂ��򳸫�k�Iik��0`��l� }>��i)��󫧚��`��pձ5���x�C9}��1�d:��|5�k%����G�K_ctB����f�[�I��nHڰe=h�V�\�>ھ�&)��i����3K�!�������*�~W�6.A��3����.���F2�{�+���鹒u,a5��W�s���hʘy�<J�j�]��r��]G;�pS�*�?{�J�^� D<R�R	�tܐ�^��g<�g����j�b$&�:J_�����T�MUܴ�Y+t��J2����ak��X���R	SH��Y.7��Tܜݬ0w���#�$y��\�v�q� ���:p�m��1�OϲD(�ݭ~�J8+�&��+l<I6C��$�t��O_jf�')�M%Bł�-�yb̥-^���;ٱ�sѐ���շ����UyW�K�h��n�>�hf'S��G尬��pLqίZ�p;2�E|$�c����UH�Q5<9��Y2�i����-�g�re9�7/^iij�3j3�Lc6,��R�>�d�S����Ra?�=�v~�)�z�"l�m[�x�-e��;��N-�No.]h�)��_J���&����v�<89�����(�����L�`Ѷ=C@1����v��:<y*Tǂ���"�C���&��B�giS�Z%��)
��g�N�j�C���њ/�0~�M�vm.,� @��#1��7����Z�Y�ԙ}�:-�i��qߵ�Kd!頚�$�҂��a�t�R�e����!�]��:��Tge>�\E�v�x�,h�	lcmi�1-DC�b��N�>��jl;�:)���_m�� �����,D��`x�{�o����IxytN��Z)zs}>:��>��KkKDF'����	s`���#�ޒ���`�=���2��\�u�鐩"���aT: �8�쾦K��,pn\��{�p3���R��QR�"�X�Z7zMKXd�A�vx>�=isX�^�e�u� �����P�bS�&�|]��Do�B{$������/~�!��=��)�d%�|�$���nvu'g8��f��n�1�-Kۋ������"0�d��w�S��	�<g{��gΌ�$O�)Y��9ziυ.�2�~����Q8�8S�.��i�.(�[�F3�Et�����|���f�3���.�5[��o~�����K�mI��~��pCw�BQ���߄��咊��o��޽�H��t�L���ϵ̢R�/p��z̴�Y��v��|��7��Yu���u�A�5����J��|.iL���C_ų5Im�{];%Ɂ�u#a����"(M���Wd�Rx������L�-+�#�jEU��%���y�R��U3�T���&(�U��b�E�`A�KJ{7�B��S����?�cx5y�Jl���r�(���BH�bz�V�ܙа�t����?I�U{�+�cשG���*Y5mT����ښ����c��*c��Zdv��ޱ�"��V�z��v O���j�M6��/͐�їΔ�����t*|V�s�<�"�J��=[P�i��������ݍ��PGp�!3f���4�W;@f��z*��vx��O߄޿s=�N.>�t�tOU|S�Z�n�́,��o�O+դZ��4���lA��5��R���c*Na�3�ڻ�j�Z�Q2���+�u(7�9�@�
��[� QѤ�B������7�nײt8�HK|�'�{=dKi��V��$�B�g���+%�!�M�jQ��y�ud0�'��m�+�kQș�
�#K@�,`�ߑ��GD�g���|����V����(����8�E{M eOv����3` Cp�m� ~:�jhh�ꎭGa�{�����*i�f�=+�qŒ���܈�K�9�b���e��H$W��|4]�Ʀ2��d��δe� \(�=����Pω�Ln5-���@n�j�D����P��Z�G.�9D.�\O+{o��j��՝֘�Fd`��%���a�Tk�'ڸ�¡�ȹ )�%�YXs;�.-х�ݷ��J�ΡUr<�н��$��E�P"\!�[��(F��pt�v*A��:
�����$R�<�,�� ��G���9��1YzN��/�L��*�\yi{2t��0�-DCpv[C$F�'y"ϦJX	�N�`Y�x@��z�uZ`��3�����%J^h�S!��N����.`� Rȉ�JPYh���B�}~�9a7���׃'n��b�� ������g�㌘�C�D�,��3���up�D�u���޳T�l����/��U�Y�P'���m~�B�.6�"Ze��!�g��������o��g7t�C�l��I�QvԴa߼|-2=B+�����վ^� �_��1nKRAZ�4��#y{9[ʖ��d0�&`�ԏ��D�1�+�4J0И��<u1ˬ@a��$'(�j��sߞ� ����v�fRe�1ACb���@6A������.?_� ;��\Th�Q��I���e��a&��\� \oV�Sj�iT�qA�mz�������A�W��T�vK�j�A��A�A��	5`;h���`�yx���N�F(qX��PpZ�Nsӎϔ���4L|���
�f��	����B�
-�Un�qc��;:;�	��k����v���EogkWq���Q��;Zpľr>+ë���۷*�{�l�g#y$@��|�w�<}f��k�ja�P��,Y� M8�H�  ���S��u�G�j5]�k�=&�y6�@Y�2�c�~��:{���|d�o`�e�Өcf�����Zv��%��'ak��(��P�+`f�#�k�����|;$�Yf	`�(ZrWb����_)hj[��-+'���3��琟������UHW���������u�'�fF���	gA��>Cgw�GHp>˶Z� ��{�	s�J��ԑ˛��qb�x�&
E��Pр��Sw3c�W�!2*�:F"#K�n�������^��ucg4l���6L� 	@���l���O�v��J� t�HR���t��Q<	I�ۇ��;{��C̕s�v6�:��*`O���*��N�u��:�֠+� ��>vsKN���.3{�璑�z�����M+ըp`kV�9�Y�)(�g�pq�i#LW	:%,��ܻ}K��-Pc'�\�r2=;��G�����p����4{j���H���c=�(����Nض=8���j�� �+�}^�|�={�}�k���oép.󈼖 �,ko(��=��;�q_��ES�/�ކ�$%u��:'u����_?��b��3���p<��=W��3�R-��^�ϭ�dI��?��_Y�m�
�Ge�� I��l����ɓprr$> �~�B�+r)�W�錚�L<�\�*"���MWR�rK��sH�SQ�-k�;v=���ҌvZm[�`�-Z�<%HY��1C
nV�K���d���/��Y�[�TX������k�r&R�TbR�mA�ὼ�"���`g�)ITF<�p������O4�H��A�y�:=
��^�#����Gt�\��p���<<����%�e�0�M�2�����<357��D
D�
n��-B�|A��uo����_+��`U;G��r��.Њ,J�������������	�� �<"0$@$w�"{&h
�t��,¡�
_�x�u�������q�m.���pH�bv8��R�@�`ږaԙ��*
�̍�d>-J��tY�Z(�~ߪ��*&8��~[�^8�Ϸ'�H*xP�Q��vpr�wl�m�ڀ�B�*L)-Z�.�s��Xձ��Y���*��~��65ݪ�M[�[o���0�X3׵˝��w���D޵����]�g�&aN�ˮ�vl�"���vm��U�HRI�r��2��CO����g3�\ �@����c����R*��]������,���O�P#�؋��i��4(X�<O�>���N8y�TU৳S�ک�F/J;/B� Ep��ٰ ��to]33fWFq\�9/��`|�4�JR�}��²�V.�	.k��EjZ9�,�e{a!��2
�=	�B��73]�+�21��5��`��	>�db[��v�mu� �Rus.��k�ٳ�e��/.d�އ5�cgסT�v6����I����������뿩��,C�}J`p�~���
�K��oW�K[W���z���0�k��^w�g��6�ON�y�^֒:��6�l'�M'Dݐ4*��^������jҽj�e�����H���U�Z±�� �*[�9ٔ^_�|e7�f#������������`�I�\־i؜d��
jU�~���Uq8�핫ah�am��wqۮ��©=X�}�9x0�e��i�m>�0������J��%�_Z�����o��v0���*�hep1�*���Y˃���&.|N;|i���߉z���,|����y�hJ�&;?;��C�k�M��r� ��������)�.�D�Q�)"jQ�B�\n8��f��]�k<��=�B%f��^Ӟ�I�\+-WZB\�{-���l'�d�^!y9�;U�?(:����2͡ܖ.Q��,���9�y�Tk#$��"U�Qs�P�A-�'Ǉ�7�^)4kR�%����6jA �Ё�������.�beۨ���͵��5��.W t&�}L3� �}�_�5 ؞eE��t.d.�0ޛ�d\���E.)�xI=�
�қ�`ڪ��o��s��w�$�@-Î�é���LHcR�#
��%m^$j�2&aN��b�E"l����9M�*ղ�׳�s`��J�E�/�x��F��֧�m��eAjU��>\Ye9^;n�	�,>��&�:F%G�#���Wm��t��gZ`�쫐�|T3��G�Tr��nB^ՠ��V�} ��F����["�F>��c���wVY����N1�:[�]��V�6�,D7����Ȥ��n� ���Q�F���\'����k���|fφjN]8���4���V�0K_���������L�+�����ވ\h��J�EK�q�$�(�7����N����#�c���?�	� ֤O�4!�l�Y��ٍ
[��T�B\�Տ�����V��`'`��3����|�]���p۝�Ot^�1��=��>�^��~�s��I,O���g@ߔ�3��zM��~Q0lh��#�����}ˮ�R̲�o�?�)����ZM{����͍T�lʹ@_��������H�n�u���o���s���>˴JK��t� )IB�š�Ni`�B%<Y�E�`�qUS[8�%����e���m��2����-��=ǱeB��%��!0��wgCz�R���bBk�9��NB	���a;�p˿�{e��	:����â���	�g��e���V�BmYf��8WD�/m+@4����ZY�E݀
�Vl�|�W��a��#߇2E�DB��պ��X�Z�D�[1Z&��+�2I�%��Z����2�Ϥ�q�ϒ	��&��6�$�3}>���Uv|�|�cױT�[ʠ]n5j�%�������2�t�Kˠ���6�M=��X��)��f�r_�T*I�l@����:4�0^;M^���z�KlPc�:.�m��x�t'[2:��f1�X��ծdL1I�yG�����9W�Lr�Z��BK�'
Av0oZB�0�RgZI	��'H{�,��ꬎ��e��=�c���}O-c�ݬ�����M(l����]���]�S��"�Ҷ8��0kW�
ہXfbU�*�%�����A���GH"R=ʾ�]�s;�l����0���Xj���-J�^�� H�d�@�'�I��`(��y��fV5�Tc�A3v����/���
E�����0�ɇϏ�,�~O�Q:Si�H'z`a�2���{J�~h{p��M4����Z-f)��xj�N���X�1��vVT{}��4!uŵ���v�G��v�]!����Ϙ_��ѐ�HJ�HU�d�6�źV� �[�3�=L�>���	��{�w�z��T3�/s�{���t4��u�k)�\H-x�эS@\7�ItV��:$>SU�
��Sv¶ �-[���g{N`..?+Ѧ# �e��A�I��w}�e�B��2MbG3D�/<��R�9Ͳ�:���O�D~Ư�]	7��'-�M�J����.�nڵU|5�04�kGV"�O����e>�L�Ü�!ܸ''G�hz�ٯ�z����)IfC�(���/ʥ�HY�9+	��z�U]�����V�B���\(�l�Û��¿����ɳ�.I'�w�����Y�p�)�����7m�2fRh��__�{���o�t��v����A��F�
 �
����D �R����X(�R�E�.TY1C�WtP����m�݉�p�Ro1�~IJ��
��.�,r)�P�=T �j�no�Vr��-¿2��b�X�|v�"�4���;:���{��2U�z�	�b�p��%���i�h��U���ԩa��'0D)Jb�:R֒�Or�&��Q]� �w\���kw�UK�X�0�)�pT�&����
}����+��sn&�K���q-��]Ჩ���g����в$e��5�\L(QK�@9K�����C0��D4\��D!fS���7D�O �,�ܝ�*F��[j���X�ހ;�ɪ��{��[��:\�A��{���Ī���%\v�aׂ-3��3$�T�HF�J'G�2��嶺a�pg�/�R�e� Bb���Y4:���@t�K�"��+I`0ؙу�	����Hc�>q $��@L�/)����y׸k�}$���6�c�i-6�I��Ʊ(��|�ϸ�|����GJUvn�v����w5ݪ�5܊Z��C$��Ԥ*�\��G�O��Cw�X��T|��w�I�!�e4��=��r��'m���:�tq ˲J�$&�ݮ�r�$���Aa��O�4q[C�ڍ$8O���W_Y���d���!tÙP�SL�������l�{�-�N?]���g�c@_��|x�V�Bk;�^�h�ʖ�ל}3B+я�8|��>}<M��?n��x�G#���l�Εբ5�g`���a[ϩw��,�+�9�_/��s�Ҳ��Û�+W�ܹ�<���{TB��������'G{a���M/���i�4�+�A��B�{
0"���eIT���͟��\���E�P⒝�^�%�s�R���*������uOL\k�*�í�x�@ �(d�����\����/�B-t��b���n�9-��ӕ&���K�pD'�R�)�&:�@���i'�d�g�o~�k�<�j͊�"�@��"9hY�+5ӈ�ڟ���Z�qa��sv�Ҍ�D�Z�DN��,���,FZ��O�t@�w�ނK�`�77W���:,�<wr��9/>�Pܖ2P-`Dd����ծ���������KP	���W%y�4+�@�-T����2��l�T�M��h��3J�6���FN�C����L*1�9�>���+Y�*�_3y��)3����m��Y5���\��D�h��7R�JK�Y7	f��Ү�+mM��h�-Y�ߊ��^��Z�tX���dR~�z�}�����;{ngP>�A7��uiIO:	�5(���k���X���ڲ�y��ŠM;�
��Q���V�"���gn��s,���:��Z��D`I�Z�
>�!�|  �N��̡�;���_������?C�Q2L�&�.1�slTIz�����b-�6,
��U.���FҪ�%*c���V�@�p;�&���/:JT�7w#u�&h�[0�6߻�M;� PC�iT�d�h��>�`�svt@��ψ�1
�om�;�X{G��*<{mL��qC�὘�f�FP���Z�k��@�A��,�g��J�_���P(�*��y��߷s��2}���U@�ىz�ͬ���<�+�F�p��s���3]�or:pT��_2�!�Z�~f�Z��fI�Q�T����V��ʎ�	�g���F��T�4��q\����zP̈́Y��EɂW�F�Is!:��#���n=�dZP+��������Ӆ~����pa#��\ }��Ү*M�2N rF�ޗ�/��~�
��qS�*d�J��۩�d��fɴ~o��͋��ѓ0�)e[>�<0h��S/�Ga�U�{�;NXeݱ�����2�c�9����̖����eJA�	��2� �R�j)���U��~@�xY؝V���Ơ�|I|�hZ/^	#�Њϣ� �Y�p�oF��� ��OE7x?�u�.?[0����v/�PD��ZA�q�ʥH��3JrOl���4؁�؄��oe��Xղ�ӡR��Q�ǌ�%<��q���CEϪ�7h9j��1P�~M\�����(� ����T� U(Jkt_ �(�Ϻ��3�B���L�(�+����`���v��IH���P��4z���
�&s�xݨ�U�f�q碌��E��+&�H R]r���k���ځ] Y)��4\���ե�ѳ5�ϩ��Nͯ�����`Uh���8���Ԫ�"&"��ŵ�OՂ�6���X(*����|��z)f#�N��m����{r��Cow[.Jl�uE��Ee�똤��;�����m_��J4���sYD����!��$5h�#��rz�\���3;���D���:����7v�#{���$�����,�s��U�5mp�%��ۚ��~_b�H�5^wt�$
kW�#��-�@vO��f�w*����e��o�c�9Z�e^;�@V�Y^�q˞���X�$��k�c"��r6S����ý�ؒ8����ؤq8���e�$]i��&)�=b	l���	�x�a�d�S�]fq�Hf�Ɗ��������;(���3�ռh��v���dÌ�#O��~T!��	֍?���ˣ&yZe�_H��=-�b���P�m�.���Ȇlok�~�ۿQ%�	�������͑t���%&	�����n��o0�([X��J���	���|fE���#�Ptd������]��pG@��	�s�`�{��F%-eg�fa�r1
34��-��E��5Tf^d�H���^X�v���[Y�t[.�A�E������b`�U'� �Q�S����a�8X�i��ZVЉ��M�&�/�_��Q��)W�%u����}��/j��j�����Yx�x.��7wd�5����Wz�.8���V�h5(혊N��ع�Ӊx�M^E�t0���,*�r�)����y2�r(�Y����M�?���&�q�
?s��r�1��4Q�WT��[�� �k�j'�i�M><�U�k\'z� 	1��-�l5���k/�NB�=����K�Jm�9(���8��g�뇳խ 6����
v A�B��n�4��p �l_Z�v�<�P`��v��--�k�[p�[�9�.Z�h�T��,q�Y��ͽr�G�v�����.t��f.L�+���Ba�~�m��( ��ݳD]x�6��8�!�����Ց�z���������(���ݝ����<�����g�l3U�E�N��*kq�[ҭ�m�o�%��h,]�/��R�QZ ��`��p�S=�m��.���w�S��m��#ǝ��\��Y���I�dw���fwg7�X ��.�~t��p=��� �x`�!�m�.*�&��"˾�����4��s)�V���JgF�!�G#98�D��?�d��l[�$&�����m�N������l��8F-�;�"����� �M{ V먡Ѝ�H�F����
�T8`9KF:Y���5�~��4�����s$ɼ;�s�|!䒆����"� -<G��{�����\ER֏.����c��)3]Y����VORm��Ƃ�|���zM(�|6H��V{�Q����ě�������=q��r���p����8�	Uxz�l�����"���;�l�� ����8�f�ɑC6�?��.|�(�G8@����^wv�nض�{�u�����'Yձ���J�tt?��x��;Ӊ��2ix��yc{.hǽ<�Z�Z '!��aLe��w�Hc�T_̿�S���63���\#$e%��!��שF��QHms//�, �v �<�d9s�<y:W�vz@c���v�2�Z�lPF�B�	�i8^�7� ��K���#� fg�Ӊx��E����=���mL6�R׶r��nOA�d�k��t� /��ݍ�&�v\�U;�P�<mh��Yn� ���Ul �d��X����o��W~��3���~*2�6�%��>"`�T��+�$p��Ė�_�{N �]|�։� :.HK:��$�=���H�䑴��l�$�0 0�O*���~�8[���yD�O�| Z�0[�D��5����h����?�c:��=� �U��U���W����Q�1*�d�.� T�e<3�q�jvW�t�$�<����ݽ�b�bt�&��E��P��Yy+�� ^��$�=	-[t��1�[�ugk���s�?�5:�}6I��kd��QV�_n:T:��/$���3&�+�u��E��Q��#1G ��m�Ҧf}��.�=ܩz����h��?R����0�}P�vtOd"A۸\�z^&-G�3걯{�7_}��Ei��e��0kE�F"�eߛƾ!{� ���:�ڽ�O�%ؖ nn%Jұ}O�EiK�=]�2���2x��%�{n�9���<��>�J ɱw - [�%0\�d�($s�nAi�?�5�7Y�$1H��ȭ���]Z�h������72솿����	�y�={���q���w��- �@ ��Bd���HJ0d�F����)E���{OᚲX�-< Ӧ& �(��(��H��l��V���_O)i�QJY�W����3̭����_��͛p����ٺ��
��X$��iю���Wj׬w��k���a8����%�:�ZF�/5��C0_�B~���ւ�fvR�F����>if��)/c�Ʉ���^"ص�Dϼ��KI��Փ����������
�H���;���E>���m��q�a�
?���(вۘ� ��ɛw1U�H.#�S���t�+}��bk���g��3U���%^�H7:��BtW� �/T\k[sX9�u!��o��o¯��a�n�pS+K�j�IëՁ"I�m�`
��T�y�I��taz�j�A)��9e���	/��e�[o,:��HoH3��"��
���8��QjQ'{��w<��k��K�s�2Q���C��BO�QQ�h��������Sun����  ���H��ɡ��S�-��P�p�˕���3�[�����:�=��
nc��.$R�k�g][�p�z�{��O����Q��>D����$I#:=�z+�k�1� �.��C��L�V�O.�V;��a�3P��L���7��$ni�_-Ƿ� �����Z{ z�̆9(6dC7 �?�Z�$���̤u3��޴�zҕ�>&Y?�8��1v�[��:�w��{)�U��-�B.S�R��,����DzI�+u]��^z'�5��lB��+�݀�tD�./��M��]��oFu���2��
<�P���F��>�D��$�6��y������p��'V�$�hX7nl|n�XWH��.��/H+/��	�}�%��7�F�C������j�ˍ&t�n䎿DE�k3/&������XR�?^L���"�9������7\Mڐ���jv�*���������$*���<3���T���r P흜H��iV(g�I-U*�?��&Ӆ`�۱��id�}m������즚��_# Ӂ'�Tcpn�=�������b)���}�'��������$<�9�����ܓ��?^ڡ���"���>ugs�j��������Vao-cA���d�l�`V�gcv� B�r�O�eI�R�݁�ʫdC�w�����B!�LCmLة:��q���iGц����F-�+�= M7zr~��VS�U��E�|,��4qj�Z��#�jЬ�6�x�"���֏\�F�5��R&���\m8i��Zvx�����wk�'Y>���Й���}���5c��c��2lF�w�i��vv�?���K�����ۈ�	$����
ĦUqp�q�:�<��%o�7�]��to{���GZG�� G�hfν.�'���ԓ�v��n��:޶ 2mw�cg��x՚9ZU�N5�f�[���R&����m�0����A�σ��"�.�|�M�t���S@p���[CKF�����H�X�P�"@2���  @e�E��}^��c�N��q�}�<������i�͜.������g���XF�S�)X'v��R����е��-۷�8�~v��v�*r0'�:1�z����m\�V�Y���g�a�ˍ&��1{���@Փ󁳸�9~��ݐ�Q%M��S��Vf���o�lr�X;w�[K轛UiĆ�B�;�vt�b�u&ҧ�G�G��4Di���:�N�v�v{�з�-�0Ѻ�Ol?]�H�R<f�o0��w���c>�����8���C8��vk禨RY�erOi���k4�Q[�(�x�#C�~�ٙp7���}��<b�� z*.�-��\wm-��&'¨x2sG{��9p�?�OK��N�_~��J�V����p�guc��\��@�����L���Y���_i�thA	� ��ZB�k��CHΙ��xza7�n�rV}m���,�8-�_}������]�T��h�����AS�\\^�?����_���pwu�Co��5�& 5�8��Ç���7����n(�����M(Kͱ{�*��ZB2���Q���߄��'��w-�TvP��� - �ɤ���#K"�'y�����������������o��+A�*h�� � N�� ����u��ҭ��r**���&�����j��,���t[��Z�� 'Jk��8�2b�PON��7�E�pc�� u���: Xs܄��w�5;S�jj�
A�%������*4z�Y�i�D�}�R��X ]�J��#thI���\B@=�}�����ݭ=;�ÛɁ(�=!)��GG����\�Q��s�+ſ���L�=�,ZoC�*���+�|��\��/�F/�K�?3_H��p�1OU��'��4�*�&��Ƈv@�(f͑m����?8�[�s$�TK������XI)3�F���j]yDy��7�^�g#K |~^F�f��ݠ�ݩL�-ͬ����]5�Ċ���9�|k��D����栴���7�'�a��Ӱ��$�,a�`D�	g[T�O+W�kp!�;�Y+��EN��|&����Ju8�t>���c˘��N��?��bh�R�r���ħ��\��K)߭�61m�)}�� ף��k�o�3T���"@���7�W��1#v��kfommӖ�
%i\LJ����?�^�[�F�J�� ��� �#�8�`�w�62�>#��R�����V�3���D�DnF��	�}�����4|����yd���5������fT,��R���J�{v7����7��sh�PRa�{;��]��Ϟ*U1H6�x��L��>�I}��F����:�k�E�)ی�����Z�>[k�r���tߟGQ�W󥂈���H�j�lc����W��=۽���ѹ6�Z���|��h�0���B"�����.pu+��g/����oÿ���ݨ��Q7�p(Y�w���Ls�O��=�m�S�D�%��g'����E���L>�'O�Ë�t��r4�<�Gޢ��Yf�1[5}��m��p���4���Ѻ�_�H��������'����m�c%�J߮���}��w�M6�jڬd�d�t��1oYq��Ix~�4���]Q^��m|9�� LR���n<��o����Lq������ح����w��ZG������gw��d�������	���F�D�S��<!�F�%��t�Sr<��E���j�S+��;���F:=�/W�;��'��֒���1)4�H��IKZ�;���˵z�eej���a(���QEI��[���b����hE g�25�pt܃������p�G�Β����ٳJ���!��}r��WE=�k�����|Zj^�C5!H$��¤$��I��R|'KS�J�
UK�2����ZPI�Ö
8�f8���R.�V�X�'Q��]-ML(;��][Ç{�w�Ϟ( �-�U@���޺'�r�5G�
4m8㾞X#���)M�3�������{�M�U��Fr�����_i�S�Rz��k�Q���nFk�a���9Tڳ���皟�n@�����|�$u�6�SzaC�O�̺��+��J�O�hO�uGG�s�X�0 ����eQ%���c��M�FY~^0��3�"��|G�b��Ii�X�㜓W�YX��S��m��TN_�]�3?P��s0�t�X�̈:�A�>p��@��S�2��;�Ԩ݁'���JgUd���|�"�?"���u}����������֏�y�[���:��$��\2�?�,s��-+a�0ȿ�|��jv>��۶�	a{ڞ�$Y�\]��t��n��kjײ�ON4���	"�h?[d�:�|L��,U�Wu�B7F� 15GD�*����V%_k�7��U�x(j�܊vBe�Hڛ�ji�p*�m7�V-�.~}7�v�?L��=`�FU�h��!��B�s'ٶ���{�֚[���=��~��߄�����e	K��+*M����婪Ƿ�3v� d�����o���C5#�_�K{�,��YВ.���9����Xﭲ�]XE�<��\K�����\d�9v�ȯ+�9����И���jS��ti�A��>O�6Yn5	>[S/��}��]Ue�ϮUѳ�X7�G��`-(��������h!�� ��e�܆�K��(��0��-��=o�)r�t;��r�����Bԋ�s.Ւf��Z���\���m@�d��|j|�bz^V�
���U/sgw7��Y@��˻�|�*|�mU=��>V{>^��A���D!�{ۃ�i�t�����+U����*ߥ�T��W����s;�Z�;!�å�
���>���eߞ��>ײ��M(����L��Ē���V����A�[%�o�p��7{"�����j����Ҁ5,=Y !s��J[-�,�Z��^���_�������<J�֏szZ��G��|/�Zt��[�ݯ4}�l	��� ��6��y����Y@1C��\M���_��fe����LZ�X !24��I���e:��|!S N��N۴�z����f�$�lYm���:D�N��SW����"CYFi̲~��7:̲�����tB�V�=�U��VU�Do_�>�yE���7��4�ȢkEL��F?Of���c[���_Rm�i\��%���([�(~7J�`�DQQ�Y�Z�2�p�Elm�����!e�!9�P��!��N���ت_w��])��o[�I��v��<P���r�*��M�^���e��+Ѫ����U]+�.Ve�{���"q?RK�V�h�۹X{���+k|�����$�u�dIx���Y��j����܂�]w��C���aw+�8\�[��F��P���q%&Z��[[��T�U��c���5[�̃��D����+����}8{�ђ�;u��2<����|3K���k(KMK�<]���v�$(qFS2����F�����>˷������Nv���K���ʒ�����e,��~��&܀�S!�� ��	{6NEYWխ'���<*.�5M+�.Q���giv=�l%e5Z��0Y����و�Q�P����^F�@�r��.���u����A@�����X��V�%G��%�����fO|F�՚x�k���i���hm�Q_<Υբ&���R���p���G_9�[_X�ٮ�i��Pӟl���o�
�R{�2_��mک���u�qkI�U�=�l&0�q�]Mҷ�QŊ�t��Qj���z�g������k[K��'���Z�>� �}|��lo��-U���/8�����-�-v �Z�>��ܪ��A��q�@&%-O��^����,��+)N�����{x�8��V�z�lk�(	4T~�	���(&l�� K��<��ε��D��C�K�(]��[�Y�lf���U�.��{	�a�����^S���l��"U��[U��@j����πv���\�&;CKbe8Q9�E����Ԏ'<vR}?���To��S�Y�޳ts�K-L�L�E�y��2�����!G�!����C���X�ؕx��״ޅ�o�:+I��u����K]�ʿ$�ׂ%�Y��LΒV����m���G%�Pi��)�x��,����C(�5��J��U�̼������!|<��jT� \f��Љ.7�Ў`�Y)H�*-m�
�	%Ȕ�@�r|/t��ý6���tzV��-����}�#9=�8�B5i9�PC��n+\M�ʮ������ý}���!�l�.NHv��wmQ�xa��U�ĥ^��I;�f�U,���G;a���i_~�:�g'��
��`��Ֆ�τ�;��H��>�*
���A��K���a����u�R8*d#�Q5�]���*K��`����'�O�ʞ,Z�KqGqUW2�s���-�VO�B�.l�l��5����x���Or���(��AG�S?"בD`V�fm[�Qƨ�BhV�V�	���A�jcQ���m^+9 ,��`*�r�b����F`Nc�&�I�C<]��}�s�:�v�&���R�⁸�槢�b�O׆ �|):I��P����'	�	����
iSƓ<Cl+$f��a(�fJ�4VYH�b��,��w-�� ���C���e;�^gaj�;�%�@����÷;�|:s���ي& }w�����V�v��C�-*�"�i'{2נ�^��&Q�4Z�!˃�vEO�묿!����+o����%[�$���Z֏�Q<��K(�Dj�h�ps6�'	=m�>ɭf��S�b{�`�(�1[���ʞ�Q�R>ʼ������n�u�k�<���
� ���� Q���YVў�}F D=�fF9�բ� ��Љ���ֶ����C�xw�MW֢`P!~��t$�Vӹ�	Ŗ�śynQǪw]D%�J�q@��F�3{/�% +��N�FYͦ{AqՊIUy���?��;���u�Ȟ� ����(QϞ,��|�"-��|��J��ȱ�괨�_���6M*nFc�L�Gi1U>j]�U��� �m�G�U���ݏo���Z���vφJ����K�.�)�̒�����f%r@�(�*|���~�1|�|��s�3�|�1<X�t��t3���HEzs��0�\�t������]=X�9�1"�W�@&�C�f:<�؝٫��q��Z���3­0���g�������o4���DHy���j����\��Pm���B>h)ؼ~�Jg-��I�,:���g�%�\��z�箕U"d�N����QG.�LK�@i��J.���C�k�RJu,t�he➳��7���Ҍ/��e�[�ݗ�"ӲC��T�R��#�${�QZ*=��b�nt^l��>��KZJR�՗,%c�|a�,	Ӊ��;[
|�.�~�����Y����`��.�Z��	�����YqV���j��6I�8\$������>]���c�XߋAߞ�4̸�Á��q��A�ծ%�:�@w���{��6�'B���$�^��(A��뿾��|��<���#��=%�t�=I��x��յ����+K��,�r7��"�N��Ҟ��1�>���N�^"�D�]�hY���-D9,Pp�g[ �i�N�� lw�m�o�ilb�)�/x̥`�i�~V�
��3�%j�>6Z�����2��Qǣ�ƍڼȄ�1�홆�}?���N���{����lHK7ᬛΧ
r�R	L���^�����r��G �s�)KhAtuV�L�ّXt&�~��\ ���]���;4�sB����{9/���ndL�.B+]�D�\j��u��#�"bN-�Tj�=�Y�����J\�u���$���^���9-Ü����7�j�̔�áaF0�v�J&!T�2�� ��tU*b@����ZG�,27�|����Y�	�y�M�F���q�1�괤;�yص�gɽ�K5-O��+E��z�A�0a�H����qB�d1(ɒ�/���?Ἢ�����I��2���d�j�k֐�0�rQ��~��f2�J�|��,hm7��"7-�>�k�+�7� ���-��>���ޝ��|\O4v��P+ui@M#��S!u,T�:��8L�mI�1oy�vT�èt���A�k���C��:�%������X���F&���rD%�;	H����X
8�F0��H	����	��[<�-�$6�m��KkoԪ$���J�d	�$(	}��OWN�hf3+���m]S��3��f�2�r����{��g���2�]}�rR���Ԁ��xD������`�z�����Ru� \����OIMN�Lݔ����G5l6�<�����|��k�������{Q8A ��|�k�/-k^��6�4*�,�vi#���륨u��O���Ŗs���4P7�t��ء�@܂�9
���JWL�4���R��"'�)A�k�ǖ|����б�Gi�ii����~��6��`!�A����N�͉-c:�o^�����vs����(�5�;�n��6v���@(3���=`Fo�Յ�	�����$30�بJ[R�c<���n
� ��"��cq�c	6��QH��(m�7
̂��TK���u"�5����-R��5b�C��8LI՚�e�z WW��z�����k�IQ�h��m2\� M�XP�B��	��,�?�J�쑆c����y���ߘm�Jų���V9֎��@M���e{�뱡�?A!��3�E�~�
�R[<sF .[P��l�ڭ4�Ё�3�3�6�Z�[;����(p7[�?\5��#_;�T/���y���+s�>��?Z�&��.�Z���A���T���E�H�Ҩv��#�e�V�	�P��u�1$�Z���؀.�d����Xi3K�Tz�%��vt��ȉ��YvsKe�.
�0$���ʕ�ߪZ��d�r5��N�G[��w�R�`b��Ր�M۴3K�&����$P�r�_���Z-��y��:�Y����#>�V)�T�}eY��6J_Rf��̻�Rv_�ʂ3!{0h�0�Θ��N~�Âp��ŕn��MI���B#��P�t�U	EX� @�H23�yS��������Ud��\T�c�Yg'�=�>[F���m$`��VAfe�O3x~��cg���! ��
8��A&N}lP��k���1;��D�m���h"ǹU�]��Z����U��j�(��PC�S��jCO'���������=�w�VUu��o|v��(b�"~��g��U1�3�5���ϼd��^s�`�@m�������!ɵ.�@�?�����ۡ�E�����击"RxȲ1B��JQ�Q�0q*�t�����ߌ,�]U7�^?l�wMm�^Z%L�|�j��DG�N(��h�ڳ<x�4�|�wl-!�Rwyҁm���`??o��ص����⾷�s?Oõ}�k�k��V(��p��	���PG�<��Pe�۞u����B�\c�L���uL�u�	�$/�Β"�-Yd�*��P�k��(H�y���H�w�_���>~�"�_rD3?|i����
���*h�.�{�O�	�
U0����-��'�O��o^���H{�3�@3��j�'�����d�e�ӏ��}���];�%4���1�@�%V����ϟ?w^;�ί/���a�Y���=�ܲ3��i�����(�%��Q�̙��;��J�3�ɯ�,�?	���֙��"ޠ����jL��
W-�/�L��7�<� �62�?�b���F���A�>c���5��5�-{dlx1�׫��o����4bI�z�݃p�=�6n�ygQ��4bn��_?��[^	���ɍ�Z��x�A+p�̥U�T�dl�>��o��^L�^�U����߳O�a�
�e[�������@�x�*]枫�C�$S7x\op��T�djH��ձ��<%�JYT�cܸ�8�^�~!��$�|V�V�=��C��@�v-�~��qqpo ��G�n�Q����c�|���*����m�XKDdB�g�wt7
�H��[�d�I�?}��D�CZa���p�<R ��V+�>t�<�Es�ҫ�E X�$>�H)g
z��JHh+ƕ=~��TPgn�8�B�B�Ƭ���"Z�e�)���B�Y+��k �e�M"��"=d�P���k[/i��ء��ׯ�o�|ƣ�pwy��$� AZ���;��ߘ�_^\���;�R�O+�JK�ɫY��d3jQ��J%�,�\M�/�z��,�u����Á���7SeVfs��T!��}Ι�I�+X��ǃ(s�����Q�l.m���]���B�d�}n,�����9z�c�J�����.��a�#�f������$���BY+HA�*��4\��=Y���1v�v��0�vaͨe׭Be!*����_n=���Dr�]]�J��Z�i��]'��3��7����;�y� ?�R�P������[վ��"�l�����������Ƿo��ŹӺ�$[Ec���^����L�f�ؽ���|��ˮU��(�߶��b-��3t;�(,�ptx��Y"���������E�2��x����X�	��ϟ�g/���?q��\��,H���
��LP����F���4j=�gK�- ��h:߅��=%5�4Ղ��up̂Č�:T��(�p�5��Fg&��oۃ���k�Ŧ���K]n�?>J웳D���S�8���FS~��,E�w%�E� �����;�t�0cɣ5aH\}/
��&9��u0��}9�jOJ=�B<�,��P���R��4K����N�!6�h|��l^�ߪ5��ٓ�w�;}���PK���[]e�+;��P�"ia�>+w��+l�,���}r*bZ>��D�;���qcьmY�'����i��Le�� ��M����@�yG�AB�:Ȧo� �
��5��"�b���%T#��KI��D&�*t�����6/���Z���&������ai�`/��0�zYE#ri
��FK�u�"^�
(#�6UYD�.���2��W�6� ~y}�C�������:����Z:��=��� G���;���	�PI��}IY��TG�j/�*��RU���%m�Y�J@�`�l)���K>�m�<����������)V����r��u�tCW�������F�>�	��\�,x�!X�R�v/���~�'Y�]^�
�z���^��i�����]�|�I
C �� ��%@�\�����S&4�l��dA��/e+�:�4fj���$?Y�=��=[�w�v�?����@-SU���G�U�m�q'��epr:��2�X���J:R�Ҟ_�C>��Y��HŧŶ��a�-�O�5��=ה���̒�Ҿ��M�T��n���Iˑ�6\�R��UȰ��]H�CSIU�x�V���>���)VU�թk��4O\�U!V�p�m�Ҋ�����þ]�WO����S��� ��7��t�Aا�����»%`���f�Ŝ�9L�<	j�}�m����Hջ�uu�8�ɫ�\�>��={�O�+�#��:ؗ��Lj���V��'���_��_�T�
�C�YU��%DU������O��r�
�A��]�N3/�ku������z�V���HO,~�fM6I��w��r/�2*�=���4f��C����$���7A��o�>T%��]7��&� \GFH3�8�@|�iR��ݫiQ��KY�N�(��]�����Z�M'%]�R���{��i��FߓlK6u������{�f����󒝝�p��E�����^����~�] ��[y�vUQ%(�H�0�G��jj��ř{R&�.��{�¯�0?�%�Z�ˈ �#|NhF�� ���0�L���F������(F+���,`�
�Ӫ�6��<���9��y��b����M�<|ba��aߪyt֥�B<�&�<�3�1SD�������(��E�f�M�:�^=}��n�Gq���W��f�J�a��cB�D�- �b��B�����p-æB�d�V����hgف���3*,Z����9`kK��W��kq$�?=������R���Ύ֟�㑱��h�!�e����Ax��e���_Kp�.h�F��k�t;� ��L"��3Sk��:^}�}D�p���*�;[��}�hl����ɤ�Q8RYs2S[���<�ϼ=����h��V?��b*[��z6�J��Z��&����S���%K����H������QD�a�(�XBw����+�[�gV��u\2��JL���RK@B�﵀CP�ʉU2v��/�&���l~�J��h.��M����B�JD[���:J��k�3u\��J4s(�v�P��k;�T�|�-YC��`��}�'Z�������JƵ�]��=~���%�N[������������n�]�h>�$��%a��! Ȍq����ӧ���_���}�oh�$:��Τ'�+�!�*`��ϟ?��?|'Q�@�> �D��"r���"���G��w�Yb� �������[r�.2B"�+v-����_�3V��COy�}�i8P��D��_{���]y�f�yb ؛]��������-�C+�aBӊ�r�ETDk�d~�M�F��[?����
?����vY=&Hގ��zD��Ts�5�8���	�ZNi.�Bkzf�w�P-jT����W(k�.�k-�������k�ח��ga��K�嗕��g��A�c��J��1��v���p�Ï?(��û�0�*�2h�j��*��A�ǌ�I<��z�������NO/$��!�.|���ܥV#�fz��� F��;���'���t��ζ"變�l�Y7�o��C���0��CE'��X�d�9
7�� �d�U����o$�`0�@.l��j��e���ԥ��#Y�1^Zu|{/z
Vi�GG����pp�/�13$�1�Ev�.#p,�y���3��W�D{�{�&tum�!c�Ks������ˆG����1F�2�Cw�t��G��[����v5�:�xx0�;!�"Z�d��k.O��**UӅ�^��㳟ݵ
�����T�s t�D��b�E%�X o��F��OG7�>K$�0�
F���A��A'�T�A7b���D��ڛ%cT��^_���K��@�6U�x�($v��\� zhWnϧ�x��h��4�B&޲�0��5��a!�a�Ug��Vi���v����'���]���'��]����~O���,
Kۀ`↧�-�}�[�s0	X�K:�v�� ��Be�;����a��pϱ��:G��@�����ӧI�*>��T����$�UҔ��=����}�|wc	�HV��U�� �$:1Ӌ��NY�;�@?}�.ܾ;յ%��Ǜ��Q����l��]���E�������������_�:/�/¥%�nz�R���F�
��`g�量
ƬK��+�͢��Z�ȼڽ����o��J�t�Q����΁�"?=f��]x��4���*,���s���Dv�[�@{>v^�z��Z��.�Jw %��h5	7�u�*]�����~��U��5�"�Ơ�(���$c[?Γ�o���Z�X8�U�Bu���3�8��'-im����c.܏<Q�0�B�G0�񖺅�p�,�Ì	�eC�jb�ƿ���­ZZ1U���i��թ�ĮJo�+� �(�}�+��[��{���2=�_��w2 �eV'8�"T�)E�B�����B�E���
	�����>3R�c�.��#�ڑ���zT{i���	�DU�������y����doW6hg�w}g{�UT�x��J��.2�I�Hɑ�v]��C(,�8� 5�bq��.�@�߀�A�{O� �N��|���I8><����v�P�l�q�cj���A��#K��(>���3�q�����3K��Rm\�a��u�. '�*A���ж��V]ׂ��{4��q����i���a���W�r��MD�j�?[�-H9PO��NO<R�3eLD��N��������p���ݶg�Zb 1p��V���y߾O`�(��ª�{[��v��C�%r�%p3O"hˉ�.��Z"��Z�q)�m<o�����XC����@��V�M^�]�s�<��8�I� ���� �T��4��Ձ����6G�ߏ�@?�`�~�p�W�piA����y+<�zr`�Ӫ���в ��y��e�I��%Ѫ`�1��=���<������lW���ّ��n�tw/����Y�+E-h:ܛ~�6��3^�n� [��B�^Jn�tE'&*eL2P��������9!0(�)\G
��3},��o�ُ?���$���G�Q�1m��#�����8:��г����c����#��z#%?�0��uh7����E�1�:�3K�y/��.�"wv��g�4�+�����|����	�$�--]����25`��??���>>����A�ŧ��D�L���`1h�>�ĭ���z��zu��L]�F��y����"F�we�x���w��;3:ծAW�r���o����V��EU]\7�GQ'M�1��@2��9��r�iL*��"��N����;r�"����6 �����s
�v�Ө��
I���N���W��y~������j-��d����Zw�!�n���fM(9;,|[|{=TF��Εy��﫽���\*�-�T��-�X�"��x)�P��XQiv���r��ǌQ��<���di�Dhc�EQb?7���H�Ti�H;7q}�R�)�8�.�J�O3tm��1���*]�9U�}6�����me=����YY�q��ٳ�\XKһ
;{{���H	�d�~x�}x��dSfM���mc�Q�!��)|MHPTe�����,�p�j&t�U�y��ӧ:im>�ymf�fa�#�1�%��h�w�N,젴����Ϭ�������N�l�����6/����	�"�
�F�i���&��6�4�bVЭla�>�{��a]:��9���u��89���w�n�Z���Ѻ�ܳ�1����J
�Wͳ4���Y�һ���'Yl��0�Aaj��f,D[qm����������D,���K�� ��l�$+��j�Q� d���c����ϥU�s�J(Bm˥���:�ۺ<��7W7����*[��%'t���K�NÐ`��n��ګR6��^:�Z�+�����c�M��Z��К��=��nHW�ʂ0^�IZ� �Ś���G-k�T���K,�����!\��������z[�2y��v���6R�	�O����> Tunm� �hYF1��n�u���7t�琧��إ}l����U��bl�9$�v�����p}�������������b�m�um/�^~V�3�=�["�A��4|������i8����ü�ϾՓ�P�������d.��"Õ��o��$�xo�^�/uFE��JR��^&?�@j�v�U��Ei��p�ߗ�����rb���y�%�)I�p�`�ަ���cE.�Ő���� ���u�]HΓ� w��]
)�|�V�nFJv$@��<Q�un�v�TG~� \�դ�S��3	P���N;� ��g����²��Pse��!xx�vʯV�g.��؆e��"EzΛ6.\��S�x��BPe�j�C�Е��R�A!I~��I��:j����@���=���h8f�����(s�o�tH>��ʝDԧ3>�j����c�z�Z��}tJacw�!�Z ��J\����u����~?W��=nmuT!ɣ��E-���Q��*���N�V��K��r7@�ARW�`~73�2uII��<��|�����G/^��ݝЅ/i���e�U#̞��O�]�	��*FIJ���W� �ܑ���*W!jÅdё�cމ:��?�Ujbj��_�0�)�$��l~_�Tx�R��!c���$MbL�@�B/�D4:B0��J�|N�T@f�P+��+����y��_a����:�����0Bu�H�TEXr��n�������*�d_H���p*��JkV�U�?�_S��x��M����9�I\��<��{*���PX��K^��U.l¡ɾ���m�9�
������U;:�-��h�^��B��Cb�@Y:71Qe_�3]�TIWQ�ΰ�u+�GPyJ�,RS���C��pkh2�wlC��B�x(K�A#�R�5=�3t�^nՎ���hq��{�%�0�C&���~i�:�[��z��@"�~Gi�}l�2�y�uX̑�q���m�H~�Q��~��ʖ$��E)�sn	:tK���/�(/��?�>ZR!�j.���[����CK���E�~}{���ӟ�~|�>�s;���a��cNړ�1����`t� [(�(dUѯ�A�r���oΙ:�-em�H�=�7������S+i�P�C�d%u�c����M��ԡj��$Y٨7f���q���]�
��hH"?�����-������U�M�:y�w�[���F\���2�9��W����Y+9gf�X�"�#�a�o�˫�����qU����?��ْٙ���=�)��P��&y�O����z=�E�<��L�9fj��n����yΘ�����G��NѬ�� P����{����jp�������´�*,
AJ�;�H�E������k3RÈ*�95R�������j_V�Q�Ӌ>��^ p����Z�D΋>dTL"�I*	�3�*RӹȀQ�!�$�d�'�_�vU�Bd�yԒ-�aL3���![h͝�hp� @rR���]����Y*�d�P\��x��0zE���H�u=��q�@��C�FU�j��+�}��L@�n�tA��O�D�������N�3
usw�-J�`0+yd/!�?�	�d�$h�up�J�v:�xxK�e泊:zT�f�(+I:��!��������@�>�����"���X�RsNT��-�l�)��s拷�4&2-p:�.d���Z��2�2�g�P���Z��c3Ҽ�4"�S�w����5`��;ڴ=T	]�g"b�G�}���2$k�bi�7Q�V��x(�C`A�Dw�� ��}����
@�]<�{.��U�����f�N'�pck��!�ّnr�7���̥2I[^�85r}'�N�}�1����	����v���
��j 8�6g�v
����po��}Z���ҍj�����'���3iZ�y�,�ph��\�����t���Px���c��-��Թ�,  �I���"�x���,�V����7F
�ɢ��v��LH�z�jϦ#�#�T&(��"X���'�_,s9׾٧����.��Y�rgvͻ�wtv�de��^���m����
�����U��Q����%�ro�On�&PR�?�E/��uE(����2��{v�U��IG����LY�]u_Y�#�=�2�	�5{��ԞI��e���jTƱ7��f,��Y�)�6lt�%�ԏ�pk�ny*�)Y�]�q<1D�CU��ڮ�;���!�����焛fEtt)��Z�G������7a2�8�:Gvg�"�mC.3ȣ�&N���zgs��*���ĉ�_|��VW���CT����H)8H��� Z��ֈs���"���Y�`�\��T���c��!`O��K�q���蘬XΣ�hP\<��Eą#&B��G6���J��,{*��K�M�n��c7�5q	�"��Z����hI�Q*R�f��N��ƈ�k����QXf8��A����#��fS=rL%i�jN|&��e=�Hv�2*cS�����'���?ܔ�����"9F�����!��蝉O�D�Γ���}�6E��"�{���[G�A�|��%�7�^��.���/����2d&}n (�Ygh��`qf�{) ��ȼ�b�X�
�'T������Qz�K\�1�X�Έ�D�ckS��*���:A�����V���1N5^"�bq{��`�V��ݪX�Ǽ/�A���0!Yc��-�4�i�v-3{N������7�ښ%a�ӗjSi ����>�\?�G�o W�n�^p�챽�D�(�͗��^.|L�����e�8��;�L�I�2�2�J�v� �5��{xtwy.�?����d�D��M�R5d��E�^���eO[���[ˢ[�����e���Rޅ#]YUZ��{jB�:8�	pp��S���p�l��L?ڹ���C�>��%*�l5�F����)���"�2U9:�o�aTcj��������~�S���G�!��K��r&����O�jj�4�>t�g[�����������[��=�]�	PE�F��\W��j��J>s�e�s�hĚ4*��/V�_���;80TϠ.c�~rZ=g�e�`k�~*-�ռe�f�[;��sjVHG9���.d��e���e����cx2L[;�h5�9�W�J3���R�Y�*:���oćy��_?�j�%ʊֳ\��ۡY��~�Fs{@��2�}f-eX�Ј� ��*}�:j��jBO�Q���;NE��HʱZ�����ʵv�����������ə�B��c�D����4Z9 PV�٦��R�\V�M��rX��R/��
e��k�2i��$�w��'g~{k�^[:ܔ�U�	A�(��Κ��q@�K���+��U�����*�#��ĭ��NG��9�~:���Y��g�3�Z����h�`V2#�xh���6��,֣�na�V��cd߹��5(1��-]G�R����>,|��J�����^�GC����x�[#1�tk��o�����ǰ�w�> �y(���ɡRP�rc�4g+ĵ���}��"l��#������"��9q�n�*P�	�'r𑰀��gG�p`izH*H����B.�~ �DJ� ��Ssg���h��J�N�M|꩞�K_k���s�dm�n���-���҈�y$s��z`ی:#Z�Ϟ?�W�q��e���������}lk��R�4����e�渚T��$wΑl%D��$�5��o|�>�|:���*V��\��!@%ȅ��D`=Y���mX=M�<k��0_m�]�/��'�����*V�8k۠yoh E�P��׶ F�q�����Ѩ}hDTF���-�O����v�p.c�!U�����d�?�ۻ;�p�������nh��6���am]������m�IOә=��0̝uO���l�t�7h�ý�ph���ˆ�]��G2ޭ���a)��l�+Dy9���g���qƻ���z�y�%:�8.��m�.?��g��A5��"f��Q�k����j��#�խ��7�,���|�����("�z쪓����t�vA��]\����lS;�+�x�v	DG ���.3i��&���CGwV�������SlLZ��<�Xt�A�W��(=-� ��_/��xrE�Y�T54>��Fh����D�R�ꗫ���W�s,#�@�pD��&e�
Ǩ�x\g�4�"�XE�'�XӬE�o��*�.�U�ቦ�6l��s�̧�3��ABWw��/��/�7����-h�*�{Tm��jR�3c9�F�Y��ة$1�e��V�	�ں�/���
,�vc�K`��K�-Ts�|6c1�2���g��!����=$fsq��*������+mdq���;-��%���P�hX�k{�^�k�ӝ��*���RС�%9�b(�Ѓ7CE俷{�d�A)3^�,��Ob	y���}��͝Ʃv�	�lvn�cwQ��, 8֠�y�"�ϑ]㈅�s@�����]�^����}��0j=���ê� J�0�-��� Qކn�ג�-�)�����1�2����خ����~�oB�s �'�<�=�S����wS�s�v_MF�sL+l�vm�3�/�V��/zk�k���'\��� ̶l��4'��4!��G*?�D�C��J���~m���@/O>���SD�i��QvO�}KB�_�4�9��+��́�ˮ[��tq��L�5Q0K�*�]�4i�ɨL�L��g������5�*��p��"(�gZ�Xf�=���L�4�'�i��y�Ã��}�ph�@������a��ǻ�?
�L�r�� ���8h��|�	����LA����U>c{/���~�,(�l��ߧ��&�EYYE�a��3J�c)'�WZx�۟�#��	;�g#E��|� :]�-'z	`H��h�$K��8�,�m6<����v~������4b^�(�y�)�y����j�c�7�����B%h�w-"�5͈IT�{�UI͗AXv����˄;���h��"
��Te�0���4�Xy9PE�V!��(j��W�)fy�f��*�E6!�y�ڦ�T�b�7�Ϣ���Iֽ?5����4��Aeom2[x�v!>�5� E2S��x�Sh��,S�hP%���B��*j�اH&�������*p 2�E�wy�N��|>����׿��sKe��f�3�#D� QQ����A�O��pg�β9��<��^hE�gK���xB�/�g�DY�?��Pw,b7ð	ےH*X�BC��P�悹����=��`�2l4h� q�J4CB)M�J�i�#���E��"��E6-��bo�{��,tp�������q��9J�k�J�+20��m�9;���FXX �����H���a"�/߯�8�^z�Y<�����.��;�1%@[��]��M�B��¢�s��	���?M�($�.BIY0͝�#f�A�}�2��X���7�������/d�	@�)`OZF��Đ,$pz���y\�0���1���0���X0��j{�v��2f���3���a{���a80���; ���bb�R)�4��me2�S���
�N4~�
�&�ex)5"Ҷ�]	K1{���sc�14�b���'L�<\T�9*W��:0�X۵�[ӏ�� �K��&<�ii8��D �!D���3�s��\�O-��}X���e֋�+!p�QP� ����'SU�(y�'�Z�|��������cנ�	>�6"(��*h��_{;�"יY�r�x
f��n帜���899q�x�\b�r��	������^��>'��J`D���;ܢ&Y" O#n���_��Q�<_WS�	�f�h��kL��$���H���Z��ՅȆ&j^�j�vwf?�0��h{�@/u��RS9���&i��L��Ns�UYo�&֬��w�ݢ�j�-+-=�c_��.̘Me0 �OʘJ�;[1�e��������yN�`�-sG��zq��6���8)���,q���2�F��/��k �`��|���T��a�!K�������H=�`����-�'%�*��?@�-�a"�/]��:Q��gHA�6A�ڽ3o��<*
�����=����~c��]"�4���Y����"�J=wƯ'3F�?<i'�8T�m�Z���;6�
����Y[0�)m3�d]�~:B#�E��K�v]]{%T+��]> �J��g�rǘ�R-���/c�@Q���\!G���vGcY��Z�fB9l���9���(� �Pr�:z���Q <�Yp�Zl�Ä? � �m�:E���$�kWѨR�^���mM�B�q?[��Ȱ���4'�Z)0@+�U{92��`D�����k�%���x���HA;
��ӧ*�,�l��T��h�9c�@�T��� āx�@�ư�%%y�ˌ*�ջ�;�}�;[0?�°3���ۗ���gtk��N����� ���O�vl����T��2�j�W���q|��|�vOm�|��
�j �l�ޜ���߿�漘�
���ԕ��$[[�>�4�{'����ߘ��sг���Pd�kf�]"�tJS2vQ���W�x��t	BXKz��.To?G0�c붽��`���of�9��W���@t�fK���Ӊ�x~Tͤ�]Ub;9?��/���ȡ8�ϊ��b34(AK�����EhMQC_
P4%��naY{�E����+zQb���O��"3���mP� F4sUX:���u�K>>+k�Sᙱ�F�i����8�y��0-��J���V _���G[�tđ%�Wa�"b\g88�@?��٦l"��a��ѳ�Y������]�~����=��WAk�ԩ�8�6���Ls-[O٤���4�����n�o"��Y��0�v��N�]6�VƳ�c�S�>������FG�k�Z4����ߋ�R�|]ZvV�B���uxx���=��ˮ&I�;����u�9��@�H�jA{�ۖE��ڞ��P�4�1�(��?��]٦Aƍ^Y�
4o�-�����6:�'=M��@�1f����z�Q��\W���U���ξ�:��O���e89�6�ԫU�g��pn�$Q�9g3�Q}wN�1l�vD���t���#�o��
�Lw����+&r�5w{>#��(��Ԗ�Q�BC���ENR��e�M��k�ɤ��jߟ�#�1ë9��񆔗$�$k����3�$�ڻ�dڌd%�q��d[E�**�Tr�m�}�}[%���1'1^��p�(�T�
#��e��8&6�K��dQ1�yN63�2b �	n�Z�*+�B��b�G�����ҳ��.ʥ,�3�eDf�	�x����ί���� �Z��u0��TC�C�礱=��6��k& �:;HgcG�o�q%3�v�(�n�GR����We���k�&Wg�bb������!�=�zas���)���L���	3{�����dLd<��?W@rwz��}
�gW��|���]�	�5�H	��&���1Oae�ײ�6�ad�i#s��v7�R,h́�d�5(��5=h�"%�4�[>(к}�����b�yyl��Wط�~P_�=���+?��4\S:��O�L��^��
�a��lM;ɶ�����8����p��{0&[=���p�1���;�BT�ٞ�b;!��Y�&�f陃DyB������hd[b8�}H�J-��k�S݅J��`�q|p޼<{���dR��l��H�2�K�����xd��x_e��Ӫ�m3�#���ZY��8.J�RE@-UŚcZ��HU�
oP���H�\�E ����x۶�djk��i����H`���fAa
�挥���F�I���6�#���rU��&�,K�F�71pc�����ݏo5�Z.ܐ�Z����.z�"9Ə��c|��Lc/���%��g&z��I&�D�:5��po��_����$cM�3�h��I�;ْ�+W�J�<�2ѳ;��Yq0�d�d9
7@��x��ut��XF��YY7���C�����ʚ�u�~���2�Z�N)����"���9�g##u.�R}�Q�BG�A���T�^��# +�5�����ZDA�(�F��h��!=(�Ke ���/��=uD�H�^2<��i��5=�{^��ep�e�kkc�^S��NsQ���R��=�O����Ϭ�j�3�eI%g*�M�J�)���s��0��~�����?��E��ر���C�m�vvv°�u����˩�$F���O���ť��e��Kg�j5;r$����xd���y�Y�F��c�\��o���x�{s� {n�/Uڄ�ϥ؞uEʈߎ}J��^PV���]�[�"|���3�D���YЃ��i9�b�y0�z'28�����<<A��C�"8`gZt��x����k߂ ���a��Z���B�A?�.���?���R���"�i9L��9~���c�;��\ƈhYd�<1��?獩5��Q�tf/p�#{��x�0��y�A�\X�nd�Ӽ�(nKo�$�8Ώ�HNnn�c��X����.����>L���<X�S@�[�.�c��SK6f�^��L*x0�!�B��A/[��fا�70LO�/VKi���C�"m�+(�'ס���Xm*D"���%J�mm[�r,��F����]Ά����G�W_��v����qN�*]=C_W��e�AL
#�\}��)GS�Rm�\��3	g�g�+9,D�f�Is��MB������-3ޗ�-\���Qh�����"��e� ���4�t@Y�rz�-6�Z�<�s�U�T���N�����B�:�P�5�׽"6)e��%=p���+��wEWY���H`)��r7��D
!���G=p`-s�6��Z>��	3pXt�0V�Z���U9\��	�!妅�A����� �j2���g�`{�8�V�ψF�\Eۑ@�C^|&=������"^5:xj���d�璋�<��Z�#M쀏��G��xD3��'	I6�5��!�G��󀩈��=K�O�֦��D,�����K[�,� +�D0��Ec�	
2m[�'���1�|�&v/�׿�&~y�ÞZH���^!܈k凨R�֫V>�PD'����DQ=@(��m������Pҧ�빹:o�K�:��"�vҶ��/{C�}��ٓV+hH�3��r�<#̻w�¹e���Jn��������9�˿����p)��T�#�:	v�P��Eb�:�]7�ω��4i��<D"�  �N�����ێ�y�D�C��C.4��D�˖dЊ2�k���m�``�)(��]`�*E�RHz:78Ƃ�gm��*���f�g�ƨ~��H��^�u���<��nP=J Z ��)�2J�s&��]ߜ��ӏ��y�R`�cv��L�c/o���w��ɀ��Mv�e����cG:��I��W]D�,Wa��##$�:��2�S�aX�����T~�$k��!�psy�>��ҏ�}�����k%/���k�s��6J4�v��S;����R��H��a���ӕð��3i�T��i�
F��Ո$7I�/�������x���*Uk Z��v�}Wz��`s~����?}�_«��N�i��������U�$���j�1��(���H.\,xk��,���������i�\��̌؍���J�n؉tx�������'m �� ���Y�]^p���Ch݀_��E��g>� �k�D�9K�J�N*J�g˅����~nD0;r7�SC"H��z����l"��u��
9^�2`�_�g�[�7^-�ؔ@�Ρ�,�<���2���4}DMM�Q`��,�xFR���,A1��
�ک�F��x�����r��
� �G�-��5{��t�]�>Gq+zn5�nq?��3�= �6�.E�@����߇�˟�����PX�E��4s�8Q2,"*��y��0D|�f�l�׆X�-�>_Y3RA�R� �Pj��ْ3>�@���GeP;{��`�E8x��F]K����9s�����a�q�bC*D�WJ�pb�j��z	� >{L�#�1J=E3�J�x�����,�S&#�>�n�̌w @�qJ�2wސ���*�5���/D"��"�(���dq8I�zϕ�^����ӳ6=K���o�2���-Vk ΄@~�/����J����#�"s勬l�h
}T{���˼ pa�����v�Z���t�B�lWJ���f�"�h��<�X����w$�C�|�tq�����Evn �-�:�p_�,%U��;7�l��\3�ː�s_��d�30"ֵu������>\߅�|/,;����C��7�o[�-�x�3a��- ��9z(F	�X�A��`��E�Z��IC�!-2�>*�0�h�V�lp���|f�Y.�4�)k'���'���kQQPM��K�TWro1���4�g���3)p�(%J6��k�'����]���,����9�)�r���U_A��YX�pq]�� ���_Gk���D}v�g���T�̄M�헿�8<{۟8@�D_V�wJt�Z������f7�����3ǥ���3ЕNk�*�8�W�d���Y�O����:5����aQF�g�Þ3�����=��:�'���v��3O0���H����<��K�7	)�g����3p�hj$a�n���se�h�z*W�,"fޯ}])Џ���.��zoƑ�"������t�m����sl�B�I�t['z,��(ۂ�+
G�3�1�~�V9
2�E�f�aP6�Q���/����ChX6c�Y�9��ǒJ�0�RB^:2��C�|2'0qr����F�2���e���w�ӧO곡B��W��4�,�j%Ks0�Q,��@�k��#H��4�ϡ��� ���b�_�2|��������@�*�;�#3�@�1�4#R��9ꅍ~'�ۍ0�b|왷��}~S� x�Wr>QD��������'�*܉P�����*�J��CtBI��OX2x�����-��J�U����^_X`���8 }���h�lBt��~�`xpÓ=a䫺g�3h:�D��S�7�O�O�_�9Ֆ��"��|>�g�[����T!������>�5�C�Α=3�ˎ�s�m_��� ��3��X:;������T�e���ՅO3];�N޻��2��(P�{���i�x)��(4]���e�N����{A��ٜjF?�!v����V�o�����9�9�j�q0���$;eVW�|��'�s�����eoX�O5~�ĽM(�=��ʯG\DҘ�� �>cH���wF�4fH"ј�Q����x_���b�JL��YD�c'7�m'~�4��	���g�xXΈ�\#9�L@�c+*Id	����askG���i��1c�udNX���0��%��R�P��٨d��82Z9#\���R!�z��v���^o6A�O���,\[����������}y,�'Q��Y�b$l�52��++���b�����g�U5����JX�n��z��@�[����T �r�&���k4:�C"sB��R�c��+U!�
��J��u)�R\��Ahv����?'��/L�V��1��?�F�f�a#K��-�������a�^���Ww�"	����O��
.T�^��R�R�֮-Z���^%����4�K��r���T_AJ=s��#6��Kb�3�O�%�:2�1
D�4�e޿K�j�Py�&�A��0��C�r�Z����<�>��G�^JkuT���r`�����z��8|��7aW������p��D�O)�ޤ���a˂|�,p?lY&|h�igW�i>����Z����'}��Y蒍�kl��̲,�!<�#iB��DJ.�:ʌS����> �9X)�o�=nkB6��q���&AT͈zJ��L\������I�fU��mѻKP�_��&����$p#%_Z����˰�1
��������������>��iT`|� y��ۍ(6T�=Ҍ#M/�u�'Oj��z����:`��Y��6\�b1�S ʽ�h��g��-�ɖ-�2u�e&�:��" �@��U��Z U�z~_�y�b[mW9���J�]��MHj�ѵ����83co��"�����^2�VtU��8�=:�?���;9����ޔ��>
X�>�NB�r�96H8��L�dv��	�A�����]��R��i��G��o�� ��X"�8���=]?�}_��������I���XP[�T��Z��k�>�3�!Pn9-(�c�/u�V��kUz��Ȉ	�CUTA"��F.Үg`�6���Hס3j������W�]zy5��2uX\qo볼�|�^�������P~���L���k����fn���Q����!ցXmK?_���kg9���p�{�*Խx��w�qM���!E�k]�N���P����$˕���4�/�%ؤ���J؅�=�S-i ��s��MM����v`�l�M:;�W�l�Ҳ���7}�,'<X�Y�inQ��2��*�0Uk�"X|p�=44yHd�D�d[��um!�ٯ,b����KI�	�M����&2����P�A�zZ���{'~b�N*t5��E�b/͖+���Z�j��,��kh�4�I����c=������xu���+k�W}��ō���)���65�N�u`׿��ڦ�Â�IHbs�fh��_���/��0�2z��)�-Ol�r��u~��6����ɇpws�1���=]{?
��#\,\� '��_��:�I^��Ӟ>���=۞9�'t����Y�/8�����"q=�̧�$#��gM%BH�<���CP��MUV�sWo��>�K�˞����U�\���j����D��x޷�Z�:
��0�ۚ���i&N��_]˨4Ĥ��vzy��(SS�\h�p�AEE��>�䒕��a2Ot$˘qy��~������7��kl�o����آA����zŌ=4\l^s�R�I-���N���� ��N�Oy2��g�}2<��h~őn�J��lF��Zw�rA�l��H�H�2
�Q����'kP��]����2'�Et�+U�R�VsۗWW���������ك�9��ZAg�BX3���Ps�K��i;����*d$�T���P�O�5�׶;?T��n�eP\-��Y�ph;[E�_�4���K��?��?i?��q�~��:Ro�I|p�³_0*W���֬�5U�J���y�W΁�F�]�����_' ͬ�Ԫ�6�^T�#*U�	~�BV��^{����	L���(�$&0��֠�:���iW1�M���F�Q�f�W?��*��{�v}&�W+�������?\K��?��J�y�
��Y��	V겳־��R���+�����໌Lrd��:G������ �Ͱ��n82��r�������b]�Z{6���8��&�����tZ�/��#����amG�%��!���p3���{uu!������T~��qj��F��E����Y��\�O��R�V�l�Y�!\-ܸ��2�a�ʣ��b,U��{1;��2F��g��ș>B�x��b�$�sr��aѷ�^�馈:i+l"8�iJ&����ێ��h#X�{`Yߛ/���^��;��Ks�7���'Zoл��{�8��6��@Y�ut�����QT�/_�"���&���_�@��Ȯ&v@w�i7Tz9��-ϰ��lK���#ef��I �<�^��JGWe���o�����u�JS��v����A�9�U�:J�cs'?�N%#Y�0�z��m=�N�!m�F�*�l/���Qx��u����J�Q�s2#�:�q�������(I�����z^zFzH����V3�%q[�ttv�x�M�J��_�{ ��٨g �J��S�Ԝ�t�������p�8A�����,�jv�XA�1� C$���DO&a
��q:H�NH]�����e�8&���ΞEy��zΊ�uyp ��{~��!��*U��)Μ����R��'�C�����L�EŲ8�F�'/�tا�s'Q�;��g�ߍ3��:���(O��?��?�f�ɚ$��E+�1� Ҍ���ʹ���ޤK�ܴO@DT	(ٷ�v��Y��FE�ŽՎ��1_�$��\�p��i�f'��y��M���5�ă�G#4?��d
 R�g�Ҍ�,{D����|�r��2s�c��ũD����no�@���m[;�N����SH�R�\s�L	��������������n�XLqd��	Hٯ����3U��Ib�@����c�;�^j-��|a,[פ)\�9���V�w��s�g���`�P߂4�
�㔼�_�,p���C�%,IA��O��or����r�^�����v�%Ѝ�,E�:��Y!�g�i5͕�b��������d��m�<��Ϟ����$�>|�(R���yÉ!\�;U-~fbzJl�njb3<��)Rk�⑭�S x(������Hr,£O�r]�<�U�D��3F��u,�FT5YiSs��xdx���$#���[�B�U��(;/�"��,��ʉl����-���3�2��Xd΋zp���*	�$S
y�=ܐa��\�М��Ʀ��D������~��������?�	c�^(� ��û�|#Y���s{{Kkh�)z��g�@| �6�=O��t�*�e;D/Y�ud���īqXA'����DN5��D�d0Mt��1^j���pO���`E������=�X�E)�|��W�섫����ݮ�ї�٤����������m[&�H$.��P6^��.�|�H���
P����/����k%�8�
��w�w�ʯE����[*�	��9�v� �Y���i�4�&D�\�� r�mS��r�K���$I������ΔP���1�����z�3W9ѝ���H>~6f�D��"d�*ն�2�:#8{J�������í��Z@!y�*�#)����X�\�A0�--slGo�k�S��g�d9��cFY�#�� �겱�k�|>�B[B�C���~��z��k�4�����@�9#e�h��mͿ��h!
���y��hbD?S8���v���T֕j쫧�Xy��+T�x�p�p$SU���6 �_PƉ=z�hŞGfAu�9��N3r?��i[=������m6����vU�A�|nv� `��0��C��#�([s�ɹ~�m�x�-�������0��+���O
v����۔طFJ��,��^��������i���x��;��9�����w�(��bw�����q��mP��͛�����T3��Ml��}rqs���;t�N˜My�-YIZ���U��-����)}u��v����I4�r�psuI��H�߷H-�MoF�Y9JM�`���c;���b�)筄:��[�2��Yİ������~l���9��őʄI+nRP�sWu
��g��$ν�qIW1��"��¼�+ku�~y��u��PIS��!�-�?�F�qh�S�M���z�[)C��ޘ��[t~�p�,x�;��]|<�߿�l�A�{��0�-R���:����9��)����=/���,�����tB�l��AƄQ�N�+����!�/�YPb�X[[��H�}��`��8}����ж��2R(���Yќ�/��Xz��x����X�Si��?�`ri��Pℚ望�h,����
7S�lN͈�,�j*�i��s/'�I< �N�<�P��H��$(;���>�^%�W�v�|-dl�Մ&����C��y��)7��]+���ɅӮ6��!_��b"f0N�P	�C���z�֘��5ok��j�B�| �L����.��0�̸H��M��mt�׳��7����,�pR'��L��7�(=��=Yʀq�tX�*��jJ��Z��X��:��iC$�3;N08<���bI[I�@����c[����gbn+=z��~��g��,�J����r��p����h�Z�AAE���g^��E@TN�u�r9ha)	�����9� �W$��`��"��-����PvK�6��\��P܎�H��\Z Op���,�\�w�� ���A�AשX#�lH_Z��T�l���NU�T���_H'��%����N3��HPiYz))�,�z-��:=7G��y�	���R���T����U�:��:(%�����`�6� ]�s��-$�%	Z9<�Э��������m��w6� �: ��p�zt̞���ݡJyd�������kؘ�&��J�U��f��N�I�������e]���uzR1/�l��u��o�zo�v6v��!Yب�L�ҫ�c��fRY�K�����b�*��Bk�h��L���-C�W�ʈ{��[=�[����y|B�M��pA�2��j���`e��x4���g�O��D��|T�I�@D�s�!�`��z[��m�nf��*��L�!�d:��������p`���`#��?��������ʨ�㩮�22s�d��A�l�����Bxs�>��Q� PF�b�A񧳉�Kkݛ��'ο��1��'PY�nt�3[�v� id�c����ޛ���\oZ��Ybױ2#1�y/8 A}de�p��9?�.�5���Y���d mf� K-�O��^���=8�'avo�Č��,L�'E�{���p���Jj(h��$��pr�)+s�����:��-�jV������n��|n�nm����Z��8@��!�b2�Q2M���w���Z h�(��;!�Q�"+h�1��C�41#<��>-�Hӹ�\�Y$��=ht 4eu����y�"�DQ�m���.6����R�ك�!��lf��`<�w�׆�����Ƶ�R�l)�	�Q�%4@@S:�K����=3���z4<#wX���Oo0�dk�X��w��sT��#p�3n��Dc-�e�`���/Te
�kd0sٟ����W��ʂ[�� �tQư�|��t�/+G�#H=��	�}�4�=G~��XP����۹��m����Yx�ڑ	��9��6��B�2�jK�豾}U�4A`���ɇ���^�a��e��d'����:#{�����j:sF��g�$���}���5VF���]�#-�D�tw+� �1W�~����_UW�0M;r�� �1C>�>j~�
��=���-��=�:*�SUH+��M��^:Rh?��%��%�V"�^5[��n6ZSۨy��Tۇ9(�>��L���F����q�XdL���9�f˙�0�z���J�_+fd�XnW��f:���@L�������a���<|~���p��{Epp w{Ͱ	U�8�y��1�f0��ߒ��w4rR;ID"Ǎ�T�T��EcD�axaQ%���ˣC��@�T%����E���ܣ9�;;܋ʉ�)[���H7ʝQ�gSp�&�T��p��k���>ybß}�R�,�Yq�5X�?/�΅�ꫯ��|��mx�L�@�׿��p���CG�^�x:֡����i'��?�2T��mQ6�{�����{��3��/���J�l<�M���?�g=H�� � �2�`H�x����r�W)�U��R��s�k�*E'�>�}8�.s�S[��b5�{>�����pj��c����|c�؅2��R�Y�>���^;���TW�>�A�zVeG��#�֌3۬/�BPD�$?D�s��"	y�x�����,��f��ϨW7��cPUK�B��䚉�].��S�ǽ���|����&c��X��O��LÜ9k�k07ʙZi$p������@3cF���,E��PK��q������B�|�5{���wtp^ �g��Ǹ �Џ�H�������ٔ9k=��p����6}ܦ)
�U���
g�碡�jgZk���:�f]y?��L����� TI��1H6诣����ρ3��3�����p����PU���O�*ӹ�Z�L*)��i1��Q��O������k�ᛳ�hVh�5mg"���G�JC�$'K�2�\�}Q�R-�}C+��fe��l({�q.�7d ���W��!x"sN�gnn*86i��sz����.��Ȕ�53�y$��ͯ~�j�\�uo�g�`� 1�]p�c�a/�q:��s��U�__�59�1A4��	I{� �1��B��%zPvJ�������س�͆�2�4mZF��?'̗�����xAY.azdf�p���
!�x��U���a�6�؁Tn��䳢!�೭��ճ3_���J��7��5ʯf�aa޼x:K[����� _�a��;�?Y�x��鈮�bc���F`0��S�%T�-T?u��1���{_��-���C�Ć�P�,r}�(D1���b��{o;�-2�)��S�S�Qa+e��P��R/K�Ll`4�zmSO��@	��o��z�7�Q�t%�Nֻ��+p�;��	��~�Oç�s��8��bP�9#�������砪E���&ڦ��1t)�[;�g�o1��襡 q	�,8Pm���zY��N��R%r�	�g�x�2Ld.>�T��AT��Se�K��W�E��вg�7cз5Û�s��[�c��$��Y�T��s��7�'��C*
Rx�ɠ@���F�)K@�ON�td��U�<�@��Јt�b��}� �����}BP��a��Lld�y���%�,��h�DJ>�p[y����5Ƃta�ֈ�c#
j �U��,f���У����5:�G<"
�ҿeG���)4��\h:��"�ɏ2KI�����z�Ke��<AQ��T��ަ�#yO���JU>��;��9�Ab��f�����l�uC�5#��� �O���dnY4��
[���MPەzt��zr���o߽��Z��T��zW>M�F��$��38x���F0h�z��Y�?�Q�Ԟ��O°���m�zq�^H�z��Eț�E�sN��5eӨ��0K��$���3RJ�$x_����s�L�[A��k�r�T�'y�۵���a��sM��&<�|a{}lA���M��);Ki��X�"<�܊۝�;�!_u���$Ī&���} ����eܶ5��\��N;iE���t5��x6V������l����_�MAz�aN�QEv:f/�m\U�*$�x��!m��ې-ř�'�HAbsv��2��Q�k�:�2���>Nx�X��8�H#}f�R�Z9B�7�'A��R�M�H�R,W:�_h�v�+��Y5U�b.PĒ_N��C�l���qx��R��O��)é�R���Ce��D��i2�m�tT��}19#�<�i��<n����{$�D���a�i	�E"h�)��p�?��}�c�Ȝ����.=(�E�c[��J�w#��^8��Kg�b� ��{����0���MX�;�{"��ڌm��ʁF��5٘�n�}���բ?���;Gw���޼�^=���1i�#�2��e�����X��g��҆LJe�M[	�@j�?�LB����#o��@�8�� t��L�;�ga��������G�3�ޱ=�����~C@�xF�P ���
Q W%?~�ޥ/�r_���g��>�����qJ���Z�p��D�h��O�����i�\�����<.��kx������7�Y�g"/�rX J��!Y�
1rg%�7#�}|ݍa�����k��Qq�7�C�Bũ̵jY�e�2�Щ�T�!�W�*8��l��C��!ґ�eA�Q�����q�Hf���-��':d�TU�LR%̈�pF��ȃk���3fCk���[�*!_G)��b�*<�(ml��v*�8�5Ug��RZBX��f�;�7Wᇷo������"�tk�:�`�@׈u��%�,�`�`�1�;�5�7k9]�����H�׶Q;��4����Was�ᝈ^V�������+�K�0����y��#A��pp6c(h<iSz�g�p�C�}p����l�����e`��J�����p
�݂�4�$T/h�\�&�m�	x綷!U��$���UC9'c͡?�һ�i\�./5��*�NU(q����z���(I2�d�xf��h�J�`$8K���ͭ����5���
d��[�Ȇ0S0�v ��ػs?��n�}ֈm4�L��E3�7|�l'l"�C�Գn^2{��)BEF�C$�o�¼;h#S9��N��Ă\�EM�bf7q����������9h)������jn�Ms������[e��[���o~l���`N��N�!����ц]�^(WЄ���͙ ��q��m�h�A��4�m7Т�n���F��3ޑYv������[i��?�����>�O(Ȧ�PU$&(c�C�3�B^*��YֵR���<4ˆf�PSs���kgC2�se%Y���A3��oa�bӐ�,}a�A��2z��7�on�`΢f2����F��:���c�(7����P�[/�Cw{ԂR"'+�h����H9%f<��L[�h��vp%>�=��}%L�@I,/u�(u���ͨ��-����B�]ˌ̰\߅���L����a��jL��^���B��<2��WB�yFI�8U� %�D��$�ўZ>��%�A���1(���,JW��'�g&��穌Yl]�Nb_��u7V�?����p&p_wBd�@|1ˏcR�_���a��v�D��D�2g�XW�R�R��s��@�7�{�Ou�0(���ѹz� �����:���0��ޚ�H,](�	���?�_��$h�H����룰��4�E�G~8�ic�L)����1PJ#��h)O��0����zr�V�A����e�_���F�w
0p��1i'��?54�z��z�̎�6Z�/���R���1�`Ks�C�*2��aOgˉ�c�\<����O���j[۹F"16�9ћmwa9�윘=������p���K��!��,$s;��Mi5�~���w�lk���!��������"�ˈ&E\��z&IKs�"�1[�$��k���R=��W�)�˄�=�.���I`L��A��hؾ�����~���?�P&fÀdi�p,>2G��6���=�ۑ\��6��u4�b�'�\��TF��jm B}����.@)�� ���� ��r��t{l��I�\];�Z3�A�}ЂU9�� dAB<�d��U��0�y7g���\%>�u[�CQ�����t�2��O�T+��S���2�Zv���K3��rmk��p���PyDZ�/.����X�"�� ��e�����r� �\�qi-d�5�C����Si��
������W�	��_��p�k�}���?�������z2����~��*��������Q�����Z�b��F�Ʈkck�����>�9�)�����c��d���� �rUK�u�{k)�$F���(��d4�J��vOdsP�!.A�4��)X�szM!ʠ�K���(G���=A����Ĩ��E�q�l��s|�$J�\$ݰ=42o���HN4�Y�B�Q�LHk唚� �<��U��\�T�"I���~(�5#=j%�7�p�Rsrg+����^�lz��ֆN&�
`�1:�d���G*}.#��(��U�"�2�����V��'3д@�s^�/�G��`A�g�<E}D�l��:�YiQ3�L�z�|�jBP/:�Q�R�!� �; ��^4�,s]e�b)[�~.���Iy��pĠ���w%���j1'����o���`����n����Ok�����������N�9=ֶ��=+��]��%���1�a��$ T<>�M`hl2���VN���Wֿ��pP��X(�no�÷-�
�M` 4��d'	�V�
F=�pi�:�)=*3&�Ng"�����+@�)̿����2s�~x���9
������7_j�_�\�?���j��-p�|V��S�ڟ�fG`)���n?�Z�P��Ǡ���O"�ȧ�N����}����4�k�m������\=g��Ԝ>�i��=A�
YY��s���G8��$��"���h��+�c}����:�\H>�ҕ��J�5�d#ɋ�O&�U)2�UgS��4ET��`���	Q��<���/��|̝9]n�H'��et�:���e7��P�m��/5Ξ��0����f�Ȫ�OOaǲ��08c+7��Ӊ�}.'f*gsg�*�z��!A��}g6
��V@KҔ�0�>LA��8r�1T�p3}��%���oZ�{>Ov��f��._yV糘�z��=g���cK�VtG�Ɨ�ᴏ��Gm��r.Vv�l�7���/�٩
��-�)����v!���a�^ ZmT�X:�,{?�� �������xvi�0S�
89��G�𿀏�tP�:L"ηW����a�KR~I/�iQZ����\(O�J�ՅD�}죊Ƥ}�̳��j���L��8Xz(g�Gۚ\�_�������2`J���lS�t��ͭ[\N�7P`$'[��Uπ,G�tmd��R9�P�$���N���\�ąLp�dp$>���@y��Hc?�/E����PZ�U7�6(yv8;�F�k����8��g�dN��)�,Yr4v�<ǎ�b�Ԗh��ۮ4��g�l�pe��D����6��H#Jr}ϞgvE(D;w�O)�A����u:�a*�v�E	��� �M�P��	82�V�폏�zO�����@G�!'ȱ@�}�(܋/_���~h��hH�[IßE� ,z����Z�9���7zo��ݝ�@���iv��qyqf�B��Ζe��03�v���U>�v�T������Bbcvjǲ޾=�wv��s8nD$h%���{8c�-h�փ��%.���mߟ=܆;��ω3�@8�Q���%Z[U�����c��*�o�}��u¯����ůG������s8�����e{޵��[U���Y|5�M	���I���!p�]�c(w�?�h�)H�g3Q-$�PϞ�F��jן��Ɡ]����J�ߥ�.��Z#�C�lX�z$L*́��]�����0M��CyH��R��<��]μj�v.op%p�<~�.��S9ڲ۟i�#�|pSc;F9Z���j�\��45t��7*^�2̉=���?YT��)Ά��Q8���@��l�t����1�33jw�-K��8���;s̖%__)m턮E�`J�n������7J"����_�����s���� ���;���hz�k�8=.Ɗ��9����ŊQ�A�,J4���%b<��TڰM,В�=a����n���`$w5���4��sy�G黕]��uC%��c,�\�۟��7]��'�僞J2�T�!�L���� !t�|��<6�3U����LYF�"��% [
,��IU�t��$t��I�2�2�8�R�_B	G:T�r�&A ѿS)�@�lʰ�P�@��Sb�GL�&.�O�gW��ә�)w�,�rz�Vϐ犳�Hy
G�����[��zΰ����Z۴&����-۟��l`x�;�ZV;��p0T=��*�{^�G9�����m3 X	F�	�k`�rl�9T_�8v�S/RgH�xJٹ��7�Le*'�_#f�e���a�"�)�%N\!��L�m&�UpK��F�هf�S�w�z��BV����B�d���Gn �y��W��:ե�*rٳ_
d��~�çS�\f�m]'�"�{{�5;?x! e��	�a����_�	��J*ԫd����?�:�j�YwQ\F�+�L�[/_�L��-��׿V����O���K��L}n�JƠ������
��b��YX�B�aB�Ӟ[oϜ��
�TA�Xq���#���ˁ6Q3Ui���vo3���?������a�?�Ϡ��m�_jrЙ����3gM�EUi��o�f�go,�z0����_^h�2`���$����^y��w�j�aOA�/�,~E���,P�f�T�^KZ0O�g�AM{�5��4mD܏O�h�@{,���VJ�6IS��aʚ܉� *ƿW&�&ٚ��6H�NV��a{�w���R�ʐ%Ν^���fH�!E�0�� x:U�S)��^����P���<

�H�ճ �E����o�N吼�{��6Ş�\Ur0�ʝ��5Z���ݻ��
���#�;���{/�"���WԈ�Bt����>G����������߆wWgB�,�M:��`�^9X(�T|͎S�q=�?Tr��@��ܘq8[Nm��m7�p�B9[4N����Qh�¹}٤���gd���kS6�X𓸪NM�N�"RƬ>����24F֮�ٴ�3�,���V����xaP��A(S~�?��*��Yаj.up{vp��qo��tЍm�}f��c{��Gs���abw�(\�ztR��"�4�TD��n)���e�N��z�r_�EH�ʞ��.x?S�O�+#��E|����*<�5��]#�O�ړ=_�� *T|��d�mҺ�V��[��H'�XK�Uѐe��zc��LGγ�d(�_��,AJuY�.O����{8Y�,c�
����g��-���S����F�k�8fS�/������/`g�7����S!��[�ȓ!Hj��F�Cp؞�xȫpg���oA��~<gS��v�+�O�����G�\�0"�E\ce[�8]�aj�-�EFh`o#��u|t���K��� ��'�g����^�}���Zu'�>�z9������]\����8V�8��X���(��ݖӇ�NZ��Ys���f��L[ݰh0ni��ר�06�G�,q��=Yt���)8�8>D�5�TrՈm*�/��W�� Q�P/f���=���T`�����U�ʟڪ�B�d���1�i��\$wX9��pgK	�`G(󳛫pg�ڃ�Ih���2m�3��Tf�����l��Q^E�Q.	�D��\��I$��̒Oӵ+�9_CO8�v�LW<D"=��x�E�0�eQt�rtw(	)YZ6�$�p�ƪT3"B�-S2��g,Nq����c@��Hc&�^���!��s���}JJd�g��"����h'��D+�ԛ���Y�|��ԜaS�$t�����L2GG�2�S�F���^okv����5�p�1�Ӊe떩��B��i�%�t�1��d"V�NJGxq��zð�M9ƥD�g*�(����wo�[cn��;�e�IS�JY��ʑ�2E��m���x`�k3�s��f�)�ƹ�r��[s �`��غv�MI��N�td�kk��:�V�3�A�h`M�%�Ele���m��Z��Z�\�,dZ���ߔeѕ�Yt����bl��<�N�}��C��K��X�����+�(�R"ʯ�<k��xn��c_���g=�HZ;gU��/n;�~�4��v3 ��@��*�A������]��`�ќ3��3屗G�P��i0Y��4k�q�#��2�_ZB���'Smii7��.Gא�o�����!$RhN8��:d����Oa����D��s�D���Fj�wK*>9.���&��g/�x��LXN���J-n }�߳h
a����pI!����MC٥O7@�`g����0�0�R�T�����2��hs�cMR �Z�$Ƣ 	ڷ3O������9�}A������>'��Թ�8"�dI;(d=f��x�9*���'�C�)t!
�n�P��,%����@�G�K��V���PU�n��>j���T�m�̆�N��M�	��!��s��ּ�*A�� �1s;� �I�
:�K����i�^76���}l����s�	�E��&b��t������e{������Hh�Fx��k���Κ�dE�ā���+@BX��F��W�8P��:��]�d5�T�qoQ��V''�H�F�Y�#�5o� �A�ڻ~>xt,=�ԣ`GS�ak�v�8߭��%��ҙr c�)�͈�3���p�����K�IƖ)�UV`�@����(w��=J#��� �^���B��#;4�ab�c"df.����Tܷ̙6�ME:��L��L���������&�}�.���,�e!7���e���ۓ��_��Q�20�n����x��jWOk�]p��C2/ႚ�Ԍ?f{5-�?�}�1L��̇v�����>C���^��B���{��D�K��;�$��8`
��\S�"�w:�-3�2������_3(���i�Uj/�1��e��F;�O֟�K|����T	p&V�  ��IDAT�rZ����}'�B�zow�z���^��Jg��<S��A�eX��ݪ�S�_>��Us���i����U���V�v K]�ƝY�zEa^���f��e���H�
3��Ҽ6_�;� 	@��`sG��w�N�-Z�� F��s8/�A';C��+�D�i!1�B9'.�����m�f��3h���^w��̰W��-E�O�i+�1�<�O�,;��aD�|�2�m'Q)�=*y�U�?1B�zw�ŝD�0@geO\��W^^M��hK=�`�l��=�@��P
@�9aH[��p�"�HD�I�� o<�zDAH�>:k���|�O �n�&Nv��{�9��4W���ed�,R�ӳ���\�`�\"x>��Mk��D��~��q�MQ�O\���,##W��<J��྄���k'k�ёF�4�-]fT`V {�L�P�9l�m�X����"L^>�*)\��y��}���VB����݉]<��Gl�]+\۔��<�<�;5[%�v�u���sgs?qTHY߮��-eM���}��X�
�݅��+a��N`}3����	�A"�eIц]+�yM����$<;_�^la�d2��2���dDx� ժb�-t.*;3��x���|`V��Z�V�� ��E�hȶ>�0Nn��H;F���0�UC����RGRr�ȏ+�V���T�7�B�f�!j7Ԑ��A�g��(�6��yS�r�;��mh�ᇓe?�����PNK� ,�Z��*�H2^�w���,tT��3���ۢ��]�6���0�-R�΢����Ζx�+�t�_��n�/�J�!x����BKV8(�R<�dڸb�aF.�,#�]��:�W(��*@n&'����;��Fǲ��*�|u�%�e[���l�n۵IC�s�R�A��p~^�(6b�= �@�t��J։|��T��
4d�鶖��ӣ��5��Z��H3s��U,a����=���$R�+Q�[����c���	�4�D�D���XS�)Js՞�܅�2����r�B3��9sUM�!
�2Y� U���_pN_��J�;ۡ�1��g�)=A|O�܌��|�
9�*l���=��n�u}��]YSIF����s��  ��
���m�q��F�h&D+A�'0��K��z�%p[Yp&r�T��%�.L���Z���ܳ
���P$p%q���Q ^"�C@���&@ߒ�a��J
xR�b���u��:N;Q;�L-�2��1�PkK����h�I��+�ԡ��U_Ɉ��>���j.��<+1Q!x �Z:r�U�`1f�c��2�Ǘ�q��Y7�.c�ƛ{e_������;"���*{^}{���XFp s��.�/�;4��Q<�
�hs+��|��!g�@��_́��桙�-l���R�|�]&�����hk�Q���_|<O����z�L��6���|��|�?έ�b-qh����i-���0 ���譩����}�����i�� ��x�	�mh{�Ck�ϕ��7�U��6�<Y��
zD$�bAu+)��wIX�|ΈWJ�V6�oʂ�&'�@y�>_��Ξ��E��yY�.�x�\I��KˍX�p>[!Ъ��[�5Ek�z(���q�a�yR*A��5 ��^��9�0�2��s�\A�\\����F��9Q$�[^���%�D�MW��H�!�GT����ot5��P����aN"�Ռka�Xc��s�C��5���>�G�#�v��aa�0�o��ʔ��>��j����rf!T/,".�����e������2e������=�,ɮ4���O�V�JWA��l��W�����
�k�q�F94�h��h�P(�:CG<������s�GVS��CGged���ޣ>����@��|w~�m72���������W�!�bP��Ϧvh;W����>�� c��,�����F@
�Y��\� ��=�+3���IҞ�uxC��l�nv���?W!\�d�穴�	d��E�W9������*��Ρ�ỵ@�S-A����ZլՅO��R���d�g��ݛ瀚'��#r-������|ik��UW꜔7.3H��x/.�ώg3_jg����F��.(@e<}d)Q�P� ���4�$~��i8�%(�\��^,��@�T-�H�s.�IW��(3��yDr*�s���<*�G����DA��o�v.�k���V�<���8+�y���~_��Z�u���j���7�Iˢ^*	e}�-�"h/cV�i?��G�T����jn�_��t�@Yk6lg�����huI4z��%x�R�+�ڴ�^-���:��?�Lƀ�l���>��4��������?����
�a��F���w��7ߧ��>�V%��� �0���V��P��g/S(5�LJxn�υp^7����U+�2����me�%g�֦^w�p��Z�.�^����KR�K��z��#�PZ�t08_wO����-	֠��~Ғt��v:��*�F!�{��M��E�+^�64�,��]���j�\�x�)���=~rV(�ra�ɲ�OUA�d˴%��y�+7�s��P�l������DuJ�L��ᙝM8d���9�ø��:�^�5�½��5\�q�j�<�C�I7�r�?�Of���I�����@�����N�$���8��Ȥ�L�A35�LNR\DX�PA�k���OON���+�O��;���S蔔	+�f&���-rjQ��M��7w�*��M�Jώ}����NZ�]*W!�� ���B�NU<�8.DN��>�@�#�0��woӥ}	]	
W�+Y�q�$Ȳ���$�h�Bh�����z.Cm�w�q�g:$�	N-�����
]���M���}��K*T��´�Ce��_������|��w����W_}�`��\�����-h�t�w�D���w.8@�A�Z<{�$�W����O����E���[�N��V�x��+��8�,0-aి|w��-�����{�r�`ӎ
�e�) ��VC�"��>�ˍ�1v �$�����X8/ea
� ԡY���n ���J{:W\mt 8�B�Q�֑Ǽ.�ex�-Q��Xu�I@�(��J�$r�i��$��k���L�O�j��:Hh��<���_�lI!��J9'T|�UW�E<d�^d$w�dk���U!�Z�˰�c|r��d�ѯ8O�Q�Ě��l��S�s:�$�T����$�Q�hw[�����3�׵p�i��gcݧ�Fb|nY��Z��<�'��3ivy��,�]�)Rk�
Q$�d \Ž��}�$T�B�w�~�wФ�S�pr���)f\k�N�hsO����~��ME��U��uR"��2��Y��`-P�J�$�v��<}�=�>��SKv�����W���;�p�"��v�����=�{J ��]\�[b��ma�A�˴ļ���G'*���W���j&l%��2�f�W�c�d��&@�I2��<4�;���V�'(���j)�4��)A���r�z��BҖ�����r����@oE���@���z:�J�n�}W��A3taC%�
+�6�.y�g�&,2u �a�y���5�`�!�#6@�!]Z�4�f�5ʢA���;@��,��p�t�=P��e^#o��	�e�r/�w�"^��O��A-f;(x�Q�3go����DS�����CT��@~{���X�r�=��:2{/s��2
p��ޖmr���F�~S��Q�ZXlf����	O����N��Q��J )���4s�jDY�~��F[�d{����x�z?:>M�}�yz������{�E���|s�����{ �&ȲO#A��vn~��,���b�±�	�5F�XȩR�����BF��9��w{Ko�Nή�m1JϏ�����v����3�����`�%(��%wQ�ֲ`���lXv�=} ֶ&����J��@�/G��1�h{�y��h����M�s�-D5]�jJ[�^����D{��+�+���H/�J{vH�^I����5�N�
ʟ˧fQ�����l���h�Xpw'f��t�)���s@)�ss?�i��2fռG*>h7+��|���c�Z	4�k�Ύ���?7vͥ4T�[L������S�3��Ź(7x��hC��ַ�,��~��e��uw�������|ѿ�*���c{_C�z�̲��4����3���	��:�u�KAΪj�|�墲�[�>��ҺQ��A��t������i�ۡ��_�����u W�6��lqr�<��Y�Z��Wě��Yg�;��[��dk�>#B���
�"D:H@��~��ϟ��O�>O;��p�r��BQO�:<=� �IQ����G=����kۓ�E���O�ȷ�sCkb�Ck�8�[06�B��o�]��Q~(ϗr%�|��|��ﵮ����nN�֡`�dr�&;��BӔ��r1�@ ��H���{����X��hO���A�=H�VA��N�5�V�e�}f=ᯂ������]�qKv/+�$�:<�r�b�M�G�I�N<��[���M����'�RNXhC���V� �ME�/ɹ�)���ɢaE���zc_�:ʄ�� �<�n*e�)M�I�aV7����[h���tR��u|��;>[�J�߿�z{�ꅃI<Њe�H+u&k?���V��������rU�Y��m,���W�[��.]O������Zd�PȖ�������hf�$�����g魃e�N�
��[��7�L۳�b�����X�D�IR���#mj��!s�!Y�ݛ���y �,k�'*o�u��T��[��Lp����ގf�t�b��y�<g��A���k���JZs1oŻ�B%� �t��N�'�1W8���]˶*��^��l�k��,�JKq�Z��%�3�K� 4�V��s�٥�(l��!A�׷ ���#�Z�/q����w�T�KѻQq�mqz�z��`���G�p�+@Hj��¯�AjۂF��t�-��ڂVΒ��!���Jg:�_��/��u���kU��xIl��U�_k��w��0]$,!AÓe-s_��H>�� �a�ʾ(x�_�J�,㻕�vR"E/�S��t$�\�R���~ e�Ƙj���}e�ٮS���������bѱ���Y3��E�����Ӂ��;s�D�_8��[�w��$�8�����Q�,��X�n����j��Y��,�'ѧ ��'�t0�&u�Ty�w��]�����'�S�˟����h�џ_��7�8�l��g)�X�0> RoT�&oy��L�}B%r���\5A�*�);\|Z��[;���E���o�o����;ڬT�^�������켍CG�Z$��Z��P7U��	�ҏZ���+aeDMX�X�f
���4�siF�y���t���qnAf]�!TP9�
$���%��^"e���֍�bK�<�$.�7�P�Hݩ���-���D�ڪkwP�\a�b?����	d�Uۢ����!4]/��D���6L�Ꮶ6�Z	�P�%d΀� �5��񇋢d&�us�Q�Y��x:�Ѐ��,�}�7������VG�;�	���CU\g	��u^8�Ta��l�Fz���y��"�5�
�r6
�"��ަ�w]x-����[�e���ew=�J���@|�εU�tw��N����+a^p������{Eb���Ѯ^(pֺ>��Qj�����h�q�%�.o����k x`D0�M��{)JR���Z��ʁ�;2�A1,i5��$թ�Ł��pk�Z��f;��](�R!�b�Y�>�:� �t]Fl��8)Ώ>�$����歨A�7����ltfl���dׅY���sK>fjQj�4@��Y{w��Z2Yr� no�,O�\���r���wqs+����:x58ьU#�p�b�@R�z��K�;��!�^_\����ݳS;OO����]a�U�(���0� �	t&|��]��Xf�)�QUvz|m�F
x���XK`��EG{tl���F|����R(��Ψhz)��2�	w�S7���}�>��|�TP߂��𽞺��\��u�,A��zg��%;W��,�k�Ҙ�]�$NI�Gs$�{����(	5��3?��W�l�-"+pT\�Y�	X���깪�,5����\Br�mh!��K&q�L_%�w�5�! (�B�-��_�F�3�����;�!� 6�n�/�--��"# �Y�FWv�������vT!��W���[0U]�}�H��K�y��Ӽb}Yܷ������"ra��j5K_�}�^ܜ�������IN�k�d[��%�-��T��h��o&��w�jUm�BP�1����*�4�6\I�'��.���{Oָ5�M����O[�yH�(@CY��ˑ��'E��_�,+<�C��#1?8bY�j��	�[�]��p��(�Ц� #5�ܘ�g�)�M���AnfR�6���.8�ö���N^a)a�L����I����g��9�g1�B;N��w�^J� �#k��<x;����Z� �����la�5��hߑ�O�<I~�Izz�&]`�������	-�\��]����#x���pM�{�57�6��T�K�N���+�5�����H��j�U�����:X7�k�ި�Zۚ�ɓ������v�~ש	$v1p��Z�\~&� �N��f���g�W���ע�P=yt*@��v�v��C"�)������6��qP�A߳�[v�������c�	���_�g�;^c�Tx0�PEok�ݥ[W�>H/��� q�Z�����R����m)/��vj^� P���D�	�b��KԦp��K4Rv�����6*���0�u\K�-���ɭ�j	k��C����o�������j�Ud���vI�h�W��#>�!i���\3�+t��lm�,���ߋ^�̱ƪ��a��]�%�4B@i������W��oiK��J��������I>�n�*�>T��oԎޔ2��}X�^F���ѝ�]�v 	0�Fi]�N�+dZמ~�K�Pƌ"�K
���k�qs``vtt�v�沠@��.0� +��M\0I�9��9z���l�R�p玆� С��>�x��p,<N�im ˔�b˷�1��Z��x��=��MG�@@N�z9���/�H_]�IgW��B���J.R�?���5�Ƣ-����}>����g���Y�����m�qr*��=;xWs߬�P˳�|y� �+�ؠ�=�[� k��̓0%c#?l�~L�����W�����L]s��Ѥ�)�IZ?G)x�9��?T��#���{S�^wVQ���xC��.ިtO8�n�/eb�z�j��o8/Dt�+�qb���G��ޮ�ൡ�1�~��pvy�6_��-
>Ĩ����7?�U#��BRR������L�������Cw��v��!�܅T�>�����ç���M�?�1�7-t%G��JU���z��e:�;H��'$Ϋ�8�7HZ�xm�cj�������z���:� ��-�퀞"8�W"��w�V儇���b�CE�p+L06�>Hl���#��~Vkt�	2z�Ⱦ�ş������Y�fmn|<F l�Ô���(����ѳ��-"8,r�h����z�\�����?�W��ֲ'���;�r�6��Z�B�=�����-3pʕ����&���O.ܻ�U�`5�Ŭ:<1��3��|/���n��'��R��K?~o����c�zv���Z�Et�6Eʑ���=8y�k�jZ]�l�҄�p�v����9ْQ��F��l�tQ+Z]�2�t�TE�;�t�۰<�+f�됖�|��縴sA$� ����wq&�&UD�/�{&Or�BQ4��H;��ɬ%_��h�C���ڜd���g~j�m,;+���7�w��V��������Bҏ;��T�����6H޾j̞�r�b֪��o߼J�W����Xl���0%���E��0�p ���,�gj
t �ɛt������� \�Y���G��Of{'C��-`|�⻵�?O��a��d���6��r����l�J���`�,�+o߷��&�2Y�����t���{㴾�*�o�*���lt�1�Ϲ@Q� ���9�Z���RhN�Zw�x�U�}�ϷMơ@���t��Q�i���j��7��C5j�z��q���x�k)����P�:6m�x�|�b�p�Q����T����1!��p����'}��xy�^��G��k򬷎CU�|9`�gܲ&���X7��Yr�"k����������5�~5w��﹭C��8@�d�f[�k�ʻ�ttԁ	D��`U�U�<�ONR���j_��+��U��Vii܍���EZ����Ī�k�ewW��F=i#��J^��^�Ģq��	�2��_m�`��RU7���O���Z�CF �Qd��*K �?~,`�-ISpQ����]�޹�b������I��.
v����;�ן}���=�?��~Mֲ.�n< s��zpf�f�q&�d�Q�6)���.|��O�}f�3�����<�J]ӻ{���Y��wu a�
ipT㍝{}����,9��	[���hфmӍ�<�i�7l�����￴ lI룣c��H�7��鲻vut3�A���{:R��x	I�8w23������>�l��e~�X���o~)Q���=�\8!ΛyU�V�
 k2�W�E|�L�C���0և���8?Rt�W^#�+Mvl�y��&��'�^�Yٛ�<l3x���C�����;��l@Ax֛�~�G��	���eZ�D A�Ȃ�Ֆ��6����Hawۨ�]&n2A���ŋ�����L����(Љ��=3��E�z�psiC�×-���UfT��meC
G��+W����ů?s>�}�N�ߥ���=ܖ�We�ד��td�M8�@��\����5<c�G�pG��,����4��v�tX-ڶ��h���g	2[�z.;׋,�-3�����T��� � ����=�p�Q˥t��'\jG�G�����x�Bb�T�u)�.H�N�!�ބͥ/\��0SqW���SAm�VH[���l�VU����8�cZϥ]��Q�E��a�%r;,��P�~��ߥ�w�شCkC�Ш4�^�G"���5�D�j�I·J^��7�m���ѡ����FR��pX�=�:J;�'��z�(�:x��q(q�2E��?WVh[t����"�;ܔJ7�Y�������/;N1�`P����y�.�7����×j�n���_�z1������%��2ڢI�a�Bఔ�u�z�3�tc*��	D��lt� &�)�]5��2z�[��;9<R�{xx�>��4��ق��)�����7����C2�,�}O��;�˴o{�h�@U0�pL�n���ξf�@��Tk΅l��LV��u��FhK��,�E�� n�����P��'�b@������@�O5cS����pAܫ�DAc�$�nɣ�4/ڵf��Y��Nm~��z]�F{� �y&���܍F�EW�x$n5F���Q�B.���u�BFW���:q4B-�����oI?�m
���qCm��{�ׅ�����vZJ�%�f$8�v���܅F�u̢����E�E�J��q����|���ڑ����>�o��䟹켏�.�܈��1�'�F[�,n��|۠��ƚ���P�$0��Y�B�IѶm 4H��P�:���-z;#�qH�;~/�P����d�,]^����s��W�V���ʹ��3
!iK�v��������~�Ĥ�G^����yP-� � ���U������N5�����w�v���3ٗe�AZ�S;�ok׎��-����A!9�]��D?J����婞��:^�vh&�!4/Ckۘ�j��Ո̿tKF��|�Y�4�Y��}kq#���_@=d�E�h/�q}5[m�ZI`��-�G%Q����6c)u���@�����K�@�����M�ȣ�>	A��Հ���k��|���:-ə�Qp��*Y'9��h�'�[
�z>4��F8xe��D,}����<���rJo�	!�p��6��ɡ�T���.��l��խa*:Dσ�x����Q*,8�7�YN_[��q�ͬ�,��T��^��gO5k�b^�{G�Jr��#>I�6�4]�~��YPb!�����z�4�!�@���;�����*��U�w�~��T0�lR'��+��4A+�߶��;�b���&��p�r(��a�'���JrG�D:Itȇ�- a���

{H���&�(�w5��H���C�t (��?�����*�u���H
�*��ˋk%$i����y}9�
�]Z؁����GR�R�ŉ���Y�?#�G7�5A�#��j(}l��ٞ�]L�sb���֨�,�H:
g`���d��R9R!G�<�N8q��5���ٚQ���м�!����_����W����~͞�)��$Y�����C���� �ʻ2+�%6
�`_t��nY�Fm(i�1	-��Q'TB ��ݿbk䒬�:���mic��H�R���I?��3�u��<�=Z��om�]�1�M;����|�m��y;��Ѹ�$�zr�^��O緷	;�%�{��J˖�����3��s䚻j���Ɇ�:�
�ǅ��n{�+R��{\�BN�n�L�W�~*W���~�&�]ԝ����~g��~u�bj���=��٠@��s�s��Z�{7��p$���ήԼ�	-[ݶ  kn�����T���&�k9�L{aY�v?mnW�dŎi9�0cAj����T���TN��+���H�B�YC��Md�1����3��{���r�$�hnՏ����+t���sr\c�����'<�e�&j|����+%�<SWOr�=��]��ɥ2���.L��ȍ��bc?g3ݤ���D����u0f��'�@ #�tBHָ\RH�
��Hx�sA��u�ڎ�Q��
<R�xu$w#<w�1
�����L~�4<z�>�7�J�x {�vP���i�Y�$�[��؈�����m���J���[���v�JW���.�H:p��k��i8�sD���6oS������Uz��u�Z��hf�$Q�{���JQ��Y��ӕ�/���뙤d{����+TM?[D˖ĎQ
i���q��m��{
u��� mzZ��;#������c��eYb/��X�*K(ґ��]�Z�7�kT����٨�Ჴm	9����?JǏN��In���=�@O�U�G�;�UK�����m�t��&s�P-3�CZ̸Y�6�&@��	#':���Щ��q�����.ܗC���.>�T���;�a��yTЭ��$̓�j2����Z7� K����K��#V	5�X�s�;��t90��粸WXLq���eXS��t���r�*I����{�r N��Z��r�tϮ�w���|ظ�&3i��H>7nJ�EܢcKQX�Xh�o�y�������i�=I'U�Ξ���T���.o�hI˦i�3?]��^�^��EH3�po!� 0�h�����{�ju�����s�p5	O�\�pұ�
S��"���� ����<�-������Awt��>9uA�9��,ח��/�����׿U~������E��ܺjL̃�&�������v0���VQ0<���M�{WW>��{m���7��Qq:�����,�^4�.��jǅ뒮˨������h��4��� ��E��`�c��7��E#��RW�7aYwc�9�OHd���|0ϸ��:��7�w��@ ������رѩ�c1�ƣj�Q&+�,�FZ�(���u���J�-T���N��ޫ[.&UĴU��o�ab�@�מ��0]�M�%�&�����n�ԝbv��q�G}�jmj��E��mwm��x_��&�'Mے�>h�E�	\���A:�J�|�#u�X�j���n��ͅD򡖠�utr��..u���O��T��u�X޼|����w�9�vDy³��	���r.kL�G�	�?nv'~p��]:!e-1���ܥ�k�������M��tĶp�?�ĭOroz���w���;;K����̗��r���V� AB��7NsD��v�2��H7|I��Щ���	�7VpM-���Q�B�m����u�A���Oh@-㤡U��E�T�^q��!�G�B�ܫd�gA�c�,��z��������9�.J�|t��旍�Z��o��6�~�J�[���$�Z{N���c��ѝ�Ɨ.=K�WX��^Q�K��%����ep��h:ܽwCY1���7�GU�8�\�ljԝ�F:��I'��id��
A��NaT��q�8z�f���a��1�N�"�b,
��#,�D?}��Q�髯���a�@�xG�JRJ9��YU�ζ��X�l��:@�Q���ĕ52��Dpj�rГ�2�6+���K{�;,ά��P(
��f��*����~:��6# ��U�h���
���?KG�>��7r�x��]�>���2c̈́�0�@FA�f8��&U�O 6���?+7Uz�T��x���(������6�<]\��?�������ÃG���� ��},�zm�ۢ߂G@P��3w�p$CĽp@��t�@��j�H�#kU��t�	�`Tv�2�3_Z�\آ�<���yH_�r�-V� <U�:	�לD@�c���+���a�X2[��8��@bg����v�ֱ�PFk{>�B��΂� �ЌM	��8�5��`S��������v4S��B�L2@��{0�,|�J�]|n]���K�:؏�ܰ�rP�%������`L�j̒�]���ܱxb�c��ª)I�h�Nӣ�C�1Z�h�v�h*a�د��^����[��dH���@�/��ʼE�q�d(����p��wgkW:�]�I����#�\Ҿ[�^��ڍ
�I�j�xe;��o�i�lK��*�=�d߼ycAr�잭[�b&��u��^큝�X��t$��B�6pc����-(�~�˽��� �
��g�ӓ�G�'g�<	�G�c�x�oAuI��#|7ugs'lA��9�3��;Bf�)$W�1Pʫw�Ô!3P��H�ei�����Q��3k���~Ï��W/�yF�c0x�5�M����2�\�^��2Nh��Z�;C9:��ɾ�r��hM�j!��*�Tz��U�{>?���2�{^#�Ë�/�D;c�wҳO>J��-�k�i�s���u:�ݦ���\q*ˁ߯��#_���=�Gn�c��k���>K����M�#���#� u`�zQ�h���N?���$Wj�u�ѡ�AVr�Q��X��\��h�of+ׄ�kF��X>��S�����(Zі�N�r,��N�� ؽ�H����A��y�a(�^K�N,E�ǖ�Vk������g��>�N�MR��KT� ��E����2x��tA���^�z�'�@��7������W_�Wo�t��G���)��P��V��Rm�V�Oᄱ��m>�L8/�����7�PuPUw��3�ף����M)�nb�|���X{�	jPx5��+�������&��R�hI�KoWo ����1�jD����M&M�hf���%7J��'<hM笙"���T`��C�Ͻ�>mlt:�<>=},���}��?{��������=U@�'�������!�F<�	)�ƻ7�J���	�H�{mJz�S)�*�|F��BSa�:T�21�5���d�k�+p�d��:=����}U�pCgv��g� �N�q��k���!d*��r^10jm�˹Ь��c�jìw�V7�4�l�R5�-
]�/�d���8�$(\j3�� gm��"�j��$�nDM���.�m��K�e�8���-�>:�\f��*,�P�S��]\I|��H"-��T�������?umt��wV��+Bҟ��4~��0�Z� k4{Ugr���쪭O릣�I' �P#�KЭӌH|d>Pރ���5*�j�ty-\�`�P�/Cm������\�y:�;��[1�v܇��W�H�s �ɸ�r)漲��ǱJ8�P�(%�Q]�5c��aydH�aCɄ�]�,�:/!.0��Ŋ��Ȳ�йܙ��/�����_�
��ZR�UH+F%_�m�����,�����xG�<�'�<A�(k�_zHM���fl��o������d�m�le\:x�#څztt��?��ftW�/�"LY:q}a\�È��J��JtؓU]�
t��U)H[2 �<`�$��S�<����4�J���{��k��8���9�r�*�?t�*ti����B*�l������ԍM����~aA�����EpfQ/�X�*����u��k;|ik��.���p����N�����+�w6P},����A��ls�[�u�P�9J=�
Y�t��
�b����V��=�
(~�\��RI������+�d��LP�	ʼ�ĵ��L���W���������7"UxUwT)U�V��!e�C��d��#��/q)�`�H����"�?{'ay�H/6g�!n��M:hl���4M��^\�p�x�V
F��K��q Q�5E���r@�T�옓����l�z�ܘĀu��:��֗���J�;��_%<BbbU4s^����E�ʿݹ�� V�{V*s�%��<�L;=��ǅ�y������D�%�v%�>w�ɾ��?����}�:�e�l�m'�� ����RvE+�Y�ފ,3��?蒱\U
 )H���|��+Q<�V-KU�vIȦ��
�9����ʒ�M�m�;��O*F�R6л��ӗa�?����ܣ��������7��)���ӂ$nFg���4�E�dtSDP� ��Gn�k}E�ݏj��F� K�����\��<R
ի�ݎ61ߕ����N�(w������v�x6�ɘoGW]7И�o���.��ga���z��TN�sW���X�I�q������N+d3��N����I��F��k�wڢ���ף'��s���G����=]׷V@A9ݵe���(nVR��$��x�ֽv����?���y��I鲔�I�	ylAc梱���҆�}<N�[�v ^�]�B�I�ށ)'�ӑU+��(ޯ����N��p�R.�)���U����2� k~��Uz�򕐲l,��]ۄ��9ܳ�o_l��tr��v	�}�[� �ℂ�mF,�_�
l���AS�S�u���(d�}d�E�v�����ttx,t#����
���m�E��о���6��~�n.C{�U�C{�C;��m\�fi�P�5ai�siٌ�RZG۰�D&6�x�T����d�� �r��;���EՑ�^̪�³{���8�Cg��y_	�P��������{ U5
�B�P���ֳ�C�p*a�Ch���9�P���;{�6��"d�0wA
0�=v}�:���y��t���H��pH:��bpX�6����p�U���	���W��<�ZT�u��D�(!��S�,�@5YW=w��~v�cW�7�}�wm ����reڄ{�n�Iڽ8}y�����.��x�W�]��%�fi�<�^M�m��}�*�
�Q�s�"������ByD��`�ֵ�N��ϼe��>ढ़�oHn�2p0�m�S�]�e��,�����@<��t���u7���p��2��TX�mT�hp�񾳾~v��U4{�s��$^tu���'�GN���Y9L~օ����C8�k_��L�C�~-�؍��YE*������"f���l��<��-��F��էR�ٺ����d�Pw�fqm9;�H�,2���@e�əNJ k�!�"���~ĺaV�*��v`��z`�Q�*Π:�qu���x �tU��ė��t=�U�G�u"B]0+#>�ړ����u����Ʀsݺu��ӧ�����6F�Py�q����'r�y��i*���:Ӎ��`�ù��@Ipf7�=)qfi�� t"־�n�1��L���裏���m�j�L[TrV�2W�(?�?��b�m�2�2?�Z'�KvW�>�(I��U�e�9�̮�����6�N���z���U6��8Ǎ�W�f���rI>Z��ᵓ����LW�̯���u$��X� 
��Ar F�k4'�\��-��V*�t�9E)����&�s��(c�i�e�"]ܹ��:���mY�n�yk6�浖��zE�ilI���+���N�J%�"Y���^j�+���;�c�	��[�_Z�L�����(�c{�^.F���h���Y�mВ:N|�ߜ}�v�����P��%�k�w�x��b#�b���ٳ��g��rh�y��9O���'��\1�l|.F��gvG����PDnX�_|��ڍ�^��́��:*�wgR @�ý��T|6�)�ݷיWP�r��J���� �Y,�
�h &� T�4�C���U����<�<���.j`�׻��U�Nsh��#w+cD�^9�Ǎw�h�R�P� T!�vhl�H8���ˑ%�G�sT�����e4���<ir���0��+�h%�h-^-3g�>?�-w�Ꮅ_m�����ῧ*4�\�"��(��
#�`]eQ3�F�/u��n�\���>=Oˬ��h<�dg��D9���)t~��+���̨��5�S�,���@G���Vׁ��b��I�EF��=+*a���k	��'O�3�'�K�K?Flet'�?3�b6���8���"X�6�����Шv�c��QNek�	~����]�Q_�-{9��Y�>���l�B�UQ>�z������Ya��/�p��Ͳ�7����E�����zd�v�s�z���)=:y�UJ�Z��ˬ���sd8�JD7�����T�rȶ	y�ą��޳�!�~���j��n�+�ޓ9��yᰡ�[��1b�j�7ns�jnY���Z�ld@',:�-�����{���5h��n҉������:�/ߦŰN��wiv�&,Ze�
��,�
n�xV���UrW�^�,m?{�V[��Ȭ��C�&s�_��g�KJ?��wk_�����iH�X�s��nX��kU�?�����Ȭc��3�\��,*�Q��m9̱�G7��jn�;�5*]��Z���4� o�V@�T�p�5h�=}t�� ��@��٥b�h㉂�' m�T����K�>�͊T�Q>��(ɿ�g��SʐA�n�x��Xpy�����_�:�X�6��җT��^�ח�����q�t0ZVt��<�q�ɥ�-F�y�'�w�'�^Њ��F�Z�p�z(��G�V�IE�~���T<�S[2 ��
VAv�`���S�oF�l�F����E�� ��<���;22���H�9�]:j[3�� 3� Hl*������Tctx�z ��:�KgFh�ݸ4g��N�����=9�8[LW��j(�+1�=�g�l.`��x��x>N5Qb�~�a��g��_��ݝ���uj���DuVu��Ȳ�r/Z��F6��Y����{ۊ@_m�,ԡyj������W�#�u��~�ZR��z���l�V���Ư�+�g"��W�\cփ�lm�]�!
]����:g;�=X��ڸ�<#���c� ٞ�ʘR7N*.����T�J�ƽm�������h��ίε���6x��}�"��@�s"��ߨm7�X[I�i*\<�m�ㄾ��lo���7��~H��D�밈ku�b,�<��Lo޼K#;HD��w��n���g�	i1x�Es���ʕF捖#�3d[l��i����f��8]��I�M̕��82=) y."����2�mU�jq�[hQ�8YlU��F��vlcL��٦���a��`�>}v�Jl0�J��K��ަ��U��j���P_���ե+*�,V�#xB�[Oi��R7�z_Z%U����4:��p�l!��ñ��p7̊�f:Ql�k��T/	��j\����?�o��	��snK�N�޶ÇyX�<R�mi������ ��J�kB��|4?����Y�)z��2f�w�~����s���8�>w�pmQ����2ߥU���\�����6�*@~h��5	��U�Ԥ2Ț�p�N�Ӯ��ބ;�%����O�Z2ٷ��h�0��?{_;vF��7��+��oIIH��@4���w3�R����I7v��ߝi�Hg-h�#�k���ѵс�H[�����1�z{���	��e�)�t��D�J��ҫ߭P�ۦ�����{�9���쒐nwH@!9��Rr?c8�����t�p�oR>�=�o)�_Z�B��ɷ��'i~;��oȖ�O� |���rյ��ҳ߸�R"y*�mߩ,ٟ�㑘+�IT�=W/����ۏ�������RV��/�./=�e�o���9'���c �t�����X�L��5x���-I=�������~v�v��d�::]x�_����o�Q�s3���B�W�@ɢ{�y�⅕�!��PI[!F	(�]�g���Tc;J0��s.�
v��Ҧ�ꥁ6@}ϒOT�@,�2:T�*E'$���R��9.�Fr4����Lg��iS{�����Pe�n6�u������Mm���U���|��@B�]�X�rE@ ��0���2������u��-�
O�h�$)�b7�O�F�3*~����Z�x���v��1ֶ�[-�f�6�+�D���&�H	����I�iC,Bv�����ךּ�M�yO�y3�8�B��g��`wh��L�\ڂ���(���A��G���0]]L����4�xus���`��j�(��`A��S���Zu�;��(���b<>HO��>����6�Z�V��V��Y���Y��0�6��a��a=FU��9�@���%�	��`�Z�O�Gل��xܴ�Q�j��[^U��/�YXHm�2u�Х̄������$ �9��������qk����6�Qd%�ql����B��5Z�|�y�����dA~#�����A�XA��/;��Q#�~�
�������ߴ!��ć~�<������=o^�L���&�lB�� 2x{�ZӼ7Xr�
d'�S@��Y��#�u2܎������&ڃ��5��?H[�;�d���c�4�Y0f��	���6�_�x	0P�a�I�c��m�wЙ����*�J�"�|m���Y]� ���f�4<�{��(K�<����w��W�3�!M�Z^���	X;�C���R��0<���R=:I���o���b�D����~d���������?}�^�=}���߈hW�<|�0�b��?ɨ�R�^�6�NV�u��<?�� �D\|�ׯ_*�?��Y��o~�>��s=/�<g�?����W_}���se�r��wZ�EI��*�����|��>�sN��:��A:�Ƌ��*�����	I �	�w�sz9(�jg��-�@�r�,�!��z�8�Z�Evdj�!wY�X�C��)���M�[�6��g<~rnBGOrF�j����z�0���l�9�ww��G�3�=ae�uW���|�}ڝM����Գ*M�,K����>O���*,�A�KU���(o	��� ���*��C;�M:��b7�J��1���R����	#���% �,l$ �k��,�K3����2{[�y�wM��`�}~���M�ޮ�>��W�f~����F�tk��Rϝ]K�l���Ȃqdgkc��&.�W��Ҋ�5�s*,�lq����>r�N��'K0�����4��F ��p�*z]�?���`,񥅌�8�T�K�x2�D����]��-g��cq���h�
Kq�3�6���L��-������-HUorZ����$3D�^����v0�� �!����E/����0�����vt�Ic���õH?�L;,T�J\�  �z�=�}�c��z�Z0���
�g�.� ���H��#0j6X�;F]+��pC�c-	����>�����Q��Y�Ⱦ@���<�L��X��uf����,�aK �EH�q>sn,���U����l��C�����ko:�]3"�����U^� |��4�����#���>��P]��H@@�M,S�{��ʥ��������G�����p��LR��΄ar��w�g�Q���/Ŭ�2�����P�^��x7WWbx0>���LP{r� -iG�3���:����Z<1K�=��8��+Z���#�ԹoETuШ���{��>��3��\o~���������?�o��֋� ���a]��x�L���E{6�'�~��ϵ�4(�;�sY���������G{���
��r]�����xv&���--!bT�`>*�䬗w=����>Em��/������܁���3�j�vhڥ������O�~m��^���[�34? 5y��m����/f�����!B�Iq�A�6���2�Z�vm6I�!Q���ɔ�C�`dA���\9z���K��w�4��K;��ڵ{�b�ǌ���7��a#p�*.c�����4\U6�X.&�!���M�E�Lw�*��il�}x��w�V[6zw�8��\��'2P���?���,C\��]����͕Ͳ�J��B�b��+k�aN�p������ۖɼ�N�b�l!WG��ɩ2�w��Q���L��)�KQ]��	0
����ݜ��C�rT4<W�9s8?p�)?0ĳݸ�C�����ބ�q�9�l�*G��f���9�c�*HE�o�VR�r�1khkw�*�Qw����Di�@���v��[|^�zPu���9��w=�
rKR���2������sV�=�����-C,�6�1>�v�v�r`�a� ���ۧ�Z����z��h�|]V��h�0����?l�-��A
�)zrK;��E��~(~�ؑ�n%��*��~��*r��q �KQ����N��<�q0n#'`��EtA��y���	N��U�����$PU�͵*KZ��)g�"Mh��!4�q���,�
�w5��wijׇ�A_��Nt���U}5.������RO+���#)<�M}�. +TlP�J�P�F����ܸ޼���c��3�<'�m�EA)NH���̬�{~q�}�̏�}���xg?���k�c�t�ϟ>U%��������˗/uN|y�$���Ɋ��������������$5���|�$�9�,��IF����G���B�{��(m Ȃx�rT������(�AnS��k>{'��4�u��c��Š&`O�4<���*ܳĖPY�͜��������������E�MU
�v1�L�.�U#s�@���:ZՀD���|H��`��Y�8�ݖ��=�b#3�UE����k�ւ�K7�tP�`'��R�Z�Ұց֦�|�K;�fw���t~u�>{�<�o����2D�Y��%_����|�-2;	(�UK�v�(�DF}�ô?X������t����҉U�[����Z{a����� �4��k/0o����E!4mch���D�K(2N-�]YU7F�sk��V}�Gv���vtc��z6�I�U�L���`9�V]���8\7a����k���:/��*���SP>�����5�nP8|Q�"�J�0��G�d�ڙ+�b���xR�چS�h��E�u���[��m� Zcɑ��-�����Ȯ�2��������:SM�b��gj�Dm�C����?࣑�������Լ������֮%J#U�[�ؒ����J[Tèɥ@��=��UO���hT%)v�JzҾ�D(h�e^�?�TP�޾z�F�b��?A8+�=�Go:�����Q��������`�t�Ł
���R-��bH�2|��s�k��]�<��]9e��\&��\�k�:[��6���8�FO~hA��)IS�(+�<@���T��(|�ѭ��k��B��RB?�"$Y��i�g���� ,d'�}zٗ�A�b���6+�#�n���oi���8[$���}I���v��uo�^BM�� �se�	��~�.D�r���y����/��|x_{���	���NR���ߦ����?�)�����?��_�2݈n
�S>�+�P4�l�աI�b�*����=�W�DaL�{Q!gIk��oH��B�����u?>����`7!�K��_���,4�+F�,lK�����\�d��J!�򑚨`��6Kn�?C���[���������Ę������]���?�7��H&�3	��l3 3�J��NB������sD���=�f:;�-RQ{���I���0��u���SW�L��I*9�?:N��8h�����-���h&��ki;��_���*[D��/���N���:�M�:Bw�n(U��h�2�^����>>�NOO�ӓ�=��ýt�sS��f�b'��{�^-�W�d��/�ծC+!��A�|[2i���K�6�J�:>{��|�Iz��'��䇠4�앀p���+>f>g�t��;����؄+}�� ��lB\���-���GlW�&Wȁ�Y�AN�#' wR,�)�C�>#�f��r[Eu}q�I.���꨾��2��	��=�/U���}>��U"���q����nnId`3���:���˷���7���s�8fO_9�l%e���8��� �u�{�B�l������8yr�v��.sg���(=;},o]�}���-c�%tk��x98�����ϩb�=5#h�}��5��Mw�{(�
�D�I�E�}��B)�����աԆ�Grh{�Z�}�j�5�]� \?PT��0��l���4��L��'۽<b(~̇u̇��4Ѯ�1ya�s�$�䮷5R�}L[4�Y��du]�u}�d�7I�L#�RJ\�G����E|�rO�Q�_v
X�%����[B�p_�>�s��iź#�F�O�g�	��?�r^R�c�z�D�P�V�Wu�@�g��?��*P�J)�a(:wK�ym�(��뻫4���h�[�@_�xi��Ý� �$�Ǒ��k	�8�3�@�C���U?j�7�E����^��L�D{��(IGE�C�I��a7WJ4O~��t��bǛ;��wv_-���4��\��`�ݖ�:Te�g����sM�'	�'2M B=�mm��M*��iӫ^/��:��o�*���~��n��5;�,�Ck1_kS:	�[*��dh��g��`Ó�GV�X�\ �<�E|F�j�P5[�ƅh`�4��$;↡�L$�,S;��Oӕ��v���������j�n���L��i�7����\����l�8s�p����N:��Ǐ����N:��q@��� c�k{�ۛt�����n���%(k|[jW=�p)PVۮ���)���1�I0�;�'O��g���Ps\��i�{ ���vA?���$%+�s��/ׁv�G�:����o���W��u�V�����#�u��T���^ג7��c<ApbC�	���w��*hD v�Ӂeړ|�}�,�:��\y_����В*av�dA*[�Pr ��CZ�*��D��������s3z��-��I ���.sA�g0���"��T����<7��GOғ�Z��Ez��T�ڽ` H�G���Z�Q�r	@eb�U����Շ*Or����:�kϕT%loZ��(n�1�9v=�hp�K���&�=�(Ў�����.�_�B"���^ �T�����KByk	�t����	��,}Q�lW���y�\� �G�,/π]��g�U����>���٠u�����s�N�.�V������}νa�Z�<6�{���PcI|�{�gIp�1��@�~0��m�G��pV) ֮�EВ.	siڲ*S%]��e�  ���6t���X�!�
�����\Yu	��p��[�\{0(p�E�a�O�u̮�A+�Mg�X�N�+bKB-�Z��x%1� ��u���l�:d�sU�M���l��)b��Y���G�U?	z�u{�/�ޛ���i���b�7vN�������N�nbӔ.�J����R�zsM�&�[��n����@)z��ł�b����2|��}�XZW�;!T{�[��������7H9{��C�oU�R.�F%�y�����?t�h�Pˢ�̿�ʐfl|����ȃ�����Ӝs`���W>�Y��,�b>�s̴�J3n��������V�޺έ�7�5��nʴ;�]˸?�J��'O���g�����trb�ww���Y��Ƨ˔nI|��7��o��ާ��m ��ve�W��~0��?ÿta�lm��X9��^w�v+6����!-%��z�p*\��B.BϞ?Oϟ�k��LhS�?F	q��� $ ��bm��d��)2H��Yɫ�LQ6��A�E�Cm\ܕ�|��勶)UWOM��
����*�'���K�{�]�~i�KjQJV���}�'U1��Xo�æ�J��~��4�,Ɩ�e_d����ڒ�8T�8�qjZ/�
����nE�V./�ߨ��]��V%�)��GO��_|�I:==��L��S�nو�D����V�"F��>��j�N�z���B��;�X% ��)�ñ���[F���Mݼ���GV1"�����tu}&�D�a*��A����)��Y�ME�:Q��g� �'�E a�)��b�������wlc ��L�h#�d�mT��on��V4ma�%K�Ğ�u�K��̘CiD@JKHI���g�X򩃨��2�qR���B����
�0��K�4k6gȉJ,�DE��Ų�JI�*���%�:p��ܘF�J�*7�3Way~��+��{�����k��
���ƍ��ʲ�k��-uJKɫr�YвtV�s�x���(zT�	��.q�dJ���N3'>Flt,j��w�i��N���g��$m��̂�)�l+f�^���
݇-�;;�vGv��5���F�&��X@�F����L�=�$B�y%�69�i�����2�2�ʹ����˿I;���������~i��A�zѷEdpPl%�I�h{O���G���O�Ԥx�U١p�X�E �F�ߠ�����B�Ꝧ�u������,�*�o��Vsi?k�b�`�0�>z��]^�0�^�`Ti�'�*�U��cʓ�sZ�G����p"�vc��e�����1Xϵ(S� Hc��ާ�����Hc����8}��qz�ᓴ�o7}g�vwhu�!�������6]��H/�y����Ez��,]_ݥ��*ݭ <VCz��J��~lTD�a�,���=N{V��X�-4"�����o�w��"�	�aZ�;�⏂�Z��M�P���h�G��Q�<H�Y(ì@��-�ni�'W�s�t��N� ��@Σ.vz|��?R��T6�#
:h�P����P-<��@�ݿ=�'���,�f6�8Q2���
8�BX���ǳ���! h4V�n�#H'))� U3R�ן�E����s�:�#Xռ�Ls�Y�x��R���3�eqOmQ�l�v۲����v<U�ϕʉ�;߻��쀾�I���{�s��>ɲ��7Լ�n�:������)�󃎠X����߽t	YP���qO�� &��^��+����"ߏ�V%�4G {;e6.7�#iqn�Pcֆ�t�+��5�Me{�n���)f�'@�RuUd�X�i�]9-M�8���C�V�w�nOr|�J����wI쀖H-%���L�:�Jn?Q�y��*NeH���'�����T9?\3���'�'\Ԛ�w��`�Y�9-�JLpk
�6��6�� n�֚K)�5g%P-�ܪC\H]�Bҟ�FB������{��S��Q�f�+OX]RB'�6<�֪7v�V�R�j}��/Ա�-�؁?p]�(�,纂�`ܳ��wPET -�0�4�KO�D�n܇{��Q��|�n�lO��vV`0�o�e�-ڪ�z�(���I]�6:0�ҫo����L9m���b�:�E[����m�0��ߤ������f��חgi��e��hV%g���J�eɳ�. ����ٞ�}�X���Tvw��l�#)������\�I*M=  o��8�
�C��NyH.����9�m�!l����q�_�4��
%	���G���.o5��]˖ТIb�?� �m��!�gt3�;�O�;A��R�Y۵�[Bp��<���Mz�������[Kn�`�(T�2D�����q9�T(iac�ǅ�m�׷w�u�n��R4Slҫ��t}~�n���ZO��Z������9��3�������_V�ILe!����½sMy8��8���f��&Fm*)4e]�AF���;>:N?�P3P�͗�W⌓���>�̺'�L#�}�k������������Gif����&}��;mzYY������U��
�O/�}9(4�/�����R�nk������L�����j��Uֿ�"ñt�����JN�LT6`!-����[�a.��,����+o��V��3s=��m�nN�6>Y=�'��ڽ~H ��F(i�;+q�/N��(Wj�r �
�q�� A��w�	E4�ǥ��� n�����Us�Z�3-�W�Mx�+N����eWiI;���{W�xru6��!�0�D�U��1ʮ�[��tjgM@CO�ˠʥ�[��k��r���6����D�N[Y��i��P�x��{��_��?E�%�=�wh���HL���j�#/�c�;O���u!{ۨe��s��~�9��.� �E穊R8�V�	�<��N���_T��.#y�<P�5^�Q-�(�b�k��޽��[�=R������+ݖ�^�fL�#�]�V�DYE�Y�wO��W���[��Ϟ�>�����Ox�� ��Q����"�/�R��ǇGB�Z����s�� T���b���]��& ��{���+�;�.&�7E��C�C���2�^ڱ�x~�,���Q�L��흃<�'kӐ	z��΂�D���+���v�Owd�.�%|O�N��vP^۟7	ۄ�q�*�])͜<�
k{�z㾂o�j���wo�������cz��K�~�Ց^A��;�vq��� �:�Cvu|=}��*�qٵ���*P������̪��t��>��=����t���ٵ}��)����U�Ӆ��v0��ּ� L]��g5Ңn�/��'�0T<P%u47� � �Ȃ0V�|!5	{�z�B�*{r�v��
�$`O���?���G�}�6����7�_��i~�M���!�OCO������%�� �B k&g���f���/�j�z��8�;�:��[G�r�<� dV_�N���~`�����B��v���f݁bR�r�:f�{|t�����A�"[h����Ks��f�Ve�mˋ�!ߛ,���w�����R��p4�*�v�Y���P�Ď�ġ�<@��9�*~+w����$��ȓB�܀���"悅������HJd�!9TG����+G_OEXe�o��J�U�;�Uц���"�;��E˝u��0#�v��`Y�_^*P�	A�NG���4!��d��Hb2Xͥ|��:4�$d�;~B�V~]S�/A�}Ѯ>0�h"�1w�"��,ٛ�i���ѯh2�?f�J��_/ј�[IIYv�;V�-R��֓G�4Vʞkĸq˪�a��d{���<�+��P�eu�^��v�2�.��q�2�3傁����=�-T6{��9��'Y�)Λ���b�w�_?ZWM�S�0�1KfӴ��Պ���)��g��>�Ԫ�;�N[��	�X8/�Ѹn$�ѵ��ܫ'�G�RES��t���ic�מoa��qa��mZ,dT�B�G��}�Ɯl�s3w��ݾ���-�
9�Xv��hs�{;��Z�aZ���-��H�����% �A��������x7=~r�,Ck)�JN�!-�߽}�ξ�!���������j��.��o��&agW�r�؇W�� �V�7�����s ٷ�\®��H�%z o��Y�������*o*�T�v��.n���~����>88I�<Q[��7J���;���y�*]Mo�B�P��z$���U��Ъ�:d�b�EX|i�遮�^�Z���S���m�h�,-8IN18߹E%n1�J�n'�G���>d�|p��B�d'��H�
)2���Fy�o�?<8���`{W�
�5��Nn�_::U+JS(�}��ג�$�l�F�6�����!���j�g�Yv�u8���&�W�g�SNT�<ߩ�����x���Ik�c�G�� �j��C�a��u�ܶv��B���#��������~��4��YwJ] S�g�^����~/��$'%J��(C)�籬)��s͏���sDɸ��r��z��!�~큫߳R�?t�6�#��:yW�����&�qG���� m� ���=��W�z����`�͸wK�����?���)����Q����^��u��R��q�B�~kԵ{ݏ����tM:>�F<�46)(���޸D�TH�%]��{*�Q��et5K�����:��I��q)at�Zd�cB�d�?w�J{m�24?������Ǔ�%�=;����Kk[w���Xܮ+�L��;*��~�?�G]B�k ��:�9� ���B��b�3���W��Rf���?+/Z;�����$��U��2�Y�ju���!AK�9+��#����� |���A��V&%ZKO�ע���V�">�Y� �Z����$�]�8�u
�'�L�Rƿ^I��v�݇ZJ\�,�P��*lՂ&�Z�ʅ�ygϽ����ݭ�U*�n��0��K�Тc��i�݋�������^�����;{}��F{�9��`+ 	��m��h��]܄j����0�K4v?�:�Mg�Zoդ�RϦ+{�UsJ+p����j�>?}����_�FA(����G���Gi��ߥo�����oP�cJ[(x�~f���d�3`.D���iA���ޤG�,��{2�h����1efUe�Y�fsC������pC�pA�h W�^pI�$��:�YY�{�ln���"�߹��ZdsQ@�&,���LU��{w<��lx6UPֱ�)��v,�ەӕ�h�6����9��c���j��*�V��zED�K�Q#^8�;���������G�/���38w8��wG�*��2�@lvZH;�2�O�?I�N��T��4�����N-�3��.�%{����T!ݷ��,F���%�"�C�b{��@���u���ۃ#��{G����^/_�F�It�;v�f�6t��:1�o�h�YZ5���w6���3q~�B "�9����=Pթ�H�b\�����=�J}�u8c���֜dC)#ܫ#sK��	=�����x+wu�,�:��{�y	9�v�b�h��W��Y4~"JЍs��r;: >),E�W�J�s�����}��=ʙ��ߺR�N�n88��ө�:���OH�O�YV0#�c&;�S�ϕ���Y*9�&�u-!�^ �n�a[2p��;�P��C���b��|�׮�im$z�/��W�e��n���.�)����-~EJ�_xe
GhpI�Z@����tbw9ǩ�����Au�i�#�Җ+a�XƑ�7r���`o(��z���hTi�w�n�u,��� �����
w��+�j����(�UZi\na���H���4��������YN�,zӪ�_1�d�rP�!l՟�$%��W*�8��Q, ��d�8̑��(A4�+�E�l��rn?kN�|��R[s��+�������Ekc(01h"(��1��\^�H��T����Pg���.}�IK�llӖ���\�ڜ�NZ�{��x͡Y6�%��@@�t3QY���<���������}�:]�]�f�C����l���2H���U+!�5��ި'��^��7�@`v1׈}��f P�do��'���č�r�vۥ��`�l?����7_�E��Ͼ��n_�2�у#��k�YJ�� �ױ]�t�7��_�Ȓ�����Q.�]s��wD<��}�3Ƒ���`$)U��ɂ���Q<��R�؞=s�̐;�pٕ����\b�kC��֥��\آ��/�2���̡��9�Е�pXu�Qd0��uA$c�5��y���H=i��[�
u���`��Tzb��YPJ��pj���+�*��6[�M�^�XuBtw�<�|k�u߲�	��yܘE��e�ʘq�� �!��x0��Z�A��!=�ss}s�F���)I�#�������f^���#�-�ѢI�=���mV,i��
���:�C�ȓ���G����ޭ���pN�R�S��!:O�*@���g0Ҵ*��Pu�:�65�.ef7�Ugx3/7Z�p[k\Ezȕ�|��J���s!,~�R0k�4Hv�����FN�3��c�R外���^�
�{�x�=z�>y�Dr��O���:�i�5�^k�b+�.���db�0�����(�K�,z�Y}�(�$]n+��t=r����c�˘�Ȝ�1��d�:�~nk��#5+�fT#69��=WB?��2�ҁ��%y&� ���`v�fa�"�J[�"6l�"����:�Yt@�"�`Ϊ�͂�g�{��j�ivS{��q�;������ݼ_\��eIK���&F��ʀ[��B�gY`�n�Eg,}>"F��Y~�`wY81A)�q���91��v�Y\�wu�^Yƹ���eh�K���:]L�͹oҞE�=�}�<c��aPyz�@�f�w9XC��{i#'�_�&��������3�Ŭ�!��,h�*�4���&���1���+��('������Ʌe�ש�n����?	tun�py������a:����݃��*9a���|�N>�j�^\�(���6�玕%Å�j�v��6���	��~�o��_|�E������
z8�B!�QB��/-c��ߘS�_�����7�G��ѫ���+饁���zAK�B�Ly�`gOz�d�88 W ߠ��A�����1��#'�`�$#9�{c�6��20Sz�E�$ ��a ��Q��g�#o0[Y��	�ʌ�(QR�n��L)����je���F��F���5pg&]jx���=��se����2�"��M��#C"JE=t���}��V., �{T���۞%���j)��� �"���]��Bp��d}s���_�_��W��.;�D��9@�q5�l|F�B���Sy��F�zN:��٩4^΅��n^���-�C0Ȑ[��[�@�h���6�\����\�y�=;U@4/*ȏ��r#3�TP��?N�8Ȃ�w��G�̎dR��ŉ���N`���#�gW�H,���W�]�Y�]�q�C�e�í`��:��az �����j5��̮���6�P�2�c�p2w�鹂P�ш��X�W�=k�F�*},d�e���:����ή�C����-�{�ZI�ĥ�(T���un��?��@w�9�u��d{�%0���&�6����V��Tu��;c���?h=<иӮ����Ƕs�x?��ck���'��,'��sps���������(�(���J�ήn�2�3�c W󵢡Z���ڸ�U+�vᚥ=���-��ۢ�-������=P_�>\s���A�ަd��60�@��6õo&��G���=��k�A��z�3�T�����{���O-s@ǗL��+�f�&�o�� IZ�K�\]Y�l_�ʠ@\�:w�{�G������!�`T�C����J$�m�`lRO�6�M�?����K1wM��ZIͩ��cF bq���o�A:^zI0�Dṵ�3����_�_��eV��/�Od�eїS�@F�ϟ<S����Ԝ��H�kXpڶ-�(d"Z�Vr�1������JV��|@9��2���`����\�Dׁ��u����L��� 0B��L�h"�1h:K�'������ZUz���1'ȿS2�y6@��鸝
Pد��0Ӡ�cx�o�罼ް�/g��$Ve����P�q#.�<�M��`)T=�L��]�&!r��u�م\Uv���:�Rpm�;Zʙh>���
�E�\
fv]dՏ?y"L��_wFi���pz�����P��}[�t2"g����}��9��:��n旑�]f}r͒���*V�p$�T]> @bTs��"$S��n2 +�7�4�Y���g�j���������~���{y�z����V&�����؞6ݙh�M��#�ء�۾�>���Q�>�ǟY�G��:�n ����y������(1:'��=�=e�Ͷ'��/U�Ы��M���ߖ?<uY��)*�� �Q�N�	G;�o�|V�3�f�6�L5�uoV�#y=�3�;�%ߙϢ#���h[<����%.S����`+��I[�+��o7����~�4���gN��M��Ʉ-�]�WgkJo@. �y��m�2�#��f�tܒiNS=Y$�S�f�ƃqj7�D��8\'8���G�r�D��O������ˆO�D@�<�Qې��Pj��?����?6���Q�5ú�zWo�s�J��8���-��&'��ۓt{r���4
%���9�f�E��$��3�}�s��w 7􃴇&�9c@N���X��6��Ӟ�O��"=}�Lt�cʓ�4��:_N՟�4����3�f����w`�P�+R
:�BzUNi�X{�@v�|�<z����/��O�I��/��;�qݤ���HЇ�:����&}�٧�����U�?�����\� i9����� �@RP_�Ҟ����s��sk��GeS�����J�d����M��p�=�� ܨj����Q���U�ә�tc�1�v@�� w+����,]|<M_��b'[�3A @迠�C{xx G24�F������=9���ҋ��0;��R�E���x�}��R�ɢ�~�T�B����/͙}�씹o�=%g�$���=�p}��s��~������[��1z��R�
��x��22�A'v�g�������/��n1M��h[�������1h��t�߽�^U�O?�,�v�Ƈtg<��=�0	CI�Y���ن .��nׅ3��<V�u�*~d,	���;tF���δv�R!�E*nϾV@[�U�@T�8�&H,�,���0�A�с��]���{�|߲8exH�I!h�}L��8a��[{���*�����y��o�ԋi�Θ�k�	PT&�\�snA��zV�^6`O���͔��]=��3N�,9B��./��}�M��g��lӶ��_[E�qG��(�����tG��x�ۘ:�X~V�L/��H���
����ގ�,f
�q�s���߱h1��
�P8�6��w�J9^���%���*x{�S9�̽�>���Ev�W�� �-F�J�M�0�-`��bҝQ��S�����(f�Q�^��U5�Lز/����P;ˀ���ض���C�Y�^��P��͏r3��%�ҙL�����(���\-�)\O������?L��7����9��s#F�a=4�����B�W�Frp�y�J�\x��0}��ߧw/_�����{�C������f����`�}*�lc�j\�39���(���V��d�1�/�?M�|�<� �;L}?"�l��σG��N�w߽M�~�6��BQ���Ŏ��_B���`Ha�Y	�j�(��s���������e�8h� �ߗ�tJ�ܬ�eM�ѯ�RF�~x�V�7�	u�n�09�ѡ�8բ�ꊌ�t�z2w�^d�d\�F1vq��QpZ��8�e��Hy�G��}�wЙ��B�qm��v�a���FY�b���23} ci�����8�7��H��Yn��������>��g��知g�?p�}
�3�� �NP�8fڼћ�,J˂*��3S���7_�����w/_�j��w�����B˕���˟=��㥴9G`9���/m��������޾9����Ϟ���Ŝ����c��O�=M��_��n'm�� �,a߲@( a!��C��5��>v�\͎Wv�(k�Dx�H\@2dbA���:eИD��w�`�Q &�WϳDZT�A�T�6!�P�xI�E��o��>�Nﲽ3Ǜ%T3�1���~UT;�$� +��S�K�4/��t��/^�y\Ɂd���_oS���@�:�	y=��P~ݭdgݍ5�M׵;�����$"ɒ���&;hi7�K魢�vX�V����>�']f{�A��u�����9r��2@W)E�7eA�����#Ӎ����]��*?.?gg|7K��^�~6��ν�u��.���Ẏ�4��}��@��� �ٹ�&ŝ璱U ���^��&�	���W�۞E~#�o���|`/1':�k������ߛ��)�j�}Jon�RO&��eN����(G�y'$
9 ��@��̵&}N��fuo����>X�y+Y@z��dlv3�k�R�,���辄O*Csb��ߧ��^��o�.����t��+�Ɣ9g�"t�v/xE!�چ_�x7Ʀmz��K۰��)w��ݵ�~��Qڻ�>���ز���C���]\���o���,�}''���*��#`?�sCq�z��Ԑ\�	.����Q ����<�໎�n,��x�6��w}��P��	ӿ�숳E�͹��"��/�p�sdk�Oo�W4!�%��s h��䥡6��E�:��	�|Y��*��*��ld ��什�]����Z�r����������Azo����e����p�v �s8�6#"U�� �o��ݍp(̦3e�#�p(ہ:�������!��ߎv�bWs��@�j�q�ފ��1�dǰ`���:ؗ����Ǵ0G����SϜ���G�,7Ǩl%�Ѯ�@>������ڲ�����=%��ʊ���X��A�y	nj�׭>�r��A�I[3�GHl3��
y�ɬvn��Ց��k��e\���E&�	܌���y�VKw��#�SdbYW�
�2N� ,Ix})2������I��d3}�����d�,a�~<��j�e�f+3��R�?+'���u��|�L8o�Y�u��b
k�߳U8ɞ�UE{E�FD����&2a�j"�,���v�����vn==g�?e�)���(��k���<=����������Gi`�c���3)�/<}���)%�Z�����x�l�~��6��,����|>�u�]��JHTeo�_�\����|v�iL�E�}L�,�pIU���"`��9z�Zpg����F��ʹ����Y��L,SǇ�_��������QZ,no';��� զ�;ܵhg�2���1�lf�m�j�S�uEGS�b�*����;3�1�N�����d�2e[��q��pm̠�xc�fc�g�6Fo���y�0��X�8y�!��?H�ތ̻�o��������1?�{/ɿA[k�6�}K�ϭ��5��ڌs΄��p@4�轶�6t<�'�?KO��4�{|����-C�Ӧ�}y���}H_���O�����?|��/�0�#{���`�@QWޮ�!�Lrf���c���G�=w��aA�A�������͑�$����޷l�7�7��g�,����Mzp�a���ӕ��Uy��,` ���ʓ�3h�1�M��E��V�+n�/�2�ABw�� �>%��]�Ke�q2�#ڱ=Bf��w����B�N>x�������a���,�Ҝ+��0�H%)9�@�O�\�@
#�~e��7��,��N���;rm�j��fD	�_P�R*�C�.;��|���h��Uz�.y�F�kƟjG��]_	�Μ�ۗ����yz����Am��u!HR�I�T>�5��W )��B����s�`�]^��oΜ3{B� w���K���S��H�����S{&'u�j�\u�"ƋJO�6?����-�T.G�=�����Z&eE��,-og
��JW�����(q�s�(S��X퐯w@Q)uWAu���r���5�ke��w�F���]V���g��.�R&��&3��e6�����yvZ[��*�6��y_֑�>�U�l�ȩYC,���n<X�F{#�,2P�������T�o�����c����jS�����ҥ ��=��{��&���	ב���V����+�N!I%!m�n-�w���$�c��\�|L���D�����_w�#�|Ǹ�Ֆ���{��r��*��❞}G&��Joi����r�9�ۘm~��z�&�{E�Yi�*��$ݮ
�ؑ��JQ-�5?(~|���!��^C$`���t)�Z�(e��ŹJ�{v�����4[ߤj5�e��V\�-ЕeM�������ٰ��������ͫ�ތ����e�� <�To�,��8��D��$S�����Q�����/����>J�����^�`5B���im������|�Cz��1u��4��-��o̱��=�ü�hkǲ���x=I@e4wv���ޡ2��7L7�O�!���h_i�	��JB0NQRCp���؜ N�ܥ�g�����������ܞ3�bGi<Ļ+�-�WuN��2����tߜ&���i�{�ae����/,AB�"�<J�Q�����^��S��������R�̮3}Q,�>2'[y��ޣE�q���H�5Hz��k{��=��]{^0�h��L��Ҳ���D9�A79J�ߩ��$k�w^z6E�E;d�X�p��(�����*2��ߦwoމ�_�=c�i2+@gD�c2yw���p�\W���?y�>y��2�t��D"��L��2�~ y,S4}�`�W��gz�ひb�E�S�� O��nA
��֌~��J�0�������xw?=~�XY{K�Μ0*g�{�	�n�l��}�ֶ^��s�ṂSZ�k8#�˨)T�Yh��3�fˊE��j��Yz/K�4�_�S�ց�`�5P_�>=�O��I���3�3���N�������lb�H�H�=t֭ �i<��ћ�H��g��'VB {T:�L��M�fF��A�*,Q�i}�ׯ����3�*��"i{C��m0L�0J��u<HR(#��]�X5I�X� '{��� ����8��Ɓa������c_*�r?�^�'gm7[6A�g��G@$9�z�T� ������u��Ѩ���0�m2�Z|wZ~��۱y��O��?�	_��y�&�]%�s�;�v;�gp?z� q �, !A1� J(M�5���62���0;fF���=�i�D�ٹTfv��=�,f�>���Ň�Ԙ1����7� ��E���޲�w����$]]���	J�M��@[��v�/���qh�`�1���j���/��/�����Gi|o��I8_���w���"]�=M�^���ٛS��EfBy�Nxa_��q��C��i�df���!�����>�3'���f��R���<8�N�#jI���d��Q��z����g�ʈ98ȽQ���u��_�Helk�lSdP�C�YC��Q%��4�d����?=hթ��_�O���>cT}���=|�����W��,�##��6ٜ�|���\*O2����3�����%{��kʾ/%-i{���������� kȖm��	�%m��Rv�{_{Y��Ih
1p�.wIɻ��G\[�yn�:ҷ��]4�5����5eT����J���]Y��r��!��@��f����ˆ�1#N���+9�j�&6��)���T>ND0�`:JL �v��m��y�՛���`�jNT�(�3����\m�c�k��?zdϫ�X�k�g�{d.�o�ԂG���@���FT E�؊�-l�r��<��Ѿj����F2�nP32���lcT"@I�,h�YP�`](�C���֕kW+���i�r�9�s��؜�v�)���رu���-"�
��H��G èGۉ��@?����z�����܄`B�U���y�L������5΁h%T c]��ށ�s�n;����K`��ޡ�0 	}��.E����.�({�`HkM��<�xi��!i�B��z�>�Ys��&�7�?��a��wC֟<+�Řʨ˪��y`{y�~����V.��|1/A�B,?�\�Ҟer���,��1/�ke���C��B=�u��gXDLj����Ԩ�D�?q�>HJfȉHS�:�������w���O��0�ڳ<c���<���2�����\�^��7��,�e]ƨ� �w+�
������'��˿�E��/>O����TZ����#�-㞟���7'�������ߧ�녜o���j�~nO�G�L&���޸/�0���K��vB;�TF�Ӥ쿼��L��ft��0�m���S�c."�p0ZƔ,?|<Q�����F}�woߊ|��+jQh"�1�3{��B��2FU4oG:J���@��� nG{�*%b����g��w���Rs����2��A��^?R9GM���p�W*Je`���?:<�SB�=�\"F�4�,���ýc�B(���������C�XɱҧjD�����S�R,��Sgn\f����^�E�UY[-{��`�(]�5ã͜��Ѯ>���[����U�����d"�����W�o��G�X�y��F�P�{��@��E��3�d!XOw8=�*i��g�e�c�q���7|�M[�ȱt +�`KMI���ɳ���C[ӕ��6�q�	_�~�����|(�-�����b��K�O�����yn��1���W�)5��*Xk�{�U4��) n���O�.��`��
 *�#���3O��G��lJ��D���\9%c�yc���5")i�� i[�|9�Z�{��|�]Y�x^&��{�&�5��TT�v�@I[���e��.Dq��7\T!�w�	�GY��{����ܗ���%~+4� �Ψ��̾߬T-�K	�_wG�2S������1��f��ߗ����3n�y�q|Y*_�,؇���Er�A�r�� �?�wOHֻi��<N���M��I���D��N��p��-���"�
��G?�008!vw��rN�B�!?� �(#�*#U�͔��̘����^LJg�ަڌ��2O�`�Z��g����2*�_ͮ]�X��}ў��]�06�`P�5��ož��7�LF��{���{��O��_<�L}��4��_yY����,��y�����Y��1�ϧ��]X�b�6�lوx�`��Pn[/E�0��()l����H{o(4/���?�"��T!���gfP8��¨�ތI����~��B�.So�T����ZH^;�Hg��,'�9���}�7�x\yn�G��ɵ��nb�BQ�ʥzÈo|��H��uH��/�*������gi�������i��,ҫ�o���˗/�?��.-C����R�27�X�g4�u!F$������@ٚJsW��9�ɍ�@�7d�YW�ݛ�K��)�4������@c��Ӷ�~�P�(I
��(��r�C���1Y�d�N�9�z�e��}0[\z����(�g"V�r��*�[�K��)�q�L�,����A�`��`f�B �/p�=�^�g��p��fJ��d��0��c����B�۩�Sš��^����o�Np�G� ��y`�5l�\25X�����,@AT���L��z��m �ե$�xǑ�џ�]f5*�뺺#n���<g}Ĉ߃GilAc��/0���x/�AY@���B��J%��v���l۔�zD��
vr�ڻ��k���W����_9I���;�
��ĳ	��7�2n=����4�6����=PzI<�U�i�sR�F�:s»#�}im
e�U���n��6ۏ�K�	�}o�H���X�&S{z�
}W����rzݱ�I�������[�y+�� �9�{h����i�\?ϝ�-R��L��Fޜ �-=4(6}�C���O��x�v����-ǌ�1�i� v,����-�ihv�vE��Έ�S3֫t���As1s4������զ���X6�Z���p�˛˫4�����Ej�.�ʾ��ޘac���ReE@c��Xfu�N,>��Q�SU
���ϐq`9��'=$������	R��kS�3`�,����`3G69o��e�˙6,h؋w'iI���is3O�t�vʑʑ"ఏ���(�R���'BG1�
1܋��\m�F��Zu=�wf;�����aDA=E3gvoQ(],"G�d�d��[�?X��9��b��/�����E��쉭�N {VB�沨k62,�Ԇ���2����]�}��"����W��5|pd���в�&���7��7�4:��/<ϽC]?�ۼ���Ȭ�*��Md�^�?� ��������̐b
�h��LԦ��rcY(��
A	�fl�a8i��L�o2�y^�f !D�@J�h�����֣򠃒i�ڌM�c�ږ��:�i5����R� ��e�R)� ��R{n��N&�����^����F>�e_ � ^QQ�u��i�^�w��*h�ch�|�>� R�h
�+=w~ґRlQe�F��֜�R��[��m}A��1Me�`����Rlq�L��|nA��#7�5� 8ۏ������]1Epz�f�E�	=�s�����:�Z�{��]ẽk�ft��c�qIo)��i>�5�ʤ���8���ޞb"u�o��ƙ�؋Ȭ���uJ.�[٧�H�rK���W�B���Ȯh��:�P쇭���%e���;	�vo����c\��~�2�=#��[���W���(�J*�o\������1L+�l�s��6�Қ����@K ��U���3j��J\mZ;	tl���5U��|�*��K{F�0G�ts�(���q7�������)7�Ғ�s��^����$�=�#K�S��N.�zT�\��q'�6�A>��o{1u�R�l��yz�kt���#� c�:��"��f�ʅ����hpc�B��D�j�W�h��Q�����?�w�S�p�Y� S/�G��ۃ��/	�Y������ߧ3s�g���q�v��F��?8�x�� �%CS(+j{�����^����~��_#k���Jeę9Cp9[�G;H#����1�8�a�m.8]/o@���E�v�0�8�#s���ӓ��c����i:?��4��sp%4�0 2es�Hy��f���7f07�o�eK���Js������^!��7�k�b1fQ���v8+����B�P���ze��c�o���}���WZ����Wi��q��Н�\�o�	�!`M���$���[}�� �'�HI탵��&V1��|��CFx%�z�irq%�-�a5��k�N,0������ ����I ���kϨUwtmG�FV��&D;c�Si���3KE�#C����E	���hRj$���{�8i���̛�;�@�{y�T�����A��g<*P��5�C�akެ�:m�z+������Z����;ʆ]z/&b�H3�u#�[�eY�߻2�R,z��^_�	�����E�;JQlp`$9X�v{{��~��Zi*  J���%��ҏ2a��lT���2�(-�E&�*��V��C
�}�z�},�W�cTT12w����u��w=#�q�r�һ8�c,'g�9P�Ylv�~}���/�Y�+���̝��28������\/�M�$KZ��H�@�y�S��;1�5]0�~h��������l�+Wi��S;a�
�`�����5ќx�(�����jiY�w`�L�gA)����v�.H�Ђ�~^z֨]�h�%�&M��^���!�5TB�
���q�<2��b�2C�i�?O&l�@���|G� �-FA��X�3����P����kQu�n��5E��,�?*��)p���S����)OU�3|5m\3@��\]\j��/�M�ӌ$�B�V�έ]�'M^���7X:�g��"&ߌ3��������]��5w�wl\���,�E�Cѥy��L뚬#O	�2�'�~�������r��A�oN�($g��tbY�(O�������_�4D��o���DiӜ[9<�-&�"q\��:��Fpy�f�qfp�#Q }��� d�N*sJ��m��>L���U�r�f������'m���2����ؽ�ꅞ�ei�?h���9��@g�T-�Y�x�J�{n����R���cS9��:�`8��Y�a�.�\ Dq�������3��cϓ'Od`nfv��t��W�e�T�j|6W=��L;�0h�֝�TU�L�e� ���3�&�]�M���ɝV٣g;����#{�YQ�ӵ�8LՍ}qH[�H���Rg�φ�#\�NU�Z�f�(Ȭ�]JF��"H��z�	P�@in�9��;9kRѺ!%�)����}@VQ�	�c��]8ӏz���2z���ص�_��~�e��!;��m��w�ɯ�iSV ���'�j��"o��1˞�1����u ��CA.QYU���:�h/D.\a�����O:�q-=��W���*f��]���[ם]l���,<��FW���G�	�Jr�+'SaT�{���J��P��hX{�q��j��7���k-�BZ��X�-P �Vߣ���G�2��M[ �Nn�;��
���4�7҈�d�Y��3z�c�OO�ʜ�e�δ�����fKҭ�'�l�u�Ӯ�w��*�>$A�~�M�j׃��6�?�%���';���m�������զbјIÙR��7��0���m��S�rdX�攭��}.��#��E�f�0���ƃ�RP�k(�Z<��d��j�/'>��׭eXҿ�6(]�p���o�u�)SW��{P������+�]g+�`[40'SQ`���v�!��4��g��P�-(�0eYu�`GD�{�����ã���ͫ�Z��\ڈ8 �y��Mz����e���jz$�&� �wx�q\d�d�+	�\G�:�^FP^����,O�D�{'��,�q�4���V�@^�stg�v�)�;�0�]��g�K�g���2�����0S�@2�����r�����u(��ɬ�d,7�d�`�����zJ1�K(Bb �&�A��Ԛ�'ѻ� �&���W�]��=��{G�zD�����U���p��s̍_]��?��Ho�H��:,\��@ H����2�|s���sm2t?��2������\_=���<��q��@�A��>�1�l^OՄ��J=O���,�Ly,$2���9������;�^��=��юO#���̄=�x	7����P��a�1�Z�~�[g�����U��S#��c{y];0���Ν�]����kd]���펆�ݞ���ы�r�v��w7�7�9��6C�R}���	��n�
gr�E:�^!Ѽ�]��-�@=��y��1n�ݺI�0?���@>lK-�1o_�����@(��y�{*7��f�c\GZ��>�.�X*J��⬦�I���\��\2�.?�ai)�I��3f61�m_�>J?r4����������l�4��s�l��2k�7N�hWm�VcmI�ە��x&�E��E�,_ܸ�K-�ɦ2��lv13s��*\�Y�������	k1�%,O'Z�e0��϶N{0D�a�ƍxXUV+f閞�4�E�,6�GDt�E��i41ԾR�k��l#�E3�϶υ_��O0��Bt�(�ƙVF�>�[S>�(��Ԛ,��ӏM�A�`WѦ�:!:}�
z86���-�UKQq2��=0c~`��
"f�J9�i�\��$���~�i��?����>O���a��M.��lj*]^��������ߦ߿J/~x�&�˾9[Ѕi|pd���J��;)�3�������ԉD,R�Ӻ�/@��'�)�{����0���i�#��T�x������i< Xcrd��n>�}L��\��+��\�4*��s���P��U9ej�ڜ��z�^��N�Ҕ�#b��V��՗
���2�/��o�j�.�-�����"~�����2$���g�8g�)KЅ�N��-��Ǵb� ԙ���������O�9Л#�؀����Sm�!#0*��4��2I��Lԙ� �!��v���rN�Y+0#��!����웲��Ⱦe�%��P�3T�̋�v	ə���	��ҾZU*�J�t�P8[��m��CƧv>���W�8]�:>��t��K(���t����l��n��z���W���<�*5�<W^&�Ve�6� ��Tw_[�:)��r�� ���y��(���q4�M�;"J��*��Y�щ7no&�,)B�%�M�x6���6��pK]b���|�`� �2;~t�/t�g�E[���B{*��/��b��oo޹�X �`@�=�q舲=�V;���D����Yd��P��.�3_|�yz��~�rr�ޟ}P��Dan��tA�}ފ��@נ=',���rv�����ղ�)�ބwa��ۮW�5U�N�J�2�]�?���3�h���?,{�~�"Rʤ�v�*�|��(���/�CBi����O�ԽN��G�J�CE)E�JR�5y ��R�P�1��63���2��2�92��q~h���C�ܦ�Zmӑ��&�$��M�?��N^����r����7d��q9��/j�q����� d��+�NO��nz������O���O�ѳ���O���{�.� Jfrq�.ߝ��/ߦ�~�>�>I��f$'" ����Q���{idka'K��)�j�*	v��C���1��bp���g��Xמ�;����]�\`�"���n7�H>���J�����L0��[yu�j��Am�e-��;#M_y�a�.ҥE�(���Y�ZwlE�?�ܦ�16�yiT�����P:��JB��y� ������3���������/5���ǻ�'� �-�f�BOXd�mP
nBUH{�ea� 7k��1����h��R�7�6[*�彆�]��LOGB�����X�8��:�/���)_(���l,=���@�ʌ�ƒz"����y�/��'�gE9W:[��P~�7��]���}[�A� Z��ь����y�WQ�X��!�i;��=�<�l5�+JP ZAa%t9��3/].W�4��L��He$s;�y;Z�˺|1j����^����)�挅���[�gF|��Ld���x|�?�iݕ��p.���k\kl��?��V$9�7�� f��_]�l'm(����LA���A�/f��T4Zz�>g�y�Y�C��%�dբ��pCSt�U�������X��uv�&y>��JH�����!p��b��

Q��FqR��fNՖ��	P�j��F�-Q����K4f��D%��TǋW?(8���o�s6�F{�������\v��T	��Z�T5�"QJ��E I���N82��U(1�p�=ZE ��+O` ,��'ё�H����Y�0�O�S��Um_=J��К"��[u�oEõ���{d͐{� �(Ɂ�%� [��TO�@<��Yb0�� l&����!���U:���-#7*SØD_@���5��{���J�7@ۗ��	���AnX�(��#F>�2zEDd��Ҳ��Qڻw��?��~�4�8>y��O�Eu���ί&���<����޼x�^}�*�{s�&��2��I옑�3ݷM�s�Jˆ���-r��;��yZ� D��@�ͮԂ� �ء��#�-�J�u���j�Ԫ,�A����Z��6�Y]�0=}-��
;]����:m���2ɞYS���%��ɲR����刻�3�*�&��8��hD��]�,����̻�|��aG�W�}��z潭{�8K3rj��y�Re��g�`2�П8ae��8���9!�Z���
�lo|:��-; ��7�h�u�"�$�;�\����R�S�q�d25C��Z�S�5\��qv�[i�2&_e�L0��ٲ=�k�5m�<��u ���8���� � ���)��ѱ�n�����e }s�3�0����}7	Po?y�r:�TJ@��۫�P�z���D�S`���V8�NN�{d�v9�3 �x>Ig�jY�`��:(z=w���O��Q5c<�`�	2z.a����9���~P}��y��3#y���)�b����t��m�����W���� ]���S%�"�]do�nj=��\���\7�3;�<7�U�B�4W�:���V���Ν�{�s6��\��^�X���L���n�����'��t#nX��a�c-��,᪖3Mb��������9-����u�ݠǯɘ,��=�'S�:	�X���XUW��t�����^��2$��,�dS�agT��[�����pz�oɳyrĕ�r�B_B�ƀm��ڴR�
�I����͵�J%d���灢#R��� �o�n��Cx�Ʋ�����wv5bA`/2� ��N�������L�R9�""یY���ޠ��~w��$}��_�g�x�|�IJ�f���e#lZ��S�t���e����?�I�/-�`�n��fwv0���G�y�U�X�e�X\[�O�������'�o��
�>�"���HFKtG���NAV����J�@=xi� l{��z����|�|/c��qg�C ���|a9Z�b��:8d�"Qq>,:��
�Ta
�B�U���1�V�Z�c�%,���gs��Z����}`P~x�.�띦K��!�>%��3�,~����xGG{槔� �u!s��������#��fv�՛E������ջ�ރ���<�Yõ�ѩA�Ч{���e���;N�řZe�1Ⱦ6^&�wpNs6 �L�t�%�I�L�'	}�� }��iKy=���h��R��\��z�D�N�9_�! �\��u65N왰��c2��*0]�	�&�RY����N��a���v�=K.�q��7�{]����x%��1\����;<����].s�~ �� A�Kh�qd�:����ϒ��!�(CC��{B��0[q y]*k�����t�Kh�������΃��K�U4"x�kyw}� �������Tkw¼����۳^Jp�g���i֡�S.���X����y.���"�H�+G���u\˕%�=�[a�s2Џߗg�8Z��a;"sY��[�5�z������m��� ^�A �x���V�虉Of��Z	[�@=��?)�yR������p�<�w/�,�Zϝϗ��xB����0��<���#����1�ѦUͽr�-�*]�z�[E��:�d�{x;Ĕ�F��%�d�p��j]�m�ׯ���H9�/���d��Q1R���!�+2���z	u���q��Ɉ��ね7"�}�$'|���˯>M�}�,=��Y�{l�lZ��,���F,F8ߓ�ߤ�w����v(-5�Z�;i���"�4��2t߲���wvO�[]����j$qp�2�B�7�����.��T�]���]D�9@D5 H1"Wu�؛'�r61g51��j�Q�9�b;�N���3�IK���(˰� +\�4�G�ל!>�֕|���h�,��B�uO#P�L!�t�{� 1��M�L3�g���}"��]�����2$�[g��!��F���M��ץsJI�p��^[u4���񅲉�g��G�_�Wo^w�ګ}�kFL3� a�v�s1��۳ ��O�+��@�*�t��" K |r9�
@�J �0,0��<p��<�м�M��>(s����L	x0D����ܩG����R	�����«KK�L'3m��$�����k������g����$���d�z����/7���,w�������![yӁi�3aGO�I�rds.�V�Q�C�bM�ˮ�犋0��NU���K����֕�f��'?�zVA9*�}Qv�+_�iس��X;_����2}�'ټ��o����q�>���u �̫IPH���=a>G6�>wr����=�_Pf����y��yr^�����uhv���گ��RU�k~U$]M`5��e=`Y�5t:��1>h�si��ū��g�#~ZzUc7z�����ˊ��������;��ή�Z���yw�%�(���8�[7��r<�0��=��*l$�~tC��"���JdV8d�}����cgi��� ̨/��似7|W/cӋY.	) !rp����!�M9���[I������L�|Ak�`���/��U�Ui�B�gl|�u��
V/���x� ;w�ۆ���-6i�V2��c��6|�0}e��g��Ѿ��L)8�R�������ߤ������@�gN�^-���#����M߀�5'|k����k��kttgi�j�p�x	�j�R�Y�<���Ă!X�2 ���l{��R�4P+��H��L)�*�b����^~�e&���!�Pc�<ku2K�O��z��h��N���|d�l�����@�U�	��+Rr���s<�w?�{�(���O��o��C�5`� �U��܎�L��Շf�HQ��R��� �Q��	j>��:�K�	PUF�R�3�K�0�Iլ
Y�RA�h�5�30�1j��6���w����>u>pШ)���Z��������Q�k�H�a̦��h$�t�޻�Ի|�y���(_s�����~�h�N�c�L�e.�{�����A���C����C�`T�v���hI�����ha?e�`�b���Q	�^} �x?��U��
΁����S>�q��;�r�{"J�t����F�QM[h�;X��p����^��]8k�9IaI9�ه��(��x���X���@�U~oG�IAV��Vq��(g��������W�jC6������<��g00���@��f)H��Q�\FQ��j���n�B�h�Mt}�5�:''�Im��������0>����탡�-U ����C�ە��4�X@����g�$X�4�����ɥhpm�){��Ʊ���̯*��˲�ty�O����y�hfvx��,�E�H�\~�F��C���%	9��q��ʔ(�p8镥�����!4�>�x+*��LLTp��4�ۦޚdޒ�M��U:�x��u:}�F%h/����#e_�6����-�o�-ՋbQv�"�v. �;D����!ޞi��BO�=I�}�L>�����N.g:�8�^�H���k�f�ROZǻG�Ҟ9�j� -!��%���<�.��/.��ĳ6��ٚ���i��4h��h��SXj��iˑ�� ��t�G���v5��A��aF.P��=��k��p�UL|έd�2�럒�w�vm������m�a��ؒ���� @ￃ�&��㰐9p�z��R��Q0ƃ8��dxvo]�y+��A�eF+�08PȍB�v����@{3��;#��(S��MLZ�����!���T� ���;�Q(n2efU� 9i�n�c<����O~������S!_SP��4׎���*;a�93�.��-X]��h?Fx��B���n���v+�Wn�Ǉ�.�`�n�L
���#(�@�g�Rld1S.f'��֩;���@D��e�۪ߕ��&u�~$gb�{�2�<�|������U=L�}/Se�S�e6q$�o<�,k���b٬��5���i�W�}�.2`ߴr�ō6�yz��2�rt<�^�x��ظj�� �ϳ�#^�����U�ApL���y>��b.��޹��Gz�j̥���ĝ�>�����Yy�m#u��%��0p�`�������t�UP�EF-��;y�H��*������:�҅0��I��Lv6�
!�yd6������z�_k���V�#�97M���:a��**�uu�]Sf��l�D!B�I@z�������'v�d'l���o���(�G,�f�H��G{�K6%>X�,�^^(�B<���=S'��4�Yo�d좘��c�X_�`�7��"m��|��5/5��D+i��6ҍ��nl#�  �Bgu�P��t�N/.���uIy�������N732�n 5���} 6&M�ADv׮}w�W�cB����̎"�0��A�~��+�9���X&��z̛�ע7�Lw��͐\�}�	�V��%t('{}ט]���
2���DP��Y�I�=S�h�twd�o\�������n����k�E�����,�J8�u�*���3N��	p���4n\�P��r��?fDw�U���O�sL>>��,!��<zO�t�Y*���<|�0��?�O!|��Yb�������e��}@���;"6����v��w�bTnѹ�ep���-wr�Yޓ�a��c���g����i��VxcY±���ɧO;���`�`4Dah��qµv���I�ý�Yi�(�T�2�W����@�^��-�Z%�M̀p�E|>�A�?@>�f2wF=�r\ �/!W�)C��MV%	8�Ֆ�R�7$1�˾���J�� �No4#�,���ѝ%��<�����[�k��)�rL+��.�~��3x��g�0��
�����ێ�t@:{���\f��3~�s^��s����m(ze��~82��2�(@0��)��:�r��Z��\�ЇnCब���c���f�7HE� ����8�h��hd����tC���P��Ɯ�՞�h�s[�e#@���_xk��4l"��@���A��j'n"x�_��E�*�m;�y��RcM����k�ef+b��(���	�Y
��B4M+$���P��cT{ �A��+	W�����$���2��2��>���<�E�X��>���C8���e%��G�Fh���\Ra�����O�d�\�VT�����Zgi�t]�y�I{�9-���Y�x�>M/�EWx��Q:��O�<��2���2�k�.�:  �0|U�?���W沄����<4-w�^D�of���:a2Գ��A֮g��l:�dg� �ӹ6�ph���q�H���6�Ԃ�+s���uz;���0�A	��Y�~(��K�����Y�>['��$UZws���F��e�9��R��ZF�7�Xf�"RTi����#uQչwXJ��ޯS���pu�B��)�=�Q.]�2kP�񴂧��s
��,����ZQs�%ߢ�P2��֨)?~�$����>��3�G4�% q�����F�GU�T��۾��������Hu'{Ɇc13�8F���'�{.�������sp�����`�X ���;R]���qL���q@���cl��O�A=E���l�r�P��8�޾Q�HAX��1^�"H�,9
Z��Hhv[�jWw�B;Gg1�5�T� �f��҈�w��z�Uٕl�O_�8�ܣ��lЕ�y6[!`�p�,*��b*LK|�f�$�^�5�����rr>�*8�W�g��	�A��c�3�
�nɮRY{�t6�w��GjҀ��v��"?O6n[�NF
�Z�pO���l���u���	�M?�]�������L�2e��g�H�I��P�WuZ'�*��Rxߜr8�`����c|�1�=�����3am�iM����xy?��i�.�1c  /����'����/M� E����C<#�Գ������u�O�q�`�;*�����V�A#��a�ߗ���p�:�'7V�Z�a{�?,0�S��<_5��.�Q\�CD���Z����!����ǏB�7v��@��A���8�|�T`=����y~~iQ�sH�阡,8�k�-\]���F�[z����ϐ��Jejܜ#`����˾#W1{鈾T
�|�F|!>�R$0_��wAvi��3�����2���D��̗j$��J��POk`�����txx��X$ψ���m:��x����%"�RbV[����8�	�X2���C�(/��ZǘH�������y�q�MR;u%�Fi���V_�p�Q�N����:j7�����(φ�P�rG�)Tى�є���^j��a�(�����xS���PJ*E>P���T*��i�/���쓧)S
�SW�2Y@7ZEyu�z����d$j��~8a���Ȁ�l�t3�@<�G#/����;̜b�G�b*?)�|5�t0I�����/�� �:~��Ș�>CYC[�tlD�,o��^}A�R�Ʌ�m"k�8�Z���H��W�3W���F\�K�M�_�
!U���>�[Z11�%S$ 4D�R`���9ud�ͦjM
�4�2����n�^o&W�rD{��i�ZU�J .�l8$�ـ	��Oa�W�Z��dv&R��BPi��9�_~�<rU<�[���A�F>~�vec�`��I�Q�}R$�+r0G��2�og��X(l9��:��x��_�QA�^�8�q��.���^���.��j�֓�����?svc]9k�����絁��ŝ\y;嵑���%���t�>�-�I^��V1�B�Ku��g|JB��7W&<w����W���j�52m��Ğ?v����]�J��*�x-��}l\��,��r�Vǝ��{�#��V���p M2p����z�7�?�������R��m*��.^}�#޻�Jd�`��l��4��lrJ�G�e�vvFi�;J���~�r��ܒ��5S� ��!�`n�'7�6PbV#1����#��=������k�W>�t~�rH{d}����Xգ���н��ފ�S���X�(Go,���{�#d�@+6�8��eTf�����o�Y�(���@�xzj�{���;����y�<[��<�]���R�*h�����;\�rhN�^�c��~vNP�V�l� �y�R�W)s�آ�E����+�Yu#4��^�,��B4�=i9��9��,�t���.E��"���KvϣRnh�vY=e���Բ�K�*��)K��l3�h'd򈎰a2Qf���Ud��)��n��6��W.�i�������G�J�1ّ�z���D�v����e3j'9�ǫ�t��Z�6��<�2li�6M���Ĩ �x��2�S�W�pE�f+^½�a�Ħ��!R���wo#�o��2p��՚�n�K��D�� �m=���#/:�f1�c��#6��+�l�ό^�@kG)~�e��;:8@Hyi�B��>:׋{R���k�ɫ���r�,�,���]-�E�쐰"� klr6��Q@�cj"��g.����>�$c`,\d��V����F/����ҵ���I=B��G�dA���s?҆^0�,���ޗ��2���(=g�x޳��xY�V�$\P����u7�-�G��={!���_�2Y��j֖��rKaنC��6�+ <�K_�t4t~f��x�l?lyGfg��"���&겛X��X�'	Һ�{NA4RfF���Q{�tv3����f��A����գ����oz�����ԟ��Ԗ��G�����f�ΑEk�^��2���BFjH2Df,Q�!�{)�,?��tog7�ȏ�z��l���qp��(G�@���
�|xp��-�E�'�YcT���z��*�eQJ�� �z�{	_/90ԭ���� 6*UZ�V�l�nў�2T�@#�#^�C�%�E���
�cv�����o-��[	34B��U�F^nf-Kw���mZ'&mc��rٸ�HU�]�2פ�(�S��F���B7�+s�#'�"�D�ʄ��J��QxD�)E7^�7j/�fi�쾉�p��H@U	B
��c�����G��)�Z�}�z�a���A>H޿�@B=������1�� m�Jd�J]d�p�6Q��r����	����3���� ��x��lN?s[��Ξ:��K�:�������D9��+��s�6v�7(;�fg;�����G#����\�"��(�z��%h�þ������ڱH��<��"#n�Z1�7ٰ�����f�8@\Rx��b� 1�����T>��0��x���mctD=�;�f<��͖$F��2/t��{ 7e�w�Ÿ́<WJȦ3�Z=��P�{�^u{_��t쁏[��_��%���N�w��" I�������[ttqn��[�d�8Z2S�$>1 ̇���c+n,����MG��j���({�+�`��3��]GU��	!Eh��~��g.�:�A�z��y���c�^��U��{��B�BF�ti|�����;ͺ�WGak#��Im���R�s;-�J�K8�W����\��˦��%*{eh	t#�Ag|�.��뱵gs��g{��w�u��/�����ӟ��.�vi�1�;�Ŷb�� ���M-e�6��(Q�X�#<������w�P�UGI`�����C���ig��&��鶲M<�Ų���4&sC0a�0��˴��(�v���T�M;����qk�yc�Ԝ�z�v��0Fep��񆈑�ٺ~�z�����9���7�W�<�م���2��RgW*Gs;���?�J�Nӹ�[s��~�<�=w?�ے�Ty�����%ן�(P�-�&��)P����x��|����,�m*���dw�"�24sW*�:n����!�2�k� ��FV�@��V8ϰ�h
W�!���?ġo�(?��lX�������8ۖ�j'����7	8Ѝ��x�J��K�aL�0J�ާ��"�f�]�x��?;��g��J�nJB�o��+�	�gcΫ�'GyN���ֱx	2��"�n�'�� �6�M,�����j���BC��̟���<^Aٶp$.��z^!�ː��[����~�z� 1%��h���}lA.�{5�����lz-�aF���d��\�+Q�G��I
&�/0I�ie�j���3�fnt�e��y޴}�ʵ#�W��@4����N�N�����4�:Zg�s�;1���B	��V�k�Guyѳ�����97pk�j��|.le>�s�Ǣ
��2��Yk�a���<�/���,z�k�
N�)�D���-^<��a�}6����z�<����r�&�^���z��_w�#��v���H�9V��n���X
r�]�!s��_��_|�E�m�ϗ���Q	LE�8s��ɂ���e�Z��ǻb���"X�K}��ߥ����r�V!����Znu�	����,V�d0�ۯ���4s˄/,���9������S��Ov¿O���Ŀh��M]�S�(�J���o�7K�4��nӎ�+�(Q|�^�| �2g�!h[�����=�]
��J��EZ�{���i�����q/�������Ã�C�0r����h�Mcƶ0�:[vQ��L�P�a]G�|q�V>�!V���]f��%� +���{;��A�C�'�f���۳�tv}��' ���7e� J���^�m��T�I��Nb�)��D��kT�	}�b��t��;	3��g/lzG�{�VEiX�՘�TϪ͚��4��{�!��3b�U�iØdV-�����a(�+0״y�i��P���2�o.��?/�r��:YY�w�1��������%C�󬐠i#w�q���ro2Ӧj����L� wؕ�(��w<��'^����J/8���s���G�R�jU���TI
�y�����׻Q	!F�l���8�ֶٲ.��� ��11��6;u"���N̑��A��W��B�SLzrb����,j윏ځP�^h���" @�Ĝ�es��F����y��u<�< ����K�Aڼ*�S{�8�,vm�%������&�WULX�(M§�����@��6<8-"ku�V�΢�QL'����=�x�!*θ���	p�>��Yf=���y�F>�����s��ΫWoӕUױ�d�v/f���n^�2��ZP.��[�9
�zgvs�&3$VT%�K�Jh�����c#k3AI�m�^e��VF���e�k�71���\si�����&z/�}�Qmbn�(疽���ZVV.�3��5�u��/���o99�vM�V���>���w�s��q��������?��#�~�����/֖�4d�Uꉅh�|&�s0���`�I��a�v�V����a@��h�ym�Tn�i�8�W�\��tb9|p�z��{i=�.�����.)���ў�8
���و�R$}s뜣gW.� �m�.�T���x$r�|S��B橧�	�t�[�9f'j�3�n���2`"����<���;;K��^�ȑaH ��NT���Q�1���B�%R� �P�{H�|6ZM�%�Ȇ�T�������TWڋr�z=u�o镶�J�T�RuN)Y#�3ҹ���w�X_(�%�T�Y�xS�<qxWʎ3�L6�?�Ӄl��O�uB@d�!d ��J��z5s#P��)���fhI����P����{�N�������K��� ���{�e�}��q�޹3CEZ�-�T2;h��n�6E5r Ԝ�� I�Eп�?<F_i���� ��GQWpK��-�Vb�Ҙ���	��R(ˢ(����ܹ���g��}���>whɑhy������{�>��g�������$�ny�(>a6�G!�$dT#��f~ܴ��[<t���d��9��&�E�	�`8�����h;|^�w�H�uI�R�t���|���0窹䀈��O�����'Η�h�J&A斯!��>]o����{JO�^�'w�s��dol�� ��D,�ᇤw��e�H΅�B�Q�L�*Fǈ�ҨPU������5�P�/���ϣ��mS�,�ɽE,��t�5�i�I����C瞏D�ȇ��p%J`����܉wC:=�{a�1�wS��)�MQ�9wߧ}�|���i����E7�k���wm�C^�ͷ � @���Qr�BD�Gwܩ����v����,��{�����Z°���H��SL��WK��~�n���('�س�uSpy�zqL���SG�.X|SȲ�o)L3a?,\]���V���,n<��oo+M��hCu:�l:t�A�)hw��c=H�
ׯ<G�ܩ�'?��[�Z�&zenbw��t�C���kDċ�{�^0�se�Nh�{� ��r����N�QѺ:��(���#��k_ǧ�x �<��U"ｐ����M"O�����ˠ�t>�"�����Q�E
dѬٮ說�*�-��iN�~z��b� ���I9&��j1H/c )� ��>����¶�A�O��n��*�nD�)���'_Nk��PS�yOn�R�KW�_��Zgw86�T"�䞋��P������W1��"uY��(&�[r'���z\�D�`8�ijκ�]t<��p���'b��"GӐ�Tr���8�Ni0K�߃�'��;^E��ls(�W�������%g���k7�x�lٱ���j��t��Y�D���p�����(l�#��D6P��4jO j��|Șa��I?w6��ߑ<��ufk��ҍ{�ɇݥ���9+eq���: m��V��Փ��7e!Z�Q��m���~��o谥��V@0��@���dG"a̩6��ݺ�kq&9`}�|�=��*�soE����<6�v�>O2����l\�j��G�]jCt�T{JM��~l��W���,�\��XV2�0H���}7��L������1P�nk�cc�5(Ņ�[7�gR��5<v�Bv��]߿Z����]��>�Qh�^iK�sj���������@yʅ�p���NZ��������jA��1�*���Y�bA�I[�O�*G6ۊJz��U3�ۍYM���~��^ʷl��x[$L&�y�G� "9��̡Nًn"�����Q�^N�b��!&D�����CD�h
gV4`�]v�Z���j!�(RFg$�ק+13GE��x�jŪ4�塸�����#�7�o��8�s�m��4��� 7�Z��l1��D6F�6-�,A�w�!m�3�7�I#���:���������1�O����p5�
�>��u�#B}p��["�.�(��bc�-x1�!��i��gUe|�(��dWJnVB�j�C!��1qr�T(~_Hw:20Y�LgT�a�k�(����{{"Bz�~&A�"E��E�:����$��v�he�����(���ύN��v��T<5��7�]ٽ�[v/:�`��}�vH��bN��9�G*� ��G>F}�����\�S~[�N�wy����	�.�/\.l�<]_}nO5`&�K)>Ά���_��DVaZ!��m��lJ립���"iNUr'^��5/&� �sx��3( �L���ӡ$ú�W�5�/[�at����07:��l�c9Aǿ�eE߄��FzT���o�^ǿ
�H���ӡn]��rV��t���Q��D��C�͍�i�"����@|����14����h<HmEA4;��}�3��ʛ�P�/�_���pMzYӽG��1�B��1�s�<*91CTO�5=������(~t��H�*dJp��uއ�W{	��oQ��213G��}���Z�.�w|r��ޘ_���j��;�.|��!��)�>��_���v�M�uS9�0��
t�~5[��+|StvCOԜ�?;<4wNO��.�7n���#�b\��HX�S,R;�z�"ʄ��aԽh�8��c�~͡/���"z��|���4�oD/-w�Ņ�uD����+�qb�F�74��F����X�)m3����~8�����D�~玸}tħJ�ͧ�2�06�)E�8�!=�Z����{ts��Ɔ�3j�!�[o;��^��o1~��84]���ke�==��3��Zo��(�Vn�PaT 6��U0fg�XO��Z�*F;EL�%�'�;}MRɱ^(bt�hva˼(���Qh�g?a46�Z�ϨB��0dxq'A�P���mA�.50�t�<wbN�c�}L�Aae���Ĥ�A�H&5шDԩz�
�N��@j)beq�Cl���Rި%�����6��nX�<m��|��;޷Ή�P���E8D�Ʌ�oA�@oYy���Q��RF��)���BNb�`�(�u�eh2I�O��rEb{Qz������CtSء~/�=g|�����e~.�(��m�XN34:mk�X|D��Y	��h��z��(U�j�u��u�#$IE�Y|P3� E�#5E�9���QD%H���i�!f�Y�%@
��fH�n�.���!�|��U"�W:�]�hҿ⬾J����<H�$�[k�ނ��N�8{[���鹤���0��"�|�ѯ�N&���PTK�{7�5g(�^q%-�C��y���M��&ȍ^��z����X�>ۛ�_���to�@��:t��|����6�l&�Ch����"(:�TJ*��4�tߝuZ�b�����Si������GM��f�ҕ��w̪��W�'_x�#����>���:�R��6����#�oi�&�����E´5��i�L��4��V�s�q@rE/��Ն�Q�{Hc��i�}���*���9�Qv�>Hq��f���F�-��":�/�f�2}M+fHMC"��'�+���v���z��x��e���Lƍ�<;e�5��	cd)��K�������G��+Wy�*Y{5���+�����	��@�k�������)��R1�Vr�$XD�+�o�f����7}�l	pU��1^|C�#+�;QC$4�D"1��9�8�BZM&�Z�b ��M���,cm9j�o��X�Io���������=)�1
��-	�t����CLz�!'��pJ�
1||H�����8�^Vq9Dܚ��9~�L��1"��e�7d�ˠ�-�9EHuƚ�1%*8m��^��"V8.v��p���c��H����P6����mD�ΕJ -����zч�Q��`O`��ްʺ�V:ۇ�Ql�8���UaA�)��Ί�2�E�L�b������{�L(�Ъ-�����-~=�
�A��Z#��8Ս⨙wAX���6C8$�kp>Ӂ���!(D�\pa���#��r�n���a�O2�*�w^�e}�b���>�!�D�C��KD�Aڶ3�̚�"�c��[�0�tJ�^���rRx?�Eq�������9Ş���ډ7��ޢ��=��G���y=��C�E�rʚ����r�����4�}���Szɩ���P��ͥ=-
?CW��n������vՍ\�����t��E߫UUQ�,��dR��U���e�����/��x=*�s6[)Xt�#;�{���e�������}�[>�x��E��"aڂ�4�+>z1�|��zS2�B�( �!���ێ��lt�*m�nH���~�ĄjDˁqZ�Y����^�s�A\��b�o�����B~���k���\\���`Vs��u�v~� @J�@=�c5�Wf�+���ࠞ��q/N֜��2�����ڄ�\	[<nZ� B6��0��zKr�s�qHu���������|B�*Jq��R�"�r�b��C��v��1	�p�Ӌ�G�Ǹ�D�:�M
�% �;�f�iȉ�J�q��w��0��̈BU��K�A!�e71h�o���"_74�p#N<�n-Hy�[�t����u��M��n�mB-6>O,���HRTzߨ��vS��f���ﱐH��XpDE�x/�z����2=�9�R��O's����d����
�����*�IY8o�_�=e��gS�.{Z��@
mo��6�?sK�l!��A/m�+m`�I�qG_�q�p2�J�ɘ����"��fu�l�3���ֻR���3�?^8��������ɂػ�3�g��P���G��O�@��w�S�������y����~�u�"�S��''G'2� {"������7{3n�d��8�;z��Pj��8]��.�����q<��ӈA�s�=оI���`��c���1ESת.K�Z�%ݯu�ԡ�?5���h��Vl��֗^SU���rM���M&�~�����+&�ݻ�,�������۴�5��8�v�\j���QML�L�lo�o��窼sy6?-M��}��0/	u.�cuN7,��x�!���L߇S���Pb������E����4�ឈ#B�&G����ҍ�4�����3N[|�r�w��%�N�b��郛���ꇛ#uP��M/X����)��3ނ���\��,-�+�ר��Aa���6�/t�,9�wQU�Eq��T�G ΋)���4~�U?ՉBgo�%�)��a�pR�u�[��ЌU�>� �tf��"�Y�9�P�
c)��:����i��$e��#FQ6R�"�CA����mrº�M�L�?X EEq>]��[�.�1�s)��{�1��<��*�|9Ԡ+���8#����n"Ig���h����G�\ߵ�"�v�X��mmk:��=�od�,
r��L����O?�"�G��c�úveU�B+[U5$Zеb%x��5��c�tT��W�v{�t	y�Bc��K'�Մ�'��o�`:cL��o�X�&�S�nWM�6gD�m]k�-�ɦ<�J:Ѫ��k���^��:+7R;S9�u}okJ�t�v��xL��>�~��o�J"�l6v)eמ�uto��f��.���J��A��ӗfs���̊aD�H�x��ᑻ��n�l}�]���j=���f���V�-v���z1]�(B�cE��K�埣`�E��-z��=�>')rܛ������
Ob$�d'��GDf�|�~��^���EnD�ߒla�/����>���#?r���t;�E:�q4�m^���&�����Y�����o�W��t^�U�+�) �mb/t�yt�,d]O����[�Y�N��"�=��];���Cg��r:+�Q��"A]"ކQ�7T�s��n�9w҆)��A�*<�Ȳ��v��&� B�a�	�0#�� ?m��_���GP �K
ft7�VAH�)T*N����3	#\�\���%�Hpi��D�g�U���Ë�T�pכ�;+머.�t��7�����aJp�f6��A$���Pq��ڜ9GС1)��LN�Z'm^�(!�P��@��B�4 �5�Lp�4Wj��)��Jn�)�^3ꋸ�,(9�(���d��RǦ��>[N�f �����?���P�Ed4 �~�x��+@7�������8G��{�{-}L�v���H��'����i�S(�j�e�jM�۾����7����p��SZ:�w����t�:��>]~me6gm��X�.аT!���J~X�zZ���RGσ�C���Dj��shS�Vw~�i�qS���1�Nz�P���<�_��ž+�S_��ݹ�'��b!���w��6	`$�~�~h�Y.�o��?X7˲��ǚn�:�De��-��׋3q|t¯Ϡ��
n����=�c.vq�ɵ
�]NC��-����W��>�6�smݞݼy�Iꆸ���s�?J��;��������ihY;g��c��T�y��"˷����x��_���]ۭ���^�`�Ilց��h*�CC��{l���,��9���t�5�c&��D���=d����	_z�=��������ͦ{=�U�$-l���b�qv��5kDr�I�\��b��iJ���І�m�`�r|�Q�.~1KN�h������8 f͞�>������_Q�=ԣP�`M�.y���;w�/����$�
���k��zC7�z����2�lW"8��f
!����j:�Q���a`�)�s]ͣ�F_�!q˧K�/S���[���:���Ns����]�:3����	�����v~C|�ژ��ўk�ߢ�\�Z�t6�����G/��+�9UP7dB�{�,��z:q!2��SD�"4ZK��`1�5�u�'%Nݕ���v�^���~m�혅�n����t�Ƙ~��x �uXӹM�����Җ�ѷ���龀c3��Im�(�3�u����XWYZ�˶���"�j2�˥{eo�_���b�7
|�����'�3�k;� �E�/��(�����O�x�{��Vz=\�������fM��p����7,�+{�[��l�W� ��� ��W������+�ݛDT��5�f[�߸���ܜ_��{�~�k�R{���7� �� ��u �����}�����H�ƍ�g�Y���B���-��.M�!�a�C�.�{���k��!d��&(R � ��u.����M;2+��m���'�w��g?Aw�"����nz���B��u��� �f�cD%��bghJS��p(���lp�I��(��@�0|�Ά#A:a��ŻBj�7�^E��(v6��=1C�t�]�s�2���d&���>�������K���V��Z�2"[UO��C�O_߯i���*�� �{uIUb�^���8)�h���!��H�S���4��n�\��:�4��S����W,�Aux�������)G�q[�-_i����_k̦�W&���t:���8x2�W@b��;��'ĨsA?���ͺ9^o�;ĝw�oj�Lr�"7�Dn�g�zZ���(�,z](ԛ֥�k"H#i��􅑴����!,��-ץߛͤ���@���J+Tׅ����(�{g���[�1޹�>��M7���>�'�����Ki�SP,��������'�Ղm��ߨ��X�a�̯:��S��%cj#Qܬ����4��71aӵ_����6E����0D��|��;���ފU��j��6���ȶ�'�x�?��x7�M�Ⱦ�g�l8�����Xv���}d�w�ǲPZk���֣7��d~{~��}����O?�����
��k���(��F'�+һ+��t|���s���p
��Y�����jV���uHf{;@�����]Y�1$}ʴZQ�Uy>�J4n�Mgl�i���۴�({�^���l�S����|�=ХE;���Fe�Y�	��<��%7}��kq�\���rmWDMt\������EQ�.�������ʕr���\ �S��Έ�ά�Z�m��:2���=fʋ�Ġ9E`ҕ�+�i��_ӣ"�\"e�XxD����MGD�ߨk�am[����E��|������XX���x�i��;��[������n|i�Yܣ����<*��S�����1E�k��>��xSd�	EӶ't�kR9+� 6ɀn�i���	���ԥ��V&���:��u�W��ț�
�o��Ț���G@�{�k���m��D�������{����ݐ�(�`�h1z*��Ѫk�	z�K�qND�F�bD�P#fGЬַ��'�V��PKc��#t)%�0��m2	�Q��'���a�|�Ƨ?]�_{��z?�7���Z����F�vϮi7�8L����<6bC/��E���>���8���X����}��eE�ra��(� mJ!��rSn6�m�6��Qz��I��%�K<GW�ܥ�j�h.X#�e�D��,�����x�>���Ѣ�nyU�B��[�k��rq�����g����x�7����F��3Hcŷ��u>v��}�N�7�{F���}_���?�s^��ԗ���j��5�$��Y%�?~����ϧ�ɤ�R׵����\�����˴�?�� ��%�*���h�A��[��7�M�zQ}�_�6ә�-�����}�yR��(���@�H@E��Ƨ9k��I��o�)���w˱����t��f���-�0KI%�? D+\ﴙ).8�H$|Q;��x0p����'����o���g�UZ	[�������Mi!��뎎Oo/��/�����j�ot�~�[}�n�g�~��@gFF��It�sfc{.W��6Ϭc��q4�]]	��W����BUZ��E�.��U��	��]�"Z]aޕ"�/�V뛛��T�/���^���_�6_�e�{
�[�n7�:����8fVW5-AM	:�I�@ktFı�s�g�(�q�;0�{pg>-Z�}���|�2"a��Iܯ<��j_a�Fϴ�ؾ��qПT|G_����M��|�������Z���,^���nu���֛w���ѽ���-c�_��߽'ަJKFF�T-��l����r�dm&/X���VE�5��ѬǶ�~�H�{ꪺF�C�����✊R��us�i7�t�^��vS������V|h���Y�6�Cf���8��͕~��Lʒ	�=��|S?��4C}�	�Vid"<M+�ܻ��m�x���o���/�=f����l�'bZ�c֪�(Jݶ�;Z|�c���K��m�X�5W��N��%
�o�h|���W��=�қG'�_������o԰�����R�Gcd5�S,_�W,F�G�TY/i�֛�[ߣ�zќ�Y}��o�VM�����kEW�u�#������v�y��������7�~+k����U�Z4��m�Y1�U!zY�Sq�����zR��}?�ZS���EA���_�����e�b'�0-���nܸ�����Y����z�u��e�@	a�N!thq��M������{����GO���D'���^]�����Wˣ{w�f��7#c<(t���Gz�N� �"�v8�t+4�h�<q���Q��O?�ϖ''wh���������B�"�S����D���_����Y��/�l��d��� +F�S}3����]�*�Q#����.
4��u�\  $#IDAT�+�q]��~�g#�O�q�����&��q�����}��E�yŅ��������x�;����2)���z1�Ȱ4$�$L��օ��1�{�9��)>��@J��_�X�M�T���a���o�t:��:I ��(��*{t���ES4��H�p�K��m�eo�0�A�N���w!H8=Yu\���UJ��C@@@rIa��\���YBJ���k%w�ZJX@����NiPx������|���9gΙ��y�Kh�e��JeF����m�Vi,(:M���n�ﰴ�#C~Z⯩�l��%���6:9��Y�°NC ���J�pJ���7� <�Qɰ�����8{ƭ�ZČl�[.�O�_����u�!mN8pNrE_�Rpƾ�%wpZ^J�]��p��o>,��q��OR5|��L��X�In���g���
Y�C�g��Y$<�'m1=4�����U��s�3���*�eɌ����}6wf�d�0|?#Xҙ��ܮ�Ga[r�D?�.h���z�Uȋ��aV_�`�%�I��;����hy����ټ5�$2�̂x�a��_��3�S�=�,gOnv������������!�{���J�=�;�Xҿ� î�}T]Zd�TWj������.��|Cl�"|*����x�	������S8���*%�m�RjƎy-�������Ə$�
{�q�wVؖ�����-�p[ ���<�ӆlS�%��nk"*��$�Y"9 ?��V����d'{�(f�<�{߱�g/��%6}ElA֦ǺR&*��
��פ�Q�e�,n�dV��M�10"������J);���;���x����ѿ���,"��.�S�i r�>%�Rw���x��Jt�:��Pa}?U+p�j�Ç֭��<�!�>	�.�4<;����\��b�=l�(�iP��U���|����b��֢�%�/O�5���_W�7W'z,Fjl4��{V��k8<��.�ɣ4*b Z���ɷ"��
E�^�$}�������ۧ���q����O1_�g�d���=�	v�c�8�N��`��e���6�O�@���V��(Iz.�wӚ��Z	��|,�҃��я�[�߬|�P}J/��3�j�d2M�z:��H�8�W
W�h���O��%�>�e�w����>ȡ}�=�ԵI*mP�������`o/�$����N6��ߺ_�x�P�W����"e�=dC9E�@�*�8Z�f����i�? h������M�����A�Sm�����qSݨ�&�jy�]14��1�t��]�*G)T���io�^���o����f��3"E�:�k-t*Ⱥ�� ��5j�!�g^i�ʡ�֚f�y/�Z~5�"��λg�#?����x� ���~E��<��RZO�g��r�<�����S�X�r�d���8��G>^��͛�CL��"!5?���ed��d�l���f&����t[��C������w
$�)�1S?�CG�X��Z}�^�0$���6�}$���[���Է׳��Ș�X��'�hm��Փ~v/[�ɚT�����f���C�+�L�_U<;��BR'�R?��52�p�^��d��IdCz�ͻ����!���Qi�L�A|���"T�X���a3M�&�'��X��>^� ���>
��#ɪ�[�Ȃ�_a�.�W�9��[-5�ɮ@B'7����xe�ro�.3_ i��ܔsX�z�D&{@M���$�j��8�ش�1�M	>�c���1Z4j�|��5��0n��cUI�6���k䮽��!�7�#�7�!��+�N��\G]3�]����U=O�wǎ�.h0uYo"m� ~BC�5*�"h���-1�[6�\N5�k";#��M�����eUώ-�\="��B��%�j�U�Uf�% GN77D�	ih��>�d�A{��j2�i=�X�y��!���k��_z� _����'�l�*�\Z���CX��<���}���2A�a&�l`�2�������{��p2�V�Ϊ i4�B%â��8qI/N��_K��(��D$1[�}G�uon^�k|��6;ʱ�%��/�|�-;�Pq���	�<"ΪF*wy�Y�*@G�?"u��B
��6�Y(&J�J~��_�(k^�7�D�0*/Z1ȢQ]��n�5���~���9�FB��T�k�X,�/+J.�����[ ��n�9&t_:���Ïa�i���g�5Q�0ߎM!�wߐ�\���B���/�]��/p�B�>�P|Oz�?����/����i�N�� ���We7#i�g�xR��h��>nȱ��k�<ΐ��㋐�2��0M�W&������q3�;Z�����h1�d³a�
-<Ղ萬�QۺݾVￌ.��e�-��>��|��1n���w�w�V�������7
U4�Ll��w��M�Y,?S�l�6����P���[�&.�]%��u\$�A��=G$/7
�K13�;i���A�Π�J��L똻+1F�.z���:�����G�+h����j���F�3��+����l!� ���W��̃2���٠�rU�칏�D\�ι`{�d?n�[z��5~�ީ���~�~� #y����M/�$s�u��MyXˉ-�w�X&�=(V	l��}]�j�qvVVT�W�x��`�F�EpyQ�:,{����gР)�9�'��;�lЎ�rU�7���Úѷ�wE��-\y��n�;f�u<�w��N��P5��)}�����Y�d�|��y� �1�ᵈ�&Dm�Vm?��%��(�Z�;�N4Y��T�";C�u�C�E��MAf�1�?��aI�p�ɬ2wu�װ9V�4p�+|�_Ev����A�iugy,ߛ��_�]n�m_�HZ^��,d�lN������<���ӵ̃�����!p��.ܚQ=���dEWh�
�y��%�<��}�D<�^����f��"<%E$6?R����X�m�!�!��*��2�ZJ-�L$tq�aοo�n����(��#rhT6��.ZJK�{>���I�i���q��ܞ��Ԃ}��(�c������Ѩl�|M-O�y�Lk;()q̦���ǅs�9�j�^���7*6��e.Q�������Q|���I�l+0�bp��n�{i�8�HFm�f��p4<qq4���8����MS��mv�<���k�Y�:�U�#�-�I�?���!P߅���7�����O��=�(,_�ͷ�SY���ꍫC@C����M��i�rs9�z�{	�2�P~3�z�Q��:�X��!���fh�^����a�Etoi�.�/Ue�$n� `!�J��+���|-q$��6"�[�e�����#ccr=v���Dn�`��w��N��` pBO�q����	 ��o���U�q-��|�Fh�!���j@]w]�ŏ�'h$���	�
��)��/W�)�*�;%���k3��i�"p�WOU��f���iUR�Y��+��J˶$ζ� �3_J�"7R����a�8Y	�V��P8d5�P�����g5-��|oR<�汔&�.��ZGn�Y4���}�����VUw�������Y���Kv����|͐dY�I�S7��a7��%m�s a���m�D��qK���H���YW�X2ـkv<�80�-�@��dۉ�s}����"��%�ԉ�5�����=� �m�I���,�=�5����Z2���D��y�#՝��X^�	�냅Mg˥N�Y��I��y�>d�VgFS<� w,혍G��X��3$���Iۭ�����p�.���%�
=!���8[�_����Q0��t��VLAt�뵧a���L�L�Ϣ��N�A���I_��ǰP�v����H���FHタ��.�_��
�~$��T�5�#��� x�K�D庝��<�x��K��)�ص|/�ShM)g��Ek�M��o~"4~�)���m7t�{�gXD�-��j%�%��Oi��WΎ���O���]�5���7A�nB����y�������E��,�ڶ��x,O��x�dZH:*����#���Tr`�Zw�b�g?}�r*5ҙ�}��|��jL�ZhV��`[4�⪙�w��l'��I�Y^z�d u����2��Rj~����Q-Q���ZJP�F��A�鿌<.�`��߷��-
ܥ�����m�*[���g�M�vi(����5!�N���}p�}�lnv^���fl]R���n���ݓrH�b��uG�mۨ��M����O�j�|�]z����rX�c̳ _]\)�?���rL�$!��@�0U��
���:TW���Z��5��=e�5mj�+�0�������LlL*U��|�w�:]D��/'ڹ�<��*�aH(lN�l�%��$LG�N��s��������I=׊|�����W�	E�(6��J�zis|����b������ńVDP��,雗���T?1y��fP�1Y��v*��%��N�Φ!�/{X�	ί��|�4�󜶟_�ۘ[.���0��}��e�,z,�c��VU�����iGQf)J{��ʈ�Y�f�]��C��$�b��:"|���U��l©��{lZ�Z���^���2*Ǿ����aF�C�����~?��iIuS=��('���ѹ�N,�{�r��s竍U
�/��x�8���DH���p�+��ū�1��
)�&+��o���K�n�u�w
$���G ��� �ڬAC���|<�\G䫼D�ߜ�)��+�N�<ڋJ�+pcTg������`��I���|$�`n�k.H�4}��o5����L�0���FoT�%T^ԥ�E{������K�b��������&��~w� L9Y�]�5��Un�����D6m�9o��4/;�D��)�R�/p�;F��q|'â<9��bϣ'��E�{��҉����c��m<y,�;S�U�ٞvE���o��f��&��-
ۮ�(��eR'_	[��������|őֶ�����e�X�p��Դ�R*63÷,�.Є�|n�S� NË$�Q�it��c����*mO�W�4(����+0�Jm�я�a�tA�^��kkg��92��ʳ�5si��X�IO�nvQH�R���?�%߄���ϖ;[Zo9��U>�i�=��-L$��<̤���:�O���ES����c9YȤu����a��+��T���s�W�?�T�+o��Ǡ2rZ� ���=����P���"�%,��Cu:AJ�U��6�&��5��r�h���*@����{G����
����׮���&Z���)�d曗��5;�����<6�H�|�d\�u5r��r*˞���܈e���2���.��wV��Vw�a������\VƆ%*�7�0�2�o��LI�U��U䖌���
	O��Q��a�ۑ8_=����Y>Q��x�$\M��ET͸@�~^��z.o����Fmud��&�!�0�H(�d�c�S*-h���pMQ�7��+�,���ה������0���Ί�D����)���l���õ����&V�k3��Al���A���ϱ¿��܁��6��>:��c3�w|R�(���xYո���W�P�-'mÒ����O+�eq�U��.~,�����n��a��c~���X��4�bLYq*�DB\�o�t�K�k1_�yRt�"_��6M�%�-oI~��Tp��$)��������&)$��JeCú������Z�5EU�,"V|qO�u�����Ά�U�#w��0�(��������>�����Ѿn~a��O!U� ?{��\��i�G�S�5hN���O�J��=yn)����?I����#�Y�L�0�y"�tț����b��v(��v���~Y���:��aT�d!*Q��������~�~O��^��}X7[o#��1�j��4!7��#���Z!��p�#��ĝ=9r�剛��/��3��q���7��f,�b�O���DU�fM}(�7t�3\H><E��+��Wl���@~DiR�P4�Q��6�G�yi�ሙ��AGS���A�*��@���lzYf��yʂ��W��Byiq�3OJ��� ��V��#<�>�ڢ�������OŨ�i�N$+��]~��VQƓ\���((�M��\�%�2nA�����/��fM�[�h�Z�^.t��M��"�#�n��ӫU�Hm;ׅ*P(j���L���>�ȲӺ6���ˌ��Oݔ7/I���(T
02���`�[�O�O���	�u�u?f�}�C/������DX��N>\Z��v�/��lCA�.�+6%	���0�ޭ��>� 9�y^-N4��V&��ޤ<U��6+Px��A�Q-\�7KV�9mcp-�����K�H�I��t���W���v<2-��e�A�A�RW*�n�/V�.�sz����0J8�HB|70���]E����̸��9���5w!ww�+4�����`��<h�p���{����0����K��{�e����M߽;m\(OvsW{~�{!�O��\l@K=�2�bՈXFBt�Ҋ�k�33�'DW 8��b�����Ɍ�b�︎fV�a}�	%�a�ȶ��Ul���v\|�Z:z�	����� ��3�D��i�E�b�z��T��d��Z3�U8�gۛ��M����W/�~ͥj��k���ކ�i���o1������>�4���Y��I�)2Ɂ`}��x�(�$\��A�[�E�H��ǤDS��D�HB�2��$����/(��+�j��jNP�3�[e�4E�I�SS:����h�U�6c���:���JQ 	M�wE߻+K%�,Z��0Q��UEP�;⠵J�f�Y9v��BGF �!lB��2�]!C���b��C�M�WεN���ў`r��Ue3��s�d���K�1��>R��BXӓ.�:�ҋ�,X�Zu����]c�h�"�s��r8��DR3\8�=*WI���
cJz;�'r﫠�eH�u����A�83��,^㮢���\Y����u��ws�Nt�i����Q���U	Pn�P��1)�.��D��mY���B�#�.Xm,�q�.A�4�ڟY�SLJ��K^fK>8�r+BrP�AB��K���5�1�S�O4_
۳�=��ًt����m= {bX^�.� ��rH}\�uwf��z�a�[:%䪯�[RJe�KǀU�jVǵ��\g�X�bbCrk '�)�
`���	~�kC���n\
�+��ִ
�⃘:7�&�V��t���	,��V.x&cOra����s��;9.�W�C�� N�Ò��U�5�'`,�G�x�9��E��B0\�=B �|id�G<m��D�l�&1}�Ze%T�F���N��!�FR��3Ol}����f�H	/:~=;c��PY�_K8}Ѡi�y�㓈x�oƶ���@�ǴL��21�ꂣϞɴg���9mT^Y��{=�m���t����(<�2���ڑF�;L�}�L��g�o&�����g�d<����EGw��ΰ���0iA��8Hb��6��J���dE���=��_mBrS4� |M\M��n|0�*?fG�W��@1�z�9�̶�I��*��e��� G%�@-}�t�V�[f���4S����7)���������g��t�zt6}�L�O�
�w� 'ۂ���y\(/�d���l��D]l{n�gЖ��(��ڛ?g�\[|�{�G*bO��v�}��t���c�J��z�^Lsj����D,��}|���-���a�����kj�mG�	9�S�HVxl��"}(�iM�g{�A�QC &$�]����͟[3u=<�ؐs��?g;j��G�j��N�(&��a�Pqn�o���C'Oi
04%ck�3���ĭ�_�F����Ť��sď�W�jA .�T��Mb�k�~'�����g{��4/��o��			�
�g��&N_I� �d�^�fB�_�$��Es�#ݘ�3L�t��4�帀Ƚ�}U�q����f2Qʹ
��-���u��=Z[OJC3�= P�8���:������ͯ�����K���V>�~���w�]K&+y؊~���O�?H/+m����D�1-�� �C*��h"XL����r|�B=���CyY�zW;�&�8jU���1�Qb��|�*���������Y>� �ͨ/5�Vt%�ʙ��cd��QmtO$��s�+:A�Wcb|�����Y�aϲ7��)s���`L&�̠�ީ��r	J/��+�8�1Ɔ9��QW[�}�666��I�Y��/�H�FX#)ӻ��sI���Y��k���<T̽�m����V�&�������B3�`$��B@���`�>�}��x1����{�ݕ��Z}��襰N�����NC�u�y��<c�M{fbM��6'ޙ|ʹ�Z��ϯ��ٗ0R}�_�,�#�q|�����}�����a���>tѯ�.]�j^����p���v��[@oD2�vVG�{��u��^YM��QǙ�cGἀ��N���'[�LBow��!{��Wm?gH=��6,�E�Uם^��E�"����V;�{�ȭN�u�n>Mt�9sW���� g��&�bh����7�jn4��>^>?;{�\���w��N~����d�[��y��ǣN�P�f��I��t�&�z��(rr^?1��� �p��������H�l���7mk9ޛ�����O�[I�4�R"sߖ�:;�s4s��ϱ �}�j�;�t����v��֒���3?�gq�h����7�W�=R�%�&�������GS)T5��!K�'E�ܖ2*����޾�d�А��QN�J�����L��:1-��:������\M6�ͪ_����T���~�߮OV_}
�S@8���~�a�?��Y��j��k�<���_���EE���G��Ⱦ����߭vԡ��������1�	�烷�����v���s�es0�����3?[�ߵ��G��Ȉ[��Be�~�3�gm����Uq�7wuD��A�i6w�%95 R���� PK   Ŧ�X4�:Eg L! /   images/840d763d-d5af-4e15-a65d-aa66cb855cc5.png�z�W�[�6R� ) C#�����0�tK7� �1tw��=t345�p���}��w֚5{͇}�~W�}��*�`a�a   `��J�#  �! <@{��O#3����^V�����lr��G9IqM��ö�=�WW������ٽ�¾�ƾ�L���]/߸w�b��t>�7#�^ex���q���qj�qz��������=��G�`0k͗
y_�3�j��er���[l�P�-���q�5)E�&V�?Lr]�5��v/�{�V�?���na�/�N����I�V���)8i�h�m�Y��'���ïo�o�v���o�w�?~�(�q��9B�1�<�=x?ҽ��~��,��^W��WhH�;�s��(��[\��_�����O�[S��ۑP��`q����(ǥ4���.���vﻫ��n���������#΂�k�k��v�=7씁�)�� S����ܼ�T|��w���?��?˘����C��ɼ{�j�ׯ��z�6S��C��Wi��­�Q��0�7o���r�2=�n��{���t��)������b��ڎ ��g���:�!�4B�� T5����� Q���l�_)� 
Gj���Wqu� 'K�}d�C�u�k~$����JIl�8�î����dt8�/�l��|��<�WN��(_ۯ:&lW�/�c?��@p�٤�8����܂\�d��\	�K>*~vHh?��<._|7�+)��֛p�����՛���4؂R�Z�Mgy@$z�����ѳ����x�݋dB���z>�� ��v<�j�ҋ$��H�7dL��.��2�9A�2�=���� #�KE�y9��B�����l�_¢jq\�D}�e{���,�vrC���Ԯ���R��u�+]�dS���*[��울�-��ϴZ�8�]���^��9y�~C�J@���^wWИ��ɦ�&O��:���M]�_n/�.onn��_+ڢ��n�{u��玻����9ZK��Yɤ�_���Y��55����n�Z�ϥ_�)s4�Uƙ���v࣌�/r��u���C�NF�	�,�0'��b�;�ʜ�W�����f*��T����=�*�7>��yz�ԾHwkw1�]t�zѧ����FDC)�qž	-�%g��u�� ���5��ִ���Ԝka�����i+с�ȱ�r��뷐���pqi{�^1���A���(jy������8��taI~%�S�[���3]��=
e˨�*�f��)qtw�0�p�3��srz��9#��u��AB������ث���fXu��O����]��DCɈ$����@ಲ,���;
yUN�� �eg��a��7�h9����N��gDD�'�n��D���?|��!�\L�l5�srv��M���)�����j�V!�䵉8|�Y�_-�u�F'j��H�<ݨ����jp�ߖ��V��OI��u��{�/x6�bA3ç����p��:�A#�SM�D�>7m�'�#�`�)a���o���ݝ4�n~p�Q�������6C}?����x5��9Oʮ@{����%�^]�TːER�j[�g9ǋt�b�ܼ}w��6���=����4G�$_�h�%
>�!?�!�6`0�|�N-�;Fi���&�w����>��t �s+�T�yi�����~h(?�I�EՏE�ǣh��C^��z@�ܖ��.#����z�$�0���T���G���[�6i&O��͠;رI��f {n��"qY\�*7v�KU=����\B�%����9'w��hn�-�)4p�	ܝTPò��́:�t���m���s�_}�xm��Z;�NS8-E:������щ��)N�@�6�'<��{.�۬�fŶmZl�o��:M7��27��d���'-�.^��[�б҈����9(rG*4[�4	[yǈ0"?=/�gw]��Ɂ�lAߒ���i����C��������Q�U3��ߣzt����Z��c;;�Gpl��Q�jK���o�W?�o���iF�Y���L;l�q��+Iȷ�ov���Jݷ��[I���T� ����\<�c1�PQ��%�v�����3��_�����������F�����B��e���&�ӯK��0Iz�E$|niJj[4o�*����L8��M'z�1JY���E�UԀ\���"����߼1Qd���~d�4�;\t�y�������Ɵ�Z:=Q%/ؤ�A%r� pW=�m��°Q˗�иgQ���_�z�ƶ�2���wȣ���}�|��t�.�V�u��@sKo��^'D^���5��N�ۚ[[�[��?d��),ۥ�����]�p�>Y#N�'U�� 
.g5U˫%ٜS��n �>hd�!�]G�!��C�l��O�yg�d���1�@�'�cH�!�����R��c*(����pD�~.��55�L��e{�eIĤ�.ꏬ��լ�M�ƴ������.N�Pu�O�W)U	o��򥥇��݁ǡ�������nq�k�m��`S���g� ��	�i&&����F�޷N��~�Rۊ���#��T�FW%���8�D��Fyk�%�(-jkf}%x��Ԉq/�0t�h����`bx�S؝Ľ��Ig.��p}Xޭ�����k
�V�k������L�k�^���WHsہ�׮��(����$��������>-�Q>W^Y蜔unp�d�Z)�����&�����k�^���~Q��h�/j�o�����m�����t���4���59��Rw����`6�!��T��i�
�	��<9�šN��׵1:Xx�,�Yq���I�V��wp��v4#'d�D��,r�DF��u�~�O���
R�(�;|=����j���3Έ
��%qP>�O�0����¦I@"������5����3�0�����A1IU�����cG��������E}�q;���gRNoo_�;�d�����SS��N�	a8�w�à�D�SR����p2s�+W�}<�>�@f��9N�ΐ.�� ��52wPш���#���c�\&�mƁo����zU\�,�S�xK���8�M:]7��k�~;	�A=��~v�bD.O8��XCQ}X��W.��\�,�N���Y�VqsEj�5އ���Xu]��f"qqX���`�񆧟It��i���L�4�>�O�@���X���8�ǌ6�JΤ�>���>�K��*�_m��(�*�Z��9Z��Ч0Rr�k���u�ި.�Gj��ǂ��Dd�i�?;1�J;�Ϧu���k���xe�s��,3!mz�#Y���m����N�eAZP��姛a�j���g�?E��B�D57D��@72le-���)c���L��,g�+��V|׽[q�W
iKM����[����M�sD��D�ٹ�\�iy?�ov4�*��4	�}Zw��FAt4��y$�}[W^dMň%�����q���v�E
�?F�h2en�EաGh�E�"+tE���Dm2��Q�f|x�;84�w�.���(1sX��tN�y�غR��~�s��0,�	�O���Zj�t�|��6�6��&����tww�.59pZ�
I�'�1MG���R$�Œ`��[�)�-t!�Η@�_�Q�k��`�$������{��P���&�9���,�#���G����9TZ�ҺW(�����P�P�a������g,,,17:�ҏ�g>y6R��d�'v�`n#�֐����[&<�o��HBY�1� �\�
��UԵ�B�h�U|T�x�|���+!8��
 
I���̉�=_ٓ�q�G��xG�"o��
�7�]��3�Z&q�W�jx��[%�B�s�ª��<dz{D��j%���d˫"Zx�<Z-����䩉�ȤL�/���B?�Q�E��%�b�$�Ӵ���|��j	B�5�����1��c��j�ob�+>췜3x�d�K.�h{Q��x�L�-#��C_�Q�0�
�����]����$Σ���{���b: ���U~�������H���a|����T�6�B��"I��A���˭�3sV���y �[����Z$j"�oݥ?2�<���9�A9W"nGa�M��XZ���a��πm�+���m�1���/��ő&ن(��=��<����Xn!��\L��<�Sb���{��������\v�Z�������$�P:��Rk�6z�N���m���O�<#�>�B+^S����Y�4+Fom�Փ�'.􄼮\R�i{kBŘ�b TӚ�2�30� ڹ�r�+��fQ��V����������B��u��O)��\�l4Cx��ADT����Ѳ���O����cc@��n$X�pQ�82�2���#����d��-��3U��3�Q\��'y�������灡ȓ,�"m��7"�'�_Ti��BKD�ND*�	on��z6����}��*�m��!�k�ht���; ''�<N8^�p�#?�[E1ǡűX�$f�c��E��S�.j�/�a X�+��N_0�m�g)�g%�R{o�x�
��L�x	�h���nm0pcv����jcE)��Tl�U�Z�B�ͧ�[iG�+���Կ)�m~��Bc��Ŭ���6	ˢ_�}|3����\�㨢��{�{g�E鸁p� �w;�u~�����x�ge���/q�o���6&�[ �)��~�R+�f!�<�����k2�)�ke^��v�<i��|�-i3���s'"Q�@�����zE4&Wi�Lv��"o�4c��@�C��-V�Ҁ}�"�г�+$%.���i���n��R�{Σ����9�9j�Ë0���#bđe������Yg�Ƌ'�B)�E0�
�.�/
S�3p2��|^���W�=qY��=��4����n��;�*����]h�-^��������+%�p�m�zfB�����f����*�3�5T��#���v5X��C�[m�� M`�y�N���r��
��d�-����0Kˌ�|(�Y4�Ь
P���5�ܺ{0���
3��"D��4�G$��u`�1�g؜�9�z�ܽ]��7�֢�vI�&�h���f�?lB
�fs��L^KD�-���=E�Y�U���%���ѩ�.�Z��0r�:"�%H���:oɯ���jk/�}v\}vޚx��- I�q}\��Ux�w�?+�ҴMG~_� JW��,�Ct��q�b���d��DK��Q����/tK��uHqr��L��>k�k|ٚ�o�ޤU����[�q��������X�3;�xu����T7��.X��~�!�C]Qsٙ˯0t��}|*�}n���N��;���&�R,������~i~��q�SZZ��
�i3��3�ԤoD`���ތW�}/;�@��5��̥)�O�f�\7Tw��IX�E��4���*����m�M%hR_���aI,=m����ƞ�+����9�9�g�0:H<"�p<]�31���R��`�ߟ_���Xڙ�y8����y}���g�z�y�;�p|�P��᧰2uϮ�ٸ�V=(��݇�ꋒȫk�)ZL�M�:�_��(e�"�+���x��\�Q����Vn	]� ����Ce�a�k7��L��v��z�8�> ~�4|���X)W.s�R�����e���^Oo�L����y֣Y����s/��A��F��Ƣ��3,��x�'���Ɍ�u{.0��Ѿ�CY�0,D'R}������L�ۀ̛n���E��,�U�(���Dj�cj� �>8�������;fƂ.:Ng�b$�L��k�\i<�f�㗊�퇟`;;��-�Ev��DP�>�=d$�ΰ�~��5�i�ɢ;>�_Zhrܙ9�x��R�/:K��Pp���{]�0��E�wscFI�=����&�O�kbfffR�ʸ��z�f��r��TH�b�� ��$�화�m�Qm1�a�V\q�1�����	�,r�o�אӇ6���'�L#�U����59�>r'B'U�G-�M���5ظ_r:����l47��_�����e�<�x�f���
���n�,j� _�~sN�
P�ٔ�^c%�3`�np:��&%%erVC�Z\GCGH=m�˴��.�٥�W��0e� }݂���޺X�e�35�C	"s3��U��>f���%cJN�!�2qw��#�U}�[X�wρsGI�J��ψ�b1�ү��� %%�o��X�P���U���J!7��7�o��u�j�lگ�@�6��-���7���*����ym;��ߵ�׻,����&���WB�]��W1��J�:-�ut�}�[G���m($]�r�b��z[l�@�U��^rOک��mP4N(A~M)j=��\�ΨV�KK���[,sq ��~�d�e�����]�;��-ֽ���N���:��ߏ���-@�X�����4�n難}���+++mgy�n�E,�'&�_9�*�D��[�`��ʭ��1�(>�c~ddD����=��V�ϧ�g�s���`R�Ek?3:fccc��K\�c�e�*�I�^ꞔgN�p�|=f(��]0��O���Ʈ��������r��*��Z�h��
2���= /�&�?-���abP��M�f�c?a%����i���	����ّ�����א)r�����~v�g��
*:[Ϳ��!�U�R�D��\x��b<����mI�	}��΋e���O�k�bȼ8;;#w��6u���T��{4hQ�s�5�:?���6���K?ʣm�S�_ϝ�K��L����'�Y�
`p.@W��f�ƌ=���ߞ�`���Ӄ%���&"�a~ޜ75�0�ҢHo�tSS�q��`L���R��}�/��_����z�d%mJ�x���� �!~��șw�5c�jX�?dfA����e^�;e~~�T+�Q�(�~��[����_��;�4�')ֶjs��<;�(�X����R�ߍ[-������	g�;U��Z���Ʊ+��͜��|
2����'��=<y�6����4��&!Y��
LaM��玽���_L�t|�=~���Ķw�̔�~6?�����7Z#�����S�k�伔��F?M�'VZ��kJN:�8TIm�_����
S��;�J-0�@8�;�K8!��Ә����M�S�TA9zX[|>>��$�����2��=�ߐ_�l}�XL�j����	z�:��.��� ���#6nt?ߎh�[y��n77_ӻ������J��)RUi鑞������B�+P`�����<��r�|��Nĝ,1�t�����g\�P@,�B}TE�����GI��g�A�VV{o�&�0����
�=�fL�ӎOI���߽��}�_�]y�y�����w�ۼsi������~����Z�G��%�6����>�(�:�°���+w�l����������b=�*]�w�@�TJ���;C)���9,�5���,\��x��L��ʼ��Jް���ņ�D�W�?��_̮ܞ����z]�ː$;x��Īe,��)�p�ѓu�hhf-iY���c[&V1T���T����V���K����r�����rbc�5b�RZ��?���B�&8'�p����-�W�͐7�Fb��y^�p�(��L�����tc����$�;)
�7^7!4;�wچ��F��(.��&�%d�߯e1���F��!|���Z�%�-�N܌�/>Fm=i�ǨqTy�)��K��'`(�l��)�\�[�(�0|�5�ĳ�9X��_$N�Q`����R ,Cr-	4���Hr��y��:������0A�X���i�F�l��_�gҮ|�^>��q�P̢p��l�Tl�H����t��X���/2�Z��#D�I�F�S�N�Xkr�lym�3��wh�]B^��k���a�	�<�D@*�+bs*	�Zk���#��7I:�
��Ӏ�֤��h�k�GS���(}W��k[]$x���b���u"��bQkk��H��_�i�K���Ud:�ȘR�����W���RȬ����'nGr��^AU-(ܪ�_�=���3��2%tА�K���d�����lZ���	KEOr o/~�6�ٝV+�v���N���i8�a����;�ِ$���E��]}�
�����o�T㕇H�F=~���q<�1��N6�kM���[��1`�%�E�fu�,�3�6�dZܴ�/��Ek}�S��R\d$�o`BUS��x^�"�3G�Y_�ktH�_�;����ae�)��s��й�Lp����5�9�$9�+�^̚É��գ� �� �I"�W+V\b��@"}���� `�O�x��]��}r�����=��]���q#UZ~&*�ƱI1]@V����
S;��k�~|%K�mld
����5�+$������Z��q�؉&O�z:^���-IIjZ����Ï������|�z�h��IѕQ���-f�p(U5�iʏ[��% 9:n+�N�ն���|��\!�'�iv<�E��Hg�0Cb���ɰ�g���)_���e�*�ffK�;�+o�M�Z�吿�v9����X�r!��/�^�+�gt����;7�Ɩ��,}�,pD�+�p.�{�t���>f]��6h峸�U[�t3Y�O�O�h�Eh�A�Ȓd�'<�[$�r��E���*�÷�T�����$�M\�A��d���-����N��]8��lƭ|��;��O�vݫ	cY�|E'%�c�hm)Ц���{Y���h��3���S�5R�JE=�V���DsG�z�-�Yo��;���o�.unbġV��c������w��|���Tq�$W�+-Le��٠|��9�}��-<����}����y���h�����n/����ӽy�h���Cߡ���?�nw|�0�{�'S�5��K �y�K�z*�Ѥv������r���T��9Y3�1�
�a������B4�ۖ��B��X���O�1$�i�,).�JQ���c
�u��MS2��/7�2��G������Y6��Nd:�y���r���<�W�i>/��UJP��%w�5�2��L����6�1(U�e� �y�tak�T��3�/-t�h=ߊ�>B�q8YG�&��9�ݠc`E���$+����v���Cy:�w?�ݧ2߾�#�*{縪����q
��6w�� ��&�h�zv��G�DmK�
ε�<�/J���'@_�P���R���bE� �R�X�G���%n��k���_T>���:�'�x'BHE�k���ؖϴ�`,1���M�e�I7��0��x)IS��r��^_�B�0�2^��ːz����)��%���h�=�X�ѐ̐�T�D��G�M��t�Ԋ��##p�^��'"i���\�q��B�
 B���q�3����E�]�4Y^���B��]�p�nZQU��Y�h�& �O�;�]�E�Z��+�q�j~�K��

�b�
��F��M#BWcS<�ޡ���&��:�`Y���u�7ZF���hI�Q��K������w�>���{���&�l~m4�|�5y�o~��t�qb�c:�$6��""��o�k��$.�&�����=g�����?{�p�9�B��+ߔ�B��J�:�9#F}��PX���,ak�|���1ǝ���� �%��ت�ΏnC�J�M�82��O�U�ﾦ>�٨�շ��O}��q�%sԵ��	�M���I1:�v��<�?��"���v%�};Y�`0�4/ɻ>m����	KR�h�/�
˨�[Uk���q{X�:*�����zy�7Y��s�xW�.-�7s����~j�;��?�w�]����.ǵ��ߵ�7n[o�?�_ոP�ZD	u.3
�E���ϧv῏�S�`��}��D���0KK�V����X��cs�7�Q�ә�kʘdBa�I��!c$Ug����X��=��[{�����9"������Dᰋa��)�O�T+�ަ���Z���G�.U�u�£��emaQ��F�t�b��o�0p^��p��m���`yx�z#l7�t�>{Hыm��X\�5� �,P�:��N��<N����޼��\�0�Q///�ʣ�Uܳ�L]�"��R�sb/��Hy�bj4
�FQ�7�.XQ��M}G.��/cJ��V)����#�F~-��HP��*�zN.��?�MLP����Y&w?�'�8)����ڨ���ʡ����v����v.����iM�myx+����L �S�i�/�ض	6L4H�Bl��'��0é)�����wSa�ýn���g8>��NƦ;��PL\��O�~��`dv�B�w��w�J���c	���)�)�Cyy��/5-��d�G��ޛԾ���\f[mQ�`n�bo�;���.)OR��(h��֥E\@7�W��{�	��MO�H�=;��=������x�v0��[X;z/e^��]�YA�i�so���h��CИI�w�����f�6��������Yɪt�y4_�T?��Li.���B�ղw�H��<��V=d�Q�Nn�'���Do���%���LBr���%x�q
"��B�P��\k Odd_0��܉�nv	av��t���1�T �r���.��N&�~n!|�fk<D�#x��l�,�;)�7mTŐ���-Tf�X��ZqN<�v�~ʶ
.K��j�����X�83�B\	�MNs��ZS;��g'��i���sbS�oU��ʥ��;�;└��gK�K�İ�	�=�A=��9�,f�����{�<�X_Z��8W֚�{w0Y:��!A7l��D��q��� ?�㋤�z����y�w��QlTzUgO��P�_yFV��S�}���(V=��I:��U��'�!A�c�M����U0���ૹˌ����y.B'�c������ix�i;�������y%U�hz��[J^��x��v�JalL���M�]
5w,&��f�>�h������oE��*Gr2��+R����s�g"R����.�`��;�Uv{ӌ �Cl�ϲ�Ѭeߩ1v;���4cڄY��7/��y|7��+�)Z���:�M,L@�Љ�>�(�ĉ�5C�ϭCq>m�(u��-���m��Mg����lgTL�ޟ�SUhPTfX�'C�-셷)�W�O�?��9��5����ݷ��]�͍UUϾ<'�Ox*����yR��!��֎]Z]�C-�0�{T��j1�S���J��΄�ֱ��Z>U,w3ޛ`��Bṟ����)'S&Cy��#�4�)֒���Ր��^�DDD<%Ү������1�����"5>���^�k��Q��,���c�/�d�{?~c�ҽ���^a�������a��GY(�-��@̴�4��n�[���2H��l��3�3"����`&I��X����[R[���WEs����+�	̻jKҁ�:S�~�o/M�˭��$3�6W&�ԓ�8EEWpE_�f�N`l}lw�k�Vj����3�(�¶��Y�����PT���3zc�T�7�l��Gv_^^Z�2�o�9�E#�su��˨�;���m�U]���+\�3�#�����R7E[���٥/�P�eJ�Ƙ�%�|���C%V��&��7���'��3h�*TL�Κ��Q'Z�����=��!�!V�T��1�����27Q�2�~��l�qEݼ"�=x�����Ê��F�Z�i,��Y�#�j�H�X���Ϸ�z�P^(w�)h���f��:xNp������\��2��K[(h�r�}J�k$*wuy.��[�:]v�Э��7Zv���J���,b,��M�o0�_Ah���� �	:[h�+��1�uB��Lڔ{��{��"1�#�G6S�Q�d��=0�m��s�_��������b̀�+(�brM�U�L�9��i�y��u�H:�œN�G�XY�B; J0��1i����t!»��\�F}s:�m���"�{V�_�~����b�^;�G�T�ߤ��}���/��K�8	���(y�U�+gȔ����W��H�e��eoU���  ��!ۅ�\dg��):6�P��ERf?ro��j2�u��{)XޠM���E&CD[�ʿ��W�w�aK��h[�����$�"ɶ�&CN
�qsR��4�j3a�u/Io.,%O8|T|Ѽzf1Wڢ.�W2*�sk����j��f9f]Ìa��p!�$���Sq�fT)U:���bY	����)��7�";j��9�2�p;ː����U�4[�T�#
j����d�����9u|�*\�]�Z3�{v�GY���a�D���w���K����
��;�jLŚFa��Hv�g����վ&��M���o_��۵�jr��2u�$��] ��)))�4��$ʮo�?�̱�^��V�Oz*�
o|CD2�y%��)�����g�����Z��api�8Af�ש��.t�y	S��;އ��x�S�ڡ��-ߪ���Tw^�p|+����&Č#��D 䱏�f���|qd7i�_;�GȢht�9Lz-�x��QcR�2-�ϊƬ��-��w���'�����{a���`JC�~���?g��N���kO9���FZ��
�7%I��,6BZf�E��T%o�s"o>���7+��9M��4�AԖ7 ���&�ez����j쾮�h��_	������=��������W�����;�����5r4�������ɠk�{�I\�_��`Z�"^���?����=*�lrFmql�C��L���$����Y-��!B
�e~��&��UF������U��
Y J�f�4r�t�m�킬��@�J�7�����B�&�FĚ�?�Y8��$�mz��#�kgJF`����|3��s�K]ǝ��kdJ�7�g�®�i?=���Q����O��FxB�{hy5��+w�û����;�%���^�2]M�ӌ�	~Cp%�L:v� di�7����SF������-������׹�ӜQ���SNtU8�i�<���똼視`j(����i���	�좔�u3�%�	s�%�x�,M��1��8\�Ҹ� �[�e
7�ȥ��s�� 	A̬p.�UI���g#�v񑅰���gzYrV�����X���	����/jHq	�cT�*�>����A���b��a����j�Z�Wt���pJ1��'�1����V%s��S���Xi4'+�듯�C��3=��`��Q�'Y��7�c����T����A��b���A�^%C��>	z[����zYBu�lOR��x��q��X��%x���X@Z�QD��Y#EN����G��x o��u��)M����'��v7�N�TU �D�)A��z�7G��sq"ݜ���r��X}�^�!?�̓�n�ےpssc��/C(�	f���QlG1����T0+/+����B����\jlQ�ѹ'l�߾�����+�� Z�6m�p�L�UP�ۓũr6"g��B�r:_�"wȢ��7��	hL�Y\p�3PH��^?7+���l��q�Q)q�P�X�f�5%5��o�>���
��D�{���3�L�����#﯍��(D�K����ҙf�Lҩf��
9�*�o�t>v"[l��DK�ϣ���u2� c�K=x�C�0S�܈�1��s�]�q6���}Ьs�Xi��G���](R����@{k�^��L�U՟;���h=�\�<v����q��|���n������8ܼ.�c��Ϟ��NcH�0~
zv�T�ۚ�-Mپ�"�m�\t�|�[&�����2�rYWa��=3W��ƗG̙r�Yz�7l�bI0��|W�r'�e���5����ayc�X�.�>}�w���uй��Y.�|�3Z����{�&�>�C/��wF�cΧډlU����=�)���R�ܼ����\��(�m�[K�쬒f�>8TA��:/�ڠ�4\��2���R�k`�"�]&�KS���H�\�E�}q�\���>��w�R�9�q^z�bi�Aݸ�˵��ޔ�.�j�PK�/��@��8�^ސ�g�3��m��(1�P�2ƹ܈ɍ����&3?�]�o\\X@|�T{�C����!��V�!$��&�ut�� �	�ҳ�����l����!�[�\���u�<��w"�E�u�7)��ɴU�.�q�S�]���B��f���kRnw9�C�%�=���f�HYc.C�����	�P���)��(�����'��`����T1�K�Ĥ��C
�v�A�"[m>S�?�� Đ���}��������GͼJ���?��t�4�����M�g#��
�ɢY�oۦB��W�A.?E5՟|4���(��;�(Zam��ZۏQD�&d�J����Pw�g\h���#���>���C��z�s�����=�:bK6-���xpHYg�B��'�8'?ً��$�GE!��(ܹ��NNȤ���9������/^�5�|rԗN�tH)mX��׈�yA��'�S��X���4~�n��'o^�i'd��7 �g��#���kH��jV��w�ڲ�e���&+���O�b%��G�������9�J8bM�^�2�tx�<����[r�>>F�*3շF�3�n	���и�=;����8��;yw��̖^�P�O��M�Wp���:K�i <�v���F��bO��,�)�ú�Z��d������[�wm�v���dzx�}uuE�"b��}��n��[�q�>���������
����$�{E"�A��X;I%SK��:RC���JG�qy4k����,٬�����r	ˍbO�0I�)搊��^[�NV�_����nEBF.��E����Ee^�J���@���mE�נ��m+N������5�F��gWeЪ���
��+.���
�i5���PZy#�0Z껇Y���/�.tg.[k�-'L@�p/�Z��H��m��y*��B�6Ȋ�KV�0�oFr�8!Gp'��0;��:��i%D+|�%"�~�Uq �Ɇ*	�$kҺ����(���M흸�xz��WF��<��dY���k�b��1�ض����Db�&�h2��C���%��qފ>6��W�8���W_��/Ϊoo#�-�
���PS��h�U�\
�S�q7M�"x�L>�N�y0u��<u\�k����	��L��������<�z����<��(��S���$f��|{l���I�o<|@ ��t��J�x>E��Gf�_:���w�j���↫�Lz�@u�Y[��(:P�!׿��,�eQzX^���O���w,� ?�gKL����ԗ�>+<C@��L������ `��j��.��b]��1+�Y%���M�[�y7hI"q�f�=���Cq�>��R�_����h���ejX1 ��;zDHC�4�$����;�q��))*˻#�ÿ�2|�_�u+}v-c�Ufq��C����Ȭˇ��_��z&f��(�=yh����]Gpɇ�ˍ`��5.�8mB��}���J�=�5�d�����X⠁N�j��@�����X�zd%��ڊB�m&�o���P~e6$߿AT��U��f�}��~�V��#�Su=ر]8 ��g���7ڶOZ�6�]���s�]wq�������q�f�Q�ޛ9l̫�Y��E`|�����k�Q����B��n��qT�x:���¾Cv��e3�[=YC����E��1o&|��Or�ih��{p�W��*pު�IM/v��*>�6�`�U"i��UC����p̑{;�/���t�?-�{��;,w�z�^6�eK_H�+e�#ӣ~�-��wz��h�T_fy#E
O�QV��Ob����(���q�����AV��Tj����UΕ<�@�QO9���s�;^p�:zЄu��X)��)*��`NA'2���X�B��n�2�b�������%���&-��kA�!#/]]�F�_V��x����*��x���ƈD`��"�`j�P>Cޡ>ߎ0Rެ�����g��DL������d�F|M:�w�jR����0D�4<���������$��&����-{��k��]:nV����V�����W�#�7$�s�ܜ��1 "���/>�CAACe :@J�y��ɺ�٣�gwz��^��,�x�~Q�O�k���gV,#��r�Nٜ����!�x���A-��.[��N{�^� 5���^�n�.�
�EhEM��k*>��H���]@�ZB�&U�qq�V��\�{�X6�*B_'C�������<��)�p��G>V:�����xע_�~5��̡W{I�@���j���r�(�h��m�0�cI������'���W��^��ƛ�Xۜ�nױ�A�TT6f7��x?9"v��BV�����ǍD��������$�B�PcDz��W�$WHgD�q~֗��`w�$g���{�m}��L��|G�0�dV�4��.�.�6�[��е�J�������_H��!��	i�v�����эw����&����T�Uv�F�^���cc�R"'���U��r-1� Y=��-�P��s���:�OH���E+�)�����T���ǆ��LI���������\�ߌTR-��jn�:ݧ[N���//?]mFｉ- s8�3������A$FZ޿�
^)�(g��(�=D���o��F{h�<88�'\�t=zc�h ���ش���ʘ4�$rTU
�KW��u�n��CJi��))$DZ�n�n^�K�����k�\`����|��̝{�9�3wZ��A��H��x�fϷPG}GV�~������@z[�S\tH�Z�m�_�;���]�<W�;���T<(S��6q�]\m/�d��tUc�M4�Ѯ��9z}�呟D��򘭭�2-�`A�*uj!tB��Mr����w̓� Y���S����̔�bC���)^����z�׼C@8�����;�$Zw��v��\��S���3z���@���ڴ�73��|���~K���m���鈽���w��h��*v�uv;�c�#��� e�*���OR��*�m�Y��?Z|�FF������Ə�N�H�Ia����5�PO\��'o�q�8D`T��5]�42�ᴝZ-}��#tH���b3\�=ĈeH��k�8��FoV�,�Ӥ�K��MyqWu q������������Jb�3�a���Ϛ�����1��2�-��k���c&�Ϧ�� ��M55q�k>=��@Z��Q��@�8�v�^�M�(�Nk�L��	�����\��(�+���� ����p���ٔ��ȸc�q�Vo]��]�
���7rW `�oI��O��Q4q&�����DHvrܯ<\��6*�����s�:���⸑�ݐ4t�C�e[0!DU�ͧ��<112l/���TjO/��4��O�3k�E��b���������5���2*��s�Z�JVy�"�;�y_�L=��G��/mw��N�Bd����Z�e�jr2Qe������d�^�#�Fr'&���<�k��Z��;��{�NU�D����^�u���!R(4I8����h��s�32�ҭ
sd�щ��l>T������������:T�^˪���Iw��te�뻤uIp	�G�G���^i[5�?�]�==q�.�P�Ѽj.��՜�5�k׳]�E�(Ze���:��@�om����$�Ru��A>�|����}'�	��)�3���Yjܸ��x	(r��4LMC���E,�H���0���}Sn�������-�'�-58;��~?�!q8����4���m܎c£��3������2�U ��d�>}7B}(h^P7r������p�?������t$��9+1119�L�y������8�&��@�qM��"���eE�$掳���T5�o�	@�_���c�'�4s� ,�������e�����<H�g�o���MS]�=�Rޞ���T���Y�5ir��!iֹ��)O�??D5o�CŧO���i��3�-�ж��z�/Y������pYMn�,��k�"��H�ʞ$�e�Ո����'Ո	�����|g��J�(ˎ_9�EN`R��dH��q}��{R�܎L+����P(l�`���U�Pe�|ǒ�֊�Sɿ�44,�}$��LPdj���s��À�#]>Iށc�����w�?�r��Ə-���K�3���G������픒��^�NO]:A����\�o��n�����mSv����?ϐ���4W-<*ݤ8Y��"�(��2ӻ��Ł[2v�F ԟA̡�����r(����m����Y��KY��E@�9%1��G�C�˱ZA�.j�Q8Ճ��PND9��'��R�r9�,~�2�b+�_C�.���5�(U�5y�d�P�8�n��*��m
���D�}���c�G�X��z�Q���K��Yց�ĠO�?7�?�~����ӹُ�(ڟQ����n"����{�_x�5i�?�c���nN8�����2�O��M�f��zs��X�axδ�T�p;Q�E���e=��W�E1�W� iZ���v��m��|ˋO��/���:��qF苀���^�0����dQ�vU����t�\�+{���������ߜN��g4�=n���2�)~��F�J'���f��a6(��$z�H������	(e�&;��\�,�V�8BcC`�l�#�	��h{A
ˀ��eL'��~:Q�]n�.n`�L2�Ql饃��9�#���ߪ�Zh�є��W���	29MZ�=���Z�l�0Q*�d�m��xֽǰ�@
,3�e�,�B'n5��3�;�n��r5�#��L�:�=8�_jE}��X؅'[�^�(Z�v��|�Zg̵eA"�O�D���?����>k�-Fgݣ�x`Ჶ2�"{�Q��i���w�[�KG�����0��v7O� �|�e߮��Z�Sēh�&��l��U�y��񖟪t�9�Ĕ8'�J���в��Y�����]D����9��2�b���\W��#Hd��qM_�k5,��L���d4�uG��d����I���@�R�9(�.u&�k��

Cy{���r��rĔݘ0�g?Q�p�X͖4՛zI��me25e�}K|G�����r�z���yC�~0	y��
+���7���3����(�4�r�_�,�N��B�|{ ӯ�p���
FEL�9͢���jZ�{㠜��}'장�����ad��~nSO�K�Ǌ?[�OKrpގފ�ϫ���H�f(��8^�(h��!>r�/��%��$M�Q��TS
������zb�~.�(n��o[�忁)ɤ�j��3>����~�����͗�.u��h�y�=�(2<�ʡ���>��b��5w�[ 1��Z�n*"��vyw)�3C��������$���*��]�QLF�I���o�|U�1��߀&g������Z�8������]�f&D�C;�}3��k,M�|�N&�Y��.5�4+��.��t�Uo5�x6��0������CQ��#�m����N���q/2���¨�QM�;�@gh���,��D:�*����5��#�jn�.u�tUb�Pe9G��A�C�t5�Eywi��8n�_�]��Ve��j"~������$q;�U��9��j���ܚ���
�v�۳bL��zS��%M�OO#P��1�mX�z�����O�*�������6�A�+�<������^Sz��qT<O����:�2 ]��U�����	���@@�gV��H=Y�D�����YQ��0@]�Q�:�9����,��Wc���WE��᜛��4�z���_�O㼁qa5t^�Q@���۩���o�2<��7OwY�š]��Ev������g_�������� (�k��"x��Ҽ��Ŕ�����d$ݾv�])�id� 9Z��^�p��Y�δ��	~�b�
<� �`Joʿq5�ro,">�9��HGy0����נ�ql�4�dY߂� i�s�b��*�yN���'���o�����ogF*Wr��Ssw��z�~����V���C�����?F/K��=-*m���ݚ�_����8x���2r���Б��l���z�Ke�����f8�ϩ��� ��,(h������w2�ou���Ѿ���.=z/ݿB���A5�B?�~2��*6�2�>y�!b]����I���Nz�V��g8ePJ��}�
	�p�_N����:�����>_]�<���b��o>1��1�sR~�U��*э�XDU��"|I9��{+dd����ȓ��7Y�;�v�������N6P���0���T%�ď��ig��`��U���r���w��?}X�~s�P
}h��6S|��qp�{��>zd|��@�U�7�����!r�OiQ�/)�����#�`IO,3E�k������`��H�����l���aL"k������z]�;Y�q�wÝ'bM������<h�kG_���������=�$eV��v��2*�7XR�:���;�J^�W[7�QV�B�^�[6R>�Bi�5[��\I�oٗ�֨GB��25��GI�4�Rj�ڤT�/�v"�(=�����~��٢b��d-c�0��� �1A�]�ՠV�m�B�����`��2��8��M��э��#���V9����~�4��؞���)Ѿ��td����f_C�wՔv��6ʈ��WOt>]��X�^��g^�D�{�i}���VR��`=D� �W��*+_ju���~�A���Cn
�\����Va��D&󾿄G�6�ph;����Gd�u\�_(����	�~-9�+1ݍ�
���z��/0u���a�#�e*�����:�Dsv�p�qil��>{ܺ"� �|�J�M���ZO��]��0�Z(�&���p����.�O�`�<�Ȯ�ϪҦ0h�od�H��:�Q�\��߰4��7�]��ee������RN���s�=�/�)�i����=��nlA�5nҲc@������KB��z,^�w�!�l�AX��f8�������p$�#zjq)���D)?Jk1姓xa���"������G���SN�N����&VH�3��B9��c���)Pu2�6氾Vc�s{����D�����1�ؖq4%#Ur�5�r_x����oo�U]�a��G�����l�����A�Ky/)����D���>�
c���L�<��G���n��������2�Ìvv�IN��h�~#0�'v&w7�\0�+����!���j���UO�F{W�OT��v�[3,�܍<�A��J��_�>f6a@!�vF�+���IDH�
8��T?��{��p�		�3h��r�5�1�P�ې����Z8HP�w(Q������������-ь�S0(U�u�K��ģ����ʋ�>��p��Õ8牰���(&+� v�CI;��hP��$�����`̹ߐ��_N�y�yE�9�^Yu�D�Wԝ�u/8|O�~+*:{��1&�V��y�m:���S�A;*��&�X!�8B�?pd�,�(L�=n����Q�]�R��=��K�LU}_ߌ�ӛG�l�����j�B�e��>��K�0�l�~)�*V-�8A��G;�
�j-���I뢑[:Uj8�t/1��Cs2���t���d��	�m��xQ������>+g�
gp�:����q�\#�W�P�w��&{���Ğ#��B� H&1S�N��3ㇼ�(���B�.�Z�j!W����K
�	I7�}��m��)��_	M>��;s��by������ɓ���ɏi��]�p��	z?o�x�S���c�,lSx�E϶��~�㙦r�)*W�_��(�D���z]6���l�`?�J�ؽ����[(��kP�������f}�lm����7�P��f>��ō��c�.�Ң3�R�vYt/�+�n^ٯ���4��1`A�1�.�j���0��g���Qp�S���
��q �n^�$x������ҷ�R���̰񼶋�����Z4c4C����a<�]��qA����ϖ��d��]&�~������<��h�H-���7dj枃�����y�d�OI2�Z����a.x������^������0���g̽���ɿMK��h~�6�n���s�:e�����/�X��[�=��[��{/��C�{֕���x*���]��&'���]1B�s��M��]��*��٫���ػ���)�F|ƺQb�cċ�-�|-m� %�L��Q���y~���(�o�"���coo��z��A���q��}��2�$(�5��iݍ7d�� ��O�[�-�A�̮^������k�Q��
<<v&,F�5yUt�o�t��Ӄ��[޷�V��j��4��1>o<�$���)Nu������6_}msV$4��\���4�6�$�j�$F`�t��/J*�����B�!�Z�?Xٱ�b����N�Í��dt
�D���v`���o'��Z���JU�9n:D Z���L����`~t)����Ҏ��&���7���
�ctoX���v	����{���Y�]��N�M��.@\����� L�3S��bݓ��?�(�3E�����P���K��Ϻ�^�;1W_�A�b�z��t[����Qv�J�������\���}�ȅ��	�AW�/���1�-�G�R�Z3�h����=�F���M��DO�U-�@mA6%ȴ!��|���
C
���� ��a��l��M��<��Ī��`��U������n�i ��L�����y)�	͝�D[�C�cM����ɪ�v�k�u�^7�J9�a���3Fw1�R%�=�$���zl{Ѻ<��&svdE�~E�^)�ɋ(��܀���X�������k�I�N ��G����v��m���S�ֲ�)q#W��b3S4`�tz;RlXN�ژy%Kī* *�󫼖��k�*�]���a�2e��x�t�`����z܉87��,6��W~|qx�춑�}���H�I�(�Sv9��0��g-�5�/��d�D7[�l}�A�6G�:OXT��������\���an3Y��:D�j�=����L�z{���x��	S����8��ʦ�2/�� ����<HO��=��˯�q:3�X2u�I�<������j�m��ބ�~O�~B��ӾK�^�:E��w�g���\�o�<L!��[��4���#�2��1��퐱��^j����؃��8��+s��-�	����z��'��}�^�$Q{q�~f�¾�"��a{[��siG[�g��F֨O�����!�2��¯^!l�rjm)�	v����e7��,�.at�xQ�]�_d��'�0��<?I9�R���@�gY��|�%]­�T��򩢞�[�*-	�*`X����0�C�R�.��.y �ס�|g63���,�!AQq�3��/�������O)mu�j�۝�( �H�l�w�|�"����^4����_4��i�m#���]��T���M��2���w�2Y��n1�3!F�L���g�E��]Ԗͩ�2������lq�1փ���)�
�o���a��R���B�e���ܽ��-C��t䎊���O4�4���߷V�������Rf��eg�P�륧�.U7��_iX^i?��jΆ/�j��٦k-��#8�z\�q�l��������琔�v����Ml�c�>��ҽ���))�i$��o+��~Qװ�_h�Ѯу��L �P��<�缹����z!ѻ�* �2:�3!JMTP���kŤ�;��?����}׫�m�K�>�<̈́Yh;u�� �����u�ڝ������/}�%k��	�*����_�|כ�'�A���'�'������0�hug���&O�n6x݇ɍe�q�|4�*IDk���ܓ��j�o�{W ����Q�iqZ��3�GٔT�|A��e-^��(��JӅ�̔ɝc'�����Y90vMs�݄�˒�)pqm,��������xtX���:iK�u�T�����#��2�6L?jb�S��w�7�2Q0��K�9�7�f��2�"�����d��?b�)��O]Ū�"�"��r�L��,�����s��1rJo4��Ơ~��w@�ڣ	��c��ႛ��*m�����C�L7zJ�j߆��l�$��"�rF]����\�����7��.��tzm��ݏ�V2���XCk���M��P�[l �S���q	����C��Kí�ۄ�b\H"�w�{��*�uUc�5뱆��=}��L)�Ko��uYЁ�b�g�^�2�Enz�Р:�A\4�/I�!�{���#�֫t쿧��Pl�<G���a%�"q4c ��[�3�Ӟd&}Ou�D��P�����r~�Ru�}8'�.'{�N�a�t��;��p<�+����:IT%8J*���,��B�鳑��T���k�cHǶ�.����Z��J�K󗚪3~ ;�}
��gt7�=�3�2�ߎ�P)^��g��/�6�;גR�H�l��r�z
ҝs�W�{�P0�hz��������b�+ŉW��;f.���0�nY����K6�&e�E��K���m�a����3�?�G��}G"l������HuS�j{���]�9o�9�"�P�{8Q���gdmm���5D���<i<�P�戳䟪��n�w�:�h��i���F��ɇOP#%��@����qY���b\M˻5@�lM<T�7�;�0�T���G,}��*u��n�J��+�������?�B�r�u>������	������"��DĪ��$2��:�P��i1��:�m��EM��Z�+XURkŶ�ykf�����"��Qw(v)�|k��ݾ�9͇T��v89T1,+%�7�����c��U554��o�X��i��� 5�(:F�����B�S����G���z3zSծ��A{�D�t��y�+�>�V�3΃�M9kV'�u�#�u3� 9��� �F���z��.KެG��{[�ӕʆۣ�p�9������A�ڣV�R��褥T��﫹х\ N���ut{*[�I����T�)�!�\�0��c�_�:��p�����4�w�p٬o�}��^������)�y;��;;�F1�cy��\�����m��|򑡏1<�d��9��5J��O�Ͻ$E	$���D�75�hՊ��������6j�My>���W�sHV�!��.�a��T[��e���Y<M���ؼF
ЅjG��h{�(1��{n���M�h�R���i��V�O�0$X������ں��6l��?!�y8]�D���DqQ�_�~0�j1�f�C����+����ʯ�_����a�䥵׮rS��|��ƂLH@�׍ce�j�,=�s�*~�"���Iu����W%�J���qV�����b�V����7���̚�<�����G��d���&5��L�-������2D�
I��cb��ή`Z�k���q�G��/��7F���n&��L�k��"]����6]D~$�SP��w�^I��G|�o=��!�NFa��L88�Y~I���B�i2�y�v��l�=�c�8\�d�o�q~���k�@�;i�\t�t�4���C|)�"�ם3�|��$�e��'��j�eES�o��"���
X��(Y����K���	�,�*~Ib_�:��$�6?�̠+=pr�6m���v_�k�yZd�É!����_h8/?�#���>ɱ3�ңõS=�x�c��ݚ�����4����&�ԓ�
OGB�H�OA���W`}�������ȥ�"e����N���î�#���ZB΄�}\���b�(:V�[,�K-�~�q1�4�#+�QBQ	#���P\$\ ӂ��	#�qR��]��"��M�f�n$����I�O�ҍ��D*����oBZ������D�߸�
���������!��1��%�V�)�N����ᱩ&Rb�^��O.��
v���7�'���{X[c'��)� F+(����?�QZ,�Q/|�ǒ*�I`�Fl
_�7R��ֆ[%�Y?�0Ы�0�ISE)�ӕ�KAw�>fG��ϒ�P�j��vp�rO�P���H;k�Y��^�(��}%\>j�y�o�9[�
Y;�{??+2�+Ֆ8Өr����(I�=ၩ�^��jl�3��FF�>W��M�摨�
��t�K%��s�J�un��f,�mޞ�D����F����<\�$*�ScT""q"���p���R��0�B���%'Vs- �/o;��n��P����S��#<o�Z�OSC<�Kؗ>���B��n���i���\W��=�A��)�ջ�W�_18�� � ��g
7I>��D7���Fm�c��d�E�_�2p������`��Ȁ�JJ�����=A���P�|�������l>��!�)i��(�#5hNz��3�鬗���l�ǯ�m#T|�`�羯��ؿp���j{��.�m��j6����#��4��g�[ ��+�ϴb!�W2�l��(J[�F�O;�/a��o�|��Þ�	x�A�F���*q((��=T7\�7�g�ي�w]�oN���<����V����91�:i-�����:	�.G�����es)�j_��E�\JŽ��G�6��L���������2��e9�uWčm��z?�U��+�xdR��Y�Pb���S�e�bq��0��e�5VnF�V�)o?#4)@O��(�Ϋ4s��"�L�gD�HF�ld3m���c/  �'�sv'O�ƕȕ]0<w(^K�R���� %ِ�l��1�������s�|��yi��)���l�L�%f ��W'ј��d�;�E��6�{���qn���+뇝�����!�m.�_�j��y��V��u�*��Ï�w��/���bH��H���rV�vSϪX}�R��m4���^������������I������4�b������6�[��/�����~�����@Ij9E�yE�P�Ҥfp�з��������=*-�3"���h䇚�j�fE�dE��&�z��v6�xWQ>�{,�,��(��:��J��,yqT�)ϧK���Q<鹯H]4�������p�op�O�������d��w�f�:���s��ݦö��V��o��i=�_k�휮���)Z�Y#l����-n?	�L�A6���85�NN;��6xb�]���(~hC	�
̌�,������x1�9��v���^P����˷��љ��p�����c�5@�W�2U��_�|<)�W�������
��y��m}��an�R��p�o���lA �G��0CM�ߵ,845�����ٽ�!�Hn��qUS�Ln�� 69�9�+-Ӗ*�F����_��zk�X�1�R��}�1;,t�n��')\Ɵ�t���a�Ǡ��/��{����Х�)�~����[o�ul�o�Y�9��,����cnjyZa'���">Y۟[a�<mA�����hT��҃�*x2�_����gSP���g�`��!8�3u��|oVf��It�*y�66zt�����reJ�P��(�۵]ZN}����q�O�MDUs�HQ���AE���"v1o/���z�;������6�;��9|�i-V��C(��n13)U����Y�b�O�4����c�v�b�D��ҿ��w�� 12PC�4�>�9D��M �Y{D©��.�&��|b}�S"�U:��l�);]
-s�r�|[{�v�W�d��e^��m����0ȾCc�b��Y �fD�&P	s*��Y|�9�+3Jއ�`���=(�ҋJ���q����[<Kp�4�p��B^�'��h�l����$���\]P�!�΋��p�>�g@�̚GG�8U{��ܥ�'#���� 	>�N����؃��)<|O_�ߧ"s�^�i���"nG5���:V��O�m:T�=	�]x�)Z���fNN�FWy���/q"��;`w=/V�Sw�	�<"!`�i�Y@���V&��uM���*�i]7�U25'�M3�:�C{^ �*��|ն�p��fX�Ax�֞� �A�����n��քE�:����/%V��Y�cj�j'���{�c��(���M1���	�P�}����H������[`��󉴝�k�o �a���/z��b���t�����f�X�d����W�X��y�]��祝ح_d2o�)a��\�W/_�I�c��i:UJc�焏�xql��y�f�!�þn�r:��
l�	�J�ꃁ#��Hz�3�,!	#ƺ5IPra���@=�goo/���)o/�'��X��(�Fp�X4���8�Y���dj�Fn�O����T�x$������C�Zැ��'JY�r!��$�>-��7��IroK���a� ���5��v�e���7p�����CP��^	,:j�����$W�����Ӑ|��Ϡv�����:	N�sϗ6�ߺ����͗�^����...�B��xe�g	>�>�ż�/�׿���U0Cv�J�#�@����U�{����@˳��dn�ٌ8{"TK�&��Y`A,8�a�ޣW��=�uAUdph��䁡P�KAK�i���B]GX�.=Jy�o�Z�>0�/uK:����8�v��h����=�!��������cx|;I|Y�Bo�Ē�
�+���w�Q�p	'>8�^�GXw�A�Ą4�~�yCy?1V�����CqE�n�m��8~q���T�5�c���.��s7�%Y�M�ycH[��?y^�챦X��-{/�M�����e�M�������+)ua�/ؿ�qV�G�t�wu�5鎕�J�Ӟ���n��~St�� ,�������~������o��d[w���ES�1ϴ���F����(�C��$��VN'���	U��":��?� �Wˮ��Kv92�89e�������'M�/6����{}�h�b�U����LH��;��o=����~-�5�6,/ QX�*�>'!?�>,(Q��ɑD�~�C��ΊFF���I�B�ܻ>O�R3��p9����N*�T��(�(�Eq�p�Z�/)oa����j�0�h���A�:�q�V�����^K�� �F��|ָT��M��6/�x�Bڼ�if��������ύ��U�3����U�2�������1<j���>Q +���,+޺���	ﱐB�Nq�|6x݆������&�p!����bFX^Ic>��7��ʖ.��z����^/rW���	9�y�h�����o����DT�غ��\u�Ƕ.����n�'Uj}}��(	���ĊN��Al��
Z�}0����h=X�P�H[(M�
��������a�j��־�.�]�y�1�����iKے������gb�R%����0�P�q3��	Ρ����m	�Ҥ��]�������bɼON���s�=g�Q$��pĕ6���㰜ԄS_L��y����W	L¿��0�܅� ��|�:��~�;�M����P���^X�ڹcE[#*�L&�?�}����"p�"ɫ�Î�@��+�~K0�j%�9��-�1�����Ȫ@,C��ܬG<c�<oy��>�sCN�g+M��d}��?fw.H�����������t���2�q2tc�I�;�}[n�
3Pz���d2=��#�
"@�P���C��4�� ���4ʤ��+(���`×�b��O��V�6�hj��b~/vr9��ߥT�����\"Օ�P����O�I
XO�!��:]�Mb�G��ՂH66���ۦ�ȁ�9�!Ռ��5E�vPs�H��}(P6��?���.�L�d�6�kH�F��`�xw	0�ҿ�`�����}��&B�R�qv�%�d�rç�R[	"��k�o���g�7�ϳ@�ӎ����2�qJ�Ӧ���#�ˡ��S�j��Vq^�5�AD��v���x��W�_	M�X�����He`"^��H{3����:![�����M4�D/-/�Nl��f;��~S	���u�EO�`�K>��?�S�4F�	�G�:J.$2 �=���7��D$�b"�^!���@ɳg�����!ER
�G�kF��� 
9T���{�(?��jzR_��>Pjo�� ����>FM��Ǝ���f���s�ݫ�XҔj
��'��T����z�G��m�0�iud��U�4
rł_B#0����b��@h��2ؿ���V����4�������\%�·�(P"|�o⧰����(aHF�B�|xnL Wa�AI�V��6dWu�lQ����oOjɦ�%��;�e��q%ؙ��J#G����n�gZ\ �ǈv6L���:���~w��.-�9�<S��؈,�k�c�v ���^MFw,m�C��Hֆޛ�B�&�X���}�f���>��01��S��Г|[*�>�+0G׫)Z�S)�V�r����ϲ���y���1#�5SyLvQf6���҆��P&����t�M���HU��_�m���(E|���������w��z1���]i��b�:{9�P$)��n~�r�+�gǚ�֫�B��ӳ���K��iEN�� �+^5ptD�ԟk���6�B��Cn�8�"�O �y�4D�
�#a�%
!�(3=�s���гNE�q��ֿ�7�ِ��������/�'�ء�~y9��ިsh��A&$*ӄ�Q�Iޡ<[�8ҬƦ�/��<Ʌ`H�1�_���2��4��� wN���ޫ;9t������_��灑iyNT�SBx���"{c-"]}��כ�����	��6����5oyV�a����ݳ���w Ʒ2�������R����æ�~)�-ڇU�g�D�=i���c�E&U5����M�g��ìz������sķ�n<�Tc�c.Z X����1{Z]�}_���j\���n����U6���E�6�F�(�ج���'�\�T�Z�����m��}�?e�+eKK�<d�x8I4Ɔ�K����x��SK�7n�$��jOS�7��>���N)��Dȗ�����`�ktHO�8>jeĆy����=��<�ħ���޽�nn���2��@�Y��\e����Vu��]�� X��E�J�A��B�TZ�%���]��O��.���y��]��;8�%��TTwx/hZ�j�~��E���)(!�b�yK� 9!�
�M~�"1�V[Cj���A^�^ˈ�R���y�B�Jލ�������2�?!��t]�/�)��#O�p�v�0��T� �
*����u��sx%�yL�WOI_1+�p��#f/��(��:�^O����}���/}a|��^IT[���8EWnN_���*�hk�;��2=�bO;[���M��������������z�\w�a����Ί�U4��jv= ���;1��WF�����M�DL�О��N�bJP�t��cLxb��[Ì,`O�t"�;�
{3��#�gZв��a��rw0���U���W�O��3�����^�(�=�ʖ�a/�$�t���,�$��7?
��ŗ#�9q	���Z���f�R�D?��y~5��뇻5YOuħ3������|`@���j뮻fA�⣉���	]�\�s�.dV8��.��K��F;��t��-�2���y���a��=��I���X�tK�©�J����թ�`�B��}%��r�=n���G?bp��8}D���B��9;�8v�YVξ�.$� �2��>k}(C�t[,>��p*A+�/
�?�W=�ֈ������z��#t��o�]8��:[���킼�� ���*�����:�Y4���R{M*"k�+%��7*\?�r9��\d(������.� �l��|0HB����J�Y�v0ORDsg����O�ε�Ƭq/x�.2��g�|�j�r`� �?�i��8 K&H�����g��p#mi#���CU�H5�XySB8�_��k���2�/O�>o��xht˻�eL�����~�O��_y�����^vqM��Ǽl�
$~`��i�����lb�>=Lv�6��G3�1wV��[Aϟ�|�{[]��uGPb%�|O9'_0�L���'G�Bq,���,*��t���h�{o$�̍������b��<��)o^���|g	4�n� ��� ,|�D�m�c�{� ��Bh�Nϫ���Zz���@/j�~x�]/���&�׃Uc�?Va6�}�@~щ�=FY6$%I���%}E��#U��2�����*+<a��f&?�3'ک�e�qa�@����B�{n�	�6��^���5�C^�y�u&�y~��`��t�z`C�V}Y��T/��N�#C%���[g�S?vU,Rʖ�P<ʸ�!�,U�E�paɅk��x8r�d?⎎�1�WE���D��*Ȅ�d�ח��~��4�̦,|�`�oMT��Lf����ZK ���9�x ��
xN)�<P���ګ��_����?��DW�>�����:<�a���۝(��rI�� hs� K�^�QÇ�Te�� ������z���������7q��_�D<����"�2x����]��� LB�Ǖ� 	ؠ��r��f�8�c�g~�7(��]K��~Z7��$T9�,�ߞ��~��փ�$��(�:(Ȕa�_��HO4=���s��4���c�N���I�Xy��a��EIP2X���tC��g�̤�%�m�'�
'�� ��3����Ƀ������-e��'�d�0��E��u*�s�6�`� *O���jD�Վ2}U��?��߷%�2�L�:BĢ.�r^�b��TeWs�_�lg���4�M��ȓ
9>sxrx�\IsEv�QM^s]ˇĺ���p=Dv�vZ�����cۘ�ۙ�9����V*����n�*b�:������_�x��A�cp�q�K|��Y��̜mE�����ȑ	�q�[Rt�=�1ͩX���z,�ˏly����!VE������s`��ep��\NM1��;G�O�^N^BI\�����^6.��"�ȟ;���D���`RJ�"��V}�N�u�m��"�����AF,u);B�+i�ak��r�!$0{: 
JC�Ti��Ҡ/���r�d�2~;5˃��}b��#�6�GtY=��ﱯ���3�P�ZS~�&lD����:�JI������� r@��*L���L�Zx'�y��1Ӳx'^]�P�
�����w�}�by�<���� =�����[�ĉE�ۍ<�gߢʘ�p���6��(�bL���\$�u�Ʊ�	�5}Wq���L��>w��5�}��Zϱ,�[���r��꘲k\��8��d�9�����V�8gN��\��%�[�q�R�:/C�]ۈw��0x{.��A����!\Jz�?����쩍���r��j%Î��e����$����5���4�T'w��VD?:���p ���QD��������vj����ҋ`WUn�P�'�m�gI��\�3�k����I�mT�Ҿ�*�*p�S���={�. �}���1�"�̙3�Gy��F+���,���ނa!s�a� ���I����]��}�>��Ϸ~������������h�;w�[O0���P��)C��*�Fb�w\�����;G�|�����q�`��NU�\@p��k�V��j=��Sq���H�ȱ\~�j�V�؆�hq5�z�Ҟ�����w��Y�uլ��u����k#�����J:�t�=�}�Ҥ�����7�K��i�Y 8P��UURܩ�1\���e4
s��P����Ť�pݎDW����SV�-�����߹���}��Ώ{�d���M�S�Y��	����v��� ��:�8h儀炸[(l*=��>�<vdT�1R���Ȕ�P6rd����[��[���:�f��o<�g�X�/ӰL<�. 7������^x�(�MX.�~���W,��tq����i��+��R0�p���g?��&7�w{#|>e�������o>2M4����
�;�5�5_|���>�!r��pE�8�t:�򉘰�>��n������X��t�RV_�#�U-��~�����>�u�v)']��Ȟ˾x�������^{�B�\0�` ��#c�fXL@�3���Y��RWKʦp��
;X��0��3�0)b2��nE;��D���W;�v�u�N���U��B��A�ρ �C�yQm���
�L&:g8;��mՕm��ώ�/ ��jB��$��0�퓎�>3o����L"�q��y晢M�Ɋ�mP��F����D��+z%R=�>�6�1�=~8!=�4�!"����3?�3]6����w��C ��hO�F�{ ���6�-�Q����-����o~�xO���-�+g"�����_���]�Yg.�Pb:�.�K	�x�����{���1�A��Hk���t�	����B����/���%ꋔx�1wz��"O�̃���ra�h�q\pq��5��;�c�g�����x�7��_� \�{����E<뮪zıM�N�\j5��o ^z�n�����|�:�ä��fK_Bt(Ln�UWcu���^�$��)B|�t�N��W�ʦi���ٙ;)�9I���^Y��� ��s"E7���y`b� S�+���s��g�����G�
2��G�������ԋ��gp�	����G�T�lW�������/���կ9ʇ�)�"�����-�~��_�eH绅<�����=�g���4y��Pr�������H����H�q C�f�E�¸7����q���@��v/����c�X�}T�ilP�<ϝ*W����w_�t�,u1J�� OA���8T'�hqi���hm���t�uf,#�I�d_��&lou0�_.��c*�	H�}��m�� (�@t����د��.�[I��J��iA� �; ��A���q���L��O��: �`�I6��rUݎ�/.UL���
V���,�12T�Ⱥ�)[u��ީrރR��?��ƺ�/wo޹]t`��l#�L�K���H����ڍ��Q��X�<]�-�������jy�9�$��2�{߮hP_ڳ��®�����������E����>y��� �B��{�{�I��\��2ڦd����!����~��=��hwIFZ�&: n���:\͝�9��}ÿ����U�q����Gh3G�M n�sۚ6��©
��1�n-x
:��.b����A�,mϜ�ȋ�p��4Iᘣ��w�}��D�+�������;�h^�<�8_4h� ��@���B��\O��-..~1���ӵM��; �
���4�=�^�_O?'�.���#юVG���P��� 4果̴�G���LZθU�s����+�(�N*��T�^~gc[��bP�S&0yP��8��b��~��~T�i�Cga˞U����3BY8QU�T�(۠�|�Dh�!��?���8 �9'd�zD��؝��#�|px2�d����t��ꔁ�ɨ���;�} �F�G}��# ���7��� A����6��
�|A�t:&�����C��_<7ƣ���ݩ�U�LW��:J�%pul��AK�/F�w�E��t�s�z�d��u�u"�����3H;�.���������?�T���'��V���4���4_��ɓ��#�� ^z����{/���i"�_����/����A�ů�ư���Eg@�$�c`$4���l��`z}@�z+舂~���Ǩ������:9)���J��8&u�����B#o\u]������:`�y�*QV2c:p�`��I������mPGL�(��6��� ��v�Gm���U�vWQ{C��<�E���W�����)�(�=�vi����TWQ|���I�ne�9N(ۣ��hX5q����=^q����;A�L���N::�F���[����Y%O���]��t.>^݉w��+������4��Ƿ����p��8�� ��޴�D~�FN�Yk\�G�Ǻ�����_�����v���s)��{i1�w�O���ٳgϵ�c�� $�
^N�+��<�^�C����Ar�rt����K��3�	��Q&��DK[4�����> ����p:)+���v�*;Dx���AS��ꪓ��I1�00a�أ&ڂ�=�mI�ę&�nF*�vԁ����V��ȇjZg3#��!8�
�w��m��D���4 �����=`"y���φ�7U{�jE�#�*����� >k�;�G�#C�z��?����/'<�hNXt�೦c�����E�O_�q��c����x'�r�"JU�[������9�8�{�z p�W����i�*����2��}���o}A�2a�S�ȑ�&�K��F:�z�C��Oi'Sҙ��0 _����Cŉ�ס��䵚��j�~%=�4���~3��<4�$댑z����<�u�ݨ��_y�����{���k�s ��S}o������47;-<�8u�Թ�.�����F���J����_�u��A'z�sA�@�E����1&H�d��Ӂ��y���B= �6C�O��I���|Άhߧ��3TgG5?�����JmC�	�BL|��@Cp��T �>U��m�2�c���� ��# ���ؒl��Ӳ��Ȝ�nd�Q�,�Ohá��l�pT�σ=d
�(��~�w�0Q�ڍ����N���� ii�{� �5Yk0v��ַ��hi� ���h��~���GA�����^�(\w?K@��H�<��\��h_�_�jWP�Z����̽/	�Ir���A��إ�*���e����m��ȣ8P�w:"%YI��si���;�F�G�4�L�6=�ƽ�)�t�f *��
>)��ԏWR����4>]Nc��tn&]��~<���D:w(�'�- ]�M��
��jv>����_��.�K� ��#=곔�A�n�za���������S_����^l5rWȾxIn��G酾���;�ot(�Y���):����U񑁢�!�BC` �@[2|TM�zz�\M�7���e��Q=V}U�k��KqF�)|�a�4�fz�&   A}i�V�!gt?Z-�̸U���b�(���:�%�c��������́�N	mlh�C�+�2[����kŶc���a�������/}�K�3�U�����34
�~����jP�N�% ONƴ���3�+�'ì O8���?�C� �?�AQ>����̙3��d-Q����Rؠ��3�5�:�:�E:�q,p'���I�����8�h~�1)Z �lm'��_���\���e��J]�'�W�=�N��Ki�gϞ�o�O��%���wFN�:u(����'�Sڢ�0���Y����V��t--�FR��x��Dz?�rF�ܥwd���xz�E>� ������{DpW�O���ͿHI����4��cIi�`��j䮓}7z��}�wޚ��;�&�3�tOQ�� `Ȃp����n�zL�
&!e<����0��cu��NΝ|@��ˍ�u���E餠1�t �U;�ա��;������;����:K�դ�7@0�M�o�e�d��0t��KP��y� e0�"@��s��!,�I�'�:6�|7�a�@nۆw��r���y|�Qw��pf��� ���p?�>�$�"+��������:�G{)�J�O��O,0 �`+��)�Ă���?�S?U�\2_�:���~�]������|5������]��d����f�6Vt:q@��.ȴ����H�Q^�'�����m� ��C�����-S�YD��ˎ�W��J������Cuv�y?���S������������^k5�HF����I�4�};M|�O�8�5&�PǞI(�hb��A� `$�GVO�%��8AF*����W�\�}l��Ț�� �+v���EnRax��P! �G�az��e�!"��V6�G��qe�/�D�?ՠd�\M��N�6��=J	�h��PW�H�n4Q�ǐip-��0!�N�Ϗ�4�w�}���{��gΜ)v�x���{B�@�&Q5�s?�s��:����c��5<��=�:r����'�0f��M���}��;�D�I���q��<�(�^��/� ����i��E}u��/Y;x޶�g�����O�k7�v5��/�����4>��G�V0O�@8�br��`�$�]E�� �	��%�+3�d{�Vc��<eʐ���t W�G�0?��V����i�>�p����������0�he^u�'#J��烉��H�B�P'Nz�}��Aa>�!<WL�j����ީ	C�1����p�:����s��O��Q���, �������wZ 3�-v���%M������ܮi � ��'~��e������`n��-���dж��F�B/E��5?}>��Q;Z�#\,�kZ�3��q�t,�#��L�]0`���/��&J��sl�>?�NQ��X�����������n	����Lj�ҽ^K��i�il��ٗ /u�ki�|=.���N��r�� E0���ʖ���
UL� 8���d�[�P5�N>�G���|��z��^��Җ�A�U@E������;Q�3>h'z�Q"k��j���J� ;�r䞗?[M��' �x�y��8�@�t��p;-,��x"�âpr�< 
�㸖f����	x��P��n�ܹsų�ze��o�fw7�A�I@ĸ{
��~©����8���P_�~�3���Q�p�~�;(�+Q�����g���?�:,Ȯ�]���:]��F��X�.n�~���=7���2F0bP�t0�|�3��ri��±Nm��>Ҏ��幜���.i���ٗ �Ʒ��R��O��a�-c���@��+�x�;)�ʌ�&ƃ��f>� B`ʲr����u�T��΁�y�(k��
������^��H�	&��?�s�����*?��~f=h��\a#�c~�i��xtl���v��'zzBr�����c K H�+���<O��-|^2�*�'�x�������uH�]Wp��g��u!#�8k rj�� � px����NP��m��Km�/��.^���:'x�>�KC���TC�����erp`��?gֵ�FZ�i;E�0�Ư�k�x�7�[9ֵ�1�v�U���΢������[��R��F�@�3���&�'/]���i���!;�4���"�:���	$9�a@�zM�8Dt0U��R���s�h��n��U���
Q��kN(�o�^	�O'N�h/n}�6�`�6� ����m�<W�N:���?�yaB���  <E��v-w'�:� �t�D��ۿ���{0��G0Fd?���Y��!�ZU�l  �[�q�=�;(��.zmD�}�q�z�*��g�6��x�8^m�v�o2�C�`qB�z�� V�M��ݥv��u���U���l�\[iy�O۔isy���(���^f�X�5��sQ���5�����]x9��w[�4�G�o^�0����Jp>H�����E<�P3ѻV�_u��O���ɘ'e�8��j��z���`Ǻ8�c�Z���*�3� O�ufZ�+�f��ʋ�����FЧ���I���r��9��eO�Fdv���l�L�Di<<�Zl'D�%U� D��������@;o���~���� h�����'����6���>4����j��k���@~ܙ[�16Ž���q��]Tv.��9'�<���A�z��}C=�^e�A�zG�����}�������G���©��*���E�\���2��<"�UV���H�R�����p����|�41I��bz?�������5�g�o$u X|#��G�cLFd00r��N��u�(Ѥ����u`'�QU��O�-K�+����7�8h`>1��T7t)�Ķ� ��UQ���ؑ}C]0��8�~`z�f���6�����<ܐ�L���ئ��G�����&s<^M@�� Rt�@�������h#,VPB��8���G3�"@�t�U�r�jD�P�?:  4�C�%��b�l��B�k���iP�s�@�����v۷�(xBہ)Ż�"��%��Ԏ.b�ܳ��*bO� ,��+|���ҳ������B���-��]Ɂ;�wZt܇�A��};���ұ����=�}�\:z����|��_N��$�:'kL�0�m�����P������K���"����,G|�DJPp��p0z<�r�̐�S�ُt�MV����4`��<V�c><�-��� ���?m�	���+����+W�TwLr�ͅ/�V��s;F�
����I��5d	õD �e��2!H"���
�k50����O��O��^z���$�j��� �P�� ��M���l�G��F`��Q� �z�|wT	�gL��mE�K�|1���g?��ʃck��8Uֺ #;�gp���}��7U�j#�!e����\�����1^����ŝ_��۪ڌ �����o@]���Ei)��[������s�=|hW�wD�.�9��7��W�"�Q�6����^��.�N�\�@�O�I2���`."�Z�๔���nz<b�~z���:V���[�y}ԋ�e���h��Hw#[�h��M*d�x1$ 	 ]4IVI���A����D@ �t��G&82e;"+��7ʆ�/��/����`��8 ����>������*� ?x�������C_A�HKO��R���e=(
�tw65'ȱ|��E`���sT���K�@M$zLA��D{�:H�yzM�G��\x�DLb�O����o����ksR��(�k@vB�6�'_4���Ѕ4�=��]��mdOe_��y���V�_�x����ElO��C�&�heX��Ǣ�� [5�3@V�E
J�n���y�	Ru�(����nme-�}]���)\K���3X<z$����C�8�u�������l���]�: d��U�S�N�(�v� f���}`q��E-�&nA��ܨ3X�_��_)���о��L4� i'Y���>���#�0��T���7ʓ�=v+��c��[�V���~
� 
�4����Q:?��UU�Y_�O�x��ˀf�F�{��y�v䱍��1���ڬ��(-���ܕV#���k���>O�I�N�줯��XyP�AAB� T�{;�G4x�>9�J!*�i6���-��cw�nmi7��JVA��;gy�q ��3 
 �=7�5m���<�������cw {��h4�*l#��s`���&2�1�G�?y�Pw�Z�O,&"��_��_(�3�é�yEc�ᯇ����}o��A5/�
��w���d�p�*Wơc�qޣ���vF��ޫ�S��>���W�
��*�)[ F߫+�_F��=T�-c�� �h��L��3�
R�Fk�k��A�w�id�e��Թ������=��[���1���Ѡv���}N�I ����Ii<|K�w0�c��S��u ����*��VŪ�*4gE#�G�ȉOA��=�B#{-�w��*�=��F ^�LiH��T{b���S5�����_���ZU��(m�|��B�
{=0s0�4W�w F]�ӕl�T��H��S��vx|�-͘��#�c�
 �-��t1�{`�BaWz�Se�� �����)@�;������ko_DㄲO�=�KM���]7�ˠ��(�	Q�����~���8�ŧS���j��=�}� ���o�ғi��c���p��9�U��t��� ������I�2|�'������У|�/�˼�ֻ�`n���;�ǉFm�
�:��Zw��K�2Qb�i0f��G `�8�k̴��Lh�g�ی�3
���裏a7G��@�b&c�N�/4h/��%��Z7��n�U�2u�����o@����„����:�g��/�%���hY?g��E�z��eu^|y~��sj��k�@��/��+�j���^V���#|��tQuYz�^]\\�NJ��H#{,��K���i��jZ��f�9C�
>&B�H�@ZNt�Q`�6a�W���SKU�Gˊ@�zq�ʖ�ox��z늴�q�����n��S�C�m����a4�l�@���28�#WV$���~
`���w����!`��U��>��x�u���)��4��s��\��+Օ$��G�ú��R�ݣ��'�
�[��$��"��#p��7�膒A�>R����;. ܖΝ<��E�V�SU��H��*x���8=V�F���iʮ��e��{�\.MT���Ҕ��]a^�D�>���ؙ�glM�lZ���j��; ��K�j5M���/��gR��d�^���q�*��0�鳾[`ϧn]���ã����g��^��n~�^�W�C'G��4���,U��#���wƎ#�#��VZl�e��E@QA$�1�C`G�_7�g�:U�����ؐ�����1�� �iNXoz,���ڕ{�"�ta asT��3u�����}�4nת���Xv�F���c���*U��2 �;��Dd��i�ȝ w�.�t<Sͅ��N;���Sǎk�+�#rO <H�D��������4���q5�11ap����	���|Q��T��w�u��N�e{m�
��+^�UCD>�8������1�!qRe�Y���� �!Y�6d�C��
�Z���������;}>���@�z��)Aw*8~�xW��m�������M�p	�؞z/ul'�a$�	Q�1��wO'"�g9�~
}a���ρ�T֘���'��5~�9б�v�x�.�h����I��$X���{NQ;��U����L���U�<��ͩD���ڲk��sRL]"[ڨ~����N���h����Ϩ���]*����x��]N��LLL�Ky�l5���{����K_K���%u��4�M`�=�{b��ޏ�DVG��$'���j�W���*�(�,�Y������@x-�CoSW뀩�A�`T�1y�RG�Ͷ���%�԰:T��]���U�N�;%Ue\+聨�[������6r
p���v oxO���v�;`�J�6��MU�5�jWcm9��~ޞC3��i�U�H���w��)uX� �յ,m�ryE�*gU��}�N^UhU���9N鼐�ͥ�n~gvv��m��=� �>��i"�^�����㩃�1A�x_`?r��s�P��):*��V�z�~�M,�k�M�	����������Hk�����e�7��ѾD��վ�ێL�4>h��:+ �gP����H�|`k*��7�]�*C�tB ��n���� =��_�ǽ�$e\�="s�y(�V�E��	����n��1�hcI6��z���}��F&��{O;hQ�1�?y�:mc��<U �պ<��(�:�\t]�Ց����\^~���U�s�3��#�^w�G���s�c�=G컧N�8�x�6r��x���^�t�?��?�	e2M(g�1B��W^��v�Z4y�1xnk�<��v����
>9 E��n�D���T	�S�8>�.�s���0�s7��N
0r�֙�T���9Kȿe��$�5��~�"�������Ve\��6X�����Hn��ylC��yU�F�C�]�ɍ`��m�x3�6�ۿў����阮A�����4��5dP�wW�E���ھe��e��:�y��c�^����Z(x~�΂+j]��l�i[�탺�5��%~�kA8�I���=���W��ۭF�CrO<����ŷ�z����]�v������������e�A�;�2x�ݯQP7�ʺLt�g��I��`�b�L�9Wâ�� �+���-ǆx�Zw��Y֪���l��H�!A �<�*#�WRƐx:�;��:��9���&�~���|���w���!
���*�c���g�9�-X�U<o�\G F�:ʫN�u�⌚�o�<� ��U�ZFu�կ�n;5.�	�q~g�ø#��
�3��s�݉������}�j��;(���<�����u����/]������iB#H�@V��ɭ���`h�9�h�TВ�hB�z�$��埜�Z��� H KFW��d�f�q{[9��{�*��l�T�W��Qz�l�7�(���P�=�}����="=Su3�~����<z���nR&�P�	��&ۖ���9|�fx���TpHp猶�xjX,"�![qc|��9@�-�C�]��l�;]�&~M�^�3�D�瀙;yD�G�����|�Ų�u��xs�Cs���>�g;��zzg������ɓ'o�i��=	� ���۩��݋/�xczz��L��(u������#��#(��I�
���~%�B��5��`^6'�����f�B�>Km�4���?EU���8�s0�!K궓O����� xȏ���ߕ�� ��x���+��(w���q�lpq�/2���6t�#Wc�����9|�hx �����Di�<�o�@O`U?�~T~�KTۤL�w?W~t��D�\�w�v���+��R����LO���.J�wN<���k�o|�j��;,�,���'	l|'}�O��Y+��!e /7�Dߣ�:)��ګ3PF�NeY����	�y+���)�=�\k�U}����FАc�t`���ʎsP�Cŝ#�G0�oOU�u�ߎT-<�ue=2ȼr�/n����{��4(�yu�`�9�Ctb�ŁH�
!���0=���k�`���'�S��@B���G喥ɕ��� �ˣ���u��>w���u�x ����/Ly��7tBn-�w�Yx�;v�ٹ��;.�4�Ko��߾<??�n�~+u�����5��X_+jD
��n-�+@R�j\��DP���8xӁ^��"g��1-A��N�^���X����]k�usi���nu=I5^���m��W�'�2f�'~�:��1�$1�C��lTC�*C�jK���j��d#��A�b}>󻫈h@�G� : �0 X���{�`�Poܷ���}�P�����/���N�
��=���d�v � �|�]��kޟ��@���|�.�=�ϕQ��,;�{��~��I�]Sv�E�?������m]����"=�J�O�1����wZ�4r�=�  v���U��c�c�Iə$��3	Dp4�����������윳��R�s
�h0m� EP�����8��9�k���E^��ʘ����Mg	|�j��#��=�J��`{��1���Z���X��?l��$� �φ�\"= (�Ó�/U�T�r`����
�"��.�D�T�7������{U�� �n�{�u�_�xU_��}L����U��/"�|'$�	�i���v>S]S@��E��)-/�ܸ M��{�|��ƅ&4J#w��� /M&��$�Z!KPE)ݮ�Bg�T"0Q����ڎ鄥�2��+�26/w��'����9x�h{G�o�����o޼�UgPm���Rr���C�����O�e�MU���������;@�$��������F �p(�'����3U+3��܉��D�+U�t|�d�i'��� O?ڎ~N��m'�=b����9s�6֝���I]�W�ڨ\ϣhV�%���cÝ;֯x�E�N�I���<�A%íNa�q'z�?J��W�<�V��F������Ǘ���Υ�w�	<s�I%b�����
�xM�7Ze:3�y�]��=�$�^��U�Re��T�n��v� <h�3W;+P0�g����: /|Q�y[�3��R�6��{&�` _�ct�`z���4y`�g �`��}�@��Ő.�9`u�w���,L�s�mY�\m�?��m� NU�����gT}��W�]��*pW&U�.'e�k@����n -Jnl���;^�~�./�N��O�w\�F�p��(�`�+��bZ4=u����F�K�x�s�|��_�8==}�󻇑p�PG����$��)���h�ȱe��
.5^�2&��F�� jhp��e��Y^��T�K�� �W�~Oz�����?�~&m�(�5��%'��VEl����0�6�4��G=5��)KG��:����: :�92tT/�);˼��)��� NA�����c�t����{޺@a�)۬^��s��C�W���{T$sy�y꼯U�#w�<V@��:�U����U��{���}��U�ò{)��|��������h5��]$�<�����z"7��H�V��1�r�D�̒�:)���`T�~�V�>��`�
Pu5�{�5���j����@���,��x^�:o�#&O�F��� X1�֩
PA�)�y��;��^��R�e ^N(��B<� �m��W�:��NVT�+맠����2��|V9����p�e���~�N����}P߁*���u� T�5��o�y{��e���+�ktm�rsi�߃�C9Ʃ�Y]�풮_J�}gff�k'O����H#w���&������ۺe�ꀾh������Q��N8�箧��[� ���zUK�����`���{� #��J7�2R(T�����e;r�U� $ N���ZXX�9bd?���377W0�8��8�ƪ�d oȇ ������ Y:�f�꽩����iZ��Ӳ"���i�;;M�����J�;� H�\����|Y}�4U[�8�,UmWU�(}��.�,�s;R��@��/d��ɍ�ѱ�|��|Z��s��o�i�.����j9M��d��:�P�`��y>��2V���2W��/���݇3,��:RVV�ӽ�;�n�k�FOQU3�:�]J4��F /�t���:���	Di��sh���M�a��� ����0$`�py��]��jV�tt� ��2贡,�~��n����ږ;�� 0r�^A��k�K��U6|����~��Ed�c���Hr����ߪ�e�G��ԃJ���AڷN}�sOڿ|+E�G͕i���~7�o4�w�܍r  <hO�8�A���;N���:qrb��	����� ��f�(�5� �x�f�^/�M%��8'ASVE30r����2B�¡l\�ޙ��:A}�k�����&R��= �N��@���	��P���xZ�q�*��|�� r}��G�gC�}��?^C/Y�O�8Q�,��|	&��"��L���"/W��U��`I��w-����d�u��יD�aLI|�	�T��{&��b�j��X�cUm�W&u�A�S��.(4/M������.�.^�c���ՕBۀ���	��y�́��F�/޻���4�4�]#w��7??kjj����������X4�D�U�8Pa��ʍ'�&5���z��W�06ATn��vgG�{������k�+�q�Z>�^�޵�6s�em����0o�'�8	�O��S� yٰ֠K��QuͶa>Pߺ�T�1l�ίu V��l��\W�����ʎ�n���s.;�/`����s~�:26TI�<w��AE�`]��/�)�(�yL�e��|���-,���ٳMܻF�J9 �K���洛�-��(u�{>{:,
Px<��嵝���(���]�D�	s���2U�}�ix��:v�Xkl�p�V]�
���N��!��uD�U��vb,��vB������j�<M��t�7��2L�aR4 2�?�t��m��J���m�ɯ
�y�����:�M��K�E����F�R�{��5ȱ���s~��ͺ�p'��Ϯ_QP��[ݡ��������&���\��qnn��{��]+�=��C��<��'	�Ԋ��a� �����T�jC4��_��'</���P�AU��g�u�}'Z�N�l}���+/��ϋ=�:t�4-[,��l��!~�l�A�<pP� �Ֆ�Չ��쩊���XA&������y]��8Sn���~��\��ι�]�Zdyj�&U�wdj���~��l'o�� ҝ(s'��M/�� 5�0�x�Q}tl��.���|ez�蓋��W[�4r�ʁ x�î�_�� �MN~��������9h�/_�El��r)�Z'W�������( �X��z��+�	;�amĻ���(<NoܸU8����}������&�}�>�(Pr��r�@�P���v �:���G=��]���2�O���Y��i��x.Hq��v����r�U|�Ջ�"�ҽ�s ��������cK���ﵖUv�nlrt�"��ҺJ7'j�i������ɉ���gϼ�j���X�����_I�k>���:��O
��YGEK ���R5A��׻���Yv�}�q[��Z��Zة�ݾ���vb����ڔ�b�t��O���_�n��Y��[����i����W���Vgy�R;;��*�*������Q��>s96P���\�w��E���y����.e}�N9;aBЯ��m�`,Vw���7��������ݨN�1��������9��j���X�����5;;{��0(k��ݜ�}�X6xD*E/�� �y4a뱜*Z��|!1�hG��*���9��t6 P��h��ꔠL�ۘE���e�	�� jڳg��6/���ם!x��L�"b��-����E�r��2Ne[�������ޫ�'��h?�*��� \h��4�T]?h�U��� n��}���v�����r�q5�������٩i�7��� �#G�,'������j���, $b<�e{tb˩H5�v��:*]?�9	�x���&���xDo���b �������v mll�H����	�'x)9ۺ����]U��iO:Fp�GL:�i	L�Dw��=((eyd\D C�H��r��ȃ�90Wu����OU ��z/��>_W���.�\=�28���a�������S�� D{���5l|����u���N�[^YY�n�znn�ْ��}!�%Y���� u�[iҞ�j�2&g���jE�p�K�~g|.��u��`�a�6�e�4��ɑ+QU�E�>
:x�
.6��l���p@����7j��;:�\,��	�J4��۪�cU�q�zÀD��{2Gmc,5��V��������'�vt����e�ɿ;�U����;����@��ɼ��&jW=� (W����@���o���N@>1����ܪz��T-���AI�D��N��Ƒ�<����^���6��f<K\⋘�SKZ�y������7z�r�*`��{���w.-h�MNN��ѣG�u�ĉ�F�r` �������Թ4q߼u��$'e�4�I��<7PA�f���\� *��*Wf����u=C[��M�r���b�U�V���E�FG�3�ft�������nnh�B0x z�T���o4��Z]e@T��n��NI��CB�a�$?D�����jj�n������y�^{���=���^�5'k��%l�6�Vj���@AK�=)w+x�0D��5��k��B�,Qz`3��)�Xz��=r2vM��Jȧ%�V�3�hW�p�f|:�d6R�F(3��܀_"����*���k�����`��g�cdMMM)�����_;�?�],XV	b̊Y�z��D�X�x�2��7d��a��ي�76����g3_��e/�7Y���Bj�4��#=<��M�ڲ��>�:*��C�fꏄ{�LL0�����"~TƊ��+���[����o�`��<lR�B~��y���� ~���ES<��o�@�Ԏ��˪��`aRpF����a�t��D.ș���*���������b^��Y����ǆ?HߦN��ڠ��F�0�ǑX��p�O�=�N	�@���|%]A9�o�m�G�A���n=/����C��D,A"���K1&�zTY�!3d�p��QK%JÑir�n��R�<a�+�h�Cf\�I�0y���Kme�+���ʮ�ȧE��O�j{��AQ�f�P2"���K=]\]����A7w�^�KV^�OE�񪏰����L1��g�v���aJ���*Y����,�Y���:�8�|.���`2 ��N�(2����Խ�Q+�{v�c����MF���U+�t����[�N�af���A�&a�Ջ�0 "���Ԩ�e��`�x�j�X�ʑ
� ��B��ko�>;�ێrY��r��~y}0�K[D�=�Č������x��������!-����8֞5�@e��CTG���XvȈ;�[�(U���f���[�<n�����5&0a� bcc�ߞ�}�ɂ-�cE�&���2�mi�o�x=�P���	If�qN���V&pw� Bz,��{O&\����?�ə�*`�B,ْ��Y1.��%�$��B0?Vl��w5o|Z��w�<���� 0R*Փ�MY�������By��e�o
�R��b�E��q�̱2�@Cֹg%{���tM.Y�A�@\捞���-���f�)My�¢�g�{0i��b�� �'�}MD�-q�3��"�Z�V�k���xc��}��5=���x���Q�3Q��Z��8s�NԨh���<!��s�UU��ȟ��q�&Q�Ӫ�,���W,��A}".f[��ɵL���s���s6�~9���*�_n��{���|��f��\�ڇ3�^8��!��3�>w��C�;�& p��9G_���.�x[!�
�8H��a�}p��:�na��`Ku?2]��>Uh-�{������8��7ڤ)/��L�Uq#��'p����( 
�Z2}o�@��X&��{U��|�u��e��W]R*j���1x9��,|�si��1HFy�r'�&�%�$�QѴҶ����nߨ�.�ld*��i2|%�ڨ�}�٫4
.9���w���R_��p�Zj.����p¨sR0q����k��rk�C��xmX��	+Oͺ� vj����Ӯ�`�������4���@>���}h&N�<֘���i&}(�K���	Qg��+ݦŌX���Ju����huT�y	�6)����
�f��Ļ�o�>5���)K��OR5I.""��z��fB�\G��cE6��1=7��>��>����D���)�F9Q����������E�O�G`H>�2�9��Mm�䭭Ԇ��� 0$dY�C�F�a�n��Դ�L��ߍ<u�'��b�Q|�ד��s�e���۰x���^hmnUh�`yn�
��>؀�p�ϻ���߰�%2x�5`X������4R�y��5� ��"�g������A?^N4���uW}n��̦��D��f!*@� ������6�F(�}�-���ÇNd/���t�
Jo�)Z�z���f�j�m�5�E�ܔ���7s�>"��'�G��ű�~���7���@(��i��1\�R��A��[ɗ�IF�كQY�<����q7�[0�|O�x��$N��PsݘsF�>Saߋ�T�0R��&�����������@oX����^?�Dr[D���Y6�?���w[������qb�\߫l�d�%��^{N�$C�i�.�^{Iax3řd�h�i"��B7��g�b�9B��@��{ҮmS/s1`��ܖu��n�;��"��u�ʫ\�ʹg�Q>Rٶ {\��ݬ�}k�=�0������E�ؚv�\�y�l����(1!��
� �U	���79�`nH�����jjj꺗�>�X���&GO`rP������v�0t<"f�%x�s��պf�'(?"�<�t�^�{v"�PQM#�B\ ��"��d(�Vc�'����[T|�,tj���Q�ߗ{����#�_e�r�x�ղ��"�ߣ���Eq�[Kt���{q��I����/�]�w/ې�z�A~�#�����_�lL��>}qr:��	����E����zj ����a�̸e�D�F�G�`OST,Lq�����Iܞ��<k#�H��k,�-P���� ���o\���Ӥ�~�V|���G�+���i�~�0
�Ã}�Ak���u�#���\6�Y���d�N��h+Йԟ�B���,�=gB5�v��XW�Av� ���-���^0M��Ҽ�ܵ��1`[�rRἕ�_bf�rT�&n�Hߥ�Lˠz���v�[7&��Pu�gf�� ���p*������:���4P0��<���{�ԥH�n��G����
Jɂch��$i�)6�V80����"�ǈ$9
6?@=���]�.qB�縤�I����m�7X|��5q�x 1�n�$Du��"On�
�3+��t������3��,�$~�t�F�"Fko����{��ɪ�g�`�mRGҷ����zz�gAc㙁v��[�g�����t���n��C��;I)���>�\?�3��P�m�窣�rD�C�lԦ+ǥ'1W�X;�ɻw��T�8ήa��m��	���qUh��#._�^7��'��+�#\5˔������wfF��O��*0>,��������1 �ɴ�E��ٵ'&��oe�)��+��H�3�5�*4n䪎L�TT����֮�i�.���Q]FF�0��������a z��Q`rrrN����RzI�i�M¸^������J�a��P��К�Q��~y���~K�B&�ͥ@xI@@���y�������7��$��VX1�~����/�.
�hp$DYk��v$�S����e\��|(�GZ�!�DH���xIe3�ih�!�&�[�S>�gB�L�n�8H�e��vm�q�w��v������I~�懞��BV��J����\��"h~�b�����>��v��\N�A�I��~���`���~�I�|U^*��#�],uf� �~9�j#�ؓ-,g�D~�����tp�#�1�����D��n��պ�Ny4:��R:�t����[q�#$��o���w��l�.��Ap��?�
�,�*�H�����f��L[�j����]�Y��[c�˚����2_����K:��|��yY�ʊ�8k%�+� ,㗌|tn4R;ڪךks�W>�2��i24�7]�Rډ�F�̠@���U�*���O�:`?j\��}�4E��)[���s��ڠwr]|I/j֍9�j��3͢ʺ��$"
Z�&m�a��F:�8���)�t�2LŁ��ht�%�#z�M�kx4�� E��2.�Wfn��$+�$$��H�w�F���V9�RO���mG�C+ʥi\��m��j3�wm��$�����Z�U �4�A���`�	_[J��S���䤻�"ˢ�@k��i@ǉ�N���� ���۵�xY�6��6 f���ӷ�z�.m�$�.ᬬ(��L�n���ɉ\v�Wl��c��F�t�n��`D6�8�ڨ�o,�g��P�_g��v���WkJX�`�u�Jo%�	�םH/��j~��vm�r4J4�
�	v��|*�65ƈ��^Ss��N�4=�.7� ����I��� V.(G�AB�lB����!�Eo̗�T5�}��Eȹzg�d ����4�E�y�̪��XEEA����]���+�
M(��]G�C:�����E��ZQV��"XM�[a����䎟�ֈ��l�9�D��;7+���~��S�I����~qƅ��_���t��P�༵y|X��~M�����Og�3��EjO`�CsX����<��ٽ��BIB�w�[��E�����}SWJ�'�5����&Ǻ��@	/��{ͥT�,S��wg��m4`7Q�Ƨ�ِbJ���9�`'�}�Д��f,5*���I@w�6=���a�)���>�׺�URw�����b͉	j"�b���o���TG0
e���%N�9�R�����&ߗ�&6�~x"��Ɇ^��!�m��
&YI�ۻ�X�J�ڏV�3&b�Xoe��}.:���Z[[��W������+��ԡ��㱠b���5x��Ը��]��?c���BE�E%���$"����O�%�{}ϳ<Ջg�8=��u$��^ �u���b�?��'7����L��@w�p��m<8�X8+a��wTo�!M&�RAz�X���WSR!7N�P�J�k�c����<s�NB���_�����o�^a-bW��\�-|gg�۷�'������jv辛�k��-#8��f�X��;=�3\ݝM��ddf>��;�8m�,R���F!��F���/�oqJ���Q ڐE���$�ӓ�S�O�G�!���EN"z^X5������īu�Z�k��+���V{��D�������6/3=�9�e�5�>-h�E�}R5u}��=��!E�O�t�M�C�Z��I\�Pk�4��}Xܽ[�ރς����?�M.�9���b�9�nV��::V��K9�#>�m�"H�v�Vș�����tPMu���K�źA�Bp*F0T�&I5$u�>f)� ��|� ��;y[�>:s�o�)"}=��]��=
���=�T-�ް���G�Ռ�6�P���[��qC5�(�p�aCo,��w�k'& h�3�|yW��/j�z��J�aq��GR~Ա��L���4�c����x��񹸽N�M���eKw����U�}vM���ˏ��s.k������?���T֪�mfԟ���&G�-�O�L��c��6@��}�:���ňԐ0]l��*-
M���p']g�#�-F��T�� ��1��R�ڪ(�*i2�v,Mg3��A�jw�/+uٍ݇�g�al�Ik(Ŏ0��j2>���� \4��LH���.>�K\�?�����0)���h��Vϋ�z���� ��g[m����K����T���)�;:���[ܪҮ4��/L�ʨ��.&q✊ϩ`��^��]9�bWUK&�&�� ^w�[Zy	�#��?n�SA1�^���x�>�nD?ե�f����q��lVD-�>��6s"9t�}�	-�8٘�8T�C9E�y�먗,�V�B��<^G-F�.!�tV�jh��	Z��w��bue7�U����`3b�(�r-5e��~���d7��`��>����3��;n$'��6���Y�]Fѐ;�W-|D�?!KNO��k��+�r�0�����|1.a�c��_�	�QVw1BO�J/���:;FR#nՂ�?P�ì�{9d5���K�Y��u�݇�$p�?�naX�d·�~�U�G�@j6-}��Ȼr�Q����p�A���v�W��3��c���՟9��/a�?F_��{ٻf�x.P�k������7/Yl���k����m��g����/��)����u���$��h�����_]��g7h�� �zO���e F4(޴
k-���Ȏ �{�c�N@�oE���Q/w=d u_~Y��	�9��W�L��M�X^-3�m6����B��e%'����Lf�ӷƓ<����[�0�[݊�i���D�"����y�%|w������ge)ρ�a��)�1�����e8����~��g�'�>�O��W�4wU���O+��g�a�ꐺg!%Tp����}n̑�jK
I�1<z�'6$�o��]�"�C���|u��� E�"�j�{{_jHA2v�JLm��U����v�X���m�*yp�B�qǱ�l�?N;�T³f�y�kP,��Sד���ۖ�d_G�:X��Ol���"|��=7�x%F��R����HAz~:@��#�t���~>=��?�m���O�yr\3H�v�t���6(���7�ȿ~�������^rYĚoF�c�ߴT���a���P&ܷ�
B��ƥ�PJ��ث�8R�>팗��ȡ%g��Id�'���k3�]������m�Fm�����I^-9�}���6�����Nd�_�l�O��N����iH�{d n�St��;nj�����s߻��tt�:YE#:PlL�3FB�F�;Q*���J�L�w<r����p6�i����,���Z�����8���H��ƻ����95G�s�yE,&�?�|d�x�6hkn�jӧ"�-^N���aZ�
�Z�x|�~MǊ+!;�N('�
��+���Ƅ|�:Ν����G���ꬩ��#s.c#F�:6�����yy�O�>�hjjV����ip`R ���M�ii#��Ѵ�<5�?⨹�t{�3y�1��J��}�ͦ���\�v6\h>1aE721LVО�u ��y������ށ�.h2B�T�T�L��E�n'�څ�����W�K�чC�T�g�V��_4v�o&�]�n@�-x����6u=���kO���R�]�.s�?�f�4ek48�zm�i>��iXh�%�������C:c/v�]���|-�n׵?iii��lE���ܵu5������	/��p���Ф�~���������ܡ�C,�lv�U�rS��髙p��<��D�F'x|������9���W.�����Qy�:�}�)� ~�����u&n���Z��Y>�1I�i�s�'V^�����	u^�){H�o�{�w���]���Ҁ����AS���ǯZ�l�W_��r90c�W4�Q-1�\�8�@T~�{�ø�e�6}�`''[�Y���m����h��nn�O��t?v�����r%�������� �ERVS((�v� 9h,�b3����ۄ��m���^�c�V�hU0oiݬ0`��̎w��C�������]r����2ڽQU{�r����Q#��"{�^$� }��/���/�٣2k�&J���]B�к|T�u���qE	k�.e?@��s++��4u-��G
�MwvM��-Ъ1�~w�P�z���hY)�p?� ����➐�g#�P���0�_�����Q��շ	5�v�\���Ј�7�$��\���[JaN�蒘j=��;�0�9�_N���5�g�T=\'�ߴ-���B��ĕ���9Zѩ��&�nV�e�����Dn�4k�Р�4v����ev����-��6I_Fg:�D4yW�{�9Vh��/e���Ɵ�[���'��G���b��Q�ĽL�53�i�X��%��E>:8@KJJ�)<c��=��9�}����#u��"�@�%�ƶ���aC�lT.:�s��{���R.�+����K�xkI�^��g�et�@�N�6ae"eI��ly��������� ��U�8Xjf4,��pZ$������"�9���c�����H�Biu�Iߟ�2����y(�W��^�===}j�w\vTT�9~�}~������i:���W�Z������̤w�J�8�ⷡ5�7�����J��d}]�� an70��N��jQ%,��X�p��G>l�ɅW�3�'��f�,h����}$��&�Tk��`�X1Gص3��^˱Qo�\��p����R~�@��)���j�(�5քX���[��a���	�]�����!D1K��������A{3%��Y�uϞ3���@���A�%�U}6��V�8x�\�nX��p�'��'|��K��ڭ)!̹Gyߌ�Yf�fG��5�vP���:<�3{#�2hS4������~���%�*�9:>~鰫�qҨ���mln��l�M��v	��a��C^��=�(V�,�qK��n)�����ނ��kz(�w�������aǜa�8�T �ۛ���]	))D��2Q��Eud���7���f�/1�}v�3�P�Ϫ3|������h`���^�Oi�����s�Z5hg��vytU&c�����̺�tK���$� �=k|wOб���l2V}Y�V�n�Q�p��`5��K�c�R��o�C�Ǉ���!?���bϷфFu��2ړ_~O��GB�����I-,a���M*Eix���k����L�0�y��Ң
�E����	f"����:;Sn!�I���޷cii�����t�pv=�=88h�F,}8�·��zM��߄st�@;'��W]��[�i'*��^�b� |/����x)��w�[a\�_�'�ق�3ag���� �ݕJĒ��(5^���,�{�;�L�d��.��LT�)k��5X��G@"a�(E1+���U+�0S��D���ȁ'��{
O���,�~%�B���0>�1���A?�	y��;��ްo=�q�H�*�*�o"_<�v��aQ���%'�Ot��}� ���8L;�2�L�٣9Ŝ���}S�VJ`�%�WP���]�5HA�Id��j����0t!�ӖZg�J�zX6ʽG���8��~����a#6���=3�v�B�E]'�o�#�?؟�~8f��^^�W��U �r�B(�_�!��@�m���ݰ;V�_nfyU5�V�>Z�t'݁�h������`�^��2������`-��I]��A8�m���C~����'4~5�wu~����S�2]հu�AO�O�-a.^o����s��q�-�
]��H�Dz`<&���9�����M̀4�(C�=8VO��G-}l��SY����\�*��Z/�s���{Q��~���2���r�΁��%lY鿊���Q���6�����qr5��� Cq�*�	ټ��ҕ��X���M-^g��� ������эg�hO�
�/x	���W[�@��|�I���;�6[a(�^L�a��P�
[L�_0�/Q��s��l4q�)q�r(TzR�̘}ي�8�� 8X !�e� ����H]q=K�9���Q[�`R�F�8������D�}�, �})X�(�6�0P2��k�d�>+���`t�>"�34F���d�ߕ3Zy؄Mr�z�:�t"n��t��gᑌy��Xj� 7_�3��m�.^_���>B��e!w����wcc�⹏�b;,Ҡ'!:K)�Y�:s���J�h�qv�T�D��=4��i�c�L�@>䭖K/��8���%�3� �7�Tg�b���uȀQ:���`
֎ܡ�Q��Ԋ0�ͩ1B�`:�`��MX���e�^�-���VT��CJ��fӆ~!��Y�k�N�����I�C�R�Ъ�GV���|�&�|���۩�磉�����OC������`z0����cY�E�����"��Oɟ�vA�1��Pb4����Ց�f(7��d��\op.�
t�K���B|�wr�m�U��s�
T>�T�j7�M�Mh�Y�	�D�����q�*��3'eT��y~@ݚƗ�m��Fj�ޜ��M��Wm�jL���7.�°�hฬm����ֱ x;�i�����RP��S�����X��	����8���~}qOdr�sk�Л�75���[������bg�|w�QL��[���[.*O�/:�n��khҵ���K4c��ui��M_Qq�^����@����6�-��_�(E/��c��@~��~)��g������v�Z3#�m��	��Z\�jq׿��uV�r� /���qf���?>5~�l����v���)Q��^"�?���{�MS~A�Ƨ9��+�YO��DDU����y�⷟�� k���¢"�W�T�����j`"�ɾd[�ѩry��
B=�V� ��ޖ���^�1H�{!�`��ы��P0�ʴ���}����f/Ϋ�7mC�o\$����+�@2��q�$�fI6�}��R?�2f�޺�q$g'��{�X'a�QL~RF�!�Q�Y�
}ń���o���8�*��W���$G������E��rfFF{�#�a�3c��ό���VA��A�@��i��ϱ;��E2vb�i�޾7, D#��J���^+s�f~�Jӌ&�G���#���Zl� ��|V6$U�*ȩ�̪����Ɂ�.��LD�9��� �A���y�X�ֽ�ÆH�w�'�����6G �� ��N0�nm@����$��.F�����ᣛ22�S����{�YQY����zV�֒V����z��r��e���@˄p�F���J��RXy0ГsR|�!�b��C�b�0n�A�x�����*{?�;F�4H@jt�AsC�1Sz�O�_���Dx�ߵ|��r 	�-5{}�s��"]�T1��ѭ29.�^������b`�[��DL�qE$g�5��oPO
7����Y�-�&��@�����zHW��l\���b4R��0'qv�1DIA�u�c�y�Om(>w��>�/�ݺ9��0��~�K��͔O�����b�v{�y#�M"��=�։o�t|4H����ٽa8.���JfZ��%*m���Ů*�S���s�"�ō��mQ�Ȩ=!�����Ys����C��5T֞׀�333)Z��>�S��a�)+f˫�
�dj�߿��g�[�ě����*�F��u&p.OY��Hh}K����z��R�HG�Vl�oM卥�M�p�F�j[�_���c�8�MR�Z�U��֥?�e��S�d��� rܢ��.z\ҍ��wW��]Det����YZc�z����c�悦KT���������]>�OB"���R�V�)�a�����.��;tJ��hQ��M�s��ī+I�@L�#&l����gƭ�����A�@kܒ\�%OL|��!�� 0P���I"4'���m��$��Bݏ>C,)�|R�-Q�@/��k��l����U��=Z��U&�9�p��5I�E{��[m��ǜF���T4�V�t�	l�Z|��<�g����E��L�2D=���@i;KTm��5��=�6S�	)�:R�̨�M�y��Cŵa
|����E���2�'��v�Oe.��#��5~���RF�j���c�i ���U�8�',M.����gذ�g�s�m�S�����U�[O����lsjA�X~���k�+pa�{vy��(��o��ر'��D
��^uXb0آ��C�2�ko�?RRe��>�f_V��#�� &pnn`��y}�c0��m��S��-�DasZt[)H>*�S��j#�\�D����҅Y�5{�?���i�uT�>X�hɎ\h�Oij���iH�qGX�sh2��$D��B/���u��c~�r������"V3��@%1������)߅�@��6n%#p�t���,��2�Sr�u�>���x��LՌȝ��5�|��u�j:�H� ���5�t�9����?�<�[��soa`Rɸ��{	c�Ѝ���/�0}��$�6��$TRQ�T��p�~��Ӟ�Jb�����L5m2� �2��}��4�$��@[d���d-�<O�����?�r��H��	��\��fM)�<��3C�\5�
�c�z	�<,Ur^�#e��S-�s=�
+hr�qP��M�.�����W�����n!����ok4�8������^R�D����i	��={���H�ᤪ:Q���I� ��8�v�G�	���]��n��_�3t����'l�	w0Pk�q��}��AW�2Z5^R�IO�0�)0�#�R/8�$O��B��<	Lm}��bѩ����wnjz��2Na�ݺ��AVv�E�7�ک��dn�~T`ݯ^��ݏ.���j�<m�RB��3�ii��C������z������J%CЕ?����w'�bDT$~����a�'�ڷE]y�}���ӛ�J�ߍqkYB�|h��� (�R�����ð�#��\�G�h��G� �0[m^�1N�"��I�"�S{�_l�O#M^S�u�f�]�Lh��_��~�_V��/�� p�iT9wK���ۍ���w`F�������᱊RL��P�ݲ(�`��������	MLD�b*%nw�8;Ozq������#^Fu�V����%��H��BMB���I��v,�T9����l4<SS����aY��V����C՘"2��Z1%�o��	yf�W+*�j'"}"��E(m� hq���.�#o�`tF��3+�5���l엷��`��lz.2t/$ӏ�"f� �֙~�G?�,��5�R�T�nϑ�ї_.)��cUm��!�d��sU�����,�V���y8������hm���R`��nđ@����]$�Ȥ��j0v�X��)���Ȟ!�%�RXP�^��W���u�ꛙ�v��L��:� �r?@K�V�m\e��~n�9v��[�6�t9q��j)�6V�i�c�zY�^�����jDjj��U�T��.2�=�#��V�͜̼��h�����]l�Yo����w��i*,�ow_�sP@Ĥb���D�/> M� �c���V����ڋ-���:��~)�!v-�j�{,�mB���]r�%��ѥ�]��[�6�뇭_��X=EG��_�`>Ԍ%}�T����/N����vj�=��:��j���Vv�2V�Hqi���T���ʡ�+��ᩩ��ÜKVi�p�oﳙ�4Rk�g���"غ����|"G����)�i�>]E�Y�����{y2P e�J��u:�m�V9r̐����S����$*� /�Ve(����R	_![U[���ύ���:&�n2-�.p�I��uA߬k���f���3���:0���D6�uO�7 ��7���2֦,��_7_ߣ��-q#���3����ӱ�|�wؖl=I��-�MS���Q��Ɂ����
6��d�I����dw5���(Z���+��Ն�	v������]�i���T?��!���ZsR/8Jq���t���裚��
��n���� ���I]��r�j���8eO�#��<X���y\Α�S��_�7X?�����i|.lr��p���v�H�{ڲ�y��Te6��y:���Z��1����}\�F6WC�|�ɻv�|6+�W	.�j�R�ų�ԢZ�F{
hS�_�1��X
���aC��K���������*��91��"|��]�aFa�Ha9�7o&|�+cb�2i)�$h(ng�vN�ϟ���o)}*nJ���;�ޥ3k�~bOd�����"�yG�����%�[2���c���țn��N./1i���4�96�b�4�Wc��`}����o�9�Z$gYi�+f����ڰYm�rgW�$]iY�]RH�����7��=��~������F'��ՈL�G!>-�x�\^J�����n+��w _��3ѯd�����T��=� �k_Kk����{��z��~�R��#��L4:?b���0n(3��U�[�~������0��ȏO[sڗ���g|	���O��Y���Ԥ�>����_��௘>�MMW&|`=a-]]]Njƪߎ6�\�\�-��
�;#�:��=i�yW>]�޴��AUD$y�I�TY�� �T�C*1	K�<!&�vm �G�OFUZՠǻ�3����yW+dGu}G��۳��[����C6��>���.���3���_Ġ��~K����\iFYf��q:^�J���X�QҨ��M=����`��#='4	����Ơ'�=wSj�w;�4��Kx1z>� a��m�3�����΃����:~��A>�[��.��;��i D��iq?՞XgXw�^J�^��ᛝoPk�g�_u��d�zZ�!����ƕ>ȱ� ���x��#K*�����F9N��/ڏ%Fzm�����2v��'^�qA��V'���������Ӫ-H Tz<��o����k�V���<��?:�N���]��`��G���T%����h�|��K�X���Q ���z��R35]��Z��*��/�J�_�2���E�Ӏ_�:{��(9O� ﾗƚ��yub��w��S��uO��E���S���k߀�@zwpj{�LJų_��m!���� Mi�9�f<�#}c�Kd��N.E��\q<y�c���R5�K��hd�@���,�v��޳���%�I5��t����y�����8�S�6ܦ6�{�!޴c���U�oz���U��`X�֝�pč/΀J��o.f���R�Vjߔ��З|�͡=� ]8�_���"㘄8�ە���b�B�{�JI��O�Q8��ϟ��$sA���2V66$�p����~iJ�j�Ҏ.*��4J�ޣ��O���y��Ö���W%�4O}����E9���KJ]�.���{_�\+�^],�Z��x��Ņx��uf�r�p����d�������rF����V��F��6>`|x�%ƹ��Vfg���{p�yp���sy�M�癫�Փ%y��'03��p!��:nzzډ�濃R��� эU))�U�ۓ���)S�A�>�&&���b��$�����D���A�Ω� ��ś#R�S���uvLͣ���-���-��2�_���Xz�X���zyP�ө�~tJ��%�)NA�ݮ�z���18���E(��L�����$mmmUe厩�����}Oy�:�+�gn��%��j��uR+��+�rg�-2�W'K�� ���(h�w
�$:i���yMA�/Z1ųn���5�?���Vq�m�?
3]��[�U����?<<�5��W�q(Ì���p:���
x��9���tVN��90��=~s#�%޷S^,u�'HH���.tc ��Y�zT�h��[�`z%3�rq:�ba���89�9G44�=���<[A �K|���E1������7Ë?��L���~���Q��R���%�\Q�9:�������. �������J�s�"��V��(���?b�F��P�9]'�wiR�6`\wBچ�^z�\wJo��
�%�����ER�q�`Wy)'?�{����C��O~�C���<�@��.[����Z�%�i �셔0��pwW��^�Q��Ō@�X������~wyد��u}� ��^D�ǈwm�4T�1Z�;n~�O��dd�.�^�>��Wāz��.�oo_ ��r͛tcr�r�|�r���鶿ܳ\�L2���-q��70�~���0q��[e2a�}vGO�nE���NڗRms���R^4X�p#� ;'4�*�^Q.0������s\ɟ�>�pJ�y�?;�����nݝ�@�8��_ /�fK��a�'��?i�M`I,�*蛖�x.��-�MO�J t��c�-��d
fu~���5X@^cy�sZ̈�e4�e��u�Q\B~0���UU���6vv�mC��?����@mA0)�L��~E������)ӌ��K�U������Hx<��b�d��c���]��!ບ�ćm�F]��G6n��sH���)#�$�'�m�W��R��#����Hϣ�ˊK������+S?������m�c���wn��<뇜��o�"̫�%�'�s�g��.����Z�uM��}۷�Uu��W�d�"�c��w��{-�E{��H��8#��kE	�T܎�he�,��h�]W�K_�F܂j��I(�����rc��o��iT�����3����'Q̄X����[��!,�}�Y�b�ҝ��>wӧ[ؓ����T��0��՚?���>�f_�@�\S���`Q����A4!l�,�R�['�Z[�[��@Eg����?fq %P�r�S+�PCt�����"����c�{�w��uuv$o� ýY�5	�$��[_�<f(���W�o���n����A� XWv��ճ~�߯5�ud�G y�
c�)�T��q�Ή��e�n��lu\���@��}�ߺo�vJ�� |���1!F�������*��)o5�K7f7m��k0�n�R�?�m��.c���tK�\�!��L�T��ݥ����##c$))�;[9
�zz�^ �;7��R�'~udhc�]I��I��&j�|���uds谿��mc�z��8��^�����l���޷�)Ø�:��d~!t�ٔ�2T�3�h�ڻ�C�v�1Ԩ򤍟>�{��
�ό�f�a�w���ݎ�>�-���^����(i�i	c_;סN;�t7	m��5W^�Ptr�
ws�v��֗#�G�{�/};�9UuB�Sy�:C,��]���`�Q?�d|i6Ͷ��w+�3VV�t&AR��q�w�۽���KK~_=�a?K �"J������g�����+%6�:Ć��	s7���vv�
�L��|"�����_3��z��.��o;��Q{���`pp ����x����m]g6y���]e���ni������-�.\�C/ ]"����"��Hw� 1
RRҢ����C̀�H�PC0�0C��s���?����\k���k�k��*�6k�^����DH�"�3i��S��L���e����B�������-.�y�IM~Q&'�t�ž�t��/H�(Yf����tgC��I�E~~��𰰺�	PI�v����]aX�r�9_�b��kQ��hJ�-����r(�̭ S���~�_C��{��.YG��n4�A'?���7i/2Q'p��dm��W+���x%wMdR���fp�m�@���me��pfSW��4Xo�e	د����@�~yøG�9��@�*y|�a��ŖHJ�cx}}�e���8\���Z����.c���Ufڑ�;[ջ���^	�C���T�貄S�'o��j��	<%|����BSd���9����zc�v��}�u=K�u~���Y{@���fC$��.C���9,m/��_MUn...��3����I���r3�_��`�hu�ϟ�l�&��w��Q��%�%�![|g���g%�A��LP��0?�N�����P�ܚa&� �VW/T$� �:7;��?���d\+�o��NF�FX�a%b@^/_�J�Z?��)��3_{Zǿ�8=XVu����\i�����W[�7���W�I�����D�"W�vH%M��~���s��g�����D�f�e��k2����U�cq��i� ��e#�qĜ$G�0�%�"0��׊f�7���
d	k.�e��$G���HVo�n��}w�Pp����U�� �o�PR��8����b{h}�W^@jF�8�U�0��| H.�-%���t�\9DT��&~�A���ϳ�ϐ������;�ؠ��L_01r����c�j��͓�+��,��mn�Y���U��P��p���d���܋g��f�Ї%�ӊ]�,��$!!�Mm�{'jwW�o7��u���gV��X��co$�?��x���mV�����\� |���9.ԴEEԄ�+�}kQ�H���:2�_>��jW�=B+�!���@^�|��Ā%����&BGE�"͑�"�u��9T�"��oY�G�+�;[kۉ`��bCȥ_�������XI��JgI�ᥭ����$g��b�	�۴h�}���&��,@�����)����,W4�Ѐ���D�K���I�z�4s�=S�Т9�r!ۊjFυ�Rs!j�����@��Ue��
\銹�_ws�Q|Y����0{���᳻��.e���%��z0��n)�U����8A,0|��G�n8��b�OWO����]ޠ"�Ȣ���Qa	���g&���W	#g#�����
����\f\E��ٴ7���e�|3	�)_�ó��̒���x��=rʆ��L	2fG2�������'��+S1��n��4r����l_��x�=Yb�';�5����g��f"s�Feee�T���lzzz������_M%%'gWɼ�D��oamS����� �{~����ȇB����nr�j�Ȁ�RO�Hf��;���Y��K�M����#�mv��5������d�O�j(X�"ԡ�.��^-����f;�z�p�]c�����~#�����}:�1�گoq�F{e0���~כ�����0��4[(�v�gx���
�L�"��7�/_n�v�m�CjAn'���T6|�,j"��X��IC�%��$�1<N(D��x3�6Nd�s7��b�[�TR�K�6���5�%����A�z�����=�&�b��A,����ɻ�h��FL<:`.�^WP_��>�֧ �$�t�l?�M<�$��d{��/f�UE/"%+�\>�-���0x�g���\��y���F�F��F#p�^�z������B�wC��.��@m� ^����>mϖ�K>��'��-dk|��EgR��\8�0�ÔA$q=ꌔ=��%�k���u�Gjn��p�>���l��~��}`D<y�q�;�xX TM �o�%nBPxl*��Ui�ܤ�A^�:���Ǝ�(q�Kf�~2����o<�������7��` ��f�6*0$$d.��B�V(�+��������(�
���T�q�P�f���j��5�G��:�`��g�qL�i#ư�����kj���V�	N�z>Tq#VVVOo&�X�<B�ɊX���,�Ț
��Ӊ�ʷA�
��P�ד�t�ǘ��E���_ȸ��Z�t��5-�O�Y���8kwC>��&ע�}��}Ǎ���ys���Y�8u0��&MMI�����9���im	y/'Eb��}���5'��k��l�����/�d���s�yl8d�7���Py��1ǹ�>.? �ѽ�1��'�F#�3�A�QQ^E9�����p��2}�f��~F��X]������Մ-n���R��g8����&�k�F::�Ϻ��r��X���89+Rf��˓�[l���M�C�� �v)f��+��1���Hh��4�M
��=q,D>l�����(E��/�v�7����!I���G��3*N�]�&��[�߱,�������TI��4r���OZ��*I_6�,�Sʕ��Et-Η�f'�	��E���XsfwLON��7d���al�����ܔ�x~���ֺ�hYuz��.�(b�z����b�izO�4!����b쩧��qE����Qu� �)b�*�p.����>�o�eȻ�N[_�N���pZ�~�5�\�̳"Ъf'&�ihu�	�Fp)	v� �d���gE~�3G�կ��=p~�^��:Xo��]f�E���:�z5)\jn	�5y��<�b!�_��K������{�to&X#���RxKna�+=�I];�5� 7��Y�ߟ��WH(����^j:�����a�^�o+(iii��A��2��Upw,�C%�����	B2��.��gv7������(B�	�Y�g77ޅ����O"�!��ms��aڠM��u����C_���31�������V��+���~�m�c5?�dU����#P#H��5G� �S����*��车 ��Y�MM}��~�|�յ��k/?v���6-��޷���9$L����Wp��a��-�5���3^���<��ݭΈ]��Z&��#|��a�QqpIa�&�+*�%"ٔ49i�����]v
(�󬗕eS@���^�|�����g҇���е�޲^%�K� 4�jN_:��Jz�ê$p�yI��0("��i�W����ء��d���ѩ�㳬�!�ʈ�����1�{�Ϳ�*�{�����g��y�<L�O�;088�j�u��t͑¦��܌����D t �A�ȣ��^[A����b��]���6z	�I���)Eh�����A����x�]H2K�Ic��;D��#t<�!���F�����?Bʩ�@|�"�����)�e
e���%U:�A��X�-Zݡ�XY��Ց�
���ƴ5O�  ��*�ie�O���Oy���o�|����<HWؚ�åI�/68W����y�p�9Z]���x����Zqqj���q����r>x�w�P��x��b�F9^X������혀�����B�H�ǲ�v��]4����[�%�JzES���8$Xq�g���?�8�=~�

��(R2�Y��U^
G�Z$��ȱ&�T��_�%�z<;�������1�n�}��a�>�5�_�0oc��$]�$C�Ԩ�k���(l.ٺ5���V�q�~����Ox8gҿ�R�@�l1�f���2�����cO��Μ��.�������K�L��;.�/������ 9�C��s0i]]�m��p�����l/L͚X%�N(�{� �똻�)&�N���Gu���@B�XII2�N��4�m��CLd�19B_U,cv@o�=u:r&���i���,L�iv$8o��d.bK:�����&F�W����<����*݊ۨK�>�^XX�Y:a;H&/�JVU��?@�J?��Zs;.N}��D{��~ʵS��Mr�o�ie����0\�TXrn�|���/����{�ό�8�[q�g���2J����ܭ����Q�E҉�`� ���`�+�Y��G�0͒A�W�g�r��(����v���mw��I�.�?6W9Y7H��d������~�^��K1�FU�=#���&d!��yyy4�¢�ܻ6�1����~~�ʐ�OEe��=�6S���z'��V�o8�Ai,�,���.��f+@Y�� "�c�Q�I��:/�� m�zTy8��O�����
�\�9
3��Z{�{w��,����b�HY�����6��K�wF�����pC���EHL!bּ9�
�=nX�s��V��C�щ`��`��.��K����w&V�hJf�G�l*��	��uuu�/*�o0�_q34���ɩ�����8�����gꁚo�	��R��$���Ӣ� �J&y��(��=��><�����_ʩ��\S�i)&}ƺ�wu$�t$f��ݘ� o	q+B��K��(��\�,��N�]t)�w��m�	2�}2��B�$��>��ԘDW�s��=��^K��H���;Z/~��	d�߿A�q-��n�K���^�\ZZr!��[[[;߯Ś��0�]Y.��?�����-�w�x%�8��a�����r�EL�пj&U�kgK�ژ5�ˇ8�f8�=^�!}�^��	���^������/�)�,T�>CVD��(HK�)��}�j+�֙��w0쪷��G˗�@�!SN��Ҵg��5i2a�P!l���H����L���G�v���A����=�L|��x���<.:	=.H�h?��:J�I�O;.���	_�BCgc�!��{�R�ҍ2G�{�6[$�w �>�b�brx�@0��,N)�h^^�����ҏ�V��!�{�fcē�#��v�굏!X��H�YC��.,!Tl��/8����2�}�`��@��\���1�,W��� �a!v�g˯U�?Ie�IkyA��[K�~��DW��i��v��b�~Ԕn�,��$���㊩E���Ѝ,�W�L1��
��QvB��\��]��@��p.M�X��b����W�?�: ��gFJ���ı�\����
���j ���R�6\���Z�TT�����/D�x$��m�G�؊wC_ˡ�ٌf)̇G�;�q\��1>�멁����)aaa��EKW��aZ�!j�o�����H*���:��Гwµ(/ύ�u�����L������)��I��������ZH��c��g�sc%�qAxQ~��A���b�3#�y��jl)O���&���j��V?�)�u#I�@�!�lo�Civ���6,��Qb� 1>X����[6^�j�sM�]�Eu[��dU�V>�O.�r�H~ւXEU>�_]�嗁��M8��<qpt,-�g'0Ѯ��3I�/:�%�pҊ��
�o���f�sjYr��0�={|4�k#�8ȁ}����_���Ic�qu���* �Y�?���GQ�/C�~��L/��j��#}i�@��X0������?�R~���.M�ۢ&&g�p���2+�d��*^�g�����q���'���H_�^��NIkk넺C���O,�M����*c����/n��R~�Ա�
�Ҥ��Z���������� SӼV�Y� �9� :�)ǋ�J^"|	�jL ��2��Q�ݟ'�;���T�ofpYPU�+"p��|R_|5B9�}�N��⛲q�Ò�K-�Ix�A�L�Pd�@����wC�j�Kˁ��_�Ş��"!q�B-�����0��ɔ8>2�@SZF>��Bqu�z6T~�ߚ(yd�ȃ�'�H+�*G�w��RG�����F@]�@3�sh� ����R�^;���V�`�6��"kMF�{�f�a�=��\mE\�1bs����Pƾ\��l� BB�a� � a�����C�2�k4_F�G�����[|ǱV8�F��9�Jʆ��-�N;/##���� C��NH`ߣt>����Ǵ�'���������t^�)�;��0�ް̨���*ԅ$Y���!�������0��s9�ߕ{�-��A�w�i��E�>�ݲ��.�D��iMaU ߄�y L��恢�2�\���p�B�bC�~�,�.S���_:e�&R�bU�,|���GB L���WI3_�U��I�o�0K�s 8I؎/Q�Ή�|@�&<K��x������L�?���/���&
���'�gh� �!�m]x�)�͇�E�\pS�q�9�,dcff�G�=�G�����ĄQ9Ƃ��e��X��T�tm�[Z�J��ٗ�"��2�=([+W='r[�$4Z"��Hl�RBO��L�l���甶�� �)���L���4���;�5k�R�R��������o�0-���w���Բ�4�ƺ�9x��J���BjjS�]N:aQn� TDOO�-�PE���~�X�M���ULY�_���|��F�"��FO�� ����&�{������1�5�7UW찙��4�a�L2L?��=5��՞� pnl��7��\m�[�F��0�&B����x��Ƌxv��ˢxl	����Ǵ;[[�jgu`�E9�z���*6��=%%55��a?+���e�s����Qw77��-��}��4���=<�Ni����X���k�CI5���k�^y1>�����~*��UG,�mt��Hi��Q9Y֓1kZ�	޿鄳Ӝ�g��7	�L)�n ���C����PK   l�X��� � /   images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.png���o&�����[��ֶm�v��ֶm۶m����U������I^�y'g&gf2'BQ^  �KI�*  �Y4��յ�?��^R�	 @����� � ??R�B���W=������+�O��O[���6Y��0�I��I^a����8�S���{@e�ΖxuV6Q�޸q��Mr�X�$l���$҄����vsba[!��_���%�{�����~s�ύ38������$������bz�m��x	�������^������<ý;d�ȝ�7a�����$��?$��Nu����h�Ɗ|45���IX��ˊ��>m��='*���'�_?^��<r�|��p�q@O�������f�����n����O��}P}ʯ#��y7d=t,�dE:�K~���!�����%�� �������)��q|�J&+��VKyri@]�����uQR�c�|5�{�I��au�t���Ԏ;��X.�h������K"��`�כ}e�kq�:�ŏ����a��Q��?V�~�~<Y�?
�Z�~kzH#����yZ�; ��_���������n��6���L�u���m�����DH��	�����)^J0�P8�8�cȅ;�r��y��0��o����L���{P��?<��笔���(�i���?���\r��խ�R�H9���\O	V1<���+�*�h�JY��]�6��0z[C��5�%�c�������sN�1��e��.��P��o���'e�����"������v���p
lqVh����m�[K���/��7���u�G�T&m�骦���WBԷ&��b����3Ǵ�{��^�>��	^rh-n���Ǘl��'/ė����5��C��D��@��x���"�}!���֭%�܋�el��l�J��=EQ|/�sGo�D�I%�s��� �]�+����3p~B��5�#9{^=�	�����[T΁�O�~��9Ρ���_Y��Q��$���0V̑1ˆ��M(5% x� �p�/N�,/w�@���{yDXoW�N�^��|�� =1"� ����Xª]�|uECf��O�v�)�Ȅ���
i�'
8#���P�1v���9�ٺ��͕�1y:����%��e7��5�y`��H]ݠ��LN�9�j!�ᣳҭ�V�A���t��l8ط��`��ڳ�p�����������o��' \(���P�����^���κ�����w�?��A6�iu~�Q�l��<*+�����"<��X��I�I�"������ΜR�{�^����ƭh���^l��8��3���V$_��ı��q�����k�Ke�2	�/׿e�jtO��ʅZ��D�����*oD�n)�ɉ�M��9����[/��|�W'�����N�O����e��|�s�q���!uO�U,C����a۱��\܇�c��}s��rs$$ط�A��l�,:|���;�A�Ě9�c�M����7�����tx���Uw��[m�ω�3� �^�3��Ðr(d^-dA��b�ܰ,��n�����#]���b�_V�Cn�&�V��W4 ,���J`���a�5P�R���0��/�d�o ��آ�K�Jiw5a��Y��*��)X�m���U�ZH�W���J��̇����J��g�q�j0f��E�] ��0��}�eD�	ߦ)��m`�L�xʭ&'�d��j����]\���\���[���0�t�܇����x(0ˡSC�g5�B1�V�U�f������!,����4��O$e�[���	sk�s_�"p����r�̙���|�}�`�o���]�>�gs,f�����[��n�p�GK+M��K���֞�
�E��Ɔ�Ϩ����,����`�5�y����D�Q���]�^���\��E�����H{Y�F!K�e��|���%�\)�ٵ�v� ��,?8���fK=��R!�Z��Ci��^~q����R��$��C��E����������_�l��-�df��� �S��)MG�l'� ��1�k��d{J0���������󑌽�,�X�����b���]-sg������6�Z�	b�93���n5���A}���O��2x9��%:����g*a�z��:��?�r��?�w��� �0f$�gއ��٪��
���S-����b,�#��W��Kl�����E��L������șxhV}!:�2��[��3�Tus�ke��oV���6f�(S۰���-�P�С^�$Qxy��ngp�s�>Z:�,dX�1ۧ�g��ޥ��Oa4���y���3�m���YsImS����x�sãY�
�+NJ��5�4W�q����wAyۛ����+_��q��GZ��s�#���Ǯ�'�6�J��c��P�X$��nЮO%�-���L�1��1V8�?\,�&�{W�D�ӕ�P��t��i0�3J0f�t�b
�i�p���H�R�����
ϴҭ�:v�^��֨�o,�4� ����<>l���'?���wt�=��^�����o��[��?�8g���Y/T����w��b�Gp{�������U��Y~�x�U���1|"3�AA1��d�~~*��Я��hQ���M�MpA�zY  XT~�2KR	t@�f�
��y�x�'�"���QdAn�@S6��f�����|��}QBR�ҸBN��3���ZNZ[�����S %$K�cE�_ns�x��x�X���iv���N�Mc�؋z�)���h�zA�=**.�_����K�AQ��i��pP3s�^$d��.��H}�B�ֹ���o_�@�To��!��a�h E�@L�����J�K���uL�D�<��UJ�_d�Ou@ڞ�f�H';��$�@�N�<ۺ}��no�~.gv�0Iv0��z�^m�E��"'�2PW��\oq=�<BR�ת$�u�[���p�(���6�m~Y�\�� �ʎ�(3XIo#&y[������)a�+Z(nh�qn*n@���t�Uw�B6�M���,H-,����AS�;�rc��V�o=-������1Q��&9G��w�*��i����b+%��;_�X�7>a-P��lja
a��ÂJ?G��Vro͡�l�FE�������"�=�c�[@C��Y�����Ivl�X�f�(ѡ�_�Hk�����peL)�������������Y\�h�-�x��JNF��YZ��5vx\@����^�
�F��=��������AA���Q��Q����0�^��`X<Q�[�t� ��Lk �^ސ���p�U����^��C7bZ������6���'�m�bQ	�A�l4,�@��Dq���S�t���ܶ��z�r�9��O�Û�|u�?~�>�?3~oU�X�� �|zjS���Uf�l6�]���;
It����/���E������q�1aN��շ�X�:;�%񒕞�Y�~�VcbE_�e���aGx6L�a#g�u�i�a����Be��6,���7������ਃ�j�D�Ҟ�L�����ieA*�0�Q>����a��^e�*:,��2��2�^$?���^��*3;�z����s�ky�1����r7��dB�p��q�� �@PCb�~&d <ȭ���6 �C�H&�1o�*
������~O���*(ӕ|�����>���:��̛�7�P�<}Ōi��A�v>�;d��iN�bsc������.���d!��1���K���օ��V�����=wOܼ��`��n_�h��mx����u��\=݆��w�5��댼<1]�'c��6��a��wN���+O?4܂�J�c~.����Q8N�����8�=�w�Ҵ�H��R�=\���!l[q��;��}ۑ�����ZT������H�=)4�]ؒ�����d$O�V:>�l7��V�р�@�T��A변+oǍ~Ƣ<J��T�L�R�i�A��z�R��>GI��8�� C�r PW��;t�v�~������F@�S��4�U��p��/`"c�Px���<���Xd�3�:�7�<�WTYa���}�q�����R��[L�k�*vP7/������H�S�h$��lݺ��9�^�t���b�^��
E�U5�z'�1s3b���O�g��
636o'��q^���RE�1Fo4�#V���}��'�Aq`�-�ñ��	�ev�{�78!��k#E@�L�Tp�? �b|(��q�٢��ҷ�L���b�?z�[�Y�n���v���ue[�qk�#���$9�d�����,8�T���!D��s)y��h`��V|'��6��÷���i�ZB�z�0��gW�H�3p����WV/���x*��h81���"�2�x�~�NJ�W�vg`���`����C���N1c��&/x�A��|�iRf4n�ZLvL��5��)qА�5Z39wĨ�G��;6��O�h4�J[^^��374��PPu=$n���Da�����h��� %������g͡!�����2��]�ܸ�/;�(��}Lak������_�Q&�n���R��\�~��;��y~�������4m=id� D/��,g���Ӻl�ji�]�0 ��("�.����TO�m����A�/!Zʸ�.B�J��3��X욻d�-��f�88|Vƌ�`ʹ�0�a~ݚY6�j�Eh���<vVsʫ�?�B%|Q�ЏW�e�dQ����Ʈ`ÁUXS���4* ������)� AE�P�J�tT���,�!צ=�kd�x��>��M��ӧ�Z?4�NM���r��!�,7���Vv�y*�t �����"U1�P�+���Px�,�8Y:�{,�X��c�d�W��Q��n0��E����T�����K?{u���A���B�J�p��pj�wG�r)��P[��I+9�!z��u.Zk��-A�,O,DS'���*;D77��N�(AQ@��{��H��BAV�"Φ���݊��z�?���l�b�:��U�}�#=x��0T?�1��������$�6���I��7������mlm�=T�W��)AA<4��?f���{�~�=�$.�w��n�]�eteL?�BE��&C�k8�H�ղ��5��s���"6y~��V=��[��F;{�m��|��ʘ�`�%�1�pzw�J�b>hY;D�X��!_�l̧w����hO����(N�`�XʰI�����Ȉ�7c��Z�f���#[U?����d����ǹ���n<]���5&����.굘s�7�K��_ ����Us�-.?e�e]u���]�抋bL�I&C�p�I��a�$��+��K�t���0�-��yf]� ��?#-J�]�2{�.��SI��UuЮ�(�)��z~����)�\��h�����i����,*�ܐ�e���*�~"���%XPj�U����8|�=u:#\�]�CQ{�����X��ݢ;3j���h��1��p,�h�.X�l�G@����t:Sh�`���V��2ĉ�A@C	�u�=.��B���7<��(q��2ޖ�����2��5��8�6�d��Q`�2Ŧś�̐DTһ��% 
�ڲ�tj(���d5#}kKl�J��M怣�M��A��ޝO�`�hF�t7j��;3{RÂ���(8��o�k3ғ��+����MW�z6!\�^��
u��U2�����A���x��&3��h֥?u����D��� qG�e}�9��JJ��f�ep�Dguw��0D�93�-Ջ5C��vA�~�V��4]qrw&�M^'e�Õ1��]�s���1�V�G��3����csGL[��=�o�U�Ʈxv&�R�5��g��Q��x�/��P�a+�3'9]�hlc�p�ʬQ7oؽ��ل~�֋8�5c ��E��w��[��Yq��#��v�
�:�׬�!�g�Պ��%Ng}�_b������I��+���ĺT�ߞI�qfZ��� �M
���D���j����&�J��̉I�6s��Ӓ`-ՈU]�eh��H��wĆ�5���?b88�꜕lђ;]."���"Ma�ۙu�Q���	�3���mdFc|�\c�L�y��כ�	1���,�o�m-#�S��7�ǘe�s�jCHѐ7�FA��+ơ D�Mw�=��;ѧ�Y�v�k06�������#݌�
OL�*) �F���v����Q𩇟������j��W����}Kw�'U��@���f۽�+������t�H	���Fc�$�lM�I�j��K\���o�^�e���A�}�@�3x.6�+�.7"j%� �ڭ�Et4-�Vx�UJ1唲�f�T}���#7�E5� ��l����Թ����_�Z˕%_?	�M% �q���<P9:�5:1��4m�������c���xRh|4M���|�\b$�N��>!;�����4�BZ���t,��Yg��)Ԗ̢�� �5J���f]wC�qr����T���Yʶs
�N��Z�ģ�
?)gr�s栞��[������#���"�ݖ ��D*��s�ڲh��J���/	��IL6�b4�� �!�E� b 7.CƢ��	��,~斣�#x��/�sr�Dn��#��w�w�{�
¡�8=>s�k�&�K�3ԧ��Z)��P���k����"�x�������#1�R
�+D����}L+ݾ,�ɼ��D��>���@f�wO�}�:'��~?_�1��w���U�	m3�fd i)���Ǚ����;j�%�oڧ�f��GzS�S�	m�,Ze�6��6H]sQ�c��%Nݿ�Qf-M�t�I�PU�C,?'O�?$|������W�)���"d�&:[n�9�5��#��ӀW�gQVL�1���;����-��BP���N��jJ1�ȉ�j���pǌ�������h7G��N��ȹ��U��M����)��H�t���!-�z��Kc�Lb�w��>OX�`6��O�{�V��	
٫�}��݌7��	ĸq�/> ���g���Ƕ:>�Ѝњ�_�]m�nN�b�.�� ����\���d�
<
8�:M�< X@�
#m�1QE�*#e��^�v}B B3���d����Ev��Fb�tw'l$|*��r�M9ŦR�9H�`��������2t�7WE�{��c�w0��`3�������m��:��*5?	���5�3�I�;�p,qB���{�q������ܱ[���=�Q?ٔ�_����"g�3GA���lKt�Ѻ~�-��Sxb�)��6��:.��z~�MƢd�3�]�{@oܰ_&x�%p��j�$u��G��,]�0��u|����1�H6����Vc%�����R)NΎ8���(8~���R�L�;��4�p�=lZ;觋+��S�K{�L���ʽpz@ a��~�x4Te(���C�N���Ke�r�4}�J���Q���s$J��wv@���=����:�=p��U��`��A�����!����qb�̞��U�F�x�8����˲~��җ� ��cjSŵu�b�I��X�9l�)�x���ܙ�"�ã�z�	+#���>��˼�!��2/��+q`�������H��:Z,��	%������p��yf�,�Dr����~�1�w�4GC��������%��+��X����j�E�D7����g��Ì6�5�sM³$}���I��x��8+*-�K<Ǡtɶ��	{����;�@�k��p�hH�/��B�H]
�I*�_�N��{��]߮ɑx&���x�J��]�s��R\v�ӷ�`��=!9�[�����O��A��J�����3�^��}����XK�l:��֊���B�T���t'~ą��rۙ~4��yncߥ���g�q�c�fM]�_њ�����kV���n���:K�8�Sm���e��c+���2b�\%8�[.T�GR��}^~���*��e�⢐��S�JI��S�x�\�.]�6Ӄ�ja���l)������~phQ��R���$�^=�]�*
�+*�NLI�]��z5U�F���C0�&��/�DG�RכmG��.:Q'`�Q���8��H*���F1|���:am��.ݩ��v/S�b��C;���v%gy�	��G'|��O���+�sJ�����üdn�'�e�Ry�P�Z�7N�9�80:o`�a��]�	��ICDp�m m��kW�ٖܲ��̥A�z��:�&XYMN�u����Eg}���4F\\���S�t]I��t��qI���+�C��w����"$�.ņ����[�n^�kӂSuF@zQ�Ӽ����j=�Қ�T�0.䮧@H<�ގ��_�� ����SY�C�EB��U��a�ٯ8��Z��J].�h]�,���ە}��Dӡ/�1g�E饚���Km�y�J4�5٣�4dK�rZ�y�j6sdz��a��Ԁ���
���� ���j8�o�L73�s�Y�3���i
R�g�ȥ�r����L����F(N�lx�
�����^��8�	�<���A����y�%�x1bz2l���S�5e��|R�� l�"D\���h@y�� y�RF��sSJ�H\B��lA�O/����rz^G6���>�!�����I�\Q*�@�B5Eh6�; Kˆ&�I�#��%@Q����[�s2xW�rKB-0y%���!����#�X��!#n���T�#y?%8a��6zT;��l�.��0+�#wZe9�a3G��G~N�}l%OŞ�3�w����tP5aj�.]�2$K��cˤ�=�uc�6HC�����5\�����m�F���u~JŲ3�ܢ�`��^XC..  |K[�.«�lD?��-��Z�z.W���p;�}${Tsk�ƺQ�P��{��qgV�����Ҏ��H�w1u/�g$hŖ�AܩC	��p�&vW��A}QkZ'D���d�%�a�LV��:���������iW���_���%���]$�N$�y넳 ŧ+�u����Q[��^󞠦��=�Y�˗!�bQ�d��8��z�֢%M"	O��˷j���z� ��?GSELg,�h��V���Y�-��X��5�ݳ�FU��Y�SUW�-4c�����0p�!3V_T	�!�fu�0�4Q^��g�?��/)��B�1���֛��P\���P]IOgN9d�A�Y�:i����,5� ���gw�%c�{Ư)<u�b��ψ���lf|�f��$ ���ꃄ�R�<����g���3=s�Lq)T��D<�k�l|�O��ˍsiF�c�t)b9��ԑ,����CO��a@W���l�4q$՞^���M��5�][ЬJ����������I(T�.D�'ڑ1{��qIg)�/A/G��
��B¿X7�?��w�;�o�����T�"�1^�� �n4Jg��/�~�U
�A�@?�[�JO�*��{������e��\�x/w�q!�~<=-��X�E���qCb�\Mg�m�<R:�|�ˬ��[�K�[��i��xO�᝹'Vq��������[}����UO��5�ꃘn���� ���_��nEfj4]χt�{m'�}��D���?>���հ`��S%�V$]W|��B�����[��H��_��iYO��H�_+��|#���ɕΓV�A�i��W�I��h��k���9��v�Ӄ�t6Sj�08� .i���I�9�ܢ���t��n����."d�]Tg��<�jK
���\�/F��yJJъ,Vy���+2%���oD'W4�h��f��2�l�>p�R|���9�L.��x�/Λ{�:(05�����S�qeG�Rl����iHo,����7��ϱI�i�m�����#�9uPz��>�c�O��n��G�@>J�E�ʴ�]�R�2R/jU@k��ƌ+��:07=�|�]�@�R�N������~		OLٴ�WYUu��S/W�a�JLnRxg�$��;d^�U�J�x�;�,�vBi��7ٖVw��i�O(Sbcۢ��}n��E�Ol���������u��>�վ[�0�Uk��&I��\�ZBMe�&WS�rbY��Kn?Ş�����#8�%Mn�O$��<BR&��wU�$���lG�
T�%|u �����*{`�\`�w�^ S�G�J+�
|�����G�l�d���ʜ�
z�&��ɷ�!�i��B�qztG~�U��w��x����\vߥ?�j|�X�|n;��� M#�&FT�I�`B}5;��Wgh{`�p���Y��?��wv���Tip��j*�CA�xPS��?������������|�bg䱡�V	����9�;�p:�9i_9�����I<�>�9'��(���4��N%|�V��s?Olo��61����1��2����*�rN�X�Ӫ�@�:N���M�|_�=)Q�$nu
�A��O4w9ĉF����P��|ϴ�V�׹��ҋָڶ��Ͻ(�*�9�ҜK��ʭe\m�����'W]�J�F\����>d�!�T(!��`��A��b���I��JoeH8k�q��N����-�����ԍ<��NB��-�E����yt0��Ի�+��;ӄ"e�0y*Nd#�3����>ꗾ�l� v�;i�?D�����T�3��9	h�xB���9�:'�d^�4���b�~`�~����j�GD�p,
�j\���]&����Ԣ�x�{����%�y'�Y�ypf�Y<R��@��
��:t%#L��j�L�\)�u�(��V߶
���c٢�>�ME�e�jFV� �
��y��tJ���B�!� Mg�h�X�bMe->0d�a��c��%?����I^ �$[�ǃ86�ڙ%<��{r*�be|�H?�O����6VT
��;���Y6[����c�*���B��fk9J&�pp�@>ߋ\�q(��>�*W�Sr�c�s���r�7���L�/�@g�,ŕ����6��[�Oe&���A��hNM+��V-f���A,���QRV�_?�cY�
��
�#��y�]	�x��-2M�w��F�p��0�}�JP�R)�B���&�xP񨡧���}E+p��l�pvT�.L���Lǆ�b�n[v�����!'=�p���N�޻Yr0a��,,��lvs��i�޾f��i6H��b���3��h`�p=�]zZ.v�6���:Z���=dB��4�4��4���r����q�j��s֐k�eZ��0'kh�>���YG*W����?\��l.b5�H~�:+;&:S����yG;*@B�_A����V�8mK�5
�@C�K�����ۯ;�rF��i��+��Y�#��3������=C����84�Ą|
�Y���:<Mi�+������`��o�	�u�E{5��+n�g��	A�L(��v��+�;�� .�����-M�ݦkI=shra�9�^�(x�;i�2P'�y��Rt����;�W�cC��K�,��{�ƚ4�X5
�>�Y|Dh\�'X􅙆�s��s|���i�|�����x�����VFH�
��c�㎪���1F� n��ͩ���V��OYV��{x�2
���L��y����_��G�@|<�GZ���&a{�rv�=��6G�o�&�*�[�m鱰X��[^�Ld��!���js��{�" ���5��W��͐����4�ر�rf�f�O<�����O'�}�� ��D|�l����Ee�scg�\C��S��.�YAI��I�i���c;��p�RZ0���ɕ��z��~
M�1�u�#�b��w�"�Q$;^M�L�l����S�����BD�Yު�$B�;��E^�1��O�4���.�q
G����Ɂ��8�y��EL��O�4SO�z��%�Z�LI�	�'*ln3gR���S�S�6�=Ň �a��rTIF���Q~��"� >���'���r���QcˁX���S�sc�y�v�����UcAex2�	2�_y�h��Mf�������Sb��&�����6Kx��6�9g�Kґ�%`��؆m���.5sR�L�D x������7���Qb骭��b���*<�����V)�9����Ԓ�	���Y��1���.�/1(,f�p�U�Z��ջ��@!���3s��P{1��'rf�w}�)o�&����3��u7ϝ��#w]<�]Z��1¦�O)m-Km���+�� �.�p�!�\���;ݠ17��@�0�A��ܒ�9aXy�dA9�w��4?�!�#�v�_+vGkudt��I�ۤ-�&=eޣ�Z���2B5M�j+x��V�%�C��U�� ɠ^1KS;h��ϧ��F���G2�ss���N�Q�{�s�Y�f����ȺÄ����k�Mt'e36���6	pg ޮ�Z��"<�1����:�_��1���9���}�ETM���o2��GE���:	N)��_�e@䝾���`;<����(0���hqQ��T[����>���')U�'����d<\��K���}��R���fm������qL*j|&ZX��ie̸
���p�~Y��I�w-�O�`N u�I�Gu�uװ��h�ȗZr
�Q�/�j��u�
�VT����gt-h������p������=.ܡRQ�Y�k��G��f5~P�	�U�����4F�x���5��H��n���v����kt-T��u��5���݋@���cy|�wa��G���v�.D�'��� �����W��ιּ�=�޺ؠق����77Ej�Ts��ϱ6ȅDΡ���rlȷt�y�e��d�X��RyO$W�,�q5�%������������� ��7�ŏw9�}�z=���j����`+I�B���~�3ԧ2�x�~���K@��u[s�?�2Tuy�|^�8S�$����u>���a���:ņ�i�
�-��U�tj�,()�]O8����唎㪣��L��M��ִ���;D�69��>O6�5fm/�4�?c�H��`�oħ`fg�<k0��~�l	����jfiA���հ>��L�2��VS�J�����ݖ�=�*�Pwt��QU�'=�
�r��(qqf��-��H(�m
�a�ENS[wt}L�A�%B��Y4v,����8�O�K΅�a�.u�ЀoI�>�j�v�ky�F chލVTx��2RoW��D��d�߮N���oi�圎ow�6D���2��� K��I�S+8+� %� =��T�{I_ڛ�]���z�}_#��b�5&?��h�Q1窛5(�;v���։M���Y�>qّ��h��l��r�^l�c�g'�Fٞ��ZX
��Y�߮�?��U���A*@��=f�H��Hlƈ�����\=8�w���txj��D3��p�(B'�$��Q�S�,iE"���T�ČM7/�A�ƴ�f��8�u(j<w�5%9يE�#��u�9,�7�e���Q��ׂ�����@�*=��i����C�:@���>�Ǭ;�������Ҙ�x�N�}��E�ّ2<s�=�s-��q��]��ܫ멏ut�%E�5i��vU�������SI����h4������Mh�%{J"�7�Y*�\bs'� ��7$��b�;��*^J}0[����WP>� ˶k"�vy�j�x�A��m��GG��_+m�����I�s#!�ƞ��~�E��1��ZvxA��O1�9��fN�B'�Jn�z���M,?s���AR~u����0�-C���M��x*Ӱp\�Aq�E0������c^y�r$�9i\~��p�zdEJyܾ�>�ء5���G}?�#<JO.�����:�.4c��t�Q������yɹ���ޤ�;��KM�6/+��Wz�IUZ��)lѐ���o�I�x���l�=��L���#��n�ڂ�^�9O��QDL�Axv��u��2�d��R��0&ri�O�.sjí�������<������F����gL�̲�!E[O֮l���U�HEA�Cp�
oIͳ�t��!� ���jW���.V[p��h�߿�3�KrV����f���$��7Ym��[�nɭe�W���XQLcCt�Cc��A��sU�jK�@�Ƽ�]Oק����P{O�n+����Z9��B��r��0�ӧOT�����闚4F�]#P��G��Rʠq���r�k	�EW� �Om�*��j�Z�~������7Y{�%��q׏�h�N/y���r���[{ڕ��5Z�ŀpFe�s�UQ��^�2��N���� N�N��)z�-�0e��>7'{��ST�qZ�߱E��X�J��x���"7?�ْ���rC�d�C�ٹNa�#0M��}�,3��Q�T�Rr��]Fl�-��pl1��Z��0���X��<��ؙz{� ]��VT����GE�������T(��bH�C���?�ۯ��?U�=���׈U���q npp���4��:����I$_��΅?�w�q?s,�Q�� 8����c�x�r�{͉Hn��[4*�ϻ�퓄r����{��M{};�*`ls������ă �y.��qIZ�ҍϳ�I	���C�Ͱ��ZX��;(�
�~����C�Ϭ�@�ܩB����N:��?K]@���g�Ɲnŉ�b�F܆�El�o�A���b�S��ܣ���ΰ(:mQg�����y�����2t�h���Kzy�T��5>S�b"���c
+t�:G��p�������0�(I-/)�Ė;�6Ab\5�Ś�oNg�B��%W3e,4�8->� �� ��όƒ�?y������c[�k�7T�;D�k��V�� �E.H�!!�Ǩ�� r]��~�~z�|Xi8�`���Kk3��l��Q�{��Kkm3�]J/�
�~�+������u*�a0�J�����T/�3�H۲w�~�Q�ZZ����^����+ͺ�4�0�Nh �Ǘx�r�w{�ʯ���N��ǧq�Qly�])�wm���ޝ<&��$""b-�Ji��n}���sѝn'��u���F�w����Gn�6�(�K�k�������WB�z�W����?��D����JY����1��)w�s���	�6�#�~~�G�p�\��Ž8��X�X��W�������p�b�E��w J����^/;T]R��C���'�j/�T�7M��e�g�y��;���O��-����B���>q[��v͙n`+OP��[����yS���Ļ��,�y�D�:����7�T��G��S���t�����}m��&�0{��+�2������$Ojc9dj��	U���w)�V�K�&7��;�^�6ւ�)t�9w�AQI"���y��s���\�-L��P~359�k�<�hwч��N�^PM�d��S��z5�r0"�'��y��
_6yל�ڜ0��p_�%6��3�L|�lO4��^@�I��]ă�+�xyz,dV	�
0,3�����&C/'>��^߿U��>����"Xe��XNKC4V��87�����V�>˶��ϑ֦훐j7�Ԉ��<y�s���|��c���͖n�,�++��y����j���!�3��_k���15�-7K�d�x����Ŀ�sVܖ9�fZysQ"��d��5/u0�'�M�mqef"��� �<H�.4�z\h�뤰� s#�z���"��bF�qA��;S������d�g-���|<�)\9%H����V�ёK� <:�r��s����iDr��@�l����k���r'"<ۀ#��'� ����:��dnb�ǟ�+�ȃ$I�j�"}�rb����>�)ጯ�F�m��b��Xu�G�}� (�R	�7�G7�9��!=���at�>��(3���I���*w�9r�2I���7�4HSՅ�J����p����j��[E���ֻ�2�A�kh�2jN�ZB�m�1�Ě	��N������7)q���4^L���I��$���Q/4:�����:�:�W(����9]�/��m���w<�@c5���sh�ʎ߯�h�	�M�L�ɷ��lz\d�������O�w�~+Zm�FX1\�j{��:�]))Z�]�t�|z7�6/幕�ਝ���:$2A!U�,���eL��.��E�N�l�(��MZ���?0����v~�R�Lp#mn^��t���Zsݠ����Z8:�N����%��*|�'|���9�����H�#D�p3^-S��ra[��{��%g�~F[��=xA��}���X�~bzR�}��I<ࡢ&����6�s/�V�Mn��|�X�uR�$]�͖�zy�`�9K�����h�:Iʜ�	�)_1B�+�7o�T�������?b�O�>X$m�����T��VT��g=�� �&	��_ɒ�>�l� f���ˉ������:~��ǝ���<�?���:�k7�!b\����U��� @���!\��A��w��΁풉xkevp+��"	��dq�^��5.��4�����NÍ���D���~������8n���O�C����e� ��yB�/���n�j����V��a ;f}�+y<Y�TVQS�GZ�`5�:�y���vε��	�Y@̑�{]_ �<��qM�W��I�:"�_�s��أ�m_&�il�g("�CϮҳ���<��%f2�abSc*�ɂ+��bKn֍���	ٻ��N�!#�jebW&v�,Ԗ�@���R6��}��`S4g�sy����٘�g@o��S�lOV�,���^��R]�������k�Pt��[g�8t� `n�.���h;�a��p�����֮�<TJ��i����{a��(�n�u�a���I�͝T���C�H�����G]D`��\$"���*`�Jt�CnR_\�W�pE/89�]�y���߫��(��i�s���;G&Ғ��^�uG[K��u��)���8����JJ.�xz<��ǌn0�G�V��l�����fm�e�D�bϋ�����Q�0�qR�j��`�ώ5�ʒ&gj�.�%�Y,���ȏ
Z`m`Sh�cԍ��w?�ɪ�[eV
>�Q1&L��

a
\��:�A����� �ӍQ������J�'�G|Lz����
E߶6xi����`_m6���������w-#<��Χk5�?��ɕ���z�{5T���qi��C�i� [�OV���K�m�3����_߭��g���bśU�Q���'����J��V�B:�A�Yf���eS~e/�����/���a����h,�5�b����}���2��2��LfV��z�iU�fk���o��-���`����:�o_KӞ��Z�cg�\l������k��l�����A�i{��{�U^u�x��@�9JUC���O�M�M�-V��tFc?� �e�#.c�72H��<����0����+���^�2e��X%td݊�ZX���oq�S��l�T?�.@n�\_��`j��eǈ�>�-�^@-����c������*)��da�٫Z���|ر���X0>�5z��"�*	���L8Bz�l�
���}k'��UW�G�@�����Χ멆���Z��e�kem��\�Ϗ؎R��L�;�0�����>��;�k7�F��;3���لm�{��7�	����Y,P\��G�m��]�)�ޯϤ�l1�۰0^�VSj���XuiƊ����u�T��6݇�R-�ՈM�ثP�l�qh�o&̈́���*w?��Ƕ�=�.j�g�s�n��:Uk����¢(�������jKO������:��j�o��jK�0�7��1�ꨖ�>[�=��AU�k�:Z+0,V&(�A+��i���z܏LC6h��s��UYbZȂ՗�L��Y��9[k+@b
z�n���\���w��k@�Y�cfQ���L�
��6��]*s�֜���+<�T��gU�L��Zb<�
e	���q72�[+$�0Ȋq�r��vKA4�	n%7��������:�I�{��XL}2�9�pŻѓ��}��\^�3S��*D�^�	�R!�����k�b�wZ��$f�	�k���>C8 U@�d�e���bw�V ���T:���;u�w5Sx��C+mJ��yE����G�ڨ�e�w�_c֘�mF�D �^=�eRF�.�w��{�Ge�[7L��n]���	ƍ�?����!m@��|�GQ�IuO5�Yg����=l;O��0B�1gcb�{����*O$׀�=*�+{a�m�[�$ �2A�D�녺��=��o�zcPZ��!Z�W 2�Io�>��h�4�8¨GK"b��V����G٩ׄD51����s�v�g�jb�3�xգ;׸W6}M��AZY\:�.;�V0�	��ES@&����@,�%8����
��I�=�z˰�o��x�%[A�҃�u�e�$��͘�D����}����O�Qp ���~e%4X�p�	"����o��Z������+���Q'>bheBbOh~2ʷCYl�19B.�a��_���^�rr1W�E�Ƴɕ2�'���d�@>_ks�ҤVR{븢�{1:�;���h�u�K̶��;��1>�L�
��`�mQ{z�0;���"��l�g�Gl�`;��?>2��V��`���^��;�#X��+�`�2�����c6�Z���Ⱦ�Q8 �սC��3v;t��p^�;��9QN��@�e݌�J�*�<���~j�	5�keL�bRl��؀�^��F@�n�>� ��s,�៬�1���1/&#J��e3�F�֩���2��Z6ױ�V��3�l�ِ�5�F�w�Y�V��Mq<�Mc��P]�� -YSX&:��+���k��>p�a��[5�����d���w����4<^�an��_�-�L�Lk6I"���� 
�1ȯ�0����ٽ5���kNNU��n-bn!�:i����]6
�=sڗ���eX+��{���`�������~�V�b�X��?��I���Ý�_�ɍ�����-�Y���D���lw�^_˭�c6����MV1���t73�\�
r�� ��o{Z�DVcT���.�g}�Y'-+�C�z���b��
l�������(C��XSP�Q;�b��H����I�O��]T ���-dpV|���������0���:�6�s=X1�^ �.{� ��>����-�`(q��g\#���0E����}c��F�^�����B���W��K�@�花�d�#�7��3)�\_I_X�+3>hSZ2�m^�B�
H�H���tc�60p� �����(�-U;ۖd�K<�����XOr����0�/�/��S��|���5W:t��d���o=�^St��B�b�G
*�Ω$
��@6�6�*#>9�����!&�� �Ί�4)6z��F�vf'�2;;e<���Z~ү��v�=xH��k=���#-��R����-v;�4�J�صn�([��1���%���[$���"�ϟ`d5ݵle�v��ǁ2 �w~앵5�6�l98�g2����t4��єeIY�b���?�I�ƅ>��W�
���P�[��K̯���h������)m��3cR`�c0E�p)���1"���2�d���a�(�ؓ�7��1#+BaX��� ?3�Њ�� ��e�<��2`F��D�)�u��fw��K{�A7k����E��i��ى���Q�G���ʬ,�X���4�`��J��+�+`l��Y���HCjT��j�'��Gv�I ��-6+i�E�1�_%�5e��on��D'��ϲ�����٘�F����� do���?�z몂�~ce�����,w�~��4��e<���"��]�"�|q�*�@˚*���(c��K�� Y�&յF�/�s��K��t��5�Tй�w����,�zez��ɜ�F��x���FxV8%��4J`����ۿ����{�V���F�ʺ��n��"�%2l�H�$n����lp{�^��6q�8TA�˧�c�5X9<���t^�<CE���>���gv/-����l�y�mVr�md�*6>�� �bM����|�:�8�v����n9U-��L�v���<�}T�")����@wL �:2&�{�X���šNq�^���������K$<!�=&�Xti
�Р�ި<j"���M,h��[Ϟ�!���`0J�P$>g�B��aѰ)8��Y*�����5v�j�����~#��s� Ys��;��z:ޯ՘,��^�-�7�� �Ǖ�j�s �h>�s5:(����Fb�Fw�8.�lF����R�o�~��(�:�cPɲ�Y�׼�k�[�vDGcS6b+	,�;?�hu<��0ϏS&ǌkhQ%O	�q����^��:�w������k�_��hp/J�"���챋3��k��g��`-�N������S�H��h���y�F�������V����浯.e����d#��a����zA7`3e�1t?S��ÿ�W)����OV���<yX��P?;A�A�61�ٽ��`}���l����El���QۦoX#c�ɇ�bA��\���^F�6��Ɔ���0X�t��e�<\ 
!"Ļ�K;�""��m����4��J� ��ũ衵��x�i�v�'���䢗z�=�D��am��<��Q$s�R`���{��!V֌����욲� ����(BM�6�x=?gK%�ù��374!�+�0/g�0 �Ѽx������ ��N��FY���ZCun��PU#�^m���d��e�ǥ��s����n��<���j���!X!`q�ݵM�`u;}�eS���H!r���d�,��$R2���uU{�#�� �Jr�[�����d��$��>q�v�Th<���y�k���]���d+�3-X�o��%ť��������:��a����� P���:�ҧ���Bqy] �Y�V��j���[3�N	4`�(�����|��������3$Iӥ25�(� ���|����'}�����?���Q�l�f�K�*�EH�7\T���z��)�Gl�n��<�ҏ:6��jŅ)!���ʉ��7��\���}xJ>��9����8&R؞��U<@t� e�(�fg*jL����т���t7L-�&��H-̫J�ji���?�n���քV���B��KtQ�8B\����k��:Y��Gl����y7���R�Fj��o~V�7o��)�� Gd_��tq�ȶA��]I�ݖ.P��6xQ��z���� �V,�B��;�~�K}�_|�+�[pX��Z[�)$xnɌFM��cRBB�u�
2(}S&�s����jbٿ�	�����)R� ���e}{'�?����(�z��3t����[�Z+��(��~��Z�k�3
��~yJA(�	{%B_:~x�<�]�Anp�^Z�8X�u	��a۶s�c�c�F��k�}�ƈF��'�E���G��5��ve�ʑZ�c����'��
��N.[M����7����Q+�1���+#-��<H�Ǿ&�}�t��~�4�c�<j�Jr���6����O����p/?-��z�����ѹ��[�&C�(��b�u�
�	m��<��3lL~�u���*��V�FK��*���*��S�|����@'���`�=�:+9Q�YיԶ���MZ�1pmq)<zX$0t:=�6���zγ�>H8���>��C��Q! �BݫW������v�x�/.�"n�]����Z?����J~���'�@��p Nv�P��%X�m­yL�Y=ȏ�k�_<�d7e���s�j�����֛�/tQ���R��F�TA���yzfȖj]7	�Bk9W�6����X�%��ۡŵZӇՒɓY�����1�n���q�Gs��a�y��t7z���@�\�R�����:P�ʐ�+�Sp���w���c?0E0�ӳ�\���D�[E�)b3�Ģ��Q��lD�&�L��I�秮P�s��Q`�RZ��Z���>�Lg��ց�d0!��Y	�C��{�"�~�x.̔�K\vZ��kǔ�$�ŷ	�&�+\�d:�x=�mc���"v'E�]ڞ��-��ҳ���R�������1���vk;�A�./�F�H��Kit�L�n�B���	�&�6D�[l�������N�'�cc솪7���ӡ�go�&�<n�ֱ����h��uN�^R���T�y*�V`�r?(�p+$eo`(R�B��!�sR� T@��}�M��n �>P5[��Ko8�O��CA�T�h���!�l�Ԗ4�z�ߨ�y�	5z���阌�Zj���v�L`���!�c���������e�t�3lBw��y�l�����ޭ�����h��.Vo.��:�3Jg�e�
���v)�o:l�Tw��N#�]=��pe����e�uFb��ny/WՅ���%v�X�
j+����L@kne�jPv��ѫ�e���Ο1�7�����㹮���Vr���앭)J)��Xneį�^�]>Ah�k3�W̙����umn���ѥB��!י���y�0>��k.�C��:	���.�~��k. �,o��.�����~�zH��8�\:��m�$�V�K>�}9���i<͈D: �'��4�g�6�m��lL�9�L�������j��� ��s�H�RvZ�܂�qk�PX#��nа,:c�#�妎Buek�f�m�0b��VΘ�Z=�'���f�(0�Ȥ��E�-嘸�u�9m4W�p_|v9<l��/{S���{�vj*1��D2u��u=�B*ix��P"�Q%���U����Ԏ������zA��o��m'�O��Z(!pK������k.(D����t�bU��G��[((���a�Hw,��]=��U
x�_��r1�31f}E�R:~����o>Ȼ�k�е#��J�x��) ���.zkI`;n��*[�̏�G��F�x�o�R7/}d���w�brn�f�߅/<�k�4�w�������J���J����V'c8?��nAa�XeV+<zC�����-������ K�E�g�\���l��2�tMQP{�����ה��ul�ܚ�Ȝ�Ţd���L.�����G��~T�Hٜ��[�1���٫+�Q���$��dG�S��?��޽��C���U���^܍�74.,셉?'�Ltp����.�'�XWa��1�y��woso�țk��%��HK�L���R�1㙅t	��]�q�m�i�=tF�o�E�L�z'�U�u�)���_J�FVŰ� ��s	�%�H@԰a�0{��;��۟L/�����r2��(�?m���K�-���-=��9���A$<��[ñ�:(̓�&{�e�
}��=��a���C7k�Z��w��rC
d:�yă���H2�@�%0 Pe0��oj7����ڞ?�Y*����?Y��L�M���ƁUAl�M�ƞ�ȧ�[@~Z?��v,
��MJ��td�%;J���
,�4��%ܕ���7�NG���K�����wj!�=���D���ƑUm�F����Uw#�-.��FhI�����ݘ�����,t�vˁ��xʓ�w���A�z�`��}�p8�NX������+�T0��çz-���}�����o�g/�Ե�W�����R�x���B8�~Q���~���q�E�D�N�;�'��O����������%�H)1��1<Tz�!co�>]oMܻ^��+�h��]�!AV�,�gB�J��.p��|V�c&g���Z��۟2�!.:�Is�{O�0=S�FK�lA� �y�<�fе%EVH�`S�d�Z�*6i�M��W6�8�V�s�̟�w<l�o�Lp��� �_��_���毕����|Jŏ�p������taC�a�X	(�Q<XUn<��K�+��,���tf�L�-�؈	'Q� �(�x�1�=�#�^F
tu����%`���VL��{U���{{�gL��]�
4+n,����C�:���xE���mh�'�u:�S��*Y�F�#۠�h��ܮ�V�Q�#�� l�v���� ~ j5����^��kT|�4V[���AA�����P��­�����]�$iQ���'|>��/� M�����B�Z#��.��2&6eޭ�hnt��,�zP�C��͛��g�|-/�.����{���S�0�\N`�8��7�d:��K}�m,�r��bAp[+�@�b5S�=�eM{siNr 67�GI��6[&C_��B�<�Q��֖0���B8*O���ۓ)O��8ؕ�ĝ�Q���䰙uʶv:�=(�r��xy��~P����|٫���'��? SgI#�m5�Hbw��Ƥf�A��:� ��}���'�gC��&�G�Ŷ촦�ѓ:>g�ťG�c�Xu���榈�z��)_ 5��Q»%;5�[�bI0���S�]�=L�
%�nY=r�7�/yѴ�u'5���[� �5���C 8��N�=i�L��V�O$Zra�	Bϸ[�]�馘� �����G�㞺2
}Q]��h�>���CG4�h�lE�;��5kSˋ�Q��ޢz]yL����"�O�+�f��2(�v�@�bg�b���LV�>�z��(cfJ��_��l ��^�CR`Y�)�����h�^� x���eG$h
��Υ��o^��+lw��[�����[�*H�WV����VX��3�v�楌fc��d\�56�QV�]��z��2�Ll|�XK����`s˥�!�w�M.�F�0]6�ʳ���h��5z2�Oſ�3�1�S�2��{����x�o��r~��D�$��g��O�'絏�59(J6(���ڴ>o���h�i�E�Nx4�ʰf�}����{��0?�;\��SMR{� ���]$̊�_v?c���U�kz����;򘙢Xט��'<N���3���,��f)����q&K��:۟n�~צ'J���`L����$.d=�/�w�[��Y��)�"-V��Pp�P���2�U6���E�
�f�#Q�HԔ끥+,zG�$���u�`�q���{ۼ:�n�=��:Y ��{c�;�>�Is����6QM�m��C��L��z#���Z�l�F�a�2����hx��|�:LP4E����.�N�Bn���YT��J����pn��Yt���ɍ׭^}�F�&{l\2;���٠�Aߋ,t��E52�*gj%�k�$/K)f�0�c���U	���D���N���\��g0�*Ȯ3c�,��Tdx�Y�Q/�%��:��Nr.��m#e���U��ak"�{�����j�X_M��P$ds����$ْk1�!Rg�VG�̅�A3����_��v��F#`����Ӣt���k�{DVc`�6C�P}��"#���|��>�T���a�,�"����p]�a�����ɠ�ԗ�V6ޝ�=zoqi|J��w�o��� $��or���6�-�!�kF*�/�g27�9�:�V����҆���},Fw+R�O� &��
g�[� ,{;V�?�I��W6$ۈei�ś�v]�϶͛/�X��4���v���`"��{�/B�#o�J{���;�7b�']a�w�_��jz7�6�Z##�{,ͣ��� �[�lWX�3�hH��}��Ҩa�kL���Aeaw�nS����dq|�#}p��{k}�*�*�#�XJ4?�puH��B4����|A,��~'��7�kx*MO������������>��k�/hW���gTm�4���"����#E�E�h�M��5!ѝ�0�N� �W�c�cd1B�%ڊtAbF��a�W�]���~�?���F//{a���"
����K,.�}��/Ch��#����x�w�-�S�n� pQ��#�ʍ����E�#���K㢲���H�:|�!�б|�떉��V��P@��!��4����O/Ӑ�_T3��d��e�t}�`�|9R.���"�9�*���=V_��p�YFŁ�	��+\a��e_�م���3���\I"�P��
ύ�\e_̽m*z5b���!m#" ?�|}�L
sϋ�
�il����<޶�R��4�$�X�\I���ޫ�jh~VS�j���
w��'>�[�/B�Sa�h�b��<t4<@���im(]�G�����G���r�R�g5h5X[�j�{���%I�4pA]�\�V��-��*����
����v;�])�&*�Ɇ�(@�a�b�Ë�����I6T��{�i��/��g�π7�>���q�B��<��|��x�L#�)��K/`0�2��k���4���5�r<�f�(%�\���nD��ҟ �o���@,ئ��j�;QJIh�5�Y��֠�Vz�4���ʍz�L��RIѱ\CX�z��^�F���r'��,rYJ5`��� >Y��_]/;K�F��KL��Y��V�Q��1.wɽ���hÈ@�EI'����dA��;�Qc�7q,����<n����,��:�XPё�:�����d~��)�3 ���EO�K�ɇ�qPx��ֿ�Ȉ��=��r���Y��2^b�4�	0��&u4�eQ	�q˝g�c�o�X��|e/?r�;��EA��*CX{I����?�t9���ٌ�B�h.U���gA
Fs��@�Uf��Z�i��}VC�6�f�i1�uY���Q��y����xo찖�kw���#�ɈpJ�9�β�<�|N�H��^�p�<Y@)}�lȁ���P3n�U�ٽ9dU��>����>�H��(�J������}���	��x�	�:�R�SK�J�H����nT?�iܻCgk#yBEB�6�����������v�?c��`%��N���h������&�L]��Sķ��1,s�#����0��(��{)@�S0j$|�0�����x�v�o�d'	O���4���}u�	�°�����d�P�&�'%qV�:Y��ul �Xlx �p@ �2�<�9�n����� �F趘�s�FD(ނ���J�����d�A
R���9�$Q��<����P�a��X�1�����9
�Oۍ��g:Ѓ��E�����q�t��̃C�3�����ŔY94x���vd�jP�]�r�6YAKFH�%8ܳ���4�&��A�;SFqx���i��1DK=�5��V��̰
��n�҅�������0r�e1���\�R��aL�UC����e3�*�i4�)l}��G��[2y.b�>�����°�H������.��0�����L��t&�O#�)����vŖ��fK3��M��p>����:|��3nu��\���[Y3c��ʦ�]�������)��&�y�9�lr,��	����g+y'���O��q��Q���:�����M�M����P�h����@҅.�D%�E�PFȆ���#H���w�>��7��|���$v�c�|�{ �˭�\ch��^�;�^�3Oʳanĸ9�> �!̈��syؗ�K��4���C������v���f{�O��G�Mz3H=�zjHB�5��P���L�maMC����d�X�P����޷���Qs��^��*7X���<g)(��4Q����qϵ�q|>:5!��^���ŃnNvwε�b�������r���e�Ww� #8"�HHr�\�?ֽM��<'{kC{�%�x��f�y���1�Ҽa+x�~Ș���#��]&*��4���u#�ӻq�'(�k���q�A�1*� ���㘺�Mj#���&㦳
����qS3��������|�/�Y2k.2��uI9����d��j�%n ���s���牏q��c����1��˿+"Tͣ��%hٯұ�x�>�K� ��
�X`�JisR�����|g� r�.�P�H~�.�,#�_�7��Z�9O?@���K�b�z�N^��n�[�?�`�Ы!�ACb��'KY]]�Ww��n��|$�g�ɠ_�(���\����~�7�?pfЏt�;�z�����"6C�\;�����y=V���4��2��Ƭu���)!����}��/�U�����;�ƍS�|HZ��k7I$\��{�b��r�bT���A��u�b/��"L�.ݔ<ꡎ[ʞ�3/1�ђo������XL�\H[���{(�в�>��W(����;�p�zb��M�#�-
ީ~�S�N���R����$Bp��S� �)g�'
�����+eT\�|��Ќ�����h����04�ga؊"�c�i��>�΋���t�'�k�ׯ��q�<������m��1�|z�0f�y�l,�e�<&[\8����f��4�u��2ϙ�kg����ć��Ê�wQ�C��Kc=�����i���Z�ٮ$^���h�� H��[�I�u�z	}|��ۙ,���y�R2~��;��wW�g�렶qZ���[��_��V�;l��兒�������b|G�f��͇g�,;��J����j�A��W�]W*�j6�nZrY��>*m������ׇl���u��d��H��3�f��`CÝ<���ݠٿ�+�a�AɌh��=�A�k���o*�������=��A�ϻtN"�[��SHlm4�P�F$����;���C�pѵ�Ѹu=TAt�~u���r"�cX�����i8��[r��Et8�^dH�j�E�b�����5]��b\�A,[i�M�4�v�x:�ߛ��?u���j���ar6o���q`�F��L
�� g7%R-֟;��a���r�8c��I��'�1EHM�a����#����5�<̻x�j�"L�Le��LV+�=�������;Y/�r;����kzzO��8A�K���w�Ï?����F�W�,пx��_�����%hI��	T`gSv\?�
E؅�2s�
���xd#L�!kF���6�T9��LJ�iΫ��LB89m��l^rU�����:�}�l4���9������<�9��W	��ܚ�c��:�!}�s7�_|Syeڨ[����	�_h���E5J����evx�W��u-L���
x����p/�Vg���a"��Tm8]W��ߩ�������iM\:ϕ�6�-���tÿc�.������)Ӏbą^��_����&�� ***���gj'yش�������w�Vɠ���%3�Y�聫����
��H�3���g����ϖ��t:��dO�~(�d-�Sr�/��2��^��1I!G���a��0���h�G��B����R�˕��n�"���Y�HqS��z�A��Tn~x+G$N�L�0���O��ݭ\ݼ�]n��w�ϟ��>��;������Y�f���u��k�l�«��\�"���[�aa�,?�&�����B�����v̸)ޑ),f���@ǱRK�����i�]�̚�>N:�^��ü�������0�[���x|�, OTx�0PYҨ���}�����zv�y��q�r��:>{��ݸ�6#�6�y��h��˺{	y���d���շ��j�6�\��NW�'3���uq!3�nx��6��$>J�q�a���H�Q�$ٯ�����߯��i�F\�J���0��F4����541�;`�'Y�(b�F��h8�y�8!Q?
yn�d�A�5�+Ak�ܜx�l��F�����)D~�$ǋ� wx�\��p��b!=?f��Y�/y-�F��6�.9�=�������^��f�~���j����ie��7K?���@W	� P	��~�����N����_��G����l(�3�^�q��Q��ƞϞ�8�f�s.�H�k�mM����V����Vs�=a1�j�,=�� Fi�n�|rhƼ�J?���~��.W��6{倭��p3"'�[�k�L4�k��9鼶��$�!vHڔ�
>G�+^ms��D�S�̥a�e4��#i8��q�&Cb)�Ƥ.MN��RG�9�Q_��HY`?ϭ.��,�Hw��^z.v�F{��Ɂ(׺�rxm>(1H~�����\<����	�?��!�2����&a�V��������<S�_��xJz>��TE8����dtL������nԫ�i^�H��+=�dV�iᡕ���\D���aUx���0��E�f+y,c�mm�5�C+C?չ�iX*�����/w��5�{���(�k���@M�/w���dj�lX��Q^��>??���_�|�_�R��zsK��j9�����(%��-K���)�ea���J�� Xr��%�Q����ҙnP��f�ַӊ����X�g��%�� \ЋB�_|�z7���G �������(($h�i��<SxD8�����%lx�2��N����Ȁ�����=J��qZB��%BP�;.���#��6�+�:�Lc'�Va�E�<~���V<_�r�_��&�V�Z����]D^��r1�EX�� %N��V�W�G�'�CQ����?^���{K�[���W�j�S���&��|:$�d� p�u������<|N$��h�g�r4>їr:�m�3O*�O�3��hM�q�h��[��_��>b��(m���$��z���1���Sk�c�^`v���T2���7O����T}��D���J^���&WW��r>�Y	��կcùJ&��,�ޒ,P9AU%�ݙ_g��SG����\da�j�Y�o�UQJw�=hm
�«A�$��TA��B�"�b�'RT����osg�#cPG8^Tg�2�֖0��l1�k0���=�2uxY<�`t���C/����xI����qK�A{�55�1�浡b �l�I:�s�q ��z4t�-�|��͆�qX�s��2zi����vT I�� ^Za*�qH�����������-,�a���0��C�0VA��-m��qaY(ֿ2��C�"]`7��H&D���3t��~�@9��ھ�.���ōn�p����uC5$�㳼���dJ�(�����!����Bi48�j��P�_���]��+���ƸN���l��`�ċs�1�J���!������DQ ��H}��1g���q�v��!Q�\�A�75Ps�~��� �ܪpi)5vF�md���sxU�=��=g(��a�xf�����y�¨���P1�`�60E�����m=��[	K�8o�*[���̮]�f%��RL�v���XK� b���'6�*��M�WKI���B�5�!�3f�+�x��ۡ_Y�߄���$Wϵ�vxsֳĈ��`0l�v<��L{�T���9e��8��O��ŐA����8|�c���M�!���J���iJ��p�\T��
�Y�P�꿣禋8!�7��"^Q�.�q�m`�<n>�n}��~C
Ɔ��P��D���͸���vd�F�.B��<���OD96R��XC8��w1�sO�������h+V�����Jօ)�M���~8�MUD���5ngj����n�X�޳7QS��}F�n�]��uC��0��üE����2����9�>�]x���A�,��`�C���do�a�3�徑)2�A]�{].�$3n%��d�c�g�04"�W�&ǄA���Y�D3rn�9�;K�V���{�H��S�z�%v/�r84��UE��Əʳ�WR����?S�~6�29��жe~�lT#\���ʥ��h=�	�"��������:7VѰ	�HER��Ll��C��>!�������b��I���g~}��K°8�W
矇ia�W�C����<�
!�wNR�����o2nM:�̌�����͜dld5����!��{�1(y���'#a�d���S.��WY�ˁ��ϣ����W�0f��p
�����\��C����,0ʃ�^.?o�v��bɗ3M���p�U�O�/�YZ<�o�s����W"��#\�6�ĐJ��g�
n�*��fir;x���W<��ys�{��������IYy��n"�
�F�a���^�¢�ݳ�n�ck���bcR���~^c���!є���zHJ���X��<�r~����t����g7�+y�n͎i�ɂE���{ު����([����;;��ᓤՌ\��%]x$��L����<��<�ތ�u�3�8�PB�F���ލ{f�G�/�l�@n��p	�� G#%j~�u���R�Hn���dې-��{�v��~ˬ>/8��!a����86)��u���Q��:�_���\D
ظb}��ES���5,���&N$�a�H.��L.5�?�{�3p9��:����$�&�^[�]N���;$�-��8�}��CB�Q��5e���;-�~� Y6�r`=�H�)*�˽$���F�D���O$2d�4�g��o�(M맹��R1x��4B�4��dPK��j5��p�����P6N�Q�����|�D8)����
!�[,Y�vq�W{��U��Q���������������B��=�B7|�=J��"��'���ܨg���[����߽�Q�^_��0&S9�'GY&��Ѹ���Y�7��_�g��_?�g@y��%(-�2������&� ���m�S�����Ρ���+
�
��C �3�ǗA�/����̨�ƹ��e���v&C�Dҧ���uԈ�����<�1,m�u�x����͞�,���LP��t� #]Y�����D)_�� f2��|�Δ^2��U���ԏ�[x�"� 9`fn�x�H`'� @鿿�w�����^%=J�u-�v�]�'[������&i�y<�<�������i��C�T����AW2<4��h� �����̀�.�Co��
I*q�
���+3R�m��yF����W�C��7/5 ��u�)�p������/�c��\�(�NFi�U�!�g�0@�k!J�r�ҔQx��Ϛʱf�3[� ċ�Lw�+��CU�1R/���,�Ӌ�ۓ�N�������������7+�n��z�B?������NGyz�#I�_?}���_���^����<��4������c�,�7����pt�B�����7��
��N"��R�c�(1���N �\��pY����Z���5�[�-a2��K�i���J��h�;��UZ��~(��?�a9Q�"������!�Pߩ)3^��̓Rm�\�|�a���O��������D^�����E� �� exp�q�u)'U�r�M_�������]lg��w�V6jJ+�w�f�n���<Lo=����J�N�'m�),`0-�%�VR^a+��q��P��S�Q:tA$�.��0l(��^�ΐ1n�l�a��0��P��/X�̓��J�"kZ9�"��Pz�$�v^�$�\yP��.c������Z�)֑{k2�Hq{�+�P�ڟ�y�H���u�����?��[��~����r[�%mO��ye8�Ԑ���^��IZh�:�~����������/��i����@��~s+�Ŕк=uN"7W�*P��u��l� �er��m�(�b�#��(�&��F3nT=α7l��2������mq�<'�Z�T�PE��zuu����Z;��u��/����$cȥ�)y����+�H�u"d���3��!k"���#ri���<^z�����2���v��̏�\�y4>q��J㤉�N�!���չ"��jx~#4{��7���w�Uf��1ݟ�/+N0�zQ�!(D'E!g
$",�=��g8E�iH%Q��N���W�Ie=em8��=(&�B����}�Ѱ����=J��r@��fh hZ!zg$�T��M�I^�}�,��ʚ*�Q]�l�tgWo͔��6}C
�v"QdwBjP6��2�ټl%?�d�F�7�~����'����gy�\�����v���e}Y6�9@:l+�q.�:eo8�(n4D����ӽ4z�\�9'��R������o�,��vuB����0<��rZ?����C"f�CqBI)�J�;[��J�NT�z|.�i�9���6�ͱnz�Vmc������փ٣7�͎��9%#����%�Tx�b]�V��� ���ɸM,���6�����i�b]����ݼYZd�}v�.]>���Uv˚Қv�hL��S7��5��H������Y�/|x$�hj��(1�ώ��5�Vr���c$i�?��gC}�<z$��.���x6�3�l���{��	 `��No���Yi�zϧ�z[���O��~ ��٭��e _�����(&Et��U拾�JO�=o=Nmo����K�+l�b̈[7�D���b�3D<G6�s��h���l�K5��Y`8�n��5�c�?�q淪����ҲX/ZD�5c"A����0�m]�����@}����k+y������/��������[~���}'6�Y,Wl�]�W���cɊ��r�_�56C�X���3���qK��j���֬�r,[�5l-�����^��������5�f��`�lU2,�s����z�e�/04���B��h����Sم�$��R�_]k�d�ȀAG�c͕�D���{Y�*��A��}�j�	1�����̿�q�Ӝ�mW0�m���x�C��)�<��w7�sq�x���R@♕X|"޼䫐½��t������]�{�bT8-�SR؉ǲ�&.H���R��8F�0�)&�;��R���j��;�t���� bc�#�D��2�b���w���{'x��dy�_LjYe3`��eW� �A�8��Fb��Z�!�gY�m�����b���Nu��Y� ��I'�ֆ!�0�����Q��aa��g�kا{�����kK�|�O1N�	B]Xқ�}��XGs�d ��I��b�N//�gA���o��� k݀�W�����35X'����VL٥˕y�8�ը�ԫ{�\���A�P���ey��s�s�# ]j�
x��;�I�*�z��֤eԷ��4��0�j+�
a�DI��zb�p���'/��P���Cq��T�a�0�Xc�𜖩F����D��w��K��׎bxYԣ�¡�b��8����zT� T���ϠzY�{@؟}[�T�e0��>���66$۵��X��C��eb��.N�������J^P,�\j�e\���,> -�j��Lo�+� U:�;#Z2S��G��ش\P�T�N�Z��tF���Rb?�&Eax���P/�؇X��e�j����G��r���L7����4���]MW|>�B�O�X�
f}Ox��Bd�9uf�I�<Y+D���a��s�o��C��<S�S^�M#�b9K<�����L�A+��k���4�׽+3��m3�$��%���ϱ��&���!�=�N ��{�8� �h%x��E���������r�0���^�ܩ'V�&{�����T3T��޶��r��e�X]��������1W=;}=�d_�h�Ax�KfųeD�lj��S�z�<�0�:WS��Oe�0P�9���X����}���]��o�o`Tz�q"�8��pbW��~���TO��FKT|�zr	T��ƭ,Gޫ��(�O+q<� �L.��=av���鉱��5�J��1�t��6��a��0���8������@1�s��RFn������z�!�a����T��5���H]��A����3�{���QaA �D���`f-����uk�	��K�qd|N��dYT����2��N�+�D��.�����7���.iA;���xtX��������~l���;��N��?=�[�g84Gك�_Mt�ZC]���ݤ(�b,���1��L���r����<{�O|9��s���5�.�;��G�B�ƉU4@6�1���>יִ;��0_os޻�����*R�O��0�h:��To�������3族����G6�.��rVCUV6�,{s�¹�ɋ����� /�O��������_�Goqx�v)B��R&�! �g��(��i��`m�g�)�[�P�*�?b>�RQx1���-���:�gCh/Y�3T�Ѵ�p��h�[*��������c�׈_7:W�W���hh���5��&*���skm*��v �0'op������7�s�!F4ϖ�'#9�ج�[�!��+�o�+�8�r4,�@`�M�@��a
/�Y�lӋ
O�!a��������l[Y���|���x�-��ϵE_���*	�L�G��8��s`�R>����.2:!g���r�a�ՉB{����~��%
�j/4T�/
�7��X����,L<�͒��g�͉�����Y8������%i�"��rv�FL�� {+�v%���(��u�;]���$r�,|E�Z�3맵u����E+����'0�j����P6�nx�Ȁ�PK���x�$ �44�Iv�`�'����mN��1|LrlQ�n����0"B�	G k�Ѓ}�������z���/��t� O�찅g�A���//�j|��
���&�_�y||��v+��Gyy���n��|2��0�eMl��s�[� 19�a�����`U���ߗF��W2;�d�׻��&NV����0PC����/�#��*�Z�)�r*�xV%d�Y׆����N����n���N@��ݔ�9���?���A/�6��p��N[o)�g�S&=�Zjhߑ,��]7x�}_v-X����
�m����^��1X�z ���M����^Y0��4���l�3JyR���Qv��UX�d$�8.��ƹ�4��,�B��-V���c��9�P��x��!���Y�����w�k5<�<=<����7Ǔ�2���l&+]0t���O_�><(ƂZPN����s>S�N�M�Ps���3O��`�!��U���O�6��F
'��M���x�0��}�PR�I��vl|�]���l�֙]|��k����@���L*m����K�z4�-�G�gHK�{������������*\�y�(��C�L��=�/z��<�N�1-ۖ^5����>��&��3����٤{���i8��^]��vC�����OT����j�Ow�l�Sc`��ӂ�f�^�a��F���Rm�Q#��s�����-Ԭ,�F)U�6�ֹ��6�1�wF�.#��,�YN@�d�X����0�,��W��ګ��Dn�n��Uo�H�� ��T�d�����Ŝɔ���E�{�Px�>'��P���?6�ӼIOi�G88�G�Xo6f�k۟�sn���6��r��8GC1��C�=�i y��͐ѴT�Ճi�xd%/�8�2U�ޕ+��1:1��?~�M�c���λ�D���ٔ�DÏTz+3��]!�xĀdlT(F�a�.��zd�\�Q�W˻\�ݞt�\�Gp{s#+��u�Vr��E�h'�uCSl��ޛy ���i����Ȭ7U	|>z��'�4i����
�zv�tj]p����I���5�Ȓ�@�!��M�}S/���V���=��9��
%h��EP7�gq�q��$��J�q�lDh��]P����,�*j����r��+HX���ʊ�"�
 ,-�@� ���0�=SW8�2㑹G���/��77�H=����9�N  ��ڂ"����M��p�Ǐ�~oƭo�k�`�тg
B�Վ6rF�
��z���J'$���S,Q�J��&+�Yզ��^�z�U�]��ӓ�u>n��]�4T]���Z���TKf��Hb^z�䣪0�7�������i�O���7[9?��cY����!��:���D&�%�C�l*�r*��Z�~�J���������6lMY��N[���˚�[R�I��;bnM��l��F.[�9�R~�ʞ`�N��6=�y �YO+
��W'2��8��<Q�f7�KO=�����m��b���h���t���� O^Z�p�Z��u�Kw�?�-�j(�򮜳����ZOW����Lx��#p��ky׻�H�A��XS6�$,pF3EȤF�N�����׃.�s��N l��r�1t��x5�/��ł �8�4Ԃ���B��bv��z.�l!��E}䓾w�F�<:<xt�ֳ��[��Д�$��hԯ��G��`��ֿ���;dI�k�ޢ/8����VYay��q�%�|�6גX����γ��񿽾ᚂ��A7eRc߮^ޛ)�Z���>5`8�`���u��A�Q���ƷfL�0��	��`U gf­-��/Be�^;�|������	N�U�>��:�lW��v������պ����2J��L�Vk�J`�������ck�=�w����Eԃ^�����˞��roQ4�F+Dqaܦ���5;_/��>Qe��!��1��Yg�YW2�l�V���̔��2.�M�R��ɸM�sӍ��	�r]�Õ�݀k�^"r0#�W̋+Bƨ	��7$.,c(R1���$6��Z����oo����
�#{[�xQ��%��$������	�N-�#���ɰ�ڱ�����漗+5P�+y_��'��ޖ˘u�V^	�F��'4ew�﵅��r1�`a ��u�x�A=h��F߷��gѱ�*��uwE�M�;��W��)�,�_?�V�[F�w]���	��∧!�9gy;Y�Y��;��~#O�QO{.�F+h0~4X���2fz�������%�p��u�;Y���xo���k����%��� f�P�aiL�c��r����&��ï��ԏU1�ߝA:	jjDw��ul�h�	� ��'P�R7-����pX�p4�}V�W�����0���Ğ�.H�`E	��#15T��Jƙ��<B�$5& �= w�C�*�W�dB!���:��'�����3?�x,Aҹ\�gr��(s��!T��oNj���=���L(� krA�{�k���볍щ^�u==���P=���C|5Wc:���odv�RCw%|_�t�u�*3�O$i��	��U� a�y�Fo;��7.�#�� M"O+OYG?Ğ"{�u�� ��βq�Ntv<n���?���R-E�<��{����a0c�驐$��7�%h�Zy�P���!�غ��x �R_�NW,�B��_zk��J��;��`��M԰���t8�����%�r`D���ú��L0�x,��-���xsE�EPK7��A�r��2��lʽ1��vt�(0?��FNj6�'�����ƛ',�)u=�Y	c�뵞�����G����r�A���I>nɶ��[D�w.�� �AR���<z�:� �D���A���������ȼGf�;;�B�"�e+19�����;��;&D�Fױ✕~��C+��qA�V=��z=���������x�޼�poI��^C������n�G�<롱�ɗ�/���d�|��'O��馅aQ����D	�&4�F��2���Jㄤ�̂zB��*n��ab�0O0T$HN�.�����:,i��!�B-�#����~���=��0�<5z���w|�����c�er"��Uc��ګǷ���9Jq�Qȍ>�#DB����������T��HpI������"{1��nMW��� ��(u��h�̺[�e�L�E�g貅�J��1fK��A+���<}���L��`��،O�1\�5�h졃��?~�v�_d�*Ȯ����.�4\y��B��F�~����J����j!K��ۃdu�'�^"������G���e9���
��3߽^�4�a���{֌�\>YDd-l0<+�q)y�٣��:3�B��1�5�������	�RÍ�����^�=y�]�/�72��|P���A�'0JZ�� �p��^2e�3F�3�`? � ��� T;]�����6Ι%f�0,a�}�ec��@SW��`�C����hkw	j0Md�4U�~^i8�d�����blZ��0L�@>]7�5�ww��net�O����B��/Q��u�!d�J�,�&�h���O�Dbמ���g]�B7�jL&�(2=:Te�� �Y0����{$ԒZ�Y
Qc5���H"a}��OP`rR8�d�[�_��V�9-V��i�uOL�L�k5����h)&��6zg��(;���{����X�����t�!,.����*`��
���+�)e��l,9,䡟@��b��F`_���b�4�O9�%b��^��^%H��wS����W���b��+]P��[6-��q�g�~�^�9�SG���a�Эe@=-��亞�[���M�n2W�6#�C��I���8�@�}��<�
�Kr`�5�a�+��U�dL�.����~����� 𰢹K��;�AC� ���!�4bXQO�������k=I�f�` {���T7�n���?J	=�7k����zl+]��^�<�pdQ4՝ #
��0�ʏ{u��/4�tl���J�Y�P1C���	ei�g{�&�����d���ьĺ���Bћ���{��Vu,47/x��pu2�{����]
��4�0n�x���a���6[9��̎�0w�y��A�l�C^��(�9S������z�$�j@�ׂ�]Y5B[����@�	�]���'��ٌ0b�6�6i~��bJ������)�l�7��{/��$��%+�����dD*�����%���P��e�E��W5�}�ެ"��Yߋ�G�V<'����\z���3nxQ�!W9�0!���Q�Q���[�S`�ul�^Y�G	Lz��Do�*!xOa�"qAc*𰄡#�rpB�uS,�p,Q梋e�%Z�z_�]-������]�����'=��v/�A&(�4:e��z0j0n��n���0Y��vM�����x2����J�.ƥ�~:1� �$J�BޚY��y|�n�������ɾ����X3��7���� ���[�YHK=�s�K�"=[�m���x�d���lj�ԺU��Z
�@�b�&'������_�{|�+}���R�\�%w���}�,/H8 \�{@�~�/���쬔
O��"@��'fq;��^@>�k��dU�VI=;����Aui�����m��:�H�ueee����ذ� fx,UM�8*�b�������W�x6�*ɘ3�&8l�y�r"x���
���q/�s=\?��\�����C!z�k��;���M��e�������<Y��Z^�um$5�(�_p��>��AL���=��t�����:z�a��p*]W���%6�·�D�d&�
����U��M� ;�������'��\u4jp���O���;Oz]?�j�����O���qs�κ�?[��c��"����z�W_���xS`T7Jf��i0�T�,�i����[5,0D��k��w��	
��������J'o

�n�Jnr-W
�����ƫ�'%�޷��ota"};[�B�zх|��"LR�6���4�n���jmiw�Rb�_�`�0!�'7|c�� Wh|�w��)@�I�%4 ���� �֍��ނ�tE^��A���Ga|�s=���B��?���Y6�ϒk]�7�z27r�C\ȾT�Zy��cj��%�U*L��X��D6���4�e�ĺ>	,�l�D� =���ES���eWz�Sr�v#�f���;[m%_������$��J~�}'ǻG9������ֈ�E�1ʳu�F�6�!߲NX������5�oO�Cޚ��lFϘ�x $�|��0F���4�p��{��+��6�S6�:nb��Z#��u�!�pF�"��h*/��u#"x�Cz��+ԡ����g�a���vZ�p�� �|=G낉Ʃ��s�n�N�op�@'���L&'�A��> o<��z�hE�n���h�tse���JjHȧQBh|J7ݭ.�ܡ9'(���j�F���X��L�V%�G��z-�� E���D�J͇�J~Ұ�.�_�ߒ��fE�~~#t����:��n�y���ڲK3� �iQ�:!3<ǒ�\���a��NI���9��[�Y}������I_�^(1�l���y!х�ԅ�N�%;���5�Z��>ox$�L�rx���1)�W�xk������ E,ks��4E���[]��Q�%]�E6Y�L!�i:I�v��@�\�d}{-�j��ۻo�j ����Rr�B{s�ӻ��<0//�<���H,��Jf��I'��:�X=�B�%_���ŀs�<.HF\����{,��Ի6�l�[B�H��a��_c���3���k8'�O���͛e�؛�gL�S_��:cO���=���
�':7v�\�5�[���<zA�B�{���,f�r���|�C|YMI���\5�l�c�ըmv�LO�T�z�v�����T����FB�u�0v�U㋵ Fő���q�� #�_��B8���&IUÛ'�sFCo{�m�j�ɘG*S��}���
�֍}�
�1����<[V��l)�h؂������Z�o�Gg���ʡiG4�Eh���;xna�_�H��3C�w:��Q��7�ky���;���8��=��]x���yB�w��`q��n��u���}z�\2�`3n���U�԰��m���*&�j�g�N\�"����߁��G6IM	�A0Ҡz1��-ԃ��F��g��a��A���LtN��g����J7�X�(Ga70S�b!�ą���x���5�Ԑ��n�`�����nʵn�:^��-c�U;݌��[��c�IA]4��E��s#����$���F�i�v��/,��P����^"6�T,�f�oK01��u�2�IÒ�'�����P����T%���!)ݜ�l��"*���ѹУ~ޕ����`\��Xo�������1�5��A���s�؞axO��3,F	�J�jH�nO�L��k����Z��!s�^�kV��L�J?��!�#��%�l����C�f�;����P���NwP~�x�	ɢ��ǭ���t"��߽�!p���Y��#1ɉ���A��w�`�4s�p�"=�%�V�Ђ��G�*��/���m���y΍�_z�a�"W�';	��Lo�w�-���_�~�)�i��
\��xNNzBr�Ϧ����),)���9p��cT����
Lq��?��/�@~@���3`9̚B���|rz�� X���J�	�X���Yo�7t�H§�r/'6.�ՠ�'?u�
�	-�y�.d=	�Gè��wd��!;7�`�����Jne�F����ozWเ5_V�U��(9>4�q\ϓV]�4����0-A�t�ql>l��zq�Ylܛa��'�P�dψ,S}���$�_�(�z�7K=X��{�dyX�t�'�ھ]^� �|��L��5��X�ٛZ�΢��ܻN7�n,$O,I�0C�P���2�-Ў 8�d;������J-�����:?۳\���I��O��j�xD����`�4���[�?�m�5D��E!a�]� ��)u�&f����u�W�NM(ݪ�f�_�[�����jDO��^��UT��iy�D�FG�Y�Éa�kx>�e	�L�ª@Ͳz�S��+�wY�bp����U�%�S(�Ld?��a�p^Q���8U#�A��m�Pb⇆�g@b	 �|��j�#Z`��ut�L�D���0NM����A�	���3��w��^���������+ݠ�u��8�1����C�$�dV���d�OP�d*�0~�ۼEp�\ZǺ;Y�}��_�<�9BJ���.�Z7�l��I�j�L�� gѵ<��RO��.p��B����
�0(����N �_�]+X,\��ɣv-�~CCgN�g6�&`,Z��7���E�������s���}h��L
���h����D�R��$�]/�D�«p��.C�'O�ǀ������,A�7;����H#+
�ڌ0
Y.�;6aƺ@#�0�s}���Nvj0�@��P�v�!?/�|�ֽ |��B5�A��䰈+�yZR��%/�/)�m�9�	J�����R=�j#wꝽ�Y4�}e�B�`���VȽ'�]s:�Q/�5�"����q�Z��A�-�����'�?!d=譟ڣe��_�ԋ6�a�֍x'�B�AwS�FC�	�i��:Z��?�\�պ���0Cb__�u�)�:ڽ�7�UA¨E�
4�3��B�gJr);fqX.�p���i43e�0p<�T�8B%��[��1��bz��J�6���>�����an�t�O���-慑o�00���Wt7��]�4X-EϮ8��[�y��<���0�=>���2E��p��ܳNH��6��}y~${�˗/�j��^���ݏ����,2�
��F��F	KE������o/��PL|�#{3/jL����&(	um�R�0��Q lB-�i!�X��A�Bh����P��
/���z0P�<Of2>��R26L��f4��
�5��Pǅ6Yi�E#�,ױ_���@���d���F[5�z��:޿�~�k�s/����"PM4,d�p���
Y���-m�(l��z^Qd�r�'-�b�eHM�?yØD/ tB�CK�YG0�W���,y�Њ�>�~f�gk�E��n������:���)V#	���,�Ʈ4t���p�ko����������y��Kb�E�#�{fn�T͂{]{�/|e&�ڂj"	�7Q��2���F~�{G&�"T�9x��"�7V��R+�(@�R�g�d�vf�V�����V��-�h?�OБX΃�AS��="��fFi�Yߐ=ab˴�ʚs:N}mN�����8� ˦��}��gsY|Ǆ�,��l�Ɩh��R^[L�|��'�ӡq���T��E�B`C�D���$�B�.�:.%�r�b$W2�&E�2���,t=���@���a�Dnn�X�7�5���͌�`?�$3���q�(������Z7d�A�Xܨ��&�G��fOp٠0hfZ�R��,W��[�ή�l~\�����qg�R'|ރ����є9�7��j8����G����X�cy�<5:~���µ�!��o++�A�������e�R$a���1��=���^G��2?���F�<[�:���xfu.Xĭ����(W7k�R����>��L�H̺��pHӳLk;�ȳ�Ȇ?�@��Y�V^L���LO�e����O%��f���E�.Rjq����>�Y�\�D�wI�@���D�����Nc���Χ��YQ�c�o=�Ԙ�:�' Pu�����|�nHZ�<���� <'�Kr-u�Y*G���~@��~{v�V��^�1*�j����O����[�|` ��t<z��Jz��)P�Vsd�W\S3]X�3�\ջCV}��g$��Q����{�U�_�T��L�?۸�s�ꏡb����T��Ȃ�@cj���Z'��Ȃ��ɳ�0t<��z�̲X����ΐ�a�V26>i��P�Z��4��~����I=�B>���굮`b�Pm���0 9��:�i��ߐ؈&�gd� ��0���9� ����0�˚��rC�1Jq �c�������&,E�$�������JSsF����5a�B�(�t�͓�[eQ�[iH���f�<�i�J�u=���1�ձ����7����~w-���Z��y;Ȑ�jy��}EM.��� ��'�s~ܐ=����
U�3�̌���\2��H�agR�-8h=[�;�G��{~��%|����lW�ި�R{UJ�9B�D|�g�<0�G����j���GHA�Q�,���p���SgeR��&�d��7��B�Wy�i
�b��)k ��ÞXqw6܎
"��jIN�w�m����`�a� w��ek�����![�'9�Fϒ��@���O�aqO�w;#Л�ߙU/Viҩ�WoU<�/EȈ���h�H�ݹ,�%Q�����	㻘�y����`�Y��Q�L���b"8�R8a�h�����6n�~5 �)�������`��ehXI�o�샞�X{px��H��^Ð�5���9s0Q�UO�]Q���Y*��d����9,"�BX������1غ?R���^�Y�S��j	(*��}~��:MO���¤c`dq*1s���:�ZP�x�M�!"i$���@��b�o����4f�9��"g8����www����%�In�􋅈争X���$>��u���,)B��~>�3��w8����	�����::��0$��?������^�R���X�Kc@�y���S!n����w�|�{����]�)/g/�kf�9ƺ�q+�d;_��Ê��W�/n�.Z(!:s�p��F5`�T%t�RE�* t��: Ƴ��5��#�� �b��Vg��Om:dSB#��
}N*�h ʀ�m��l)1t���'k���?�Ia�cPY��m�,-s�L�0��O�Ճ|ɮ�b:o��B��Ϊ|��j�@��a>�a���Z�1o�gSn����J+��qQ,]|��[_���-bu��=u�?��X:۞=�������3Fa)z������L%�n�݌�4��N2���N+1�Y�B�V� xD�Qț�r�'bdDM����`�׺�����P��p������G��<k�#���ŀ����(�����/���͵K�$6Å��f��	��.�3�����z��T ��zƙ��-��G5�,��yV����0d�|��1�*�c�։.�3|����===9�h;xnы��L��x8���p��>�(.���!�$��˙��{%C^�|��@O��d����:���@M~[$t���T~X_�1o5������zS�-ʞ�B���b��y̯��V7)���O�mxo�ct��0u�^��#@l ��v09l�PK�������'T> <M�93�s��z�;)�]����1<����9�h��$�q�"!p:�xh�ڢ�~�IB�I��	y��]��[G�CXZs%xJ��:v�!b= Q�5TGD�l>��U9�$f�䚗(�������0�	Z�L?��f䭖���.�ɲ��AeY�@AR'�{T��qa�k�L��a~�g��[����S��{��O���
�	��
���P�x';��
�Xɍ��g֘Lt��湯=\��^^�S�e6Y�z;���a��t1 �8S\7г�d	�g�H�L��'���.4����O?I9]qcn5��[�\�	���[�uN@s�)t�6�����V(������4�=5�s�1E�Y\�RèA��-��w��e�"�V��u�K��K��0zq��]�u� �6���G�߽Q���eCc�Ul�քI(���\k�Z=_R�ꊌ�)3|-�n�i~X_�T~O{�FQ���ck��'�m4��ֶY��\�����o������ѷjH�T��)��C���P"������Ǌ���|�<���S��\v^��R�4ަ
#���ai`ΕU? ���ۂ${:�tֵ>�V�ޙ��l�,��E��a��ؘ��
�E�9��$:(M�`��6AAJ!�a���u�35n��\7�mVԎ{�k�����Iu�d,�|�M���snd��m�:����õTY��\5�z˺^"��Hq�>FL�]h��zi��h59Y.\�	�y����Q��?Ӹu�\?r3l�x���-'-U0l������S%t=,�߻VH�dK�\����zV�T����B�k������	�̾�g=�����N>t�N�޾�w�ox�H��\���)�ȁL�^*�ۡe+}A%�e+{k��4�]�g����ֲZ�N����x{�v�����pzY��gݐ0l��"��v,�j�S��-�>jW损�X��l�ˑ$	#�ր�ya}29��	�4�H��x��>�!Ah5s�]X��V#�<B��S_m��g��T3V�d"��t�͐`I�%^�T=�:O�������`�%��uޯW���ݿ�� �ݪ�TO��w?�R��TVV�o�������&��N�e�+sbҿ�͊5��A[��	�R�8�I�N�\{���X_��ԆvOSc��O��`3�̨sqM���2i�[��o���4Ww��23Ľ	W��$c�gu�/ڐRH�^]ɭ�,�̚%n��В=;е�:�>�9���B��K�K��L,0����-�p�	�'JY�\���Z�_�!g�7˴`��9H!�6=<c�W���R$�/>�Ÿ۷�_�.Ov��#��5 K��F��3E�6���|^��t ��y��:ܥ�^����!ˁ�?�":%c�����>\���N��~���~��(���1@Tԁ.�ؼ���%�Y�&
4���&@U��U=x-�2z�r>�6����s9�����5�@��Qc$���q���yi�c�b��*jD�REAe ������y4���po����$�l֩�9� �IG0j�����!ݪ�"�ίË�g�AWkf�9�V�V�0�(�nu��	2J'�\�w�`�Q�tN<c��R����g)���!�P���O&���V�'T;9���l�y<b�Cc	,R~F�sMb_l��t��ܘy�c�s�7i/Jp!z���u�lO}���]T3��?AB���=q�U=e�-;��RQ�MQ�pN�l/�klz驅�;Cs!}�B����^��ǫI�A�5웬g�������Y�[s�޷�����afY��3�z��jY��ST��y�wv�.$������L�M$�p�!�X���]��N99u��Y
'����sWKS�R�m翽�T�[�n|���Ԩ��46�e�<[=57���ڤ��Aʮ�b�[�U��m?�L��ڵ�t�����蕞��x>��8AfH�r�$���Iz���ݫ�k=�:fY����'`.�9��"]q}  ��Z�`� ����F�]5j0hu�>.�mہ���~~���ɂ ��KS ��0T�P�Ǥ������|����^e鵽��A:�;q���,DĂ#�Kl�7�Bw�'wl���:[��
 @�C��!B"��uCLuu�c�$������Go|�#��{�����롪��ՍՀ̐}�k��?���}��j��s��Ut\7F<��'�t!+����%���e�:�s� |j�l��e�3�FxEԂ5�=ꀖL�dkx6�ɕ!S�H4��.��0h��R���#Ja�u�lE��a�Zx�ꡡl��9Vsyw���+=��3�RϸZN��r�a��߁��ʲ�$��,�G��~w��8`���F>=>�="�ѐ�nFm>���I��Hc�:��+�����nt/^���"���Y:�d��y�dk�#�9�#�����Ը(�j;*<���FxP����]�)o����G������7����m��K�z#�V�i�A[��H�L�ٽ�N��L�1��,�_D�V��ga��:	/��_�<�O?�d}���=�p³.(��t	��<3�Il��3�q��_�k{f�Gd���QC8�-�O�d6�`+���?�L���ȟ��㢶2 ��	�������;z�q�,�tx2���H$4.,:�r2&p'��7TM�^�X���4Q��F�����@2���T��KD2�t�\��2eKAh�]��E��t5��n��|���@/#dw��ҰQr9���� ��>��O4Vg4qy4���q"nC1�r�p	J$_���dYY�k�J�k8p���=)A���Q]��s����UN ��0���y�M�����~�}AR;�R����r���J��(4h�b��q �O��YrӲڢ4�t��%�%�[����3�*�o��<����nK�B�[k�5�sb}���P}w�߿<?���Z/O�q� ����@��։�p��G[�r����2a��$`z�����~�ð��4��[2���b��ɸM�7�FH�Y��'�"��S���>�8iw�A6�HS<�,B�K1+�^. O�wd�[a�e`��NQJ��t�uZ�+V��<�{:Hu����� T� �i�t��ǭ�yײ̈,j4e����c	ӧAg�jYM�X�e�0�����nff��`<#Dzx�Q�|�ʱ�����P�����_�CZ�:�٧�BLzi���΂2���H�qCb�T��`�{]jH���
E�{`q~- �xsܿ�����O�)��  'P��0��w����q��������r}=��zۛbG�Z�[�6��Ywh*S���B�e��,�ߟ��-�<��{�8��?�����;�ײZ_Y�]î#MKW�g��]�kU��N�k�!���E�u*��h�ބH�6j�1]�y8JeV����s��I����-{��Z"J�~pL�ɸdb2鬿��=.����~����=t�ZθO`�kd~Y!P0�����ߘT�}i�J�=����v��|�kL6��t9:�ف%z�"�=9��:ƱRG�s����WbB�hۊ�Ԝ/�,-���ξ�{�&���y�m�����!N,8_����	��a�~<N�G; ��Vj�G��1�t��"m��M��l�[x/+���f՘qk�wRw��B�:!���K}ӄ�mL�Ck'*?Y\/^�l�z���Pl�ݱ�
7-�DI]�0j���
��FL$������*���+[���VZ�Ɏp�5���֥�q?��� ��ˆ>��O��P��ᆘ_j��2��z{D!�m��xꂣTٸQ��x������n@�A6��p,�t��nٝn��)[�y*5����u)
2 �� �wA;�ȠGm(�n��O�~���&ơ����i�C�� �8�J��e�j�ݚA�c�vX��50l�5�yZm�;㣣β�umz�����6[)N�y]Ty4��)����3�P�َ�W�ǠNW,�Hg"X�NV��zg;}��H����Z����fR�`Ѓ��5VyU:�-O�/@	������X[��P~����GO�����J>�X{q:II%d@<0�(G��	�0x�\���VLф^{a�A��E��m����:�6��|?�N]�l�~���g�/�io2�"2~�������A0�e_Z�%���ϐ=�-�ș)k���λʎ�$�&GS߅N�Lm:5�b��f��'�|��wo?ȇ�7o�I�FL�V�N�L&$i5��f:�\0���p�3�D��y���@d�w�X�� ;��^v�����?ȧO��ݾ�齮��)zA��j��#v��p�2��&�v���}�ԕ�)u�D!c�cw�FUC��WYX��$t������u[�ۖ��i)�κ�SC���d.�J{��z�P�`�G�b��b%VȺn����k�`���Uz'K5�� >}�J���=0 w5���E��o(�OyG6��7����t�α�a�,�Op�!�� ټ-4j�����Y�2��T�S�7�<�A/�k��4[o��;u%E/	�ª�Q/�\O|���������{�
��O�+�K��~I�EeʪX��G*X�u�7=n�4r�A�M`�����{��Ǿ0�HfsY�g�εXH��4ͤҽs�{���T?O��5Y�$�K�Ӧ��i��d��`}�q[�Q{VK��q�2g5����I:�-��:n��z#��\v�z�z��8�u�4���Y�P䨨��^01E���LY3���?�8vtp�,\���;������w�����������uf�z+%Ib[(M��Æ�io��A�Y�F�����Ef��(]��g`l�����p��JLC@{�|�{ʶ{=���������W�5��
�U�}0>rA�q�7c��l���`�b	ɮ���3�j�L[�#9�%�+3�bU�[T�t"���8�"����d+;��S#��r�	 �N7g�vo�y颈h��S��� ��Ԕ�QO�9ORx�1���T�Qʑ��3[6`�qo�</p����|a����tgR̬5�u�,Qo��O���Y
��Em5���~��C�I�-��
 ��ࢉ'fr����t6sr4��+aM(
�Q�pD�&��)�U�Ƥ�� �un2�Ǯa/T���v�P�s�QV�2�^̰y��'y�):�fx��d�0~X?�:���7�"���&B)�r���t$������.Y��t;��}� ' 4e	��̊5j(M��c��8Z�c{��/�T�����z{u��֛��i� ��)x�7O:d�fݸg��.z�e�ă�<,.��80�AZ�^�o��7������F��Wj8����V����񧟙Uv��D��U����cbqƊ?��Y�3�];�\x*�Սܨ�>��tN��`�A��	��?r�FV]��Q�������lY�޷�	i�+��#�#@� ��'�yA#� B��������k҇�c�~�Z�Dd����F!qo��s��k/����No�MA1b�B����O��xd�,�ǝzW�h>��m���)�u#)��=�y/���˼���}Fw�J�=k���D;<���/ǂ΄�*�6Sj��%˕|:�q2ңKd	*c�D�m>�ƶ~��\��������ɢ�䥖7ɸ��>h�k��9�Z$o�K�yH�О���B���M���٦K2��*�DXFX0+[O^D�j���$����:�H�$nu�0�����3i��V� �y�M�C�>�V���v�2/	ܻN�m����=z�ʔR�w<k��w�er�E�AabY�Ģ�8Ⱦ�-�,P&�y���wV�C��B�I���'�F95t��XB}�O
qY�9k�*"��޸�K +�)��(����g�E��Y�pYxK q�����v��n�22in�<�U_)s���`闼D��z�R5������+e.�����>�����"S�u�:O35�>����M��3�k>����6}�<�Ϗ_Dw���ח�t�����������Nȱ2�~�!�{�N�I�#�Gm�rj��m6<'�����&c꫐��f�eh*:V��{FIa�3��ϖm�3yzq�T0�΋+yV����9+�b�ZGƤ,�i�dC~7Rl=�뜭eX��Z02�a�bK�s,�X���jѪ�L[�ѹ�SӜ����:WW)����\n�ȥz���s�%f�e��A��7}1��i�_Z��c���sjP��]�Õ��j�<*x�L�&�8��5��ѯa:{�����{��c��f%8˔�7���@��e����Û�����l@��!�E&/RX�Йޙ����������;x���(�	%aϸ�r^��	�ۅ�s�Vi�Շy_A�״�PGS-�8�.�Y��ϬV��f'0u���)������L� ��lHm�N��ѯ��$�"�LY�������Ȱ�tB1D�6�j�{�P&0����j�y���}��6�����OG�x�A��w�7�tg������Twm���b�(�6pKbZ3���v�Ho/���ޥK;M�|J���]��v�fp�W� �V>n^���Jo~�&]�b����(~��ߥ�}2�V4�G��l�p:w�F}e��G�[+E����ӓJ�I�	�/6�"��bX�k;����_��FcwRD.> "��\L�M�D�^K�K�}���O����F}��,�(]s�̀����B�̇�$9���J����W�̳�5�a��?��?>C�δ!��/���5�'Y�vT�c����W`%���u*�c�f��I�=��r3��;�>\��j!g��������}�d� ܭ���rfe��^o����@+w�N3j]@�)�yϒr�
HP&8#���}ɑe��L�"��G���g����g�Iw�]��n�]1l��>'X�:k�dNĄl�,���*�S��k�,������u�w�H?�Q�|!���{ჹ:��>���b>;�;���Rib��%b��u��y52�*̣S�>�҅ ?��x�3��B�,B@�:�h4$�$���oӇ��� i<X�%�^�P�,@8F��f~%#�o�n�;+]��$Yd��;j�z�=���>V��e1����������I���eXY5���n��A�RE����'Һ��4���:�#3ğ*L
���?���h�M�RQ�(k�tʏL�����Ґm�Z���E�s��]7�U������y ������6TfŬ��4v;����/VB��3f��9��<����l��t!���CArC]#f����>�<�'Tf�z��{��ש����>�Ab\��LyB�{�-��҂\=u��gp���ەL�V
�no4Y�y�����Y�Y�A<WAs^T
ݗ�=�!�����0=����rQ0��U�CIW��"G���wqOa�����s��k@�u�|Xs&�������R[p<��I�|���o\��>�!J��t��1�|I���~`��џ�0��T1�g���|�FIܫQ�@�4E�^�+'��5�g�H���,����G��ܾ��tm�(��"����ǩ�G��� я���m:���l	�Nm&ZPGf�&�`��e���[��������H(�RX�I1U�xXl���J�{+�Oi|{!�	8��r����,�n/nR��r��B�f�+Ed����$Z��|Q_�L D���tuycY���|&�đ�c�K�ԃ�e��� D��n��!H�R��^��yum��|k��9p�S ���\�w�s�0��d�A#yFFc[ezs�=�Tr��,]�a���G�(��f�ń���s ؈�RE���~�g¾����-�$G���������.Mn��\��%��_"�4���|l���>7v �$�d�괹���ݧ;e﷨RX����U�u��d�yVI�)@��y�ON>��v�:�$JZ�Iަ  �	?�����=*8H�ߍF��|�d1���Y�]Z�$�YL�'Y��ݑˌkY ąOm�v�=מ����h��_m? 3���S�΍���z�d�Ay�Q� :��V������v��uh�iB��6�L��"��R}Ad��#�-aU5.����W���6��ͦ���wN�q�">D𐁁h��cGYi����ǅ-(����en7�\�E�l��v��\���tm_<7��ŕD��'5�8q����(�K�~�J��zds��N*`r�A���S9���<�b>�Q�-�r�Ȝ��J���$5X��p��L��)��I�rC�`!�"�d��ܷ������呕tٰ�"G���v���e��W~�K�B���4�}%m^/����� %e�����g_3,�7gv�g����^�}�FK�<�j�b(�l�Ц�Œ� �_6��U��`V��ӟ�\�"I�]���o�h��`����Y�b�TdM�~*�e�����U?��d��D��G�~��R�������~-9����p�d�W<�i(�hT;A�ʀ���=�bM��,;�*��e��r�Lo�`}w}�?��_ν�S��lhF�6U�������}�❢�J�Zp�h��Ad�/�2@�L�q�OS�|�%��:�a�~]��K�J[��m�i{}�sM!Ћ���Z�l�C�ݧO�����ܺ8]*ɫ���Ԑ\*�F
]�4 -�������Q�i4M�(&O�ĳ�۬�yH?=}�bZ�Z����ΐJ^����
��SX�d�"j|:�i�SQ'j��;Ґ�G#R7�CWV���|��K��u�8��xO9�pq��UM������el�B�P��z"@�=���x6	��6�x� �;�|Å"�M�G�s�}�1�l��ѿyp��I���+i#�W1S�(c<a?'(C��SY���	DL9U�Y�K��v��&u�\��-B��@)���E��(���e���`�����rI�e��y+�vsi��r��k�����+��lr�<�MA|t���ʳ�7�j��Ѷ_>��x��EF�׷�����\>��^�J�����{�8ɒ�9}J2��Wt��wr%j��&}����!�}i�Ke�F��0�>�_��tx `gvPJ�LU�|�)���>c��/�O^d����WO@��I��On�+`�./,����j+��g�_O���(<�R��:�n�ұ9��m���;"	B��w�`>��|W[�Q1� �������Ϻo�����V��\�yE5�y�>��F Ք���G���e���2 R�no.���O���yI���~z��>�_t��'�\�vͦ���o���2��3�bN�k�>?�l��q��5�P��9E8�l�!'.	#;���6�M�#`6u˾t�z��蚉y��ǡ�E//�g n�QR�M���|�^dW���H�/�~��<MZs��e�$b��,�?���9��_z�9O�3��]�����5�ػa[���)C��n�g���Z�W�u��@΍+ܒq�~_�l�ٽ�ܦѲ�K�X�Ȁ�A�ݹth���V�$S��7���=�_t��Yp� �k���/��j>�C�A��N�0�����
��٪���ݧƧ��3O�ѷ,�Vn[��P���E��
ư.f㴰̔��x&�LY�S���0��Nٍxؘ9s���4^��=a�v��Ǥ��q���ah�����F�2�&7Ԏh�^�[c Wr���>���ПӾ��2��(2o�g�~��3��'z���-RI��yn!��E  ��D$�����?3L�vd)�چS�����e��Y
<=ֻ<
 өP[�W���Ս��i�����C�M��H��c+!�-�{ss+�r�:_v��[	�[:>���(��%#�����{a�� ¯�a�5����<��>e(T�F(�I:XzN����1}���5{���<�<m줲M��,����%$�A�CǢ���9#��Y����0] �5�������QX�Ss��$���gI������nP���4 ��I��������DM�&�CT����8�2͝��b��'C����W_��w)F���*}�����KQ�����(�-`0��F��g�d��R�,n�[; �>6�������©1���IĢ� V�T����3�'�@D�Ү��p;d�N���o�M��S:~yR�!���J���%@�G�1@����ɟ|fJ����-�ݯvy_&V6Zp~�{N���q6S��;_W���ɴ�l�W�R�pL��%�Qa�F�V϶酇[�<QY#ǅ�*�l��2���>d��l�4�hG�n8��~��8��;F�Vϝ�B��X;��̝��maYx5�ZPt����� ��ƭm��-��]�d<2p�m�E_�^���w�+zT�rl瘥���+���kO�{�*pЫU��a�j����x�>�.��EZ�fRcpw��y��O1���Yf�ڸ�v�g�����i��}ƻ����K*.U����a/����/O�⼔i#�ʯw� H�r��jXș͐U@��r.ys��Y��p!�=g|}VQ�~���H���X5��������͇��yv��I���vVEx>L���a�]YФ%qX��@�2�B��ͦC�ݫ!�ngj� l�D8=8K�4�`����TЛ,;G�˵cd[31�|N_��`kBs'<�.��I�w�xן�����t �X{��m����}h�@Z`#C,�!KZ�[�dlG{}��ݞ�:&1i��JbA8�T���t;�6�:�,�g"��҂�8],3��[b�m�lݺ�Vzn]�춍X[��j�:����ލcrp��:d�}x�g�u��0{��d����Bz�`��G@����Ӭ�un婵��bY��_ZL-�.oJ�z�_�-ل�)�.��Si�r��H~�L��Q�����Ý�_X�L�Pz�k6��\�O#��R\���<��5hn*;� ��}��G�L����<�)��Ǆ����$��3_�՛�_�M||N��Oµ1�lm�L���+����#b�GD@&�]��Uy�y��v'������Yw�MHjO>7�郓s"5�\�+C�F�Y�����N]��	����\�����*�vM���S	�:�ڇ~��L6k��ళl�͂i@OJ�D��3ɶ
N��þ�$z��m���+1=����͡w:V�2���(%&>Wӷ��F���=J��5|e����Q���j}��G�'W[1
�[]��)���&���H��)d}[O���v�is��Ȃ��t۝�RU(�d~){�܉I2t
��h%�=�@g�v¤��2Ԑ�$�� �����ԓ��q*�^Ӯ;O���v���~���h�S���ߣ.A��ն@�x�K��F�GɈ�u�,Ȏhg�ч��+ڮ��!�thG��2����ùI��@uT}��[y�e	�k��S�ą@6����(�>�*8gm̵����	T?�N���ʰ�X� �0��υ�T�٥�`�*�)Y^ 2qn<=#�Z�0FJ����U�L�N����T)i-�v����?����?�!=��e,�8��d�������K��3�gQX�P)��!�y����!��b�=S"(e��sw,�j�������9oT�KuB���t}�޿�{�I�t�	���s�O�9h�99����JX�g+l;�EoC-��:J ;���malW������l-����Ӛ8	�A�ƭ�dCɰ�썍I���l��m�d-��Z{.iA�|gȵJx���t�����g5�a��a�~X��+�~w���ƲL,c"\=YPK�l�����M����,�Da^>`�  ��AY���C�H%��ﴆ��o��ihZ��sL��d6���ɥ��h1qhʒ/��撫�>�Y�*?h�a����D;��_M\H�
':p��>���#A	 s��37[�V�7=��
��G-��Q�Ue���m���2=W�3���}�̋�W+�"dn�r�P�.�B/�3J3�����9�z�Ʊߟ��A��n��ۻ�R*2́�l^�?�ot�p���z���,���L� t������A9��@c�x�!R���q�	��M�Sԉ��A$�
QbR�t!C�YS+�ma�Ɠ�|��4�3 ��!pe*V�g�d���A/�\�fX�лKΦ@�k0� 
�FL��x�q=���ӕ?WU� �:�
�l��#pgd,��م�{����8���5��Z@P��\���Ɩq�6����}�!M1*%��/��e�o��JZϓT��\,�5O��Q�6�g�鬡G���C���z	�0���*���Ԛ��hj���~��y�J��8X��&n�M���?e�6���ڊS��JC�j�R	�B�W
v2j�k	��G;ZSp+�`(8�<N�Q[�
�:�*;Y�A�j��D��ZA�{IH�YJ�yT�E"�_>�5v�'v]��D��{ݹ%L� �W��ZA�h���1�������7�޻�ޤ]P��]��ұ-�pLY����.���7�-h�U�n��8�pHQ|���~��}���J.n�5#�By6O#/�	b��8[�'���#��7m�4���x��Qv	`Z�*�G�2ĩVV3����Uv�ޞ������S��AGjvͰ�s�JF�2�8au=#���*/SF�ZT=�<-c��ӿ�	m�|�߯c��
��ɛ�Ǚ\Ƥ�|�z��9���}�Y��_�'�Ge���I��K�b(d��32ZĴ�ı_�L��NϏ��(�]|9���F��'�|�&��/�J�X߿��(��c�R6:�{=��5��gv8�I�v���E�b,B��~�M/�i��Z��ϢC�bp}T�:��5#�g�9Jf	����l@î�� '5�&d��]�Q�.Y
pjwVQII'L�x]�6�9��A騁��`��"�2Lb�s���n1��Ժ��hZ����a�����IHŵ��6ɨJ��H�|�{`@�L�b)��Wj�IO~�~��[��dne��MyJF�Yz�\7�v l�%+'A7n���)��:�z~������J�;|H	\��"ρ��ڳ���FP ����̂�7�&�R����qw�*
��QC��43�U=[ֶY�h��aB���}�F�� % %.�?�������^Y[�['MK���\
	�Hʩo�pST5��Ќ!H�B�S�j�J�����^�W�z]���� �{P��$��=f��\���9�y��M0��7��mA������^�d쥛E���U&�F�\ؑM�>4�AΡ�#��F%�u�"ZG���u������^vO��~<��	B���b���bV6'�3�����M���7�ߥk��w/ϒ>��B���0�e�\vW���ػ�%�	�.F�V�Y㪁z�V��ə$TI�K ��QL��r���f�2��~ѿ�{  �҂ǒ����*�;�1,�,`�,�b<T-�ow���vr�o�����[3��ǳ�_��{k��L�?���U]�y���%�Z�?�s��8���"gLi��(0��о�l�����lK�B
�R�P��q�R4rb��}q�&.ox����%"�2�v+˵�O����Y%)��)\>)�2��RI����y��ҁ�>*n�"����O@�G;wm�OD����W�Oߕ� ��&f�N�pK�<?=��~�I��}���f��QZlC��<�:�Րiz�V�
(��ޅW��d�^����G�,i|fS�X ��)�_e��2��0�z��9��V�́�1t�L��ɟ�����!#���>�'9+~�^a�Z�c��3.Om�I!B��\T:���ٚ����Nk#ː�/�R�]�����S��������7�ٮ,ȝ+K�2Ⱥ��t����5,���Š�'���,��D�r��3�@Y�p��|x�NY�>�^\��WV�XV�����J_�F�r����	�K]�$\j�8fA��d���%A���tR+ �~`b�Ϭ�e�d6��\�O���ݡs�Jl�1X�}D4�B��i�w�2���������5������.��(R��L��7vK�3v���}��^pk7�N�Lhwq�P�d#H?zT��٭$O�s�JGw�s'�Hyn D��XP���OOǝ����:�R	EＺ+]y^q�Py�����GRr+e�nhl���� $I6��p�����KܻL'^�]��pQ��?z�?��s���:���Wui ��.��$��Xd 7����p츳>$�r��S�A=�(U�g�d��[��'�U��n�Ȯ^��Ԅ2��3'�l��Z���C	���� j6���+��+\�U	�#,PJ��d	�ᔞ���s�
�!}T�����u{YW�(����.{��{��[o^�<��P�_�A���њ�ؒ�OSe��p��^V�4ۼI��.қ�����%�1��lh>u�2���4�*d��|�}��e�:����С 3���wmZ\X�j ��m��TZ%��������6!`�ǋIzo��?�����U$��sZ_^��gX�1Y,�a������>*A��?2Z�c� ����0/ҷoo���WK
��M�˂5>-b������aׇ����]{|jw�3����y�hrl�l}t�2:�7�b� ��P�����yR~)��9t����q:G��RfI�@M'��8;Ț������6�P؜@��n")'������}ɷ�����mh'1������dA���6T�1�㴴sy}ez��v���˟e����D� 7s�Lf?�J�ESR�e��
G�3���I�gq��짘L/��##��g��Eߏ����jI���Wy���V挊�R.sphuWMw2��"�$�T�a(��
<��~3dG93�qyq=pM]�n��|���e�����Q^���b���0\,�Gb�՜�d� W;ç䞙e��iЃ�}T9�5��-�[\+2^�ͧ���� x��V������.�lwO۴�%0;lţ�ܿ�uyP�F#^�t����X�cuV.-8�pl�
Ң��b��	Ӗ����������v�jm��b*�R ���\k&ˢC�ͻZZ� �h�Ii}ܹP%�$�NsA|FQ:7R�A��+M����L�������&A�L�d�C���s��v�����"�k�:��j����%��p��*gD��ӴG�6e���vN���2������=�Y.:�'GT�k �{z|��
p���F�qiY��]����܊���h�PDvo򍻴�t}y�Ϳ}y��.#d�X�	��(Mil�0���ςI�E���:�O��y�O㶓�Li���L%�����.���GsR��f�V�
���ġ|��b�M-W-���T�>�EY��I��}I��GPxU22�\��م|�Fv� ��B����s����F2�A���~���p�z{���U���u5c���M���H���k�{l���3ȸ� �ϰQoo���d{�>��:�-��y3�5k�	�;���J�)>c6��B�@sPV0�}�K��k��r��������{I_[
��Mske���B������xP �A蓸�-��げ�����R�s���/�(g�'R�U���V���2*h�޽MvS���-��~)� �#u��1^�Ā-q��͇���ٳ��n˅��
!��K��#�?���݉�?b�S+Y��YB��a��ϓ!��Uw%fya���^V�����-_�/��Bo.*��P�]�w��U~��:C�3�h ����;�<w���|�0)ި�>����$��	��WǪ�>-�̭,kVG���=��"I�u���[+	��V�O�����/O�0�(��շn6@(Jw�i�=�E~�gBˋ	Sod�]�l��d��+SJϼ�IF���J8��*Nn�L�Hi������!Y��3�/56+ЏC蚱�x�c�7`s&2`�β7�犻}d<y��1f93�P�s���\��L��L��m�W�O̐�����à�N]Ri��d�N�lAR��,��I�T���&�^V�wח��Oݹ$S��d��>`/.jp���{�f�>h[}TtMA�Ogi�ڲ�[��"L��l�ҋ��[+wn�{].�e1kb�l��K�����>�	�ni�T�B;t7�/is�(E�_���E�����:�����Rk?�Z�G���2eA#I�2�S}�����@�Ͱ^tPr`�./�"��T2�]��ut��M��Jj4ܮ�.�Ȅ�s�T�����% ��/��a~PaG���X@!�y�����fgAm���YL��P��CR"�d�~�=-�@8i���̙���3�Ãk��C��Ju gb
�s��[5�/�M��2���q��Ke���<>Hl^�| y��5���'�����q>�$�,��d�i�+i<�iJ���Nb��t���]���|�|��S�A:]��	���p\��2��0kQ�$w)�&�p��_Ʀfa����g����W &�]����8�i�Ut��Z� T$��\W.6�Q��(r�)�4ٹ	sT1�Y��-W�I=X��޳�����7�a����)g��O9u��VkϨ�"y3��ʿ{�>U�H��!�e���|9(����U���P���N�b��I ���b�m��V^�i2N�0*$��k/��i1N/�v_>��l���*ɖ�;���O~��S�:�k� B��]�����˜ϖi7�u�vAR����C�qp.m��Y\��Y��0�/8��\��jUa��0��^��*�\�rXg]�C
��P2p�,�M+| ,���G�v�G�$ie�7eZ*|�o��~7P�T�zkS�n��9v~5a���\/�	��S�DTA���3�f��[+�/��mv�./��>&�Y`��6��k@?C` �`�Tr@�i�������ʣLp}�r0#���5�8e�ѷ�鐾֥xj���ɠ8�A	����^٢��0��{�yZj��Q̭�<�E٩���F'9���Ƃ�U)O첏湴�8�h��0����/ه�p������"c�	�I���� ��+۽Q5���S�������|�y�Ƒ����M'@&��2� 7X�@�:���{<�Yf������zdbdB<..��Xdݶzb2e��e0��|ڛ��~����}�����<?}�sm{<Y�IW��t�����:��<�ɏ�>[ ZK��|i�u-<Ze����Y
�
`Clf�#ê�n�uSI�K���p(˰����2j
��3�c�y�>�ւ|�S9�2���%W[I$�P�v��[��<�N���٭+��\8�X�R��N $���A)e\�{��ZKUy�
p��麆�j�}���>�J�=t!��}�I��m�|��������A��E	�k��|����c)12�oV�6d���;�ٕ͟��?mӯ|��̭�Z�Ȍ=�/;Ep�#�v�;��V��=byr�ƞ�l����S��G{��ЏSY
����lT*�=����b;{�	���2KG�K�h�UOp4>hQo�<�¢���f�H�.J�w�v�3�������-��/^ɡ�=��?@����r�SO���O)4#��P�������D46<�� A���߳2,?��:r�v^V�@<+*�,� ��We�̒k�4kw�Q��>�93�ku.x����E�t�-�.�������Bb��Go�dN�t�����\ۼ^�����6w*�����8]�ޤw��=�>�d�O/�e�����K���Щ�^��j���w�> K��g��j�~_��U0�wi{���l�ʂ`����û�ʬã�����zC=��e`dNR2�z$(H��F?�d�.T�g���w�T+�q��;)�tM����E,]�<d̳@��Z��EE�g�P��lX):�cY�ŝ{�R���f�9����SR&՗K���}(HJ/e�c�>N�@������3~������'����������2V���V�#�"�-B�K^#ƺ��8��*�q0\;�d�^H��"M^]^{�8 �.�5�\'0��v�.X�t5�--N�E	C�~W�S'onWڤ>�:�d��gJ���bcCP�[���l��!XfZIބ�QT��_yZX�L,�2F����ܗ��u���E��(�٫��E/����}��rN���:p'Y$�^��C���Y�){����9��������KH�9DP����SS�!�qv#�vS�9��I�)Lf��M�@�DnWV�q��p?!�_��N����ߨ�����=�Dմ  ��IDAT����V
!e��sK�c\��Zzr`6k+E�[��|4���7�
Ȼ;�D6�Ւ�A��R�!�]���X��a�0�����HT��llh_ @�GUNi}(�� S�{r�]�Ve�up�{2�^��֤ۮ�x���7a��%�\�?}��?��P���>������H�j%�D/���M$�ϫ����c�8f
�E,
���5�W$��;���Z�pA�0�'��U���m���r�m��$Ⱦ�(7��+��"y'�8�T��gy3K����\1�.̎`�M_紖�;EY8�{�-2���+ 1N��%��!Ӏ�޸����{'cS��-���&�H�<�tŏ?��'�1�*N\�S	���w��9�)0\M��뭞_����@}g��u��� c��¥б����(�(�L��3�̓L�,7��% �"�I��@���T+@�`�����$}1��u}*b|R]FpMC����\��du�8�k��x~Ѱ���8jޕ�k�<��`a�B��B���5�c��v��'��o�'�����xg�(H��J��^sz~1v`z�Z����+m�>���R=I��C�ru}�൵�0�ѩs�\&(���jJ�d��j���䛰Ɗ�ь�rV�?	��=5thQR��N�Af�F7rҺb�������)��l�~S�wI��¶/���%׼��,;�iS*����nh��&l��Z�
����9/l�ҳ�8�*'"�!	n���r�P�����(�~�ߥ��L��1��*H/E�x{M��>��έ�Dx�g"5RW�~�EӔ�m�z�1	}�K�M�_��4=�S����-`S,��r�B.��S��}��L�둸��/
$®Un�A����.t�#�i��zG��ɟ~��M_>�,$zO�*._^hڔ�`)�����{@�l�Qߜ�.�/����2;�<��~9��u3f��:G���`R����/7����=����!1�d \�yh�C��� pb���B���x��l�=��Ͻ�|m~�X;K;ܖ��6�9�	�j����ݠkН��y�f�=��
�J����R�C������H�,�[N�8/S�{�y��cz��`���;e}b�*eF�Ui��� �_�~- �����OS�A�*D�S_6<I�=dx978@i8�T���상ѵ�<)]�&�(],C�v�Q����S�K�H��)�BA�"�zfB��+�:I�ڹBuU���g�ItF��TV�QQ���G�� 	������s4.��F��1��ށ����[0�N{
�ĩ������ wί�:��)RC/5Z7�/�
'�^�U~�#�1j���f���F���C���LB����T8e %��ΐO����E�wrk�r<��ce��6\#��L8��}T9�A���.\�M��sa?�}����m�G,�����m4_=�sG"�A�zV���v�s�fCZ��8�����O9LjVP�����RD�p e6��i�C�z!! z	�A�@��P>sΆ2ؘ����{I���JϷz�P�:7�FJ�(����gPjxE� eTD^V;R>��!)����U"��Tw��d-��[73q��.˥K�H�iK{��Yښ򰚏��[��ӯw�U�>[ư�H���޼fܦ����أ�\9g�2�Z�GD���M���$���JO`"��i��f���	��c�{
.m�y�JPi/�F$Ƣ����R�Po�hv��Ҟ�N:��h�t�{�G*2��%���sG��!!KEw�d��� y�5ѯ| ����:�¨�d�n{�X����X���AG�p��+Q_A;q2�� �,���1���z��]Y��mQG0z8�,����`$iw�Bkaa����}fW��y{�;��Z�Y	Z�.wbA���2�l��,�ny��B��S3|����+��2'�1<3����;W�̆�=�IQ��P�xfdD��&�}�]�������Ч:W�8F/���id,DJM~/{�ff�����`b��2�V�<���OI����JA���ݦx�u��nvqJ�_z)d�q�����x>���g�6ׯ8)�d��4�������1iG�����/���)]]�{��uA ��#+��U��$�ͭ��|ӡ���K0*�y<��6\�*�Q���F�4�lD�ڂ��6�̟����鰲�a1IWdy�3#�b�Դ����jy�,�����.�l��Y�Cu�̔���#�Ry��#�pvm��0 a�W�Ր�l<���&�[��R�vV����� G%�l�=1OJw��Δ^�5�HS:l.�Є脘'��eLl���Č�D#Y![-��\,����r�ꂛ�=�W��2��:{p�׌�6���{.r@�^U$�P:6����W�����ƣ�]@���u���\)6xN�<ꝡ�M�7z]�f-)�7�l�j�s�-��4ѿ���h���|,\uޏˊ茉^����G��U���߹ЀUi�6�B}����D��\�L�d|��;I`����h:dA��L\S��+7��9v�b���+��
�l�㤆1��-G�/T*��4H�0j�1ܺ������+#�	��"�����i���3���[rI���<�)B������ ��=���Qӧ����I=��y���6(��e�vbH�)��[
 �<^Ǵ]��7��DV9�/�dd���m?��, �3ʗ�2���ez�@�~���2]֓����Z���tc��ś�����RL�̏�����{X!kE�< ɮSk�j}p+[���n)X�s�#�����S�?���8���������G�Ŵ;�N��l㚉9@�� �x��ߝ&�!k�D��V9�A�ރ����+r�d�͈v�T�x2Ӏpj���������)�|��t<VЇ®�]�M��hJW�C���X֎`
�n2{/�Au�>{��J��� %�N.�r�;oXk�!
��[lݶu:�#�E�v�L3�v������\�o�n&���9��`i������.����m��C/lKW��B��l=>�ۃ��u�e�V��,�M�6x��ѽ��G�-c�������(_{�����������s9���0W�i�n�,�j�Kmf����9ϱx�=�o��##̘3����NeiƤ��ʺo!d�N�&cs�։Y#��:W/�b:|>1��W>�eP�������uUk�W�D��1qS��t�שt/��-wz�֒2/��4m�/�i�|A#0��R)׻b�
�KJ���n�s�<�);��4�����=�ϖB�C��6��ڮ��&uv(τķ`3�:eǍ �U�!�x�{4�'T�ۃW;ɝ��v:�
�5�:'�I��T�4p�Qx��P��Npܤv�)��Ҵu��"�����&�D1B|5y�IS�ҡ+������d�L��H�پ�-ӷ�_+ʠ���%|2j;�n�\�w�v�!Ǵ�ؾ�Z�����٫�?��p}Ⱦ`|��[�¾ȃPo��&�DقE�'K���n,�q��d�*o�iR�����[���R�SkFdG�.��!N��Ӆ}R<Ke��s�>�X9+�k�#0f�RT���j�'D�v��)�V&��AQ�=2��\�	Xػ��γ�}�vYH�3�J���D�`�<U���v��^�qI�D�-7��#�^^�
:��~wԬ�Ѓˁ(����|o���E��:��� 0���~�!��୚�dp�f��\Y�w}kϽ�;�el6kW@ə�h:h��\i��~�yY�ۮH��4�|
���ʝj$(�K��['�saPB����(�ki����Ȣӛ�\�S������w��<Pg�s�=�GM9�R/zj�gzL/G�@�0�$�W���ޱtOR?��ʱx�J*��)���Vb6���mI3��Zr*�"#�̖�^:&��\���gyH?�1��W���Q�Z�!���Z��ԓso]I���r����]�pg��v��h[i�����>���&]��~��V�o	0�Eid#�H���y���_��J���8iW����'nQ�@�#g���L-;s�x6�{X����S:�uH�����,�FJ�v*ӣx|N��wi�?�+[D㢎f|�Sp,?��2��nn��x�V�&n�FD6�Mח.��ޮ>2����MB��s�k������O͌�:)�z?o�o`�r���<]��q����$��9Ȁ�"�䩤~7�O�Du~'CpCL ��O��+-|zZ�̨,��:��hW��>4���Nߛ�b���=V�5��d<��p&��%�n%˓�+I�c�'��� ɥ����!s�OP�?��z�� ���a7R�[=����w���>O�XV�N�?���S{�+�,����u���
Hw��>m>������lm�uY�r]�Rm̄,�]�z����Ծ���⺞I�g_�CO���g
��:q�\h��)dr�v%%Yߥ�&<Z�#�!Q�xj��(`U���&������u�8'�@!�~O�ʅ�ݪ�V�:��[1�1P�J5d��,��PT!��y��W�}E��5z�닐��]�-,��'n3��}���|����2�Cs��_p�Z7��--��Rc�sU�D<u-�J�r�H'i�<�9<H���&��SL��c�����kMGi�S��8#���	`lz ��N]�J�/�;�%����AS�4�
,���y�&��[���J��/>2�y0�B��3��=�����y]
���P�-}*�l�Ϥpl��"4k��ɲ��V��ߥ�\^.$��ͻ��ρêPA��f���n/��:K�7l���&��G�,� ����f<}��=^��}uc���r�
u��I�A�凲H2w.�������O �Bq�}��j��>%�޼7�gU,������Kr2{�Yji��|�V��,qt��S5�<KA���k�dz���c�&zo����������Ó������>�tU�ڳ�����`J�}��E����By�Oo~�!���R��?TP�saJ��aIDW)�����ߡۧ쉪âO���ó��ݫ:)T��SL<���&$T��%%���E&@7짪p�tl���/W΍`���,i�o��QwV���1㹆���i�ؿ=���3�*�zv��VE+<��J��؛�'���>��
n�ΒpK��k�i#�jK]�ߤO�'	��B�6�)�%}
�a�;�%Oq��V�Ӈ|6��&�q���F��b���|/��2��O~��H��۟����@#F�S��Mg�Te9x/Ҝ��@�E�&u��V�
[�W����z�%��s%��!@���"�\ʊ�e�6pM�s���Qf+��!o���$p�l����M2���� ��`�c7�����
FC�>��x t�{���֚�z��\B�¼yg奦�![Ł7�Ϯ�Bteb�%���_�28��T��z��-B�qR�4{�]ZНK;���.g�ց���^;���C�%��9ey�K-�z��ve�Ƈ�2��|��Y^�s�}�F@�߼��ǟ-�AtG�`��=>�d���,Ó8�ŉ���>�+�/��ot�0Y n�Q4Dn}`���`%+�vE��.��g�,��7�M�^e�	h�C�}�,�^d��3���2`^�'t���p��Ku>�uK�� ��LECn=���YT��t�b���ge�����nRFpw-U�J���~;��:�ѹ{�itͩHLo�n������f��(���<��BË�|�{i�1u�w��'�'��Fo���N9�!y#�r�)�sY�Q�9��%c�+�G�Y�k<�Ԭ�ք
Hw�y�YX&�g����`��-c�����@.�8�y���;�y��p)_^)��Kx�f��lڥ��,��E���Btdr}�x�ȸ�>@�y �� �ȡ�p�b�YFQfg�G�x�B��͟?� ���ˠ���t��ǗiV��A��wi|���yc��բ��m�L��!�� �������$K߯�o�����_���̷����}�M��ǔ��ͭ&�?|�>�łڿ���:��?���כo��7�l��{����m��5��괾	�oy���vR}�V����I���Ł�(#q�QIA-�y�8��\T8�#�k@�_�C��eq�3s]��R�Lz6�qfH1`"3���X�沸�L��y��͕����V�-,9XX%��C��N���j�'���﷝_݉��+/(H~tQ�k����"z�YJ�x'G+dW�����O�[�4!(��@Jg�5�2�{V^�ϛ�a�H���A�����}U��̿�"I�{TI��w�۠;L_?�-]S���2DKv�4�_?/���ya�k������}2�W�*�g���E��Me���t���}�����A6����̸<-ʶ{���`�E��RH�X�ʍ}�KO��D����Y����w���cy�z�'N�tⲎ���R4Ι����=G[C�& �H�(x����-X�p�M㗭�۷�;�X��0������*}��[������J�o���%���$���M�|{�^VOiG���`�}�/?�����af�=�9�ʽ��Њ�<� )���ý���i���=߿���2��[B����4=��{���0=������.N�x��Q�9c��[�I:��@�D
* ��~8߿�n���v=��*=����5����<�z��C������Ĺ�G��m����~����ZM:'\αX�q����鉜��GG�����E�BR}Nk�h�T��$��0��E�%���9Ť�+V6��([�㰙��y��9� ��c�p`��D�ss_�Q���a���� g��\z�LrF���'k"��'?���/��ֻw�`���U����y��Yj����� �����grӐJ��Tus���-��!�8��ӳ�d����rj�s�7Z��P��lO�(��@7�Z)>�C�^s��>Gm����?�Ò�eAeoץ_�sUv���F&��l�u`����ҿ���g�<���3onoӷ���.��: �`�a=p(Q�M�|��6�]�}�F�xD>���3L1�� �!��@��`'z��}��÷��ͻQ�'�bѾ��"\.EOY�~l{� ����-R�W/;�֡)�k�'����mg��O���6u���e���$�̅o޽OWon-�&-�ޤڮ�
�ƞ�uq
2oJ>0�žm~i^�#��G�6��ߪCitu�lErMuɆ���S�p�ڕ��I׏�^u==�iii���Q�`�2 �m�1m��b*���gQl A3����@��b��m�Ep;F��G랁�bE΢�Q�b�(���T4����2����!j3U� r��e9��s�Ld���mϰd����$�	7�=�ɼX��8sh�K=�����4��D2�U6�	�A�����T��L]�l�Y��N.[^>�5>응�e�/	~��N6��\�읚_��v�g.]��v��׵��a�]8��h[�u_]�P*�@p��/��FF���^��ÿ�W�:�����H?Z)�����M�����(�d����4������i� ��ڴ��Y`�?<��2֏]��C�i�t01�`�ﯡYHZB)��<�ɓ��v��<�sn��8�kD����b��59#�)?���sc���L.n��g�c06��A��e�ǡ���u�H�����9t?|�]�}�6��C��JX
h����ҨKY�w�Ԥ*�-X��W4e.��8l�"Y��P}T-�*�v��1���7~�]`C����
�i[�K8��Y���p���讗���_>i�;7���oE�B9k�ehĠ��"��k���//k��t��'��<e�A ��ڜ�S>o�
q��m.{3u+o��G�t
K�ܟ�٬JT��Ǝ�r���� ����9�<���s��uz�N4d'b89������d��=g��2�y����~��=� ���'ף��+�����r��������+^]�|Hd|`��br�#��{8� M�Nl1D�ޘ�wdQzA�6&�PWV:��β�"]�!B����?h�:��}������������SK>s�NTo"U~m�5Ss��0��Ʊ��*?U?���*ع��
��^��;�}�z�YS�FG,@{?` �-��N��o�5~�$ãZ�:Y){�,>(;�R��g_���!�F=�\�OC8��cO./��w����������	R��ԋ���hI	U1!z��G���Y�v�����kfn��*��}xIi��Φm��� 3�	�i��J$��Н$�I����Y�޼Q�\%������������m<���;+5�@{�]I��z�|�4.JIm�t*�^I�ŀ��F#|�UeU�O�";H	���ƕ4F��Й�X��}��4��?�⹴�c|F�S~�ſ�;��t�f ĝLX���9�g����Z��x�MЦ����>y�%0��\:+���p#2g=_���M�L�<���ʌ��a�r���}�s�Ã��O�&�3����n��`�3���l=�\J�����Z?��w��O�mzy~I����/u��^��U���"�'��)4���t=�I������Yغ�B�ٲ�FRݍ�����[0e8��1��Z� ���ϫgeoE� n�EТ@��mde~���0p|�]�뗂4�\��<����2L�a!'�h�ں�JW�}��Dd��B�>�lJ�T.�EX�Kd*�$��A2�\�
{�o\��\Y����.�L����qQ5>��X�����x�c۴V�*��JO2���d0 ��߻v��(����T9i�Ҿ.&����ϣ?�/S���n����X�W��t��o(Ղ���������]�OJ�!���$4��dQ��KÉ���O>������VϮ-��z��2F��Ep���M|>L��`�s<-�У�]eQH~^V��?��g�8�~���L��$��̌`�z (���7��g���A6�����b1{�� ��� u�x����R�oS��f�G��f��LCa$k��2����M���u��Vpñ�6:��f��v�N��"�y��h��<�0�&kl�1p"H�����O�������l|0�?���gA7���~0u����s 2�qn��I���HY �5�"sc�A0�y�V/��������!RNm�q��M�T���/�{m
h���ץ'�+W�
h�uڳ��K/�B�>g�j�F3\?X���@���!�%�F�71J����̋�����C�е�ߵ�H��㜑S�۳3I~���8���}�P�e���9O]ʨT^pab����A��9f�^F]r3\N5��(6 l6b�"r�c�,�sqЮ*\OJR�evti!�\�ϡӫw�U�ؚ��~�ͪMs��E�6��N����1cꆅB:eS^�ƍl`�aŹ��95����!��{ή>�{�}��{����`���)����a�ܝ5��!�����}���2=�������3M�G΢�1ȟ㗰�,F�?k.����^�������X�α�\4t�' ���Rw��m����1��?�>����a=	?t�Ni�ݯ�2P2��j��4�C�f�~	\�f�1ד:=�a`F���v�u'����jYT2`��Mҭ]��ȧ�H�H��x%}J/	�Z@���+�l�"�h?�U$�s'��fw��9��zw>�rKI	$TαF1���ڭ;��?4�z�a��P:�C��?�A�gvq)OY�F%Z��Ӈ����t��v��R�R]��I����v#�z����(��x��=�N����t��� _�S�Dzg�0�E�D�9a��)hvƂ�� 7{ܫ9���L
��m����B�7m�0}����'��
N=ɽ0ό�r/�Ap^�����נc߼�)5݉������EFf���͞-�r�JfA� ��r��Ƃ%����X�j�����!��DÒޯO���A;���y�p � _^V��t�H�]A�:wi`q��8��(��4�_^��U1[�M*�Ԑ��x�Q���tT�~X�'���d˼?��9M�/wV�>�z��i��;o4���W#�Y+l�3����f�L/�Ijոa8ЕqN_�������\[��9TY����q�n�����.�o��5i�W����Qv7���� �$@����dù��V�۝L}�i������&�<�R���d�}`�N@�s����Jnr�\�=�-/��w�����?Π/<ڮ���}�奪b(�P�uz? �3�!�������n��Q��6�|⅒C�;:j�*o�B�%3���đ��`YD1�� ��-�� ��տƞy	뙁��!����i]�A�����04���&�T����WO?�`R(SiNnV�����Ϟ�;
��C&Gvu�V�
���)/g��<ਪSV��$iH�@P)
���"�rz���\��QR��������?c�>�r����B �D��C�se���~nk�2����{t]h��|��ޣJ�f�jf����G��*���Y)����Et�欜c3m-4�$-�*�MP��G^�=��̚V�#�(im�^_,u�Q�������:���}���kJ[�dw�7�����ORߠ�Ep����Y�{��.r�aLֶ����%��p�5�8U��zy��L��]|�غ�T�����(�_�~7�8x�V]��d^�]��0��J���h ���3d��Y�ӮV��eh[�H�G����qK-E�֊~�B� K��3�e^b�GbW��.`m?3a!N���_�7:�HBh�c}����縗>���B�9N��/�拃6 c����u~��YO������v�%ET������ǖN�J�q54�	�R��NVz�P���P_X��˔,���&~H����R{_U�R���#AU��R���qVn��D)�N���/I�s�-6L���F6�s>����š��2�-��d�ݓ�C���N��\��,���g� sP�V4�ޞ�~R�
��cQ�z�ǖ�YǬ�	 #^~>@��?��[/qe��ej�[t�{'�
�UiU�*,�5��c��B����$��Ҳ��8|0�������>=�׳�zgV�.�Wj=ЄFwzdk����p&	yW�����M��m�y���&�l�����\d�����e�M�L�j�]��6DH�� �c�٪������0qe �kLgS�� �����az��72r����9�&��G�W!�G��^=Ma^��Fc>�xS��n�-�]\0��u�"��߻S�냰�3?"h"��(a�^��z���,�f����c��Jt�3^���1�,<%?�W$�6RR��TU�F}��<R���ofӶCz}�-���sy����cX;~O�ȡ��5[.;��w��`�L'�X�K�\^<��r��&ͯ�w��M%��``��5�)e�\
SBe��kf� k��� ��_��N�9��5�p���O��!5��d��L�������{�ꮣ�"�RYP*�)�t��!xqM	B≾,�C�{K�c���rk-9�-(��p��P5;���j��C��e�pv�t�µ}^��$3c��ĞI8<�[��(
�E���2 �b�#b��4���Y\_j���޸�>�o���8�@\>'���v��r�]!��hh���Z��%9	ZJ<�qni�^%"��rW7���w�*�y\�����E5�V�m�w�)�\Գ,܏#`���]����!y4���xo��;d��j)Pʩ(�N�W0��@�!��y`�X8�
�UvG�&&/;�pZ���LYB���/7�ʝ���r�!�G3[�QR8��N?��a�h�pUo��c�|0��l~?��Z�������T�S�y�0o`NnM����;?�|��r�VԖ�x�R3{s#��<���&|ؙ6�2��4Q��:ASa��r��$�j_�dD�iI8e�I�/�W�0�1�sI���r��K���ڏ��@ہR4�3�" ��K��)����{��pG��1����X�i�+!@֤�ת�z�g���G����J�>~�ݠ&��A�3q_HIfl3t�N��]����z�/fi��HW�E����s�^�U��);P"c��7�*U?a��+=�ևjEd�#Ih]+�GM��Q;��q��9�I��ڃ'(�XL^�!���{BF~
d��֮�\�o���>|󍾏�*�
��ɪ�:��>��}�<��{���w�;ږ_1�M,E�hj�H!?7� .�����*M
���p)�l|Xw�� �2&bdn���C���0���)�޻���IWKm��NNF�0S��x�%b�6Qu*Ks�4:n�E�'݅V���<r�t����,�2����4�:��>��ՃRI3l��q}��(pF����\�� ��>Qݜm1� �y����+�/�d:�h��z����^/hN�E�����5s�+U��*���/iN.�SC��f��9��G��!.�F�C�H���E[�C���XƁ����\���ļen��6tA�J��3�+e:��V�����@�Re�=���BK�+$կ WO�Q�3<��P����	���t��u�M;�E��8`	����M�T@/�3���ނr�p��+�WXGڡ�����
Ҫ�+�8�"�^,ԣ���]۽����^%��׶�T�����2.Z������0vF� ��l��I�f�>hr���SZ�!��N �B� �����f�%>���v��ґ���|��V͎@u�"Ø,���']�
C'CV�� XW��~h݃`���9�=j�A'�(���pB�:���$РUy�<��P��C���̓Y/�^&�;g���Do_%@�����ǁ�7T���j�P�t1w	8 �q����_�E1�E��K����b^0�F���l�m�4�gZ
�\rŗ+�T
��Ǧۉ��Je���v۽�ʳ@�8ZMe���r5����n�ݗWɵ�^k�ʔ�-qV�'��v�q"��y�(�"D�tp��B�[�q�F����g��>U_�&�12�l�d'���J�ɴ��JW~�P�r����Nr�XvQ��=�����F���q�:�c�g,x��zm[(H�.�^,��h�-S��C��U��l���>޾�6͖3��ia�b4����R*��ܼG�[��i�%v��ϳ�u/�.T6e�e0&�0jP<&	����Ź��Z��^@OcbkjAp����x�dl�_J��(�Wr����{[��V*
����攓(� ��W�����@�=_ٺ�3������WT�SÊ�4�l��F���J>��>=�ߥ�>'"�`�X\]㡓c�v�v�ۣJ[x�����9k�2�ɨ���W��l��~�w6�D
�þ�L+�̩��E��z0t���E�l5�h]ŕ��S����R�5r�+n.�(��bS2!̈yS����l�];^^��(3��:���׸$_�2�Nђi0��ǖaè:���y�	`H���{9@d3f�G�F}yRiȽ�\�e7)��G��,R5�d���2lf�2&�L���7/*���e�s�,���ZI�d̼��(&�F�����sw�;+k��k�jǤ�r�}Ջ́=��#�����3�Gˢ���$�۩�����a+�{!�����
����x�˰��1��a����j��֮=$VK̤Ǭ�N��²���\L|=F/�q/f��f���!m��$1����:� Tʄx_콍c����, ��7x�SX��eR�J��cZi��Bm;s:.D%C{�!	��c(��,Czg���+�v/ie�cMVb�|�n��E���×����w��J
:���7�e�K_>~J�_�|]ۺ�Y�����+�5���(��n-�R6�>����G_\;����Z���
7lYx6�nZN`O^��X�ەx�,�L���
C���nU���q[rl�A�	�{>���_h�X)������F#�V*�J"ج�v�4�s�5&G�h����~x��}�r�"�2���T �B����0kY����!#�0�� L��48 J��F�lG��)�i��g�	��@c��l7�*��� c�td%8s�!h[Y/OH������p���VJ S�_8�yz�Keqh;��Eu6��|Q'o��e�t�\|�Q����<���=qZCхaҽp.AoC��>�l\.Ǯ�q �w�.t�7�K�jn[�>+/1'X��-�6�1DW�����eS�d�H>|�b�:�|����eV��hm��#|�r>�S��-����T%dpvOX�{.(]W��:�>I}y�OO��hAy#5����C�VNC��e%�^�Rb��\�}���<][���Pݻ�8�����Ez���e��7[��a��*�e������BU��ͻ��?�'�8�Xn����C��ǟӝݧ�w_4��=�l��/��~����!��؇2�ܡ2�|]���n������qK����u����QLG�`(h�����O*�E'g @1���P��\܉�������w\} _��0J|e���ǧ����j�#I�5�Y�H EzzfeE�qE���!��d���p��5��~�nY�9�2#<��Ԕn�����i�%&t���<�T�r�6���&����?N��&��J��>�ӆ����"5���P��\0FiӦ�?�Q�R����gt�T�
qN��x9D%�M`?<x��q��L¦�ߨ��|5f������L��9Mc���G���?H��3RG��A=JY�K�2�O*O��1"Z�{�v!��B�y����s�e%�i(:vS�XgwגW�-�cJd������+7F�<hGj�d���L�_<QWse6 ��TS��f��'�˹��"�lMQIl�0L��݂ȵӫ�e�Ȣx�5�?�-�(Iw*A�&�����qj߻��Ke}hXゟ��~њ����{�LP{!3�|}���*p��ệ�\8E���>Soo���Y�4�2����w���Q���f�+C��V�%"@�~�;�<XYS�Z�p`90k�Ѫ�h��z�El�ap;5��7�Ӭ��}p H�E��=)������� �-|t, ��>�؛­�"6��B�a���Y������Α�Q)e%���m�>l�/7��I�Z�����c,�)#t'z�ޏ��X�Q{L��m���G2��@(&��`�J������iX��(ި�X���b���`�Ա�vu�$ݞ����$M��\�R��{� ��S�N��K��r6�9ȃ)��ij�������>|�둹�$&Z��;�k�D4cp��v0{A[b�<���w��a�b�?U��{��K|j���"d�<;��G��Tu.w&~�)�&��dU+ی�cٳ�#��yR
�Z#S�}���Jӳ~6��2��kˀ�oT�e�{a�hݲ���e�8��,��P�����T��ޝ�8��0-��_�����k��=�?��?�\�f� �u��Ђ����A��k%p���d�>Ђ ��`����va�}?��5�g�_������
M��n}���-�9[`�>��><�3�-c;j���ɂ��(l���S}	|�Y�QL�=�Dc�3��Я��/�����_��|��v�����H@�r�8�` ��M�X�~� �����N�~P�,Fu]u�Y}��CP��2��;`��jt��$Z��}��n�ևP��)D��[�v���8@��;N�xc����n��#1Rƕ&��k\�*k+�*��?�1!�/�~lz��n͈����{�}���A��;J��?#�I�_!�������|I2�sa�&e	l���B�z��W��G�4��d�ҽI������,3�Ч>�ϛv*u9$4���}f����}��:(3�0�4�3�Edp�0�8QN�C.���f�bmY���mZ�6��t��+FG�;8D��e�XY��ϧ�*zf��(g�FX5$��;LL%��=�^� X��O8�X ;�Tۂ ��*t;�:���Y�l��������ZmRkA9S��~~u%x	,�|�.ˎ��� i�<-,��J������͵�I���F���l�(-�T���F^�TU�I&6̫��ìP6���r�� ��z��%	�a!�uoe�*�,W���C^�~��u��+_�rp��L�/�㬇_*|Z!7�VÅp�T���;&B�D,��?m?�=L?:Q�?�Pj���JYʃ�W��)��B�r��`��zQ���f݅����l�u�� ��+�v*|rX�P%_yԲ?�ͤlc�df����=Sy��+|9k1��)IA�x<�6{W��K���_$����d}�Lmx���<T������ @�SM�4��V�T�I-�}��){���N!)}4�P�*@��A�`��"�Ɣ(p����lxv)�$���8}�Ё4���P%2�,p�m�0c�ԟ�Ϛ��ԁ+��E{'ї�w��K��v�){�������^� �$d�	,���9}�d�Ű� V��$����dzLU'�$Y�W凫��e��-���0y��a��B"0��^݄+�}�Z
��WS�ثO�^��=�ϟ­e����<����,�� ��iRd(��r�����Y����0�q�.�z'
;xv���,��^�_W�i<������5,��ۅ�+���}���vhN���__,�ެ����6���[����\��ެЦ+=@��{�Rb!H*�n��N�<@���R�G�r�',�8}��a�Q���!nzA<"�4$�ge��=g������2��n�
�����	�_SAd���������6e�˥����krRM��"���4�����!�N*��cF"L$��W���T����e �l8��̍㵤�Z�Ƣ����� (Nٛ4��� �t��U1�r����\ק��ņn�SݶI�[��Hh�Ah׾��j^���9D��|h凃�/��dl��ښ�Xִ�u8���Զ ���p����d�3%ך��W�T��<����5�R�\m'E	@>}z����ު	��שs�)�V�M�@�U!���>���,p�({��7��ւςv��I��{�
P�)NV���ꇁ��=�X:�YT�����^k�ծ}7����ýl9���0��J���xN�a�vY!��J {��J�(��(c���p��h{��~���b���1��˖��UN&���-e��;]���rM�D�m�d�jS���F%6lCx;dۦ!���K�{U��/� '�8�z��)$�'�)&*�F!�>�����N��	�N�v���	�tM �A*mA�i��?+cF�Wɒ��l�'��&�O�XB�bতSi:����r����EH���;�4|i�'�d�x� ��xj�����9��P�'�����f=�I�Sf�I���au��P&��� /�A�A���T�s���"�i�vv^��G�� ���Β*IS�{�G)x�QQVC��Z �L��ͥ�b��U��/ �:wR�9MV}>�}�4�5e��@� ���|=l-�e2o�Hن�YY�XJв�X��0_�i��?�^��v^���e�=I�l���aysnn�5�[���\����r��e�V�pw˩ ꫻+���Nx3�y.6�5�+Z$p�V3e�G��L�7�e'����,�927����Mk���fn�re�i���
p(v����ˢAL/��������\��jtŇ�{��M��E�2�
5{�+���H1յ{>��ǖ�rn�߿r@�n>E��\�W�.����7:��Y1c�L#r���2�1�9����Wj�[ �C���p.��5h(�w꼧�Ʋ��yl�;r��|�iڒ�	$l���I����*S�����m6��5��M|�n^1%N�NAM�vP�Є�{�{OR������qok^#��8�K���6bG�i�qq$�e�zʂ�����j��|�t�["��ݔ�&XI��5�G�����9ǓӁ����.NN�#�]H1e��49&t�X���׮%�:zA1�5c�î�;j��ρ<!���a�z����)x�,i��
��*�tZZ�xG��+o�}Y��ܮT�Χ�z�0
�d>i�i$���6b���觩�;��R���t�Cm�P��\5�K��,�)��\��B��͚2�Vp�	6�y�և8�7�a���u���xK�>s٨����XRh���ǘ�5�J
݋&���}�W̜$��7�������J�Ub�Ѯ�up_����n3�/���7��&s�$[5Ժ�q��"a���8ѽ��R�Z�T��ezN(80�$��i� �3O���}� [M3]͂��Cz"�m�Ž��71nN�$�OLX+"�g>`�laN$�h)�-��n+5]�W�Fƾ!AY�Y�&wt������b��5�y� ����P�����EKn���
*����,pk�}�.��.F)����:Ġ�^	x��CI��ې�M��h�<P2��E�Hte�Nq�F�X,S��O��>C�|��Jx�&I�߯>�Ѳw��m:�N�g�jf��港UZ?nh��� C��0��i".���e��/�	�ʨ�Eğ�!�����u���eQ�5dm���oa�������9���A�{����&M9&��Pz\D���ǅ������2�l����_8�q*�C�����	ٕ��dVJ.�w��%<�l�Y�z}ş��<鵧�"�R��n���Na�̠a}ڊm���x��6jd���1���JX0�a���,VL-J�e�voN�}�a�=��/��v_�%+� ���!P���!#�P���^ۿܬ�КO^�l�"�cֻ�a[؃����J�Z2+�lՂJ��ݰ8I���b�������D�����l��!�f�j'���)�&�לک&'��m;��i�2x 8,8&[�n�J#��VV�SJ�>�G�.N��F��@G���KE�N��]�r4e)�{��y���2"���(��w^�?�}�_?�7/��d�D��e=L;ǎ]�<��$���2/���Ã�gu�9��w��B���ݧ�3}�4�}���M4@H�ht��iZ�͍V��S��f�d�Y�R�d��R6��T.�1��U+(˒�&s�W��u��4��l�2+\yWX�\H�'jǗ��W3�t��LV�Z�6���[L�<�Z������_��K\N]s�F;{M~���4��e�G����S>٥���Ɛ�_�j-7VN�*��^��v�Z}�i�{$PN:���?��|>��s8l�E3��:,��tD� t��D�`#�(������7싼�E��Y6�����p#��t�'J��I����+�V4����� p]V��?>+�C��D늻�*i��v
��g�[�}��;ys9Ջ����N�+}��8au<����dh� o�u���%��I����,fpq��s0J�*A�#�����9�p/���bMHc$;�.�M��L��x�����Q�2�IXxo�"�2�ޕ�_
r1X��Oٓ8|���bF,��rȎ����Etʚ�;M]@n�"7DO���g����D�-��R M[��!B
F)�6��P��^�2��1�h����v��R5w�z#�1����:Ѹ�r@5������l��"���2}V�Ip��M1��7�{��ܒ����ʮ��K7z@���Ca��\�\�UE�k�_&�R����Z�fv?��S��޵�����>�XP��)P �\
*|0"��>�����W�>�����	�B4�%``A�����Yk�~���&���~�t�쿁L��Z��6����V�	2<MFKetMa�ik��=J&o/�:WK;Xڕ�bȰ&�B�7�WL����o.ȕl|vi���k�qb4� ��aK++w�o��;%s0G_���	��������߇���_�|�U��j�^�B�yX %˳O;g�pE[����{�=�[[�_-���/�%|�W+K__�^,��l 1���ˮ���Xt�r���P
������6<[��B9�w�ċ�EF(8�GB�[��8�+�6܅'��^���-v�d�b&�4�8��w���WM��$�5k�v�zx�tNM�15��tM�F��:2d[qg��%}�>^G�^����Ɯ�1�M������K��{��v�(��]��ߗF�#ń�?��h]����ġ�?_�L�,�c�"JPy� ��B��̣�[�:V��� N���ҿ����v��}��p���]�֨�BP+gh�Ep6ki%�v�g�7
�2G�1� �=L�'��\�\�2��V����j�	�e����d�7P�,˻����x� U��ug{�(~�n��avs��]kc	��zp�g��4U�3�\����+p���5��ƫ��U�Y�鿉��9SB�Q��#�$�pc�RW��ӷS��^�6�� I.Q�4*��t��U�>1��,���-{�X�	L�`,�!�k�j��g5�2�=��S��F��wϛ���5T�;��^�L�dtzK��v��aM�7J��&wy�rE�}.��K��{7Oa�iSEs��-��?r3�����A���C�'`7��5�T��R��
����������Qf�\I��|��dz��b�CIV(\��	���i�0�.~��|%���d��M=�DɢTM%6@P��d�Oa�ĈHS�Tަ���-2/X/I;.1Y�5\T1�t0��.��S�����H�E�g!����#�:��K�`�)gʱ׃�������U$;0K���0��'����=7L������6ac���u�oX ���w����"Њ���{�o[�v������-W��M���4\UI�%-����R�(��e�����}a�W���vX�zG@aj?_�矐 ����wYyi�f���2���+��:V�<h����5ؒlYy�d͝z R=��K��.^Д�D��nڭ�>г��p�V�o��u�$����Ӳ�ӧ���uqm8����}���p3[*�ܜ�a���ʻv�ْ
[+Ѐ�0�̍�]��YP��_���T�?g_�as؇_�=���{�vڄ����f��e+�a����E#W�xXi�蘩�7Q�=y��D��wهT���Xu6a�T����{�^���^����-٠}	t<�#�F�Oh0�.�ǅTQ��Y��G	NƚTC>/A�.)�$6A¦��u�Aύ���hА �cVF1���r.
����ڧl1���a����zp'�JN���I}֓8���-�]LC� ���?x\zI@X��c�7��FT��U�Ŋ�^�� L
��Ðk�yGjAPSg��lV���ts[w\��}|ܲ�PC�]������`�j\�ső��J�+[��:���y�2�V߷��1�b&�J�9�����ҡ����u���
C��E�8'Y��·l��a@ �P���;�6SZ�m�~�ɑL�x��r��.�B�}���j�9!_����{J\+���D6���!�,���F=m���9�k�a��~ƹpZ�F�(�-R�"d'ٗ�~�ߗ��,�R����N�b���~z�j�LQ��!��W���^n�E���R,��Y�U�Kf"?F�ix�2>f��'�p�Z��Mj�o�R�h;[8>��WY�v%�a�ng�H2�&E��)R5u|��8�1YS�Y!��s�����v�,R��
������ٚ����v}ԺBZ���Ó|v�.���N�/�,�w;[Beƛu� X<#9�E����C�F�@�*�Qb���}����i���s����5-O���2	�ީD�f1����3w.�`n���pjS
��{+�^�M���6*�n� �-2���- �p���^����m�{�-��7�hDeB�d���c8���"o���0�R�,H�Cj�S����^�RU�"~����>W�����K���װ9���k����7�˿Z��e��۰�	�'�fd�e�}l�nf�>���l�س�6���&���>�Ҫ#��wV�gK�s1���ʶ���dfdb�v�n,-���a��2�e>�_��f�Rxb�?�@8� ��i�I�O�q�;�V���+qS����"6�L��2������E�?Z�v+ua &��5d�wN'��@O��!Y!P��Ϛ>+6�2�����Y����4�}�Tv)�8���:��43�p�n���52���e�|����l�l/�!�ώ4'PM� 3��A1e�x&{PȰ<я��]���������VDx����ټ���0hpn�oJ���lz��ϟ?+�	��9�����Ի�����ڔՌ}F�ߦ����+ʭ"J6�r`��1��ƴ+�Lcjeo.�t�d��'%&}�ΠYK�ấ�{:ǌ˱p*�,����&���S���q��Ol����+{�&p��](���x��϶qNVvrMy�����$FSe$��Uՠ3����$����K'���߭w������}ƫ���|��e6T$��8갰ףW�y8��bY�u���=�q��d�!�ˍJT��gm@�����T�A圬�U�����}�H���a#��Vx;w~+��A���0���ءA��$
IL� )�>�*TM��P�����qys#&
*>��O
i� ��2�������ߙi��������e� <�)e�X	�"*xQ�K��ު ׅۄy�;%C��ڐ�I��%��D�>�/�F�Y{9[�ޯ�����<�⽻��Rބ�|�������aj���x~�m4��?sR��3;-�m�C��Us�M�<y��`�L�+�v��l����� �t��ZyF	��-p���N����-��v��z[��ɮ�t�ؔՉ�P�wB
n��P8�z:!�������hCY��H�&�p*g��_�h�4X�䩠l+��C��K�C���0�Lד�L�gMdh���T�7~N&���^��a���.��=����S�p���oK�nr���,4�2��U�>@*�9�ɓ���mX#�h�Y���el7�B��q�%O�?�u���0���LӉeʀU7˔7V�j�m��Ls(�B�:�EL�$�Z�#?W�a�3��u�U�2¦��٪�Z{��1���N?[�_�ﮎ�[�#��c�K�Tp����ͦ��܈�	j""�d���|(���1[�$x��B�X�����R��cya8�l�ĵ�.ןe�d�gy�?��:(��,ͼ��cտN�b$���}:N]M���PQ��}8��~il�=��xN�5�����J���'�<H)�N�����Qe'�f�U[HH�,M���)gO��x:�����r���<�E`��v���I�V��s�en@!��~��'��G]�8a�N.~	Q}#m��X�^9~��Xc}��>������x��(G��R��^7����2~/W�͇29��LS�~��Z
�)0�I�6Mi���.=;)��m�)��|D�KC�!@ƒZ��ާ�L����[�3��a*��5����6$e�b��C�v͠)�Y���U%�1d����J���:���������2���Lu�)�Ic�m}�^������ޝ��J�,{!��rO	\�Or�����/ANe�Nj�=�>�5w'���e�䝸lSYF-ĠRzg����^�^��ִ'���{��~'?O���i�O������詜c+�j�ue �}�b�������x3p�O�CVA��w�����������g��8��>�=Q���Q�+(����K)j��A¢\^֊3�t0�NY�w��[��Yq���>6�{tх#�;_�S��82�g̲I��/�t��y���U�n?��|���ѝJ����F��Χ�>|)���Iyު\��Kٟ��&�;�Ξ7��� G�Y	��UX�v}B)� �>~�Ӣ�EջJ�����@��c�.\)0xp��R��#/ճ�0��9�ӿ'��X�'�n�_���H�OA.)	��%�Jt��I��+��Vxa+$5�$��N�{���++�S�9�ռ_�fc8hƟ_��!A�n�<��Q���$���%��.ݻ�U����6(W�>Ŭ�>ؒx��mg�am����E�"��n>�+k+��D���@ H6k]��¼d4��6sljY���V�~}z�/knvo-�'�<0kF�T��b�����Ƃ�֓����{��ڕ/�Nʿ?~��k{�:�³p���죈����3Z/��!Tdm��VH��
��Q�ł�q�Z���B�sp_&�$����b���E�z��ăe� �9� L`#����p�!M���K�{�$��I"�G��5�D㦾�KU���$Pn��h�:#�Q�i�#O$�B�� ESs
����0�����M>����V�åC���\0ONF���]O,��M�?����|��]}6�x]fY�P�ZDw�AHK'�`(������߻��}�@��&�����S�������fr�[ҥ�iTŠz1�M�N�:�뻥��y�JR7���-ϧ 6e������2�sރ	s*Y	��,�;�M4�!���]z_�Q;���� ���ןJ�t-E\���i/��uhq00ȉ�� !	���&-�	���l��>�vSJn��U�*�{�M�]]KJ��em'[�G+��p���8E�7j%(����4�OHl�|z�����Q펒�MJ�v=v��b�O�i��7���&���g�/=;��6�}�u^�~�<���=+Q��
*�t�+ǣ1��YVH�֪�R���ޘE<�P�f>��$�'-�+�l�DJQ+e�����<+�Z�h�e��=Τ�g�V�*01x�Y��#�C�I���ic��챣�AI��wé��C��vP}�s"6��SJQ�y��y�
�0i�۰���|e�עu�&�O!��5�Dgp�O���l��ra�f����׍�Юfǰ����JM䲦-�j�oy���C)N��gR����]�=W'�t�7��� ���*�p��Y>���Ωm"��ٺ�����pOD����F:'���z�p��lM$o�jQ^N�.D����3,ʩL�}��� �d`r�cS?����s��PQ�')%;~��
�}>?z�-��K�+epcAM�<��ķ�R�:��:���
�������-�p7��>�S ��8�)R���ʂSi��:|���O{�H}�@��&�X��no��~��óZ�JS�L�-='�3��`}�,ck��e�__���.�m�x�i�^1����7-����Sk�į�Yٟ��ѽ��`HTO�a�r�&��Ӗ���,m�B�V��ճ� |�
E8X0$x,��m�:�R�OP<��������Q��H� ��
qX�l��*�γ�7�\ٝ��3�p�1�s�;6���b&ī� )��D et�RRc�c�{Ez�S��<~T�S��vt�s���lH�5R�Q�P�H�P9�֭��w���oD0�QI ����zk�����敝��� d��_^��/�����-|�oCe%��n&y����k�>`�I��DƁ�/�ē�ߥiaR�er�p��ZDHol�c	P��]����h���&z�����zl)�KƷ��J��B�;e|�Kٞ�u�D�U�%\Y�0J���9�t�2�Ϩ�͋A9E��ډ��vj@0��V���$�{�)�H�ү�<>�B�2���n��b�/�do2Pf�ù�@fzI�~�1\g��%d��8�x���%�uw�-c��ބ\�?�j	�lN^OYG#(Y�TÅ���ųel�����3~}�yCo�4����6��B!_}��	뗝��v�5�<xJ�L7�B�O�m��L�7[�t'd��8 �ΰ8P�Ҷ�ן�FC	�(f�W�� ��"�:#�y/�#qU��=�4����K�2�^��bZ���0���2L���=q� ��̠&��t�w�>?~K��|:��S_K�� i���	�)-��W��}��܇�j>�����LZ�����ׯ��5�#!���Y��$��Y���߶��y
���Sϔֶ1��� ^Z�P֮9/����
؀�f`��)��y��d
�ӟ���$;�J��A8�X���cƐ������W6�]�	*P�&�!P�BxףK&ݳTB���F����I�2����-��	��&�i���}����	�w����5��We�C$�W�KpK/�� �d+qT��D����hf�`��m�\HpQh���&&S���땤�����`��B�eFP��w�a��See�x�����1k�fɲ˨��;ze�%������ڦ�h��X����q�T9]Y����fZ*�{��:�dY���[x||�5���&����y�L����J���=`=���R�-$+w����XF <���_��Y3�c TIA��bs�b�������I�pU�P��3t��q�5;��o���R�z2�F���ت�O9?�7+���� @���ĵ2w���p�����I���^��+@�[7zn��٢�x*^�u��_4rQܬ,�#��[�@����}���*�,_�|������?�i�V�BJ�@�����}*J��@2�]cA�zi�r+OY���2Y9Da<&�խz�|�/��[=(N/~��F�	�~^F�?����_��/1��(��x$x��1�i,�=.��W�x���1�s���h>�����_{x���3e||��̇
�?d~)�%~k
�!�822W2	ț^����4�wחsz��樓V�`r��d䓘��R�O��l S�os}
���0d�������p���&T��;a�Og�ѧ�6�F��]�aK+�,�uʴ��xV>h���W���2.^[�x��Y[p��ms6�%+�Ky9��B, ��*F��&|���>��7+k�R��z�Z>I!ׁ���}�W@��^��DR�r����(c���맗��k[Ъ`�XpG�G��"
����47J���( �<�S�&v�Ww����'�u{�����Vi���ab+��		W�oW\�2@>�	FԶe�+q�Nh�u��-��Źw|��nH��&� \O5Nr7�6����"��j�Y�xs���Q���uù���χu��˗������0Fu�J�</|
����"|�=�d��[\�'�a# �Pa@�x�('��}قc���d���AL����e���d/�X��� @5�Ӿ� ��(`JN3;?O���I�"5߅�A��eY�x��+k�rZ���-܄M���$84�4�E�m�p�"���L��˟������&C�?�������Ȏ &���-q�u�ʢ�����t�K�&1�$�\�x����2��F3=�;�/�ql}�o��;��}Evg�{9W�v�K���}-�SK=c�he�Ag9�w����X3}K֞@эz�I"_rH��(��`�~����֣Ŵ�l���΂*2G�<�<��15�,�<�'�ښ�Ͳ�/pP��"��U��´v�>W&u>nãUk���.�ځN+跊���į��/__4��w?��}3�,��lxx��ӛ\�Vfc���^�B���Bwk�n���>s�ihQ�qb�R=[���;)/�!F�a9qͿ �#�y���ݨ��l�L�'�|V��W��{:2;A�.҃RM,XW�
�r3Y�ϫ��ek��o�'n��JM߷�6<[i��=�_�ïۗ�n���Fګ2�Qz�$q��LQ1�!.in�w{@�m��e&SavX\�3�8��U�F+{�����l���l:������m��G)U(ë3mt~W�Tn�{fcX�8sI},6o�Z&���[H�L���u`6�1@� &����s\�nZ��/�����
��:�|I�<y�&ǮK�6eW��*��4�F^��Mާ�WWw�0{5=�:Ρ-��mndA9�>|���Cm��6���Pm�%��S$�l=�&8���<�ۻp������7Q�%sp����CȐ1��<ׁB���<��z#��� �	��"����XS[�k�X&��>١�� q��VL�N
�����3d�_-{������~�gkM��>�q�C�fl*6}�ק��X>I�Trk���ٖ���b��<��p_�ng�$���	�x��٣퉎�B6��6�6�E$��Lb%u�Ro�Q(	WQ�����2�`��@�*�_ݬ­e�w�7v��<��_n}9ɻ�v�G?���u��*<,�ß>~�����݃2"1АW++���[�ۗ����5l�S�I�ص���D �:l�
{3�\@]J�v�꺧L��'K�1���a�K$��D�4�ɒ�$'�Oq"��d-���>��TC��w\R0	���n�h�fp��,��i)P�	����o�T�2-m���$ƃ�ԔO��k�;@P.��1l ���>d�Ț'�_
~�5��<{/6YD"�����QYT���(mӡ ���$j@ ���(��G I�&��C�4t�	eD��n�gO��8���23��Gs�ޗ�1@�/��Y-����2j$E_�Ŕ)��-�G�� �͚�Q��mO���Ꝡ���Q-!�R�lEx��~ѡ��ކ�	���O�:�jk�� ��~���߿Z�C_��KD�B̨�+Z+M�Wm���@ہ�<���G�F%}�Y��y�ځ�=h�@��$-=먢,<!�⹋���ۇނ�|z����[칃}��_4ʑ�F��Q9h��Bn��ad}�v�n8+3,8�����
n��EM{񯲨���,z%�-���[w45��v؅�^��ߟ��_ޞ���N;-کSUv��� ����eY�"\�9��I�R/x� �O���)P	]��@k�Mr>]$��Z&�
�����Y^YD*?>}��썌e���4^��Z8�o�1����n� %|�����{���Ca�?K�0��ܑJ��9�q���l���G�?�b
�L%�����o6(Ӎ4�"f�`������j���r��󚦶Mr��`��O�uo�����WOgu�~�!�\;�J��lsˈ� �~���w�v��r�9�	7>]�l�u�L��������JA&��9�x�Y �҉K��Ԭ'�e!����oည4�{�C�o��P�N27�>�k?�ϾZ����/���g�v�"]=?�N�?)����R�J��m-�#g�d�}��#i�e�>%�ڂ��U���f����=��鰣G��Q}d5PrJޫ]k�B���zvn�֮�J"3��0YDa�@'\�={&ǈ^Hb��`֮� 8�mm��]|����4�tE��s[(�6�H�����fJ[|g�Z�����翅�6�b.�s0b܈�Ng��Ɖ�PvD������'���5S9�J\�'��`�g�z�z���9���ᔶ�I�FOMp�ب&�q���
���3�d��|u�#�,Z��I1�]�A�2��#w�#�7�"�s��B��28��`V�`C�^���u���wC`��n���"x�A���Ka���I�Ә6��7ey��L�=�es/&�� ���!��)���99�^T+��ħՑ�,��<�I�+����fY��Dx������2��i8O\}��Y�1h�iCu(��@Wn[�D5I��Q�MY�7�@�0��Tx�$�@�B9s�zr>%a*$-�����'GpS9�Z	�?cM3��^��/�O���S�'��O1��>�
"�ezO/o�=vךf�1	޴m�m'3�����5 ����r��kVI�+��赶���)5q¯��,�b^�A)tY~�`����0���l��� �Zv*�7)��^�j�3L���=,����*���!TV��h~�F�2
[(;t��x<�E<�巟�_���h�RYav��r�egRPf]�q�JNգ}��"��݌�z�$�:�]J���'���*3��5�A�*�M�����e���n��ܔ�zE_A�ç�>�;�.��A������z���t聥Lk�+��&Q���N'm���SS]��)��2�=A���5�fY������X��䵽Ov��$�aʺ�n"�t��CĽ)k�.3�Y�b���Ir��Y��0D�d���-����}
�����>�,{|����V�p�k#ww&ʼs�Snт�fX���l����s��,��0x�vб��J�.����]�L)�.b�2�����
χi(
��Oڨ�{T��ޕr�;�p�n�,��[fAQ,��}$����W�^c6U)��ߓ�[�`�:h�8�uu$�����y�;9��~�C><��s�����q�Æ8�d<��d���@� �U1�l?��[��v��#k$�X����{jP�Qѩ~�T�v�\U\Kɀ-x�J�*�bb�X;��ap�˼=w�I�4w@�� ]��[��8qV�+	CΧ�z1��lľ��]�������e�>���-���?BO�O��)J�Hs���O^^v�q�W����R��2.h�l�=uj���o��I� M=2���N��~G�H?|?*N�D��R�M��P����n�q	4��J�-���R��	uT���"���Os�$�#��]�Y%i�be�8�G�UUC��AT���SoNzY�4:7w�ulT�2[Am�������Ƭt+=&�(�d�м#A�s^(qP��Qr�O&������h���ZO�� ��!XPf����{j�p���"��I;\���Y�Ķ�[B:�<f���M�A�:e``���(���d�N���W;��K� ��p��������:8��^%ӛ��s�i**vd��� ��n1 ����t����ǚ~Թ� �ğ:�+�N{�O��;�[� <W�بq�8o��Y��n�ۣ%��Y��oO�0�b���Wk��?­���XB[������׵�CxZ�Z�f�e�`S˄7��s���kKvH.a4s�ׁ��ݓ�l�������
8���6l_]��<��
��I&� =S�� [Nm;��a����V剓��wiU�F&'
a���R�t�k���ٿڃ�H�in�A��,�B���=dD��v�R���A\A���v�߶��o�C�qˉ�@3�}6vrT�\�7w���m�ia�I���5M����3$�{_�B>~�o����+z`��t8�K� {�2��U'�	m+y1�m�$�А��� ���3��Y�m�6�='���ߖ���Z�w�D�v秔!�'W��g(�Z{ax	�_�iB�^�k�/�����&L| �J��q)xp�˨+G�F)U�ݠY��k��4̿���YߋIh�W��n+�d =��䳍}�,"��6GS���T.~��,جM�ʁ*@ԁh:��Di�k�I���8i��+��l�ɫd�r��b/�w�ָ ��f#�^2Ν�7��S4ꥉ��Ȼo���_��Ƃ���vy�p������V��e�Vt����@�Hv۫'@�"ך�|�bY=@���qʒѪ��y�QԝC=�Y'��ثI�B\M��.�_�Cٸ�Ϛk��K*�38���X*s���-�J�^�n=��9�A-��z.US��Bm�'���"��ʆ��N2�	S��{��w�p�/ ��U5����������º9�����<nvk�� � ����i����\B�3�&�v#Q���E5׉ǔ�G�*��r��N�����Ox�������LAN"��m	~���_�9�����Y4����w��]v���Fʰ���ęJk]g��T�(y<�Ig3��ܹS� �>��.=7��]̏u���E�'�t�~����i���W����A��g:����J%�D$Ŵ�3M�话U6��0:��G�^���H!O�Y�s�\�Ų4�r2���CY�J&dm��P��p���a5*E�j}�'T�l>-�/�8N�E-D�D�`l�6r��3����y^㬌�����_��W��Շ>�{eҴ��l� �k�����w�:Wzϔ��]�Y� C[Q���ε��9&��c�zɺq��Ji
,��j:X�iu��s��5���������`�^��"����ǗW�E��ѭ���]x���i�]������:A87`��\i���������W��?�|s[6��<|�DO�ח������Z��E��@�on�������'Q���X^ڝ|K���=!���F���T��c��v �.��D��4�L�'驱8�F����l���iSP�7zpd���656t*q�K��S����Ry�8�*%'�qy���C�
4H�x�4�L��R|(/?��AA�yK��!�M~���!�A�k����J���Er�
I���{�� ���I�a:#���=���@��H�n���h�8�Q�X�C���^�3�)�Q�I��)@�@������B�EqY
Ǉ�k	F�gĕ��R��Z�կ���l2����yJ'�)f�yn�v��P�A����$��u��ugU1�̘�VM�z�I�Ɏ }�W��<D^ZH�t==�_���禗BU"@���]t^���X0_Z@�E��C?
��E�řU0�R�|�s�d"'�G\GgAPJ�r%m��Q �(v�۬(Y��j|AC���cҡ @��:�����.��z_�����{���~z�Ug;�&(X8a��>]�[�[�[+����(C|�.��+�G����F�W�r"�6��[����2���֘Vjs�ַ�E0pa��T���Û=��v��ŕ&��݀"�Oc�&#�=���r�`��Tds�,?S7��V�BA�f ʯ����9����fwq�� !����UXo�WSU鸴N�D���,���:L��8��̋�L.�,$a��s(���M
$ɔ�&y���)�@EJ� ��T�0r�����i8r���eG��Nz\A�y�+{�W���u��A�A�����)�=�]nk������6�A�ž`�Y�EO^� ���b�_f%�Wb+�c��(+2���˟ס�Bq�%a�Ԟ�Kv}Y6��G�,�����c�ҧ��c֣�T8�|6��%␅�V}�� +'Z3|�@"�"��r�}^��g9�嚸RZI�{� ������-����� ��9余�Hf�!Nl1��zi���:�޲:+�Eq����,��֓f��P$�#�N�V琗V�z���+�d�ә�Q/��<Bw��β���7$�W}��Fp�t"�%\ْ����p܇�ۗP~�r��M��t;_��l���\�������ه�pu�����p{/B9�+7B�oo��o?�~}~{� �z%�1ѕ�Ej�6-s����86����`ԜC���h�c[6�͖1a �/�hD�S]�a4���@K�>(����*���篏44J�Ё.��S�t�;(�҂�P#y��˼1�]E����1_S�^��.���O;���R�&E��
FY�T����E��EqN��ٺU�!����;��wp��Z�K��m�d�S�4e����5� a��b��aHe���sIf��wrNe���/�OѪ ������,C������	���X3�����Z�;M��F9n�(��fP5�&	�}�½��YK8NnF!�k�*�\�A��|��36wku8��6x�YRk�-��{.��� =9�f�J&��8�;��@�S}A�F����Z�,^[FG�Ũ�쾿j;������8�W;��(ap���,�@Y(��ZL�5F?T}@@1��2���⡓� c��̈��*��)kk��$޹>����vP�fEv���W�����a���Β�uXb�z�Q}K0��ve��흝����5<n�$U�z����`�ݡC�
���MC�ˢk�\���i���{Cd�i�,͵����1��\`�{su�����L��,=��� �&�>�~w��Q8�Ǘ'Q�$�5`��.6C@YΧ�>��i�U�qxW!����kǒAi�$aK�2�:*ݎ �c*X
�}	~z����i6�^zIRG9�����(�����KV�5��,�4�琽ϧWe����H3<�{^�
�1�8
�������Tm���_ځy�����3&���)+�l>�tϒϮ��~�f:X���k8}}	��&�N�&��z��	���ʲ�X�
3�_<5 r�@�
�����N����W�d�d��w�ƞT��3>˰����FL)��(����C/�;����	y>�RJꭡ�Q�.t�{�M�cj^��##��O���O���f� ���YZRR�7�z�!$|��q�uI-�i�5�;��V������p�R��ԝ� ����ȸ��~�cv�����{M�k���#���)&U[=���YV�5�PXz?�4�LY���^�҅�q��ܼ�
����%l�{���sB]����s�[1�=��l��T7~M��p�rx�l {�R�kKza��a-�!w%�l iX�CA�?1���_���Ls��1e�+*�:kܗ8˲�&�|M#iw��閜�\Om�܏�NeU'�m%.+������x�p�2��wK^¯]�_4�T/���]��!��T0��ˤZ|�j���1S��}q��)�;�*G�X��; �`�^]���.ј�A�6�3X�j��BnP�Ct�&��>꾌2���K��-��������$32�����p����ˤp���C�"�>n�kx���<�����#�_�:�R����]���}i	���Á`�;L$s2/e���6mL�-����.n~�eH]&[N\��e5��o(P�|~~�=>Y�;���)PM�tdm���Ya�ϸ7tF�xI���CS��{��\��y�QA�iv=�0 ��܀ay+��To��!��=�S�q�Cʴ	4�����A5u�S�����R�=7��cX�b��\��AS�eh���L},��y��������ihW.�L�����Y"�mr��W��)N���J>��!�b�t
��㐘�Y��g�v��<y`bQV�f���u��2��7��!�����u>�e�=�ݫT���Z�aDZg#	�U��۪j����IT)>E�T��y�\�$��&ҼNR�I��v�H������.,�1D��!��?y�� $���I�+;ܶ����B�w{6x���P� e��	Ы�C;-��ݡ9�I����aa����*�ȋe��E(�֗��N�_��.�X�3Rf�G�wHEi��h%�XՃm	L�ȴDh����ص��]d�d�ݸ��'�{�;D%� ��l�
����։������i}h!����'����NQ�����n#�KXo����ԕ�\\�<�t�M}�,�(� �s������ڒ��F��^9��3v�P�n���=k-�#QxS�q��/5�c
)U˭UP��=�Mxۼ���]x���,�)a_{}���TM�<�e��bc�~C(HYvy��bHc�6�4+UTe�]Y�i7z.�4|�]�n�H�t�tRFh�؜iB�Ol���޲���ߔj;
�:��H�a(\��D�?�u9N ���&w0Rߟ`�ɩ�d�@�1g����Rp���� �S���p]lN�Ys{ �.�ݫ�\?>>���d,=�=2ѭ�(u��!|�A;�t�$�c]�@f�*K��j4�����,�����ep�J��?dޣ7����G��#�%���Qooyu5x?$e�wS��j I�h�C`ui����)���r�>v��a�ԣ��pb������-l�����^�d}d%S�&���o�E��["��/PL[�&�쵯,���׭��
e��W��: D�_TY��HYv:+$1_R����lW�;5%O"��3<d��?�G�����;W���,R�
����'NO�ޟu�� '���]F5Rk�M'3i��S�XH����%z�������e��t��[=6��`�XM#y(`=dn������:jr�hR�+�@l�W=)�7nU���lo�˱��Z�\4U?�j�!�!b�a���ˠ~���ҍeN��4J��`ԲpQ��|s���l����[��^m��44�+��.[�̨�SG-��#��b�{?���[��#i�\���t�T!UЎ� 0���)<�fa�����B��c��E*� �8����no����N�ۻ����?��wW�E^���2Q
�� Ǔ?'�Av���Zܛ��iX�""(w,���.S���q�6ejͥ���A���E��oޤ�{���.FP��Ր�x�t��@��=���*�gT ���P��M�ļ����5q8�: K)�C+��dNl�	��.BI��JQz��嘤�P#QO6����`b�{{fӥ%��(�U�ѷU�j�6ZS�=,�(����7�� >��~�t�=���m�|9Z�cZ���a�@ǋ�3�O�"�-z��Y�+���G���`��0�@�T�T�=SR��5;��l�~�h����'�����R��Dy}(a;�_���a�
�da��h{��oU�5�7�`0l�#LD��r�|�>�������������H�O.����)!#vW�E�|}���?��3�nȖB#����Z���Uq��\geYb��ۛ0��_�p޾��V�ި��]�4ki>G�g��K5���(
D�T�D9
�x���,s�e--�/Y�y�~�dR����}J(�T������ p�A��������#�H'OIj��� ��b�ɣbEe2��vcSv�T_T���ܒ��!��w��o�4Dh�1!��Lk���C�&rt{ٰ����Lê���wx�&i�������U�6̣墸�t�-�'�	�F�_-�PNU�g��<j�P8�]"�� ��Q�j��J��룊p&�t�Gn����Cx��.e*A�G��o�.���/�w(ŔQ`K>$��R/4�ݾұ�����q{ �tO�x�2�v����'�������q���@ok�Z=	:��dD~:J���󎲳��~����r*qm��e��4աM�L�J�����Qy�#p1H,h-� ��C���? ?Zb�7n]!�"�;�a!�aD)n��5��Z���6�x�1|� ��-�ۆ��j��Ɔ']�2�
�۫��M�@2���WJ�t&�����l7h+3�Ȁ�A�t�2�2�^�[�!9��s+��d��&m���o�X��pc"�;ᏽh[:�#h�;���<�_��
O/�x08Ee�N�,
��(U	�X� �O&�>T�}C9/�����;(*Y����w9x6�r��->I7����,�����a*�h�Č��: ��K;��?��ݐ�)ifm^�C���]��W���eػ�t�ʖ�]�1�f�}ꁌ��?�-x%,�W��J���o�sɇK��Hlȧ^`����������v��$�,��X����@���ޠ�!mD�,Q��E�[�ķ�gbc �Y)n����)�\~ۃE�7������Et��ʳ�\����T;ʵgY�"���R��!v�>h)����B���j���M�zO"�o��9�B���ͽ��2F�TxZ}�}�����g#)��{k�(Gg0Qh��������m8�&3[D�d�m�]���b��G� �����~X^���*W���NJ�������G���B(��N�۰�����]�����J��+�W�a~{�O�/?[�l��R�IP0xI7��f�l!_N ��B�DG�SG���6�����в���?�c�'u���C^2ש�cϋEΐ �}@���I���\k�*���q*�kR�MAC�B��l��1�TH�_Reo�Ҕ�'�w2V�5q8J�����������좢ˡ�����.�Gi`�x>ꋤ��6F��-�l���bI,y"���綦��P��X0�=�������P�JW�p�ę	��P��z�l�W"ӦԷ �d1-�� wG�5� �����,�m��h�,٠��%�1��W���gC0S��8VO+%�+~��͇3�_4�)�{d�����@�ӿ��;�5�?��gRvRJ�dw�_�szN���V B���$��ϧ�@i��&X����ry�S���2�I�\�JmG�{�����	�nyQ���<���W�XZ���	�����~x�~\�;E�ٞ�5�*�O����HSѺ�-�U�*�@����J�o>�b�
��~��8��odM/�OX0��S�\��Ne)&�2�s�����hg���X�iQ,�f/,S c���!|��ѧ���K��t�S����	륖O%9�XD��V.�IY���Rϯ��*{�%���|��3UB}{�4)�*bɓN޴໨���	������w�I�lk;�޴r��[Y��$����C/*�����O�R4��_L�9�
��x
}H@C���\	���,��ώ �.�pc�w���G��S�\��U&b�q�sԫ-$�K��K�L8�3���N[�L%\���A�����HRPnUS����9y=m���ɴ�R·�ArފnU��#��9�`�8;F��_�M��8i�i����y�z2�j�$��QE�u_��4�i@�����&I�Z���`#27z�P7�^8<T�0�o1y/=��b����#�2s������ۿ��ڍ)��9p��4���+�&�--�w_۵��y}
?Yp�g�;���=I�t)r���>L� �M`ѮW��S��|�?J������~q�t��)���;%�Si����� a��n�s����F�����׏@{��؇�v����TZ��ցļ&oܶ��fSzh��zP����.ڗ������5�]�݋;�e��N&W�6\z]���>�K�R:�Ԫ��L,����w6�nV��qFy;�b�gE�/��\�K��#�@�	�!��H�k��p�k�ӟ$���y{RP8#V��go5�����ܾ��2
��G�RJ��'�L�'��ڝ;�k��-u�U�!�15
�m�]	�3���A+���
�g.]ފ�Xk"�.Um�0�q��|��� ɒ�{�<߹U9w��2�'�dВZ�z����UG%bLǽ����-{�΃�l�=ۨ��(O���V����D�����P����O��d�B����A̐d�������;���d�~�bտ���E_��Dn3'��E'��a��~/'��o$ ��j��Z$lP/�����nBѶj��H�j?�z~���+��O-<ZM�Xx��>=����)��u� ����\���s�##fp���Q��Y-�#��3zlL�l��6oZU�Z�z2]�	Äԋ�����S�H�;�<�+{��2%pSyTc�ʪ�"�Mam�B�H����`�Iy�d��0�[�����s���WYyp9C$n�y��<�ŢpdYE�o&� �!�$^�,�E�U*����U�{1��\C��Zzf�
x�n��έDZ��XL�6qu��m����0%�vvX�8��|�aI��������!C<Ἃ
,�ot�a�-��B!�L�6)�������j���S�|!~�;�O����q�٪�V9x��s.sf���d�Ro�(p}����Q^*!	�,�����2\������hBk��Cye��C�f\�,S��(e^E6�=��b&޸�h|�^�]}�Kb���)����@����o_ �����|q-����iqM\����_��(���^M��{C�y���-��lW;�v��9���E��No�]��"��X���_�Gt��g�V�.sW0)	�7�k�(˒�
��}H�\��O��ۄ/����n�L�<u�I��޿�/�:���qc`-?�1�Y�j�fV�Hf��7�3l�7���g ךXFm6ъ�Fq*Ejc����;E�:eNg���g���
�2���D�u+�;�ɝN5cE�/����k+�s}�|���40w�����RJ���q��`v�>���"
��ԋb�e���t������2e2_����{��N�!��m#��l�� ;�ҳ6��Ь(��!��WM���&x	C0��&�J��VbU�����ڏ�=˜�|�Yz-�����3%0��za\�Q�WY+������;C��2�:7���� ­-U�/#� <�0w�9�ץ����Q(��C�~ԃʽZ�$�5|�u��Y,�`��F�������@|]d>`T��5�H��A�	9��O%����Gqݷ
�z��j��z�kV)̪��hk���ev�/6���տ��72��8�gG|j�g��E��9��|9�B�b%�I���wGJ�	���7j��gz���[A�Fo/����xޅ���=�}w
��6�Y�B��k���Hե��N%j�{~���_j�ίV:=x����Yׄ�( �H�����j�P�,�e�����!���8�V'^�b:u<^l�Xp�������)y]��z%%�N�|)�D�3�X��NB�����X,v�8��[�rs{����$J���c�B-�I��_�������{]��)j*3S�3�Hmw��x��/vG�����Qr[:h� ܥed�el�}Nzh��'�F��J�`(q��6���ԃ}���2XMꢹN:hryL�/���C%�/��(H�
([���K1T��22���1�.���t3b2k*�J����.B���\�5Y�3�=���O&��"�݂e�&V.�U{�6��-�X����͑@zm�'QEG��R���.jEժ,f_��Ƃ�l�b�e��5'���:�gy�!KJ�[m�x>�k��HF����E�9��𸆼��}�
}V��$�X�؉UrS2Q�g��Je�>�O�b�HӘ �I.�T�:��է@����l�%��B�C�D�ݜ��'7��rH�%�#oz:P5D�z=+��AUp"��J*�>��$LIР*Ji���xpB�'R��(�tќ�r�$�9��\�����(����J2�Rt�p2uz�b�mqB+����HcqS��V�ci���az�~�n��Uݐ�i�EJW➦�8��M��tq����q�B��xm�=,�P��o���2�S0�DMu5�Kg��p�gB)�>��<�j���>E�Ĵ�����٦L>���؀~L,�#ր�'	���|�FA%lpY�8Y澒��N�Ke�Dx��^"	���%��	�el�k�:���9��duM����H2VY̺��ԹC?�Y�:p��)�yxN������m�/�C�(k��������(k��F�g�� ��,�=�d�h��,	���6��F��2��g�{=d��yUQ�W�g7Ϭ�M��[7ZHv'���m�v%���C;�6j�V*op�.�n7 �,C$�Z!�}g2��9[���μt9�^���Ȣx�d`�1�G�G9}2�X:H��Q��3�꺰f�������n��A��X1ݱ�1//�{��x���T��͌�����!����]�Ud���.�Z��<d7��F�9�W²������P�-, �?<8��>%!���@-jM�r-���nqr�z�
����6�%��8xӬ���Tj��E�&m,֬SƧ-�D-S�}�Qy"��<�J�����3 �?1(p�M�G��`>$_�ʧ�*K��(}LTk�����RF�ŬU�IeXA�+�K��d�K�v���R(��$/\X	�֛���uU4���v�^���T�Ƚ��1�̕��u�C�t����G�(�^fF�!x	o��~g_���d�xO��EHӴ�F��\Y[*�%��r��,e��.�Kz ��U=�r����9z �Ş�����fK�$I�����GF�uuuw�l/0���+�'�?��3?| �@�ݝ�9������������"jٵ��E�^����fj�",�,�f�[����4�H��H�r�������������#x
ɬ�x��`��[o&)z�Ӊ327������Sms�ŉ�s/�&�RHk0����ԙ���,�	n�]T	�^��jS�M"���x���"��ߜ�,��r� `|I�-�Y�Ӫ"�ɋt���w�grZD�A�����sެ��{#se@qN�Ɂ\~&���]�/��4�4�6v}�\͌�������j���\ �T�K�@:�fK���m����K\Q6�2[w[h�8���ЫW��&�혌�.#o��gt�0�Ux�&2����:Nv��X�*h��>��ls�TCOP�B��?���F<��j};�G7��Ӗ�y���[����V3m�I�ѓKWt�����&Ɇ�f��hu�ud-��z����m�E\K�G�RA�����ߺ.n޽�E��}#�>��p��5H>\MX`5�\r> �I����5��9�,�b�u+�V�YN�xoťs\7�e9`Kϑ�y<}�̍�ԧ��B; v�L��qr�0��c��0��H�K������u��iΨ֍$~LW�2gP���Gvl�$��0����gP|],��yNl*Ljb$a���ğ6��������S ��}�]=&PE��`�B���3��R��Ր�����5��L�p�`s�e���2����1��]�(k$��44��������ܝ�2:�1}]Y���Osɒe�c����������$C#�1�2�R��t���Y��z��1��D�����P� �Z�xD�7�;�b��@���	^��ѡ��5�6�3�W�p�A�� ap�`n�紣����f�;�ED���r�ԏ̌��7LV5��B�
!�Jt�b'֟�	�w���j63�pՑ�=��1<�t,rV��x������L�ח�Y4/_��߱��T���$<�04���-�~&���d3%)LO�y_I>5٩�d�����3�b4bܣ�޾�[)�jY�I�D����u^又���Е�mj:�%��fk�vv�,t�,.�ث@�ט�Y�1#[���� 쉤�A>n�͘N��W46)
��D�!��
�x��3C����\?)�+��!��j5r��S��*Q�h�`�wu~a�Ƃ�z��+��\�sr�'�go���! ��8jM��{��'��s��8��L�k�t_��e��ޟX������dn9ͳL�t���W�������gk�9�0��������@�GOx _l�9�|�V�8�^���gAPY�j(o���o���U�� ��j��=����4�7'�as��%iۻ�{5�<`�M[�A.(g��*)w:���E:��^�w���Y��rv�%i2�q1����??��t*���</��"?w��6���	�1&�����$u-��M�)�����=�\O� �4pU:� ����ؼB��Q�<�Lj���s\�jN{2=�$Y��~��J�/��tU�֑CT�55zeR��ܕ�#���a�ꍹˢ']ü[%:���Ibj3�y"EM��0�$n]�1��T�%�\�QȎ��6.�1�lp��Qt��Y�G�-;�%i�X!�V
&('��J��10��T<aS}�;��(�V�;�3ag�hݞ:�w��}p.'r{@�Y	]0��=�:6�nn^kZF��w�ʤL/Ks�$�51�R\=丙d!g��&�a��u����Q��=���hu�g�L�Y:� C]��'����B�N����L�mw����Lm�avR,�G�Qa!�\/J>��b[���e\S��sV��2�I��I%>��H�;�;�t(�����D�#�~��j�+2&eG���ɓZ�^p�_��� ʉox�]fe��>|Y_���h4@�^�>����78�u3dfxy��AvO�zb� a���i�A�I�z�����/.��������M���l8A�(Xx�cǡ��
����2_*?|v�����
�q�Z:�08Y�Q�:0���fj��v1s��R�h�̗��ƻ�~s�>AcG%w�+NH.�4R���Ld�Tk����c�يgySKU�@k������W7���3��tG�2ʃ��n���.�q�h[�h��۩.@��B�C�9�'��9W�|�w@:��y�L�$�;�V�y<���`5��x��P�M��,��?�YӨ�d��,�۸^�E��hf�����/
�-�����A�~�]}��Z\;��EP+1�$�D*�5g˭�N/�):}���
X����󨮵y�Dj��^�a�f	,��V�=�F�'M,,0}$T�t�p&q��1#��V}{���ϙ����(�D��;\�34���؃zl�����Dk�%%�m;2E_N���>=Cd�+���8��� u#~����]��o��M���4r�aäw,ϱo�=�[9<2N��[�&c�����9P���B��M�-�����Ϲ�����f<��֦��ʭ������]���\���ٖi�2sk��gr�.��̡���GP�6�jK��o��=�i��	Ǖ�8:���T�'(�lB��`�-jtZ��pz����1�,������"�L�Zwp����D�����v�0(^�&�֬5,�����6#{s�Xl�t�\̸e|�2V�KM]��u��#��Įga)/Q6��U��C5rO3n�}�l�cjA	�!۟I7o
z@j���+�f'	mV"k�i,M�IL��Ɓ��!s�#-�N����;�e�M�e&��=á>�>e+e(u~.zJ�0e���לv&u�T�5��o1���\�~{� ����mjN~BI}�յ�"�
]��3��ֿå���TJ�*B�%w�Ǽf�ܚ�p|�n�X��.���U�Z�^@��G���롑��X_O��A����w�i���@A��p\����r��cb�|{v�  -6��i<�;� �O?�r�B>&�K�*��J��h�7�����I�ғ��ȝ�P��]ۍ�Ѻ��yA>�S�=�(�Y��F�EK�x`uZ�uRP����i=PQ����G�s�Bٗ��%�Z�3�%6�B��"�']U`95�n V�[g*5�E��dZ���1�������P�|i�n�@5E�6<����Ʊ|����|<�I=C�ct�%(�PQt����;oSozȢ�9���$�v���°r+#�x2���H�0E��L�/��\h�y�p@}�LQ���@q&q��������5��:�|h���	�8fL��$z�捎��,Ae]-�)ɺ�Kƭ����}�]�(��Բ�����`B��_�� �=itaw�1ˢEz�簃��#�O��A+���q����+��IAR7��[)�fa��^��Paj8+�S�J��X�ԫ^&|Τٺ�sJ{�;!%���;����� zV�}�=@�s��.3�s:Mc����a9[��� 3;��6�bxqnc~��Me$ybVZ�~T�a��X<c��0/q�f�^�(q>Τc����I� �Xpe5*��!ȖP0�����9�	J�����27^b{���� ��Zd���'���鯘�y}��{- y:���g���22,��/?�Z\]sVkQ���f�=��<P�]ߚ��&��8�� e(��h��4�.H��L%��r�;UI��	sM*Ki�ǻ�Sn:���ȶ8r���وQsO�o�C�ה�Gh[��!���X gK�0��=�;у˯�ԟ�TE	�!)p�%���P�}�Ӫy�on���yd��Y)[��>�ߜq���Y�{{��F3m������Wp3T�z��Я4O�.��̌;SҺr�f���D���Q�<����;�4� k�y88��gord&�k4.���z��T�Z����G _���~6Ӂk��_���!�4�k�S�3�B!�.�~�)-���d2�7�(�®Z;F�S�w{J����xf�����n�2�
U�\d�X�'/Gr���i}�N��f��f@}�NmY`E$��5�T �\���*3�w�E�'	�"���@�ĂA��SY u��8K�p+wD�F\���ܸs���!�25��.(ɿ�?g�VE��Nn� ���ȵ�����fAG��D`C�;�
F�; �j�S�I�	�lf�@������^ѫ�Ό-�fd>{41���g��ѧ&Ѿ���93tgrq��tx�#�(k�����H�����W�*��I�ا��$	PE];�A@�����Y�p?�ĥu&Hտ�{{��Ng_��V[t:W�ϝ8��^�#>c�k�|�^v�n�������^o�bk�MlG���5{�I�t8��cs$������	l�}�6�\���f;l7pzd[���l���C�A��H	��:ql`Iɵ�
+�?��xn���qMr��L�&�8v�(�#�x7nt���%}靕��D��Ŏ���+Ǖ,nltKp9��*@��#��F��v1��l���t�t�"a��F_�Q�kq�A�H�+o�uA��5;��2G��y7�P2�=c�����k�(������En�Ef�3.�ˡ��w�8����O�˜\���@t7�(��Ʌ��&eV̤Pz�>F�b﵂�y�Ɍt��Kc?o6�}���Fy��Md�tA���/w2翕�?
���������	.�"�*��QY2]y�fd�|����Q<�����;��v4WD��k���Rq8�8��J�(��X�+�Np��)i�2�=�t{����p�٦��እYv��	�x1��t"�Ou	�6�ݠ/ޮ�lظ����{&\�ܢ�Np6��B�9�M��
A�P����|��]a�v�MQ��4	��v�;	�dO�D�
��s{#����������z.vRj�0�K3�^UO��ni5��+o3+��AD� �0TA��;��,�^G�D��ͥZrp�k�YD��??N)�l�eI��Sͥ�q\�T�t��L����V� 2� 1�!7(=pӣ���4dN�+(��`ef�F�����5�wS�.pL�8q�SoΒ���ٌ#i*A,@� ޅ����#B�gi��䛡�͉D*P>2P�ə${�h
c~]�3�.�919dR�8�Y]�.��7��;6��Ғ�6Bބ��7�BÂ~4�t \���)�~B[�v�F4j@w�H�2��ˍl!�yZ�w��L�<��2%�9�/	�?	�P�Y�?6:�����vG<Q^z������05wр���=f�d �c�'���&�yP�}��|��%���#���q���f�R0�	Z��Sm����H���7����� �9����l�0@	�_�E=����k��b�0�Iڣt�|�=�J��/���@�Lz��0tJ���A|1�u��lTL��č�F�ٯ��ėB�sH�V4��s8�z��2O���xl�AF����q���^q̫8�.lO��7fO)��AxOk���(+C&��[E�۝'����N򫓨)G���v��7�I��l@��x��f�?X�d��#ٌܱ�o:�\���� ����n��&��S��T�;�OY��t�nXv
��B��໒��K�)�m`���*aW��`P��s��Q:��J������`��;2s�2�Ǎ�a�Bk:Nr�.^��q�#�I��ߒ��Qjdb����(0��F�4�.i��i�AB���Ժ���%x��\�^���t����V�-�5��s�$�
��I�Q�
�cl*]O��vg7��k-��F���_=bF���햍��80g9 C>��>�M��;.P�v���A6V[f��t��=s��XF��I�%d�p��0�U���]l.��⑝]>�#��0��5�g�L���X���'�$��4"5�X�m��hrG�M�Q ަroi����/ &�SI�ZĂ�i�e���9d=��D~A���s2oZ0�$֣�8��tD���]U��Щ��c�E]G����PL��QG��M
n��*N`��-do�`uF!5��A����NA]�u'���ɛ�n�}����)�O��<���.i��'�����z���z*��'��
!�b�}r:Lav�cQ�k<�$�6#�w�'��hn�ML���]��E�ɑX���,g���d��3DGs�g�s5a̐��e��V&'ň�E�n��vu(��� fH:����푧��x���7i���ܹ��hL��&��n�M��9 ^���9q� ��h~\��6���k{{s����F�nO,�;�a<���α�pI	�B���՚�+��)���*j�N�a@��[Y��2C.8��ĵ��AY%Z;�>@���W؞���qn
����y�z�	��۪�x������Ā��^���#uk�B�����F���7�YNa�����.߅�Z�o�u+s�1ج�����%��x�,���%pJ�]�xq���rr>�e�=(1�4���vr���@]�����	J%������,�Eo,�8W ����9���Qr�^��Ar_z�����������i ܙB8�cv��#Ae��Q�(����("$��h�x�;h������2��_z��T�,� ;w�1�5���K��Ι�y�t{ח�q��:Q�	,�0pp��藇�b��TԌ D:���.��L,N��2m�7zO�x�M�M���2��:��$���-�����o޲K�Ƥ$�fZ�m�yP]�'�3�i8�U��	�3X���}�~�H`�NK!�á����f�RNJU��n�����ʅ�����P\���p�a95�=�f+�s�H8?Nui.�͝;^�4�G肺�>1��w|k�������M�������5�5����E�4��[���e�w���`sn2KNJ�-�9��+��ZS�Q��8W��{V��D,4��z&��:����m��=���!�$�Fc�(I��f���E�:W�3l��y�L:����b�B0���4Ռ��N�S\Y�ͤw�� @��N�x�%�T�3�����9gg�� p��<������$��bS#��Ӕ6�5��O��*
|'a>f�3�,������=;�:eΒ Z�8����+!��T,��Y8�ʇaGw:6}�LP2ǚ����m��	�Q�Av��'�rV���y}�������.n i�XB�C���%z��c9'�Y����Ɇ�S<O�̊�
hy{v�7�5�>�42H��7�L]4�Ҡ �j�C�;A&0�<���f��'��A�0��nI�]�<��e���Ew&vf���gk��9Q�˸V��/-�E�(nGzUb�ql��Kfn�0=8x>�(o��[��o
^67\[G�k� �	�
��|�*gp��W���ѐ�&��ÃLAn6 �c����\��1�iu�K�_��ьVH�%.fN��ݲ���%��"�jz`����Z���u��f��2+W��ۺ>7�TY�g��{ސP�U�[��6g�{�X��#��s��ś�آý���Ϭ����Xl�x_��w��2���t�&��C�Kl8Rߘw�KSZ转���l��Z��\�;娡.75S���j_�5��s���=<��p���$�{Z�'�U1Ώ`c��^ꑓ��2N�N�؄QY�9
�dlX80��Y^taJ��&�1&��h  (�L��º��v��\j��C!��s*j�����en�?EY��Z��.�>��1IzTA/2��?���̓f�:��:�2cP|�B�\����5����������ˍy�L.K�:kA��%��ݲK�X��Z̩�7)�gS�$���0��Y񛬸�K8^M�᧸Ɩ���?�ò���(��iej�+q�C���B�
@�s��V��k�����AZ����7)1�L�(;]Wf�B����V]n��iQd�h! �i"כك��(�J:(�F��9���Ö��ճ.��s{�0�4�}Sd�E� l��2��6[]��:Q�Ĝ�N��Kkv,���؍rk8բ�	+p�2X����9g"fٳK{�.�qֆO�F�	��.��6�w��Ъo��a���e��]_(v����nO$4�#/g�2Ct#V|%��-UH��~�Y�G���QW�.cY��@��'��_�t}��M��w1�5b5��@����j&�zŹ�`O&'���R{6���習�XK���	ѣLN��$edʬ�\���<����4��,]}�uo����t!��۱X�ytbq�2E���.�-�W��rO�_���2߳��K��Hʜ%�T�e/)���|�`�:�ϋ��0;bd�I3=	x׭U3�-n�;@r7h7p�鄓�c�2(���rȳ?ZO��H_q�-�X���u"�Z5�	AEy�,���b\A$��6j��yƀy"��8�D�v-�S��y�J�������}�v�]+O�k�R�$,	�V�X�#дf`.��P�]�=�L�ur8�����ɟ����p/Y����;ȹ�d�ZQ��-���!�Z65j&|�B�*��um���g6Gc˽��6��n��_�di��^�d5mnPL>����]-�{N�;E-���W��?ą�����09Z�4�7�.�ì���g�'�����A�e���y7�1�����2�wq�'��у#|��l�wY,��xY4��-Kϼ�]������g���%uGy{�&�uR��)��dE��M �:�35_���8��iY�|��ܪi66ȑݦ���c�b`S�v���nGo8�Ynw���.�5�xb۫K{����@6�a%hxt�|��YK�q��YA��ڻ�<����C[ĺ�}�n* �4�L�Rv��z�Ex��b>���D��GQ�D�620ȱ�J��]}�?���c�zJf-�L4�a��)��	s�)�Sklu�MG�d%b9)��jv5W"y����d����C3%f�whB�ƴ�bA�^5()��9#x]LF�B������J�5ЈXq�G/�v�m��䃻���t�j0��j�7���ۗ�>����!7���_��g�a��%�D4��ǔ_��O��"�h�.���N���3�1���R�d�bmW����1��n�E��qϜD���?�E)���q\��F�	�R�H8�ytB)1��J�R�����hx�G�g���c����&ޚ\��f���$8�O���q����E������C��let�$���	"�1�('t�A���ݛw��>��䃶��g���(.ף�OX�"C�_�����jH�'	�GΖն@���[���QcȄR$繩$\�DH���V&;��+R��[YPj�.~��ɚ���l]%�V=�=�</}c'Ԝ[7	�Jd�EʸQ�,'�Nf�b|����(YN0�jZ!��� ��sJ�,����Ӡ�8�ʝO�C���Q֙�t�g�4�L���)�Fr�E�����]���;ylF`D�9;���S@���$#��� '�1�浩χ%(gѺc�+��׷w��n�?޾�{��^,�9���^�6������$��&��3��e)��*�R�cE�ˁM���7��+'�a����Uf��2	zF��D��|G�Y�b�N����D���E�?�̇Sb�W�ʝ���y�ſ��KzA���4S@V�(Q��}�F~ˎ��Ϡ�����A������W�^�c敞�P�ת�~���v��2�s=nH�1�tg��?�ͳ+{|qi�Zfܲsz�����[XeY�/��!3�z��k�N�ƞ��<�dP<`Lb�s�N�6��y�y)ȍ�
�cTQgw�1��(S�=��J���I��T�n�!�g�!Gbk,Y��6&��A���Z�k�X���p�,�'|6H��N����w?� v���lM���4�!� ��斢}Ƞ:W�f))\M���k�n|����\d���t�}B\���{���5kCc����>�vU��NE%8���I����:����_�����s _�3r��z�	��`�:��gX ��ym�Lm�xIZ�	/��9�#��w��/��4S"�3yB�� �'	\����o^���⹣�r\� x��*�(�`��MH'a�z1���;���������U��f2��`�Զ4/��^�b�G���L��1����ѡ�eFi����h���>�%����v~��L�Xw�p=��{&�'��A �%6?K.�ʍ�f���$��L	�(�U�
Idc@�*p����R��w�d?E[!H�(n?6�!ƥ�҉�'���{�i���)��dۖUS`���?,�9���O���mv��7��Ec��i�M�i-+�&Y�p<8�H�Ѣ�Яxn�;eu��n�o�vwǌ%<�adn4(&������~S3y�%N�]�3��k8jsSv
��x��1nǓ�����(�!���=n=�L���Y�6�JV]7�W�<�O<~�7����#�X`j�sf^X��v�w��#-�Լ���#k�M7nP�F)��-2��%z[pю���Y��o!�E=��Bх����� b��h�L�e���0t!��!:�:�f%���M-�:ny���n�jP�{S�3��@q�����F� ��ʈp���ڃ����s���&����i�	Lǀ��j~?-2!�S뚦F�%v��F)��i��^��#�Y�� t�$R�<p��D�ۚu �ƹ9��o�v���>��G��3��	z G���w/}�� �!`T�f���nr:��+�g�IVs�-6��Y[����2�R[��<L]ɖ�2�,��'�W)aO�u�L��z/yG�w��'�q:����Xs?f��@@���a���2��
3�uQ@�Ae�,�Q���tSK��~�.���rp�z<pN��]=��g�W����ʴ�&�����y��t�-sZ�0ˋԲ)��Z��6Fw��%2�$��M���"�"���{�آ�ѳk7L���G�h
V3\/�e��sr�1�KT���='�ꈳ�y��|��
�:�-�ظN�7�2̥We1(�?��	�R��WE�q66:}���)Z�j�������yH
�(�'� �i"I�6NSG�v���4�gsqs��r�l��U�CF��wM��?7 ��D�Q��$�z �Aꎋ�sE����zc��aep5�C��8I���/�q�y��h���'�:�)���E�g�İ3��4��E%�y+lNsmy���_��y���_v)�,԰ˈ��-_�Hmz�����U/�O�O���|�bD#8I�Z����L�����O���܌l�xl2_�XǾ۲;��খ�����k�]=��
я��yU����g..l=$f۷����������@����:�>c)-	��v�x$�R�*�O�A����f�_/��d��ȎP"���R~�P���x�� :J7��
0Fw��Xl67K�����;��Klf�r�QS���F,�ZY��6I�b�-�����D��an.t�u���H�x�n8f3ѺxCWB�99.VB ��؂�3�q�P� �y)ۜ��F�י��aoID��Z�,����4�S0y^��-v�����&w5sĈ���;�z�a#���X]N���u�3��<^>z��X�;:���n1"��=�^i(c��i�q>�UŨA3�8,��F��9�:p6��ۍs�v�XZ�X���+Q�$[T9O�r6��`��Y��25�[]��p����s"��R����E'�P96�sAr��P~���l�����o�vĵ8���Y`�܍�Eb��	kt�^y��`|Ju��x
�R��R�Uk*���i���]�S��ġ́o\dlKR�dKn'��N�{�e���WmǗ����[������O)X�&�~��M 'K�Ԩ���~a�g�lM��$��r��0$J�x �%�Y�H�-z;F~u��X(eBn;=7dY�C�M]z�e�Ԡ�OeE�e��˫+��	�~&L�Z�� e�fm_������^'n4)� �U�g�U�X�]�� �;a�CL��	�_�j��E�V�#x�|�G.�eS�2k�� p��<	���"�Y`�p)�z��>o����	Ƕ��I�A	��8i;a;_��)̜�(�*�s�/$Y�R~�C2�<�U�V����_�،�%�HJ��X��s��Gk2�yTcx��hs�4"��:kͲ�,���I��4L�l�gGuB=����ڦ�{��w|����S-G/�mS�odv}�4���D�x�:��+�Ts}�!叧P�}��'U �(��k�48��l���$��V��ejI�N��,����s�0�j����)�4-K�(s����2�99}�wT�ɱ)�|E&�ٳ6b�%h(Ss6a���ɢ�G�=bf6�;��J`=�Jc�����|7~~+~��p���7���gU=�7�n���ϷW
t��N��������=}\3�z����iL�-�g7&Y��6���������n��Q`w�a=����	W�'���E �����3X��(-�yTS��K2虙%o/ӡ0=�fk��P�6���s~�}92/�GCGqTF�=�(�l��I8�1{�0i�@ީ�f�����NC�a��N~�U����������tk�ULSVxse
L/6�<k�S`��!��M��<�$�v��l�vh�{(,��B�T�I�94�����U����3c�}��I���s�P���R��Zr���z8�[̗ ��]� �@֭����8וVfd�?�{c�H��`OVΡ)K�P˦�_��n3.X"�We����<�L(	B�C⟦J/O>5v��#�O�Cq�[s�]��,s��|1�C+���O�����4Mad�Y%~�x���w!����֗U%h�ŝ�6��|���;���uA)���!�o8j,Љ8�Z��0�Pm6=�F )�E:�t��U�����|yE��������/�ps���gϞ�_|a���K���y󓬬�yrI�v}V�n~m��ojF�&��l�e�)��G�Q��KL�´�ܐ1"����m��e�oeJ�� ����9���D�e6(|��U#&G[,��݃�7
�߰�2I��G��a�))��9`s�Nta	_
������~AY��H`�����_Mĩn���k�k�/�D�Y����I��ޥh6Es)��+)��`�u�]���-;$����q����6�&ŝNj�С���C�3�2�8Aua��a�ߛO ����0gu�l��Φ~��{� ^��a���-K�R���qgW�>:�{E������/��t�d# N�(�[��##�_>O4��D�P��9�߬>h���^|��V�H����n	/�y����>x�"\$EG��<%� �4��Cb���m��M`>�d����O;�Lٹff��������,Kiit�끘I���t|Pe�1���El�24��k����r����İG��~6� �Q3��_|f�]-(j�&���ɓ'���3{�♽���fh7�_�b������8r6uY?�ӫg4*D�z�ּ�>�7�}Mu��ol7쭬4	������k3�\�yᳮ�:�h��C�h�$l����BʱE���d��Fq,߾}˹���A��S[�(��TGn��HAE	U���C�2�!^��{���?6�����Ĝ�L%1ob4h�̳z#�kY<��!Op��Q�n(���)3$�4j�y�M�C�BR�@.3=lR��#6��A�j�V_��D~&Ec�68W�zn���&�C��z͸�X�1�`��/n�d��8=z�pS�Q|r�����	ds�"�[�d������˟�Ϛ�H�H����@�xF���v^�bY���<�#.B�F�ſM�tsU�k�-�lz���D��*�� ,Jj�\F�g�� ���l���I�a���ɃhLKi~=,���%�4^j���\<���^>{n��/�q1�!ѹv�����w�={�)��N���G{smk:�${���>��S{���Q�vY���v��fP�;z�_^�	�i�f���.�o����k.��AȷG����N"�, �]l����N��>��7�;ن��7)�lr<TMNR��Ѱ[�`2�U<<szH��=)�@Hj��V���'���N�5�$��s�������Om?s ��jYܣ%����d�nZ�q+.�{��G��~��;0Xah����l�ڐ�v]��K�O��{�3m�2s
=g��>ZY���Ʈ;�7f�1ss&O�B��!0d\ ��k�8���|b��nKǀx,w;��݃�-�⇏�XZ�pX�^J��-;l�� ��E����(�37,�ز,đ�a��:�7K��2��8���/r���������x����菶��y�42��:�D�v�i1���=
O���K��W_�W_�Ʈ�����ٛ7�i}=֓�zK�����~�?�[����<޿�Og�^���4._�o~�[��~gO��p��-Agd�׵<yQ����}c������J?9{l����������|�h���ǌ���k�C=6�5�ã��Z�)2}mZ����� Ph&q�����t��i;/ͩ܌���&�ʣ0ǝ�g\�pF��}��^*���������o�c�
j�5�ȗ��5T*��<��g�)��6����ȩ��(Ɠ?����!�#$�9�O� �y��ʕ6w<Z^4�6*Ա[�ȿhbQ��Mt?0���Kؚ0�n�����'����|@L�1���Y�w	9-i\���j�<�Z��py��҇�j;���F2��(�#�u�������."���M�s���ғ������M��=w��|�R<���i-#��#6�r��M�\B<��q,��v���jC�=(�8k��2�$΂J鉊C[��P��g_|������y�.Wޮ�8�����>����_֒t��o~2{_3��~��W��_����/mU��,�.�0E|y~Uˑ�����Lv8�Wg��뗟�W���~��S��r��ښ�&���k;�Y�y����7�d��sW�fwk��}kp�!�d���Nx���Q���0���;�=���˨����p=a���u�%ů�s;q�V���4���6f�l(H^E� ɘLRg���H�5��y@N�E߮��u�4NSi��f�����g��H�#i�a$i{'��,Փ${6~�\����DH\ŉ�1 S���t����Y��� ���_<66�V���i7o����8�m�;��4�*.���r\/Yc��Y�|D�������2���4�7qr�}�A6�n��A��5'�x)#��<�Y�>�,���}z��{W��^Wȯ���l���o쬥9�]��q�������D�osPO^�S�]B�ё�GRѼP��nR��E���,9���?:�S������20�D+�����Zo/jp�w����.jv^�Dկz|m��������?�3�m.���_ٯ?�ܞ�]���X��M����<Y���v���y���f�I���z7�r���[Nu�h$��n�Y�j�]�ff�E���,�GCb����Q���wZK���͝o�gl�܍�Ԣ)5�u��@��yR�|F�y�1�:��߂_��pݤ9AG�%D4�A�F�q&�6J�F6Qr°6[Y�OĭL�AR�F��K>g�m�@19p�FFwON9?}v���󏿜
�^Mi����SK�gJ�'Or#�^�@�-�P�Ohy f��&2��ެA`)Q�x�An�{����+��Sxk�
� ���A��S�)*Sr�ߎ�4�?^RC7��X���<m<hM���^�XgLL3N�m6��z��e?���/"�&e
��q^�Q&99�/Ή���es����Hp3Ԓ��,8d9��x�G--_>������Ok������}�����1=��G5��=���}bO�<�����%���}��}��3{V۩�~��^�\3��PS����vQSK�GWW���{_��qw#���\hXʴ�\��� ���{0d:�G.^�	Na|�`?��iSY6�q�>���b�n��t}�R�Φ�?)CS��`��}=S���<�|a9[_�)��������,��\�d �_C�`=Ff�?���j=�Qd�'��'t�k�9��s��r�h`�����']��@�0��8���9����6�o<~Q�4��F��e��\�}px2���4h٥Y>?2�ef[<���������]�~wٔ�����xh�=Т����k�)vUCӟ����1��J��<8���(�3��#�QJ
*K|���l��<��ڰj� ����a.�:����k+�VM�Ґeʳ��l���Yً����ӧvwoo��ۿ������y����K;����դ2������LnS�b�1�f��ym�}�ʾy���twM[%�`������?��\K��� �,澾<�[	 ������O���JǢS��F3"��Ș�d]s},�J���~�)����u�4���DmA�=Wfy�����u>�/:���<`4����Tfj��
Pr⹎�[ 4<����̝H����[�˓rn��I��N�P�� �4`h���ᚡI���$�Kj�{�%��\|���g���/�7��aL�0�(�f����66�nh��;��&^#^��v �O?�Q�}�U��4�����JX�9^�4���.���o<���L�����>�{?n�f2�L� ��I�ߐL�Я��ÐՅeT�����V^sߛ��1�s��i� ���;JS���|,A]�X"ao���a���`����颊�[�f�ٜ�5�P��F�-�Md��5}S3���������������~S���OH+�����Ћ�����������������Ԓ���l�v��ô�g��������7�?~ϛ�ef�W�<`����R
�5y�A`6�N�KE��`�'����p��"F7h��˕���Ѹ
��?t��1��2�õF��l`�%>_hV��Q�#�k�����q��UB���<W�e��4��IW�pƅg��::Ǭ$��I�p4\�G�<�i����-
�� 	)�Pe�����T�m8;;������?���	nkݵU�
/d,�N��eP����J$�i��[R<�[�����X��K|آc�}���9�E
�SPZN��.�Ω�&�@(�{�U��9W�?��@�i��J��,��~\�.��@[aȁ�{�U��;} ����Tn��_�����[�,�����՝���[����Y�Al�#E�rn��t�����9������ˏ0,v��(��D��6\����!�����]w�o��d��}����}����I�,�4`i�#,s������G;{�31`5l"$�̾f$�bty� �\fy���:�M����0���8��UD�4N5�����1O���ݜ�k�+�]ώ̥6'�uC�F���"c���4W�h]���ZyhO��47������Y�YkjpL�W�.�K�5GXr������u>�����u*� :�d�fn��>���*��$�dq��`���9��VP�	�)J3鵔?>�X1V��_��A����SPN�n�|��� ���r��� �-�W�w�Mid��f\5���gՁ�Z�.�\,���7�%��t�gw`��mN�����\�$��(�e��/� ���	��,�v6�zF������k�vz�����9���G�Wg��
_�"Ge|������z��2��i5Յ����t�����.����)K|`1谁�^p�l4�i��S�������G+7oT�ۮ�V�l�s�Zo�b���}F]��y��2�g�)�&es��Sc�(�zE���f[e����6��t�kD��BB�c�Q���@Yj�;eP�2��Nr�Qe�k��ꛣ&�͔�1T�6qC���F΍���	�e�3W��w��N��;��L�_�g�LJ�B���6g���aN&��?���R��a��=��#}9�!��E$_\t�L�u[�������{�e�\GD�>�(C{�iQ�-�c,�F�}��c򡾱[�܋ں�� ��E)�H�Ś����-�T�K�q� ׿����(�����7��1p9|��l�Rɳ_�Z�s`/��K�9��nr2��������J��41?�����'�r��r� !�c��$T̀�IL��a��|č��͊%+V��.��Ef��4+ |I�H�ԑ3?�Rx�.θ.>�q�F�^qU�ڌbm��j8LN��~,�/-�P�t�P��n)�w���e��]Θ�+C5����S��E�l߇?�jfX�pj��� r�p,���靻Řh52��٣��)$�_��q�`��k*�\�~�m�Q.��S�c[`��÷o׏�n���_dVY?xʬ���N��)|o!�'os�Ʌi�;���s��ٖ���A��(|�k�[Yۻ��/���̙�t~
��Ǵi4E J��ͳ?S 3/�G/�3�&�lP��2�8[�A�ۙ�f�����1biI��Ì�w�E�G�N���H���_��x��F�Q�ܮ�.�q�:����=���QW��\��ʧ�p���7����C?|��k���MN��9w}��(�L�VNǅ[�`��`PɲӃ���I��D$_��s������$4O����a�8: ?�L!����3-�N�ڊ�͔���4�*����&+�'9c�6uN?��[�ײ1�A7P�1��O3J��EuZǸ�g��pɋ�i�1ɘ��I!}r��ٗ�Ϗk��>*��[!��;�m��la��	���������/��~z�3e���UN���O�S���7P8�*EH3�,m�d�����`g��g?�k/�ݥ��ߴ�g`����h�8_h��=v��ٌ�Cy��q\�M�,vn��d:N���"��_�D��?���{�Ŧ���v^b���_��^Q�ĿSPm��V>��D]����,�u����|ˁ���ޞ=N���Ǵ���̩G��y�~g��[;����>q 2�	�$@����Q$�����t�I���D��}�g�zsi�n�T���<J2
=/;�@�GI�>����� ��� �+^r��Ѱ*E�7���8�Ǥv�j~>a���f����?���Z�^^ɢ��o�h��pԌ���2���6~���{�b�(��r��oY���AA��r����1�p�{�36�ɂ�x��9�e�J�����nW{���=��J�;l�^�g׻;q�^��l��4d�>����NR ��'���dK������ Sj���.���.J�e# �H~s������Rf,`�f"���28���3�����!z��>s<��n��c������IS ���1`d&�]�z�4�l���πA���9���`6.��b��:�>�-9����
�Xx�E�����u׽�#m����~����~���x����~���٧���]4����1!��=���k�����ڤ���;��OMF��4�x�{ =c������^6:�(z9�cq��y��%69B?��lps� �D�5���T|S�	���7��\xC�|m��,&��y�LN��k�}��m�I͈֡�Z�����_ՍDλcs,Ä́i`���,��y),,��ْ��:�ͮ����T�~�l�.y>�X�n������k��'�g�v^����̮>��^߼g��nwO�ȃ��oV�IU���2�&����9��M�&�\��Kf10�)�VfH���b��ϖ��i��V�xP�I�������9޲x�ۍ�C�}�P� Ω{�1�</(x�%�ھ��^
r��l��c-߯�B�!D� �8�L�$[i.��|k�e�/a��f��r�m+�Y\v�	��*�R]�w���;{���/���%ʳ�����?������7���6����x`h�k%���G6�o��x��v�\���]]��	�[���r�J`Q�hmQ��z'bzO�-<��S�%�}�#���⚜ʢ���)@~��$Bga��&�"���XB��{Q7����A��\���?�����b�]EнĽ�T�O.Lg����v�As���`�7��Q��=ۦQf�3�p��g�a�#/?�\�,�Fj��%k���<yCe;yrIі�Y�ל[LvF�pOx����!b�Y�zsN� �dn'A f�t}m?�yMũw�ޣX����G����Ο~|N�> tY�N�z�O�!�r�O�\i�,M�O���8�XH�wm.;��#�ˎ�J�����Y�������kE��rctF�(�9,����%�/���W �R��s��3��SDi���ֱ5tm���_�F��I��=�""'�6{��޵�Ke�t�������a���Q�J��4��X=��5H|����u�]~�؞����_|eO�s{{��
��/�ԯ���<����}��[{u����E-9?�7���=�zl���K۾c��T;�� 7�/>�\Z�zc�����]��`]��w�7���v{so��{���En_}��]�xj��VJ�8���+RO8�􈛳�zP�dw�p���t$���"�zR�,�7LHi����Y��E�v����zN7��yd�8����D�6ɘ:���2�o��q�Ê���<���ļQ��x8�[�ݾ��C�W����t�|&�@o9ē�Ș�q�$A;��ʇK�o̪�䘝V�6�u�lhʮ���?���nV���O��Cg�gu���y?�{c���ov{{���L�������nz5x���,��4;���I8���mx��_PZ�w��c����"�.�Z��`���e���D&�M�V��'����Zf��O,�r����bW��Nǽ�}��s�#���7���j��֓��i���:zz�.Zɞj%�
[AGԖ��_�Yo�s46� �Ew4�����~;��V��Er�Wp4��a�]o�SMY�@�xr�Ȯj �|�E���E�y�� @c����ξ}�������[�2�8\��{�9�4�w(ek0�������=�����5S;������~�֎�����?�xd_<{I�ilD�=���������/��Փ˺�jY���^_��>�_m���L�s���-a�96��������L[2��I�a^���#V�� ��S�:6�,p�'AXw��jgӝ�������V�JxrN�S����4V�sϐ`�YN'��d��Y�g�ڊ�O�X���v�u�}�E���8I�jS�T�o��X�1\�xF��M-YߝvT�`�zN`vzB�	� }�r�����=���T���S���˗/����_ܺ��-jl�ٛV�Z��l.	Fv�Ǜ�Xk&��21yf�?�Y���{�F�������b��X����^r�F��_����x:��;��90�[�j�<��s��T��Lh��E�*�g�sT�t,��)N�s�Y#����$m�7�(�u�����%v𜖥<:�a�7"+T��1hQÀ��n��W?�P��z��L���?����k��S���pk�T������^Y��	���ƣm��|��~=(���n���lun;�s�������k�co޼a����W�$F��'��||���=���g'�������kp��+'x{�!�I�u*����$�K^���R�K�h�>�������2=R���mcg5��5p�AfpG_:��g^x�S�ٮ��,�0�����2���	I��y�x�8X�D\ead ��HV�J�A�nZ����X+��t?9�����r����X��E4�2=׎:��v�%�76*���9�M� v5�?�?�H�A��=�C���?O��맪�����O��\��>z�25����IHv����r<C?ͅ�'"�Ĵв�vs�����L02�|>c�E'�g�p��/<f�x� �w�ܰf����o����<1k �)K���H���|<�h���1�%��<��ϋ ��f��!o1�׽�)�E�/���ْnyI�Y7t͋������,����Օ_wQ�~��S���5������������y���?�1{�{����=~�=���|�� �����rc�0���޾�W�Gw�2�z̯_�fy��I���j���n�"<���ܿ����`���ݼy� �Q��;��mfa�j�P7e�����W�.n��s��xTW4��=f}!��������3�&�s,A}9�ן��ک��W$���T�c����}9D#A��J�_5'8wxd��*ɧv�wV���,�hp�7�f�\]e�u�A&f�
�f�v��uq[�_�ogo����u����=";,YkA\TبN���c�a%�����'���a��ʇ��2SX
�'Os��4�� 6Ef��f�C��d���7ϋ@D���ED�yd)���\T�	2��n���Dg�<P�G�X��&e�1{y]ڽ��w�<HM<O'� 3{���Ε�Z�����]�Ls�V�`���ZV�G������kz-���Qn�W���;�zHmJ������?����g�߾��b���=U�޽#�����dgn��"�>�@�2���޽~c?���Y27p� �T�Ⳬ��Ȃ�bt�(��лag?�������~z���I 'K"Z����D ���pm<��ܕ�����O�Mn��ǹn����(��\w�Fֆ�M�D��X7�㬆>#6l�0��˲��y#�#�>�]4":k^E���B�j>�È0��D��� k��tPe!衂Y3�9!,]���٢W�2�|�-8tJ;g:���L�_�09M	$�f�ʪ���ΆU=�^N+�z���vKw|����p w��q���o>��
s���f�byӫS�J �gP�ϰ�b���,�Y��v�1��T�#�K��/�����,4��n`a����=v�8��,P�{��b7��,cX��=ǿyr
o��r�%�)5�*�K-	�s�?:d��r�Mn��x��\-]��Qv��v�
��[���=�$�$G�et*��$<b'�f��������}��'��/[k���������3w�����3�������g�r�ן�p������L���q_3�oT`3��{bm�Z��v>�`�4�T3�׻[�����ﾶۻ��o���Ԕ  ��IDAT{:�+��\�9�}�D�q�[����@��-���\��2(d;�(�Y����b��ۮ2��<|�mFi�o59�h�'�nd�������(�~gA5a� k�46���ҿ��&X�j�o#�ztd]%O��!�} @쿳�ט&�Yۢ(�,��S����0�3�q�Nj�P��fH�c'xxkL��=��9f`�8ֵ�0fql�����GaA�g6<�r�-1jY���+>n���J�J���|�̅��e���"x���u�A`BP��C;Nn�U��8���9��������Ǡ�+�~�MS G�h����8wrwS`&%e:����i�rtn�|D7�ߕA��]��&��ߛ"�:�'~F-!^��g�@��̥w�o6-e�b�8���pm��H<6C��y_m׵�<Ыm�Fê���zo�߳�8�_����X�3�V������n#g�����\da[��#ŠS&x]��o����5�]�s3�ٹp��I�p�����}pvٲ�Ǯ
-Ӂ'�e#�s�I���y�]g	)P���H2��0D���{^��o�U;\\�=xQ�3��w�i|&�?}��=�zj;�IMm=�I�Kil�}b�+�Fc�%Ν5|�/a�!S �Z-?O�N�=�e�e-���M�fc��1����{3�͚�2ϒ��f�(�$:����Ȧ^�� $��4��Q���G��Jk�X���`�������QAF�JSL��n�V�.~� dA�����w�M��^���&S/��BV�c�̒3�s?GnR'���< wy�&P����Hcz;�ó����]|���)�#�Co懚'z.]�T���0�I'�|ɉ�97�%f�&��3 &-�p����>Sx�[d[��ye!�A�����>�뼮�{ˠJ*K�mN����1�7߱�{�F�`F���48���"�fU�I�����r[k��c��Zj�����A"����Ԟ�6��1�f;���O���@��3�׾^��?�`�w��z@�
Ru]��>�δ�42qR[9rБ�׍aE� ��AWx�9�Gg��.�e�\:�QD� ��~q(��Nן��Ts���,�"��˫�Qn8�����ގ5#=��^�C'�ų�v������Q&t\��@�	��S�6���/C[���FrBp]S�A��'ev�oj��O]��L/���~�m�Ѹ?�J�qu��m�ĽH�-g��a�	U%,����A��p�����{��'�=yl���R3<5�4S�������y�9'Ǜ7��q��F���V��돿����JǱ�zqʭ����$�����"w�51���� b�)8	�p�	��L�ewӱ+�<���vXhJ�xH���|�'b�;I>p�D�e�EV��;u��8����bb����6��QB���L���u8N^DdWuA����h���8�nTyq��ûeG���]�6*;?�T�� d��S��V�;4�,'Y�#8��7�r�^`��[;�v_of|^t!�<v��k�����
�q�eu�֟oEK(=&�k�:�[�nj������p�������ѱ�1D�o-���ݶz,c�K����� R_c���^�r�Ck��
�4����{��X��YoD4;j���5 2�;�N7'/F�<zL����]�{��i�T��}]Gh�L��-g��v#�޸?����1�	�����#��>������� ������f/?���������Ξ��������i��suyi���̞��nj�����b�~��`�']o�ݑ���^�i^֬	�	�=�$����=��P��'��̱fpw7�\��x�O����b#;�\%96E�a��dtďww
Z�z��5ڝ����Ҟ������M=ȭn��y�:�q�0ȉԣc���}����
���d�H��;�aZ���.��'s'�ق�����9؝D�P�ݽ�)���v�D�a�4�S�aс�ɛ<ͣ��5�j��fB�Mɧ��4���`�1ℯ�{T3�#>%ŒW��d���QM�d�W!�P�P��u��0	'
V��)����V3����'B����;����ʐ��j���z�s����M������Kj�	���|���z�<�ֿ��L� �b͉�42��M��k�V��'�N��>�7�xe�G���Ȉo�F�Ǒ�ӷ�k+�f���k�/d9�	G���9��9��������n��ynq�������7���[��̍�����.p�zs!�u�.j��!hj��8�Ma�#I-�kP�k���{{�����3:�؀@ƭ˩�r`_���R���3�tN�Y��\1���S���/�t��6��IL��V�\Ё����F��6�Q�78b��������/_|��}������M���r�A�F����~� !y����6�z�϶@���3{��irg����rj�YG{��qM���;�^����PM#��X��:��J!����ʤ~��'Wv������M}���n���7��bm��)��SV�N��x��O�z�����}���l:��Φ�RPA�DXR+B#� �b�\���륹�����d�!���� U�5|�N��b�8ک��;ʱ	d�B�ku������O����FQqG��[9��q�5�0/P���Dϣ+!�T`ţ9�lm�;�̀J
8h��M�����0�=���G{\���9o�c-���K|��Xք�M50M��%-�W��\���j]Iy_o&�D�Φ�cBV�F����� �R3&�}$�3X3?�H�zNj��;���[;���q�fC ���\o.d<��7�Aϳ'O�~�a@� e�-�L�D[�driB;v�Q�r�/<5hC���f�Q�:,��R�&n�+(n�q���n���C��[�x�]��w�0�5���K���yR�[h���8�;�&�5�N�O�僲�ŗ����\Šk|��޼fS���+�z��~�o~W3�������d�~���:ȿ��z6u�U���Wpx����s>}�	��o~z�n4�/dl�j)zV�'����;����z�_���
�����Φ�k��9��3�GJ�a��S-���^��;���Fϩ�E�2��zC���v���f������Z_�Hͱ�j�0�^��QZW*gR
s���y����ҝ��ރ7Xfim���ܦrK����Ж��]=e}>�"�r}*Q#���Gv)��$o1�{x���� l����ko�e���X�ǒp�#ސE�]�w����U%o�y����2�Wu�j�!�/�(//`a�'rh�ۅm���<�������]M��~S��T?�����������u-%k �wi ���_<f���Dݽb�g๯�v�n��f:�]��T3��Pb��ԃy��{ਸ਼�Z��j)�nwGg�u}��~�D	���!�C�U���O�l����m�D^]�R<�����X���
O(��odŞ�;�޾~��n� �K�<��(��8Aj���{��-�BÎ���9��(1��^�L�Vg��K�Ս.���)C�~����$y���o�F���~-u��.9|�������ԑ}��`y}Y3���u\כ�# �ۚQc=b-��^m/�/~��2x��ġ7a\���O�ۛ��MV���O��Z&�#x8���w���H�(`���̾���w S�^7�=�4�Jt����c5p!�����9���P7�}]���o�����z�j�p���}���)6�g�9����<��"�t�T���{p;!��p�g^���f��KAm�)m�Ut@#�,���fzB�$X2�b�(9h�y͞�"���m���T���f$���Ҫx�#�d���{�M	��G7@T6�)>��E�c�����a��D���"x�L��_554�A�M2hQ[����^��컛����{�����גv]��N����^K��>�E�z}]4j@@�G

�F������7%)Z���Qʠ���rcRG ��P� ��c�-3��|`w�v�!�?�rWe1剮�<kЃ�a}�D	�w����qo�:��_]���[�e�u6�\�}9�\�NUWW�I��E��� �K� ��+O�[ �� ��&��@~�	؀� B� �H�\mI�%Z"�쮮:u����5��Ƙk�jKNS�:2�=���u��k�˜c��7�O���R����*��'(��ҵd;I�O4��wf��ԠNi�#�i5_�[dȍ���<gxqh�g�>����z:�wr������_�7Vm��i^V�_H����J�g9o��,�
6��x^�MK�����0�xZ-��R��b���F��*sO�N9Wo.�8��F���#�ã"�gr�i^�ӧO���c������/����F�~t���=v��#w49f���\��ժ!�#�\C��Px��+����:��ј.=�r+�7�l��b�C�z�ܓ#V��ZtN��
�(ͩ�3�N��HگtU&"�]���n�FȌO�[#%Qk���Y�<>[�ϒՀحĴ
v�x��q�O�w�) 5�����;j*d�$�t�Ho������ܓU��آ7�y�bŇ`8*$�����p��o,�|fm[���ܖ����,�9�#	;��v���_\�R��T������|����%��X�ky�	l�+ԣ�mʞ*�<!��Ut�%�9>`��K1��a�9&����<12SٱW��,�zkY�h�O�Ȱ��s(��xJh��Q������(m���*7��,��]c�y.��Ն��`�1����G�[�y�ڞ���[V3&փx���|N�s�V�������)C.Xf�u���m��ܭ1�����22׼��pc���*�P���vc8���ӭ 8m�)�:�%,2��ps���ວ�5!?}J�uw7uc��p��bLz)`�~�ï�P�h��`��h��)�#p;�q?z����O,�c�2���ZO���q����F�����Be#ψ@�d1�ݭlXhtG�d�Q�;8
6h�bJ$UHׯ:3���k��L�4�C�-�ׁ^��qv�����-61�7����{{��f������,�E�)K�F�I�È��֔��?j�-PjG�N	<�Ukg!�A������H���)Ȩ7��ǲ���q|q������+��C㖢���p;õŶ(�����8�[���f�Q�pS61���3		+�o�5	a�97,F�P�_�v���4R{bB>�P�Bb>�b��7�F�����t:��*�x�d�K���V)^<�SH�(�!0����p�آ�-Ž�ʀ�6�n�s�)X���&�ð���)Ƒx��+O���
h!+g��s���SڿQ��jӺ����Z�����jv{���j@��W�e�;V�K%�Hݖӌ��y�?�|��o��������D����*�C]�}�0j��w-��#����]\]1��8��5J�2@!d. !$��L6����^Q*s���˅�uBQ(��G�X��}�.��C�sΨ���Y��j��Ĝ�.���������rZ��^!#�e��ԩ���g��k��mdW�?�?y7����rן�b`�؏!c���uF��5��KR�Fx:�3�sg�Ʊy^���1��ab����A?鶉|��lVՌ� e�p40m�a;F�x�u��@ZS�R�K˰,@�C����,�^�zJu�(w�!,ù`� �C�-y*����
�]��!.X*�	��u}��y	E�b�ɤ�u�x $7�=�j��}l�ǙxMHR��&Ӥ�a���y���]Є8(�����x��)�<��;-�`2��)���
�k`��dw�@*Bp[���u��p�k�F�*#�� �)0p�E������2ŴZi�����*0��,�
�~ʊ�K�
�J���n�Ua0k�/��J�/����#2�r$��<,n,֖�yV�̴	0�"�}$%(+R@�SN�f`�A^����+�3�@�80V���;���kߧN����yt���{_����������Tn�6��&����8�z\IΞx�Ԕ��E�=�~x�ȋ��p�����ڑ�G�8���d��\Z R�(ęqõPu>���+uF�չ���xeyf�d䂷]ߜ �T�a�AHD(Zkh���`Ɨ��"C�&ޅ	�!���WB��,*��1*\�ڣấ;��q�^c7��yr��#F47ԯ��Gī��c��Ҝ�d��*\����oMގR}-�Q�
�X�?5�Ͷ��@��(�BM\�&�?�5��CZ�7AoL>r,ǜ#TAn
�a�]�2���"�X����]]]�Ջ��D�1��K8�b�p��j��HK�b�V0)�l*�Dg���B�%�D�V*!�����F�B~��=�22�Eʊdkx>��:	O��r�-��P�W.2m�Au.F��6�r߱9 ?vtr�a��ً�8��z���m䂄o�\��(@3���(f������):8<C��)�%rg���FTy8��S)�Gۈ�Na�x��gh�P����l2 4���4i���4�p������T��b�'jw����i�QC���g/�k6��BBTGxϓ�Cw2<p_;��r� ���̠k!s���2(T�%e��Us���'t-�=��a��D�<Jv"H� d��(2�N=(����z�U��N�����W*7�E������H9J�l*-D���Zl��"}G97y$�����P�E�(��io���צ묈@��q��yCE <@	���;=y잝>!��#�=\�ܹWw�n-�/}N��ñ���S�lr��R�n�V�Vy���������2�z�����w���BT�|�lr�*]�����+�����X�0��xS�g�z�NF��"�e� `��b0 �:�\^�t��T]H�W��`�V͟ X�I�.Q�Oܩ\�q6�=D~gLsEZ����9}�085�0`�@N���F��H��>΅���Z	������=z������ƽ�z���$�pDm�¦Y*�"ճ���%Q��9�Q�����b�@|��
P8�����Qb��Sk	k�kbQ6=6�C��2�^[��&��K�y��"���ޕ�sE�/1~�4V��@i�Kc_i��\k�G3��Ad��h�5�n��<�h@G z���29>&�v��.^�܁�Dm)!��+ِ�S�L>|8����n3�+VN<�,l���f�ٝ�u`s>�+*�e��`TF5�_��YC nF���/�EV��!O����F����TDdi�y���jm�^���(&�W�Ż1n�B�P�d���7�������5XH��5�iQ���"��P�e�?����=s_}��v>8v��k7XW�j='6r��C�dt�"���G���<��cj6A)�����4&��f�~Փɡ;#�����nO����0}&^�d>!Ɍ^���'��~�=�s���m$�C��g��&�O>�������kF�I%����X���!�Ä^CN%{�=�G.��,�	���-�0H��t1�-��~G�ia�L���4
���w��8.�$P�B�&*N�P#y9�	P�����l=R!P?cuh��<S wD.LW�xy�����Wǉ,flH#,T��G5q���6��!�ɢ�*��i]dakLo�]d��^� �k���#Qy9�t���t�AG��3�(���"�p%#Lu�Cϔ���N�8P�+�c<۱l��a�c BɗCn*CTy�K���O��[3�v_#�&���~$�W��~]��345(�q�����:��[�d�����J0��SꢠQ�^�9b�&��U�H�hϵFw�oST�CGt�6�5ۑ���Qu��n8�	n�zA
�l�>������ФǱ����G�'?J�Q �S��N/2��ad�D�,(�>��K���X=�N�$���`�N�w �>�w��� �P\n@FĜb���!7�Q�0;�_�Z����4�C���{t<t��_z�C7�V�$�s���ʹ�����q`;�F�+�}M��\�(������.�kư���n��?���@{��A��Za	eӳ���
�V� ��*^L9[����ъ�^�z@)&8�<�!)�3z�!_C�-h�L:,��r�R�������aZ���7zD�>wZ�o���p�	�]%�[�v ���sy/���������r=w�{�ђU��H���HQ�B�*XOn41畁KN�s$��BD_'s=��$*}�l4��%*����gggntp��� ��$T��&��r��䆛��C����IP����ͽ\�rN\�)�bE	T��VF��øW𴀇{��=^6_��E���`��1� ��zْ�y�L���x��!����1G�<�M����̓��j���)�:Q��A��Y�v�k���c�=�9b�*QfcJ%aM����dS^O��P��d��ݏ?p.�Ç�wi�v��,�g�2�۶$�x!���"#WȂ�����}���10����VƂ@��`x�GC���̽��t���]��]y;���
�{:cs�Px���4�Gm���zEQ�W/_���̝H����S���_w>/��? �L@�|���B�[`$F�ā��h`?M�P��t�x>X�`�H��#0Y�j,�W=y�U�U����-�d������ڡ��x���jY�G*�N&$�!�	5�d�j[�a�a?�4�a�^�e2�3Y''G���p���J�,�HN����Yq�~F����;:;uA��������j�]<`��V�(��I�t�~]���C�da���'��i����Ʃ�z��:<<p�����ch��-��#7�0^��,rL�Ūg� �#(�::؂��f��1�nke�%[J�e-:�6�#��rw|z➼�T�Ł �3D�ڐ^��������:���fc�
jm`խmӖ�娆�x�%��z����t�U�^Ο�|��p���"�lgSzq�����Zx��>�fU��E���IC���C*�zT�n��!F����c� z��>�\�(p���jg�(<0��� t=�^�#ò&��*�.$�7������Vϟ'���l}Kn=Z�O1^^Aƅ�5��VS+&腰��	�	�ؓ��}��3�	E�&���	M*'�������yK)��x�7�\ hFN
���VN4/S�7�����K�e�pW�{z$0�>r>}�=���S���%<�2���D������^^Y��(2t�(�Ra`FrK+�� ����gt�u�B+�|�X�ͳ����Um�F����-��KO&�蝆
|Hr\�]�zG�X+-�9�g;1�i��Q�H&�x8Rqcm��}�@����D�#$��V���bHL���-�ۓ'O��~�Ξ��5e���ҽ���T �ٮ�@H�/����'	����&�I�u(=v��ɁQW�0���`������X	��4�x�f�u��V�: �dգ�,�v���IOt��a,�N�ʦ3��O�����؝����=)�dC�9ӭek6[��|��d�*c��ԑ�=�_��g����|���Pƒ����|��)L��l��x�����SLݪg�9�6CO;dک����&&ƻ����+dޏ�AE��] �[����ab�2��Lq���Y��."�a7��R�R����o�����t_ʰqݸ�a���[wc��O�P7��_�P��C��b��F��ЍT��D&�������ռ7>uc�ײ��J��i�Xn�!a��cW�u/�����?u׋)�*���3:�HP�P+��z�^JH��_|���q/��u�@<��=��}���{�O��2�VwS�`��n9�c==>3l\'�ͽ��d@9h���W≡H1[��0������}�+_��3N5�.�!����F�Ў�g����ݠp^^9�0�)rO�gs�0Ia�p�3�R��AC41Q�K �2R��MDE�pT������B&3�һ�{zl��'O�#�珤1&ށ�g�	��QX�%�<���C�vNO�zc��ěш!u�,���V>(�ȎN��o:�� �Jwz�4Jˍ;9��(E&̏���0S��
��ш�/hY���v�3,TEk# ��:e|ּ����-p��D[�x���Z�=��L���L��^��7�fSI``ۈ3D�}c�߱\?�r�iwx�PM��^!)/�֭��F(�������)ӵ<&�iY�:�7��j��,� z"�Y[�����8	<9-�;k�^h���B�N�4�j(�4}��ËN�yi8�ƺ��h��~R�Up���G�`ݍe�M��J��49z��7�[���c��ol��F2t@2C�\%|9�)U��^&ӱH=̄!���켲szx6	�}��9�h�Ah(�_��I���({#�9=>q�b�@?��t��ҽ��g���e�==gy�p0v���T��Lރ	}�������wk�Hj�'b Eb`d�Ioz#�Bd�,[�bY��G�Ne8�n�
�,ؼM"����k� A�mU�ؼ12�`p�'M,'����O� ��ʇ�<z
)!��UٴJֹ�W�xO�P�>:wK	1c�U5+�^���g��Ξu%&�ݖ�`(����������RBC���h	hw`�_���5���x1Ђ�Z֖��IR[(pS����S��.�B�3��oYŋ9���@�A��\H8<�T� �F���DKU�ЌǠfz�g�� ����'�z9�]�g<�s�'5C�������I8B�9�Yl�b��F>��Ǟ�C0t�_�v���
C�����1?�~�e:(�����1�՘V ��6���9}�^	�Y��� C�ԅ|Ϛd�����s�a+Αs�{�JG�����1s�����&��j/mzy~���~6�6X%^�yI~�:܇7�c��o���K���Y��)�c�jV����P�i��0��
�C'���QA�(!T!aM������%LIĽ��Q���|����ӫdRV1��������-�7��Zj�6�9�>��Г�;�\�Z��"�\0@e��R^��G�5�Tڴ\)�sϯk=�rM���\W�RИ�W\'���k5<�RC��8puX3���^�
���_7�Ұ����F��������he��p�Ԝ6<�Z�r6��c���t�$�?���wqqAl"&*{nb�J�k"��,�t�p��������������1��y ^�Ce��%�Z��6�mIC�`P�8U�+z����[c?�7h�SF��#0Ի^���TW��Aߪ�:Dr�MK�t"�e�7��j.�؎o'#������KH!�Z��Za9r\��ԬX�{�?٨HוAY��b�L�o��_.$
��3��o����eB�����o$D=�,�d�`j0#�L#�B�sL$�J��&}�<��Ǐ��i̦��]\�t\��ߛ�e_p�����D`̸�[q^=��:9C�FL�ຣG�1*��X���Z\����k��sM�"M��o߸U�\�ktbA��g8���#j�_��7�E��)�ෟ�BZ���t�̠M�<���YMT*~��^kw��F1т��+��"o�S�[`uBg4�ѳ�`�@s�xޘdg��gl���/nH���M�S���
T G�d���f=%�[����F��"�I��l{�Z�+�m�v[,qKpsGHL���F7L\z��!�WI|��J�r��<P�(h�BC8	0�Ĕ��կ.��]H��$>
�=�𘔘�vf���h���*�8'x� ���8q�j��_�R'a-�-�>�Vv�IdP57}$�yV4�c3Z.�U��P�c1i�q�tmU��a�>x�)'��V.?���g��<[|OS�ݰ�p(�<Z�ؾ���A���gb�h�Z����h)���T?�`�UZ��>ov?�ڃ�1���Y�{����B-����H�t\�\.���C��\��lg����;��3E�� ̽k��к��3���@�y�r�/�GT˗�kD������)vz(Y��c`���`"ψ�!��9D6��+����܆�*����=3;� ���j�wi���Hۖ"p��r��#�M�pc�`���ؼK7�H�v�����t����]O��	�Uf<�G�5�3X2y�0n(@ �7z>Ф.�1#ʹ�1�B����Q�ǁ���$��Ujs�L/�oϜ
����@��U�H'TCd;�T}�@��&dd���pF���&4d��)�D���;'�s����e0�^	
p�N��݉glx8&����H/�����a�.&|[GA���H�V�,��5,�A>d���o��hi�Z�P���m`!c�Ad�E�yT���h6=w�WW�����uƬѼA���.h�=�x�����BK�S@�o7����E�8�$4��Pq�F{��G���ح���1|E�61k���E<dc�s�2�\k���{*�zT;��;���qw]|���M7+'A�9�����x����[�ŝ��W4�h�|
��[w��%I���N�bz�b��wl[C��g�Z�F��1Mر���OgJ`�D ��Q;����Z����(�jR�N�'5��&���Bǂ�YL��w�~�b�6$�1g�v�%m�-�x�p��D��Sc�x�E�&ǃ�F����sQtl�r�f�A���cX"�7���0Y��~=;MS�����שo)l��&�t�F�,wc��ap|K,�J� �5C�V>�IRȤjY���g!`�0��Q�S�ēE�c���}���	��*+�פq�%����7O��5���*O���k&������k����Jt}۰�O����s1���oi^O�e��Ϟ-�#
�y�.��}L��	��I5$�B�&��7��kL�!Pm�U�ơ�Jwh%�g�p#���<=>$������r��bn�P�Ԙu��ځl�����$��c��y��#���xS�jƫs�h�k��a���=�g���b(=�_d��9����M9e~��(3f4_~$�'<�/��uIOo��s��P῿v�@�j$4���X��f�p��#X���Z�k���q�Z���r�.>��ymlP�De�P����Ѕ���&�1�=��긮���45+H�`}Aov"��D�!�@׳�ҫ�#��\<X�%:� �>��y_9�S[��vAm�߶q� �L�������C·~��6�A\4j;ƍkfܺ�A�T	ʜ�+e��Bw	12��V�V0ꑄ8L�w�����^�c$�w���S}r^�\�ƾi�G����4� F�)���J:���H<		�d� �O�%	���dr��ǿ����  *pf�5�kQ l�k1�k0�&S=�tp�9q�b̳�t5�U'*!���!*����b�n���ߐm[��ᭊ�
%23��� ����g�����`0bEl�0E�*?��O$\(ငs�p�5�!'ј��#|A&2x��뇧X�%VM#<�ƱSwP�>
l�(�L�'��c�X�)�g��������� ���6�N��C��C�����}T�f��� ��Y$V��:�{�ț���k��>�s~~N�m(�4�\�]�����2Wb����;��У�R�s���E)sJ"��B;p�r�n�nXd!~<۸��!���[+Q@*�>'��#u��S7}%^��k~��j��ǳ��+���'�	�w%�=)���à�0dd(����c<��
l�s����k�����p���lHz��q�����
(���#.�o��wҡ�lwۭ�o��E��L�vp;qrj�h�m@Ψ�Y��W^5��/aE*�yx�?~�)���M�&�D8?;g%	�*YW���U�~�5�%&B7p��r������=W
ptX(��$`�!d���~�'���T`A�xvp���r�2�S�e?l�|g��(H!aG��@�����p�?ǰ٧��wʎ��o����&d��)��	�5f ��3�a}�4,� �DER|��ڈYGxQ̍��Qiw	rF'�>;잞=f���z.�>��*�����+�5�1ȁ6A�z��ɺ:�'�f 
l����FJ�`�|ϗ�1�w�1�	C������b@N��ɱ�����\���D�{N�2�,9 ��3U����V��.Q�5o��NN��'�2���ўEqRC���y<РGg'�=�<{�g�|6��34E������"�A�V̈�9����c߮�+��;(��w(�b��pmLCFaceN�AF!��d+C���@��?b1���o�W�D:�t@R�)��;��Ӊ�������䇄�]c,!	[ɕ����Ȳ�������G(١��C=�"��l^�'g�@� ��>��[>�� ��}R�޾qk�M�$Q�n�<u��gV��$*��{�M%��D263ËB�0m��;**��N%��Z�ܫՔ�PLPٙ���b�5wc/�ƭQ:�����Y�9�����Ų�"��ۂw�閌�_���Q��IV\P!����X>��԰��!;R6��C�x��P-�G!s�a��8<&EJF��y��V����A�]�� 9�@�}Y0K٩���h"�!�L\W���6��-�h��F�i$�<��Ew��ȽE�ę��X�r~'G����M�ʦm���v=���6%�NŘƊz�C�CFy?�i�5+���84x|A=Mxe��Oݓ�S*�#�I���D��:o�W�=w���{yy���P����9��zLSxN��gܠ)�Z����Q��<�LÚ�U��@վ�<%�)�����7���4V��>}���o�?��'�5�;�6pm,X�;i����팻.��f6��5�b�
����k���k��4ݶ�re�T7��(�`8�q�}�yP�n�p@H�v2ə#˜IKғvD�V�kO2R5=.�oC}� 2�-[�$�#TO���b4�	��o]�!OqDʧT)�M�B����,�	+�啦�I�Ǫ��7WaA)��RLu���)�"���3��R1��&�,l�������J;�p�a2��m��ޛ߶k$���"���p��>5%�d�iddP߿�Pm*x�2hU ���F�;�X=��YΗ	��V�h��� \@� 	�à��<�MV�G�.�v�	�c�3*�Bi���xϊ�Ōy��f��!?$;4r[��&��uL�G�C+�n��
Ԑ�
Q��00-c��:5:��%ｧW�N�Ǡ��,�
�䪹Pm�,$�F|TA1.��:~�/�R����
׳�V�R;4'��X�S�/z�VG/^����NO����Z�~A�VV��X �M�>x�=:�q�������g�tD����a�u�&t�SO�a^�e�� 5����d C����RO�К�����lϋ}�!�b�k��^���ZY�Y�h����94�;��[�c�|U�Y�Pl� h�"�������$nEnӫk�o�uԳm5����k3�$��]��3m�Y���M� +M�J_�V�P%G
|F(���z�X~���q�φ�_���3��#q��s�$O�TV�r�S���ᤐ+��8 �݊ Uc�8�	$��kǕ���(�?�FN
7�2��m3Y�����cVm:w�9T��]Tqǣ��*� >2O�һ�`��U9: Vrp��kG9A�]���F�\9���dҶ�ވg�m���O�]A��'�w�Oܑ��:j@�0�)J#�r�>�y�SM���^j�>�
[��5:��S��,bfhfƽs����*`	զb��ޱ,x�n�Yb��hyE�%w�d�������'�<86L�R��,dTIs��)LdS*&����"I��R�cP?A���^��mо��@J�3#s� O�g��bˆÄF2���Z�G����Y���0H8K̟x�E�zom^
J�~D�ƾ"JRR�0���Gޤ�Mo)ϧ���3�������K��A+�RbOg}�lM�(�<���#7�
�E�p߀�k��
�n0��f.�r�+/L�b���R�P��}1$TEi4S1n���KdN�BK2M�c�����g���l7K�2��J-�ҕ��-��!!	��u��:��g��Vs��x��!���C����A�6H�I�"r� 2�5�٪�&�U��u�&^��������*jF��xR� 7����H��u�Z�
!�m�=j�� �t���=�^J��1��a @5s)u�b��B#�2 1ޏi��*]%�4њ���0�)�4�ct�m�c�'�mtl�c۶m۶m�v:��������Y�V��W��n}rX�=u�Z$�΁��-�s=c7��"}(D���'�Ή����M�z�!�y������'[i殻{i���{B0^l׈r�&�F�6��\S�Nh�T)j�F�`�(-���ʉ��� |w�Y�X6�r������c:y�uI$��1mF����y'R�e*��l��A���T��Jf!���
�>vw%Փ�� �Jw��gbFX��Kt�.i�0���2H`���2N>�z��dWq� �D�U�-�*�A͕���ç�`�8�Kڟh����6x#(�e��ty��_ڰݞwR	��}!f)�C$ĳP󗵾_V��x��PrZ�7Zp�б9������n��M|����u6�`�`�!�����ɇ/獢��WE�����<���m���Po���7�cuj���Le`�D������-���dV�d�'���tzΑiZG��`���>[�7�Io��5��c^��/���B�f,Z4,���o,�.,�C�7��`�n��aI�g���1є�jG�d��O��C��5P�"kJ�1����9��@�Z�����@��w��h����C��#��6?B��p�
�5C��}\Ļi ��:�# ���h-z҅'�Sn����28�;���	�k��~h���� �N�<�KY�r��}V;-EO�N@�؈BtsͲx��r���M��2�;g=>b4�FL|�z�_���5��� �^���x#��3b�#4|01#��;7w����m*W߉���U�Zb:�P�NJ���X���O�^Pi{RB�W^`")����3�|�vQ��y�/Hj���K��+��-�E��)x074�
�;�mbX�G���1�x�%	��4����r/�}:�����V<�/�ll�a��R*�Qr��WH�i���E�(&�0�������7�ӄ�Q�u�v�q8;��X������2���Y�㑣z�||��5��u\�#'���|^����<Q\���N+��F�l�m\�{���X��)h�(񖏏M���Fn�����Se�&���(����M��I=d�Dxy�	�@޿]5w��ڐi�U<';	`�<G*@m}<��)1��\��gD���GǛ�vr'7ڭ��ʤ�����G��v+m�zī=x�1u:����,I�#L��b2�C�Ea��EgӑuU�y��*'�H5�aL�3�6�u�;��{^����"o�Rw2u�����H��.ĸ�ѹ���B:���C��S���X�0� S���h��o�� ��nd�� �&4��"�spB��W<m �W���?���"�������s�<H:�\c0������)x.����a�[�jv�J7<�e������b�vť�E�t��U궥��u-=-j����~O�]L| @��鷤!�
��XYp�X�����"{燴-� �!����Z�"��IAYW.�O�n������]���}���4���M�>�t�~͑$#���bg�$�F������!V���~d�s$��3�.��8h�;X,n�'��w!炕O%��ZHK��G��&�4¼~f��`�}?խ�c��*_����V��y6���-S�Nť_��e�]%�M_ԃ�4�Y�*e��|�Y���g��{���0q�Kˍ����3O�~{0sz��%�������M�5x2f����s���Ef ���b�l5l��������k$��tg�&1(_�J�?F�t����'Ý��V�/w��e�>�h�_����PD7�A27}X(�����jhPU���!�O9P�Z��*sD�r\[��NfR��2O��G-�}���aw/��I�A�Bp��
'���)�xMѯ��������z��&Y��$�nN�ļ|4@�G'��CAB���o"�Z�
�nL���}��E^�$�v�|�l���6�����ÜTǜ�ţ��!״�]=�>W��I�m������j88BG���o�x��[�L�-6�Z8�1���tb=R2x��/Sn/D�7\�|ŭ;c�A
�9\9�*��<���$'`�*��$��E��m�M@|o�lݽ/������9$y#9�ڪ���#x�rZ��:Uu� ��]�۝������D/�����8����L�qF=m@�A���2)ј��Du/n���L�zq�k���&)�l�H�#���b�t���ֳ��"�e��j���u�fe9��5�-v���o����f�b�1��X�j�>�Te��1}Ϫ)�T��K��A�&�]ļRD�SE�����O�l�\Έ|�Ouoq�`@�gޯ�_I�#l�4Z�W�%�O4P�Y�����OOM��nD�D''&'���/s�J����eq�Le�ڝe(�T�v*U{D&hm�=*��Br���85�1��B۲����@�n�����x%Uz�q��G�Ke=x�*��LYLV|)���W%���Fl^14�1Z+� G�� �u���H"���a��Z��(}c�o����#�I�S7ȓ�(��q�ܹ��Fz�x��>�P;d�gm��t�M5�q�@Ցv�ܓ+�!�]HF����v��P#|�]&��D$Vw0iUT��P��6���Є�@��)<0Q|BZ���y��*��PQ�"�9���c�������em������%��'!Cأ-c�8B�`L{'�v��"'�1+�/����`�k�(1)z !9��F�q�R��l�;RKA�7J�6оjc[#a>>^�h��b���j$���~���<}�Eu���+��1�TRA�y��V��r,&�g2-U��],N���j��K���g:�q�;��Ȫ�����Lx6"�G�T��ԛ���%� ������Jwh"leeR~�sg��tm�5h�Y�k��#a��_|��H(�P�ʏ�j�@kXܹ���
s('��~@A�K����V��V����^�����XIH����IR^8�{���k(��a����@ͺ8$t����q)�{�l�b'������yԐq�&�G��.�A�F7�!��C���,�l�":��BR�5�Qx�|q��`�1�0����+�jA	1�#O�s���G�����;����#�d:gX���J� F�}���1)�眊�?n��*����UxM#�ۢ���ፑ ����e�%@�//Jn.���]���I�?�����MW�@!`?��%qQ�����]|:[����}�}�a�3�v������m����XW �OAr19B��#o��a��9�u�G�:;J�j�ي�����!V�S�Cc�*��W�)�X�zf���0�Ub��t�uۮ�.#�̐|��Ky�+�˨gI�'Bw����&d���+�wQ��u� R.5~�6_9��Mz�{$�&�#;�Uj������J�~y�@��� ox�Q"���ۼ��@;� ,xL/#�E<Y��e�Ĉ��o�Ӷb	�R_�0��i�Г�X�%dP��k���Z��O��c�6H���׈���г�'4E��Rd&�u�8��!-���)��D��`��`ZTq>8�d��B Iy��$�Ǆ�U#���wO��!�MI��\rE<��c�� b���� ��Ȍ`?zF"��5��%ܜ��!b�N�#`_zq�DF�Y��b����0�雋��y{tO�z��lȈ�a��|��-���t�k��={�y�}�俍�6Uc�4�\^�e0K1[s��L���#
��<�	[�!S0B�2S���CZAa����'�>��m����I��I�y�'Y�E��v��v��o5P>�(6S+��\��qYZh�5�U�{�2;�ŹI���,[�*#�Y^Q�&,I���E����"���;~��������h��-��F?4Z�z57��4*�`�k�0'�	���=+^�'Ƙ(�.#�ã�#��
=��t�݁c����,�ϑ<C��K��7?�
�r�PnҼ��wZ�Q ��iӬ��w������7��pbe͸��V���T%&�0F�����8WZ�8��Z���'#b����Bq��}�2WEp��݀�{�B�Q�x%_�p��P;�In6l)���Ҙ�i~HwS"Qm�_�ge�x�q�O0�5�T�M�@�3e89�8e�����?�Y5V�����0�'���	�����!;���:������@�����*��#n��R���>`
2x��	��E�S_��l�"̚c�' �oW<I��C� ɀ��t}PH�X,α��Q�Q���lMa"�!�l9>O`�p��F����v���D|# �������K1�z��tܽ^e� j$�Mv$%Q�7"�Z���P���+ .>�R�o�V�4މ~A3Z�x����vJ+D�Լ�����
�!���AQ&�]�`^���@�7���z�a�O}#��-4��>�k6v!(���Ч�R;y`�-Lt��m�_P���䰗�?L�@��U��v���X��)d�p�\���ӄJΉ4{n���J%��U��t77+,oPɶ>WrG2.J���l��$[;��W���U���=q�R��_��Aoȩ)�r��~��{�l�{�Xc�c�IS���!�� �5ґ�~bz�q� �����cDƁ�,`��{�
�@����U�0]u>Z���N��B?���,|Y���W�|[��k4> ���̘4�/��G\�<`Z�9P(�<��V����E����ϓ���U��&# ���ZLAw/D��Eض�G�B˧F,�|C����"��;šR�i��e*�(�"G�=����o��
I2�k ݎ'Y���aLm�����.@/묩�5�V��SXh:�����&�&Zê�*�X�����b�(X�W�$e;�����U�\��dEI$(ߌ�����q*J�R�I���/�Z���۠�Rk����mЩ��d�T��۔NC!,8fQ��/0��kJBh��"����z���fi���'�[,�^�?-ީG{�*��<ҷq��G�����2T�9¨�X���4�*��T9��x֡�fY3x���� 5����e�Xɫ��8������v�U�Br��PD�~	>κ�k�����/yjv\�����9����z��b����r�|�������6v��GڌFY��hdT*?�*�(�XX���+�;��;��&��Br%���l�l��JO����� F����X��R§�A»�����8������x�Lw����;�4X�Ҟ9��\B�w%n?�AE-T�^G�?���h;�nA
��_�.��F��,IrfY��؅e:l������������T ����mĸ�pxnu���ߺh�Z���Ǫ��ǫ�v�xs��UËM����3��7%�
��
�P�����!�6ȔR�c���%�.å��^�i��
�T��0A��m%�*d�|f�0�^��D�7�d&{Je�Rv�W��� �X���]ү��+��kΉ>X���ս�?�/K����'��Y#�5�B֐���ks�l����}�s��gw��9�v�e�)H�f!��Y�T�D�E�Pa2�ƫf�뱜�t���;}���Z$�q����3}�iw�(C�2]��<+?�'�;���h�cT0���l��A��IK���/���D�]�pFI�y7��i��ܸ��H;��D�(!��)���ё�!�����:�Ĥ��EY,�M
n]N��q8#�3_*��%2zPH��.�lb�N^0P���@�Q"�T]�N3��+j�G�����t�p��&����e�&�ٞ.�)�wZΌ��M�LC�h��a�7��>W����h�C;�C6B\+���MpG�.5�v���SЋ���n��V�n�GE�.�rl"Wb�|�����&?9צ�.0g	4�&�q��������i|�!�dY�b��4;�	�n�x�(Ŧw�����b��f^�yy��}�d����6�,�RJ�O����R��|%9y⥵ZOs.�D�X��`POH�W.�x
I��N6�6�+\f�	6ot�jY�����!��Ӹ��tX@;��W;K�¥�Y{��Y9h�k�[�u��j۴��a[VW�m���n�x��D'q7�)_���ǋ�]��bp|���=ޑ�^�hve��#���Bh�O���W	�1�}��|0��"�/�9}L���z�.�E��N���4"N2ľ���QT�<t��{���l*��K@��1�-(���i2���o��x��<;���Pߑ�a�'�)ޤ�t����T��Ԙ��_�=���a�QL���8����f�BB(�ݕ�P�Z�v���#�	q��{��-B	�5Wg��ĳX��c�beR�h	�]�\�t˩�����5!%�7�V*4t��&�� ��&�p���<ZwRo_�r{�]aM:9�i�0�j+��q�k '�-3B�/{��5g��(U�y	�؂�?�bA�zߛP0��6�QE����[��g*'d�D1�~6iN�W�@Kej�J��,��H���P0G-���,����U������6Ht |�AnaX�HTf���@��?WOZ� ���]߷͟G��[18�W��G>$P���|J������*nt`�opv�W�6�e�9U��SJ�W	�xĬ�Vs�Z���ri��e4��զ�9[
��b)会�����+Җ�ӿT"f�~�fKl�͌A�g�R	��J��H�d��՛Lr��n�=��(�G�8����+7���f��a��A�`Yk�-� _��R������~蠴��1���0�11�2�]c-�q�o�ȫ��g\2��j]�����d��7q�$Г~���]_� ��Hs���/a��̾nu�2H���:�[z�bU�rne��
6��`��I���/bU3�R�������;�#���l�i�G�&���b�
o�i�i�� HQ9O���b���$Y��{9�td|� BH]�u��V*��J�4F]匧zE�%5崛=,Ⱦ�a�$�����G�*[n���f�~L9��&����m���F�H���v�}�xr��AΤr�_�`���b�����]���g��&7�k|��b���2�j>�cpFj���.F�N���7�*�dzSݮ3��WX�	^� ����j|�h��$�W���l^���|v��;�[���(.�[�I@��S&U�D�.�ai�C��3�CY����y�%� �y��eM��E��Uu�~�;ب9LWe���M�3�; �S���mY�������s|��]m�RM�<]DZH-R"}�rP�l1�͉�` ��
��{�ciE���P�����wq�η����~�F�G�$qTԾ��[�2˳Ɛԩ19���=�++-��̳Ty�lo���
�!S榵-��I�F�<� [���%f��"R;�rXQS��M��$���^4�$:�>pE`&�%�����N��4�l�.-�[&�7Zf���'�b�%���D]�X��s�aPٳ�����b�@XaTk�>Є��l�� 1&�bZ]��7Vܨ(�7;b4O}?}U��]WH.M�>���`̿8)��!x�� #�9���i�i87��o�\R��&��
�p9o�����[{�����';������VM�g�ȕ�@ֻ��C�1 �T,5�����rϐ�F�(�u�V8aN�T=����d�������H�L.[�j���k������3W�~�7ic���} Y���D��"�@��/��j�6���|��$qma�
3�YIMB�
�F��ԨX��d�7Qq-mt������5��b��r

�Ds�oI�]���-f���Ӄ;tJ�E9D�����\����,ǷV��1�Z�5��ꡂBNe�ㅈ�UH"��;f5���<���~�=�ƌ<��^6m���Ϛ�v�4iHOJ�|���%x����:T�^m�j��M�8�Wޖ0��e�Wh�UP俰ίb�ێ���.x�P��W�jA��x #*�3���C�+��+�(�^�]�~�A?Wo�A���NU�t�sy,��u1f|��䷾�Q���!b%̶Cp@1�Ə�N���4��p�!�̽��u�#�S;1ʭ���J�F�Y�����[������5Gф��lج��K[��6��J�����b���G-�m[^nt �7�����w�g�q߷��?Oޞi��Si��qe�Hv��椕F�;�kaԄf*i�k�wՀ�A=N��f#�40�E쑊��`�¦�La����F.���8���(��NPT�	�"P����X��i�P�>V�x���a�HH�y���M��;*�-�&��>�?@̭(h�ᗰTx^���.�tϡ��Q�!�����":�X4V��ͪ3M���L���.+Cgn��4L�	0qR��,*X���ieҢ]�'�� ��r�e�A����`�c�\f��yk6T���]�;��<�>e�K�v��I����=�=GT���'=1�M�ab����h���O3�'��+�En���xgr���:��������SD��P�����籸�4P7���X�]Z'�E(���R����Y���:b�k�x�I퓠A���%P����z�˨4eL��	�o}���<D0�iT�vcg��q�dڻ���ғs7�&�7qrE ib
R5�)������1s�;B�K�?��ɷ'4 Y��� ��_t4�ڇ�p<�q,����z6[�j�M/����ʕv8��mAuHXZ�Y�a�9�qw�:��;��-A܈|?��=\l�㕍<fަ��Y�g��{^�!����J-�Us'��%-3�T��1���d�(�>��J�J	Z ��p��0��6v��V3����C�@�S5�JZu�Q�0m�_��U�����9L�#�J Nȍ1&Vi����i�I2fŅ#�[w)&���b�<��5ssca�7�R14 s�/E��A��w^D󺧌����:={j�J���3���� ����izq"��L-��3]���=�P#�.L|��׆w�����:e+�^�U�9
 ��'���5��a�������ŪSv9�ѡ���b�H-΢I�f!�����^��d�Lz`Cs�Ą�hg:6=��X+���D��<Y�f�&I�t@,��⠄��\cJF���I���#���A�V�)��<))��,E3��Q+�c�͋G(d|�z
>f�H��Qָ�-?u��/!D� ��.v�Ř���ԅ�&;В�%b(�)(�=�N����V��rRBIV�q5UD��R�L�0�e���V�
ycy�hV>c'���B�;���ո��jt@[p���
ue�g~���{?��LOm5���t7��=
Ԉ*�6����4�o䁰������uq*��N���7]�c5S��#�׊�}ӯ�k��%h�����c�����k����� ;�9������!�wr֞?,�]��c�%��m0*Jn����+E�-%g0sp��-���s���m�6�����˘*���A�8�S�A�n��� -����pL���^��C^�`W:����	U`f(�h��O4Y���N�t�����L�4(�(V���8|��3?��u��>6�N2e<�d�M8ҝ��1�81D��m�aBvlWM�.O�����ȑ0�"=���M"Y���T��p��J�T��2 �������*nV�}z\�8E��OI�L!�1�g��V�)F�E�j�& ��ԣ9=�l�;�4�\#!�R�5��,����v�oC>�Yd5l�UQ�H�ٜ8Lo���8��Mh5 �����5�
����3��8ր�I�.�.�����p�~۫Q��=<��E�	���=ng8������a��S빍\�DY����?lߎ�{���Ld�:�
=ј�G�,�U��;����RJ�$���~���;M �,;w|;{��%i�3Q�F�}� ��k��!�{��+��a�����j�od�������0�g����ȅ����.:�������V�a�T�([|q����a����v�A=|��^&l�e���i����������cǯ���/~�L�� ;fcp)�x6�X�n�hW7ԵZ�'f�J�$�C���c:�(W*|��i� F���Ya�&�S�J8_�OY�\?��Dd�����Q��^��w��ܙ�K_W:�����8���[�'h;,,M��&X��a�ݜb�������{��rj�v\h��[�l�4�W��hD_��!�N�}B���Ƣ���}]�ɧF�*?���V@�ʿ��-��dѹy¼���~A�����tr0�x˂Y��R�-��Fj�I���u� \���jAc�˾��g��;�ױV_���M�(�	U%��-��4�@�)J7;�����vdz�^����%�~����r�F�q}��pԇ��1Ch�kOԚ���6X+�J�#���k��Τ�~͸I��D�j>?��}W���>s��C�<�7*�����շF����x`��n[��c����z���l34'}s�R�]��=��eN�%q��	6N<���YȬ��n���e����>`�dՆ�}j�A��U�|f��4\TΘ�6 ����ϝ7�G]y2�_iw8p"n��U}��+���7̇��oZ��ēRȄ�]����귭&35~��=��|���_}/c��8_3�b��Y�>[��C��t�5�����ٱ�r���Xo�K~�������������������D؏��-X<�I��y�@*�mŔ����3X��rn���Ա)���uxh�������'S;��ň*�]R�=�%dBw��N#�J��ty[U�䯉�����2��d�'�����<�ڷ`T��*��a!��xu(걑zr�+@�d9rK��$?8��&�+�]��w����}v�B1±���'���ߕUW�W��Fb*ɽ��c�:1�$�e{,�~�#$�����c>.��Q� `����Q=#��:ִ�xC�����g�D�#'��t��֘j�΂F�/�����\��qi���Rr;ɀ�{�l
��b�5�����s!�!nbǊj<~��쫲m�x฿���x��a�n��3����*� +TY薑>�[�z��17����-P��QA�$�H�K9 M4��w��om��khJD�D�����u<Fr<�?Dq��p�ߓ�R�P�C����3��!�H/����&*+��e�QY��O�q��N.w�J.����
��ǎF� BB
���Y�{e40��	�qdNc%��3j��.��Ook2k$�c��Q��7�b��hL�߱�Q��9�?�h����ǈ�dƿ3�b{�s����ο>mxgdw1��"�{'��cP�;s-FQ#E���P��Ȳ|��u���];s��P((q��`�2��a�O� �F.�U���f��tܸ)��g��uR��a�"�T�)�HW�o�M�,�mg������t��kP���E�8�����@�Hy8�n<�#6����+|�v��	���o*�����`z�!��+N����������Ԁ�����D�Y�,p�n��vᵡ�������87���t��c�H��e_}�G���+i��0Cp�u���f�]�ң��X��j]�ĺ���?"ۃC'�����E��E��������}d@�gW���Vr�>D9�'�}���3�Q���g��z� �8q�?]��T�:����i�H��bc�dU|�s>�EY�����N�a�����f	�*�uAb+>7��S0��TW�Ji
��y��PQ��G.���hwl.�b)��q���#�V�%X@�=ڵY�V��(J�	t�R�i�y٨��Q��#�<@�4��*C�; =�C��V_A*d�B����,�����6�Ō�.��~y�5�/`Ѹe[�`��Z���"a�&&��w��;mW�a ��SQj~��T�c��AV�%�z��&D��!�p�J��ʂ@�����F<(2��~=4HBR<8���ؚ�JN�0Ƥ��7��Agd��j�SP( ��J�#��\M
]-�9�nk��Lnڹ	�'v�cCz���J�pH� �h{K�*V��OȖ��z�ݪ��Jp�}��kO�����J9NH�\��_�iO�^��I^��P�h'7��x�4Z��X�q'i�G0��fSF�ޱj{�"�C��0a�R�����~�?+)���L���]R,um�[���0�|T��=����[��V+���1�AZ�;z���Q�U\�ukk��0ij<.�ǠD��G�Tt.[�\�� 2��Dc���Ѹ�j���h�y���t����#S�l�t�76>������6=~w'��vrl��n�Lu�[����^s���Q(���
[9?v�O�k�#dTf+^���``�/��w��|�>h�O��O9˂i-c��L��ȘyB�{c�=�oq3�`�e���@�W�-��H�?�u�A�����'	�m�Ҏ3�	{7�"�� +,ZJ.��Gf�[&�A����T_�$b�v� �|	 �c��jit��_���!K3d#�],Vh6G�v�0���{����x��⸲��(�W
k����^�w/*�'�|�=rI�Їd��(�aY�����~�o�S=ϐI�V9�@ݢ�u�؎@ͭ���o|���|���l���q?G��O蚤o�˲k�R�9U�R����������d6y6m���gŋ�Fb
-��v�$5���J؟�"3���8����K�0���`F��J��R��@�3Z\���%<|�� �́_BaB�漬�;�A=P"yx �d#�>�?�?��N��>���=��hB�&��|����TZdL�JL����Gp�{:�1� ���6U�!"�;R��f�åxa�e�J<)�� 0�,fF�=���xG�kN���'5?�BYy����[[f��~�{a�#!7����������%v����A]�N�1.F�="���#�����ы��$���
�1�˩��(�q��q�l�t=�Z���I5��9EuH��}��}�no���Y�Ì��g`����=���UD�L1�fl�<k^�f�t��e̛�Ⱦ�����q�����ma��B��w3(s����'-�:��A�5T���8L�恌�l}
�R=/�7�eh���,�����<�ˇ�.�=�u�F���W=��j�V��3�u��Z3�|��n]#o���_�h�C*�o81آ:��a.N6_����=��sO0
f�o�e\�jd�W��QR�q�a��D5��b���N`�KZ9�lפ���|3�)#2-�=H�-�V�^�3I��w3��R�Eq�����V��]ԨZ_FQ�+WrC��Q���?��G�Z-$T������}�L� �b�/��.AR��m������o��=��{ ���vs�س�$'ԇ�ҁ��x���~�"�	�IE�0Č�e�c>���2j�wC��cm.
�f�	/�g�x�g���s���7�G��M6пw�Ax�����ST��?�.۬�kJ4H�$��ȸt
o___At�\6q#��T۶�l~��`�����I]�3~��+_��S����ȭ��Ն�A|I?�Ӆ�5�v��O����G�C>2�;_���}�]������z�-P���7Q?�{%	�:F� ��1�f���a�/P�%��=U��z�ŵ|���W)����7�o'�#�.�UB�5�'4Rc����ט�3����0n^H�k(x������&�]3�̜ӝ>���<�`Wj99Z�=���lr�ޓ��3�{���/��c?x�3zO[��������"�_f姅s�F=�ăA�zσW�̽���@�OJ4a�n����T�~zz
�J�M�1��\	��g��\dD�a�ڡ=�)Å�Uq����y2p��������7�߂�H�<���7���y�϶�^�Wӗ��C��
���0�U	�CaA/�fBE�6�>bB ���(���1E����$B�s��w�l���-��}�iz��\s�,�SV�X}U]t�,�,��Y]5��E�9����v�ϐ�f%�����V���Dr����~�vL������J;=Z[�����j�P(�D禍���;��=��tXX�b�+�m��f�N5p��?�갡ͪw</��~	9c���ɡ T�N�9��"��`y�������r�}7JU�����D=ح���|j�mW� �-���ui����'��@K&������{Fu��#?a�������v�����gGV�j��\��VN:�����M���CQ�`ۺ�5DVX�I^�ԕ 'gl�T�Vk� �JM�7V����WO�z�oA�s�hQ^�M�UP���!|�E��j���4ￏ(3A�lB����Ũm�%���o����w�4bh����Էұno���N�&nTpD�Ɓ��O��A����ҋx�	<ad�4c��|�����PH�3��t�/(�o�&F�>��umL,Uʲh����؅��� �͔gw	n��j���3��W	'�ͣ	��xE������^�!H��h��_o���kn��z�]a�.��P$yT�"�f�Ig����� ���l}�T�1�Uut�f��15�26ʇ�������(��)U���XLk�_w�g��S�y
�967��m}Ё^�ok`�Qi�(�l)K���]]]�DE���`�0�Jl�J��U�A�im�ଆ-V�K�5׽ٴ����D�mKo�^��Rl�Gh����� J��XM;v�E�Y�&^�(t�����@C�s�6���(�������d��(]`��T2n�K;�pb����rD�6�M�V���5�m��'�TA�-���Ҥ;�d[��i)i�낽�Z{{�	��E夣nS����>L�o{LH�c�`��~�.b���8���Y�\��n��n�0!rj�L��!����G�<-l�f�2�X�%��h'����o�����k�"(�8����j�SH��XmZ��c)���{(����D澄���S	Q�r�S��ݦU���zI����dS�h.��f6z��t0�o�C����6�+n����H4�x��c��!q4A�e��"�@�擓3XFJ��	�qC+N�E�\�fE����͕��7/=	��U��$M�/�:�vu"a��Na)��=t�M��I��� ]4��b�? 	v�0�%uu�q������tk3�"�	7F].x��}���.����?\
�$���j��D�+��}���p[C"���^6ONZuɝf�p�$�Ռ�
�w02u�A7�T�X욞�B�����W��T"��r�14��71�ǖ���XQ��pk�iC��B=��M�=�!P�.��-A
��OJ����m�F��ȚX���%^�i�ʩq�'�~�enrc�嶒v��(8�@��\����2�M������5t��S]K�t�g��ؕ�c�hMb���ԏ#�;���kR���"��S����U�a�?���W7j��#8�dY������'ŷ$�1���y�-�ʽ^��l��*Y��^|)���8�=�D!xv��q���p�p_^����O'��ͷ��YI�ʶ�U._g��Y
��lgt	k֨�X>-^�k����'��E�笑E���?��5��
Wh�K�l�Ң��C�j
���$����J�b>>�DPY��.�ǆ@�r�Ǹz8ʹ���r�ЀCH�0��@��udg'�ߗr嶅aw0�۹����U��N}n=Zx�D"�`���"�b�>|ܯ��)j�[ɤ5�yx�L�z|���|OC��_�O�y<�����5��2Lכ�.ţ�r����tG��2��
�8�P�k$$٥	��5C>ep���ӭ7���[���o�;a|�s�WRt��v��}�0����ʩ�������;���a �\qd�[t��F����7����tU�,_RNW~��p��P���lU��ѨBY�|U�5�_��R��TP�����d����d��o�����x���촶�mΩ�i=02�icQ�J4���;Yr���jE��ow����U��1�=:�f��#e�.�u��X���:1�YƩ��L�rݟo�s�Y%��] ��$�y�����s�;ۭ<�J�7V���ݔ���i�s8�X�K�V��n)�6u2��W�E: �7�Vyy�E�!�HJ���>mZ �,�2	�Y��Y��J��܁��7,Ld�s���� �E�6�˟��2LX^R����ժM�z)<���tÎE%P5��Ā����s�]��300�2<�$�{�tX7�TR�d���>Fk<fr����_���k�V��F�C��Sg��3��q���:�4�Q��`v�riB�K1��j�%�s�/C����4����b��$%Ͱ�Kr��=���������������|ߟ��v� ��PEW�aJ��xs�B#��s���� �ED;���r���WH5��yo8Z⡫S�We�/�p�m�l�eQȜ;?�	���mǀ{G����?�\����l]�y4�kʋF�j�~O|��mV<р�mO�Lِ�d-?�uy�o�1mEʑ��f�E����Ӎ��{ �
Be�{�k@�M��4��k��O����o7�~�N��ŭ"ۖJ�F��o%[��6�a軸��z�bSOtr�\�r�����F-3����XìԻ�=�������ɐ������̨�Xizȯ���N��b״[�4*�Ս8�[ȓ�ٻ{��{h-)ܓ5�q0x�9�f����:�37�y��3ﭚ���ZPM��i�5���a0[�:9�!��IU�5ə�I�^���c�Lx�$5a�m����{���\�ܵ�B�����!8��r	��ۗ`��#���!�Ꞥj`B�&	�	oU5P�����G�H��`�iL]�a�,���s���d�,RT��s�W-kn���5X��`��,�YX`oH��[i��%����-FԠ4�a�PZqH�Y�����Z5]*맱_9G`^��h��jV��e7���"%�!�N���e$��d��ܫ٬k�SP��3X�vC���O��*>��5��)$X�M�9���=�9{�۫"N�_zd�G��,��	uRL�ꁸ@�Tb%�r��4I=�ˉ>渪߈�p5���*K��������M�U)r���~����6��=��T$�#~1���z�J�=�����:)G�Zr�6e���=������8v?�"n�`uT`	uT�Wz���B�HB���ڔcb5V\A&���5)/�?H��ˉ2Ϥ��N�Ey�
�Q��l�H_Ҧ&b�0W(��$��¯�a��w���h$ش^Y׋?���>���>i�}�֥��d.�')>�X����l���_-s�'�䅍s����.
H�<x�D��|�����=d�����Xl^�2i�H��e���֞�w��ܩ�Wg����cEC�J���O�J9�C���|m����\����dr:`�T���2�m�G�ȁ��<�(;���B?����j�l@\:OqgN��֐G`|������SI��')���V�n/y_����kDs�
܇�f'Q��Z�"NV��AW�����M�C�K9$��R�w3�"c�Krp,Y�gDφu�e*��n��XqF��3]��q�a?��Um�5�ˮ��w���v��k.�� G(���	��z� u�nƗ�,qە:g�'wU'�}��z�������.AA-�0c�o)qn��_'ԅn��F22�'I��|��<�%��d[|	7v3K��ߙ��x�
���{qyd���-��Q1����K�T����!c���o��Q�?�aD�v��[eJw��d��3���������\㒁�0�p��t�G���=��։fѿ$�Xހ�ߟ.x�[(6��ݺgϋCaO��0��~��n'N@緶h��[!(�k�,��i�͎�kG����tO�{���>�F,~}B'/���
Z�z��Lw�*�������±�Ʊ'��b�U9����\��>�Ǽ �$�!}�m�Je+�c�^�#�l���ZNxWs-`V5��r����2y�����K�3 X��V~8���GDݟ���p8���կ[�[�� ~و����nnG�D��Y��C�0��3
+��8m7��P=ҕŅ5�u�?Z�������ھ��{�ŝ��ѩЩ�d˥��<pzh��l��p�U�d:�8����h��~X��	�����&/_O}�$/��͆D���^ع쨄e�S34&�-,��?O�y_UKxy����7wr'ؼ��h��6�vSd~qz� ��;�+̊�x9֏�y"��^s���h���H"lG������i3=<�0��"�0��
����H���u�����%��۟��P"�h�Pv��>�D"&
�>
	��5[�����PK   >�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   Ŧ�X!Փ;
s �x /   images/c6ed6037-c211-4162-91fa-07d26f2097ca.png�gTS]�/�P���t�*�H/"�T�A�tB��#UA�� �)��j� R0��	��J������{�y����0c��v�\s�_Yk�wښ�� V  �U{�� @�  è/���	8�.@��J��_�+  7@����Z����L��aӠ_������ҍUKB�+� u���_��Lj�Ĕ/'���d��%��N��M㥹��Zi��	�2鈫R�ɫ�@Mf$�4�6~ez��`?8����>�)(����,�)U$�#?}�}���l	TGV
����e3���s�y����syH%SF��E)�	tFo��_QLn�/�����RP܄2�u����.����߇�y�Ŧ`B����a�;W�-~y�PeV<|�G!�A4u��O�����ΐ����\���jy��:(`�����<��| ���N�]����橷su�Ut�&]$r����g�C�k�;N@v��*��;yf��t'�j���e�����Hl��0s���2xOhA���L�:���Rg�X��;\�r��1�
�c1suQ�rڶ��b��cu���'���W�ܥ5tO|����!e�eXi��M�ľ'y����ز޲��%����2�N�r���{��|Yk�AɴWB<<<��wmI����5�M���~1��j��Z"��;��[�>���s��%Î}r���������3��jt�~%��&RQ��'��5Y��C�Ϧ�n�z�_��t��lez�d �y�Ґ�w�K�m�&X����c�6��3M�]Q���.��*/�0�@�������>�h��b��X�[�Y����[�����;Z�ŏ7��6�;=L��NMM%�����7�7�6�����B/�gZn��C@��i�{{��NEX|�;�7�Y�u.�Q4����(���1�-��|�	�e�u�J)�}u&�K2c�����fOY�'726Q���z�1��b��p�z�M��`����1�b+M��8����銶�b���[��
�G��I�&hv.-ר�80�}�HA�D�0h_��z��%�۹�$ϝ?n7�܊�E��5�*�ϰ���5�o߾���D�(̾�kB
��b[��|����Pb�W�ɟ���L�\ūF������`����_*:��jWN2I�tHմx�P-�ɑq�~0��{�&�L�j�7�㬊�a��>n�YG5��6��V�Q >X	 I�[ ~�,[�v��mo˦�j \������ɫJ��(0���l���P��Z ���3��b%��j���8W	�X++����-{�`����u�_�� ���=��x��E�:�K�eU�mR����okǿ�u�g;��@כ����@�:�rnz7�7k��F׽��N�D{�8e���IHи���-|���	��C���Pb�A4��L��g���,�dp��o&�����U�Sm��c�n�9絛B�0��i�W�� Bc	�G���L˰��L�b` )�gp�F�{�����զ�-~���J�t��rtt�:��j�m��,+A�Ÿ79��e�z�lIi�'u��31�De@�d�����z�Š�u5�sy�LH4~��~��=��S��h9�BX��J���� �ox�0�E�@�l�Ѷ��YD�`_�yx
��W�YT��C"Bӭ�rRL;�;�j",����Μa����E��s��Z)9���Q�fRN;�����7��h����Ĭx�jihL���Q!������iY�Fu���H떦�H�^h�z'����8�C*i(��!�6�������7:���:��
2[q�i��5
08�1��J��p:�m���Nu6[�\�2m5%6}�<�Vƣ��T;9��b��.1��r@
�Q~~~�XZ���D���[0N��.0�B?of�?�M�� P����!��&`R
^A �|��~��z�e���+Vb��F�c
���j�C������L���+���:�$p���l ��O%�~��ڵ;*3��X޻]����2��Y�R�� �C$oߎ�C�I5�j�ޠ��B�m��݅��rJ�/(X>���&K���3] ��)?�*--�Z��7�#�D�%��C�ݯ��� ɵ��g��ӓ*�u`D���^���"�;>�l��C��z`Bq�"�����i�e��n4�&K0AZ��J��%yE\���rp.wvR����Ԓ�I^>�� #M�ݩb�v����?�S����;pttD>>>����JJ�V����HN�dIP{>xs�W?�':�|����pA�B?y`27��췱}�Y>]t$�.�O�d��џ��H�#�uF4|f���XRk�u�q^��q9��:՜*�XvnV5z�-""�Vu���9�o{�b�?�A� �N�PeAAA����#����9�P
��1@:շF���p��*�rhk+��` ��Z4�Z�Af��Z�5�c[d��fܽ����&��m�p�<idd���b�KF��妓�ܹ#|r��%2�<�P�y-�W�(P�o�`�&�...�K&J\\ܢ^:ڴ�� �E�!G�hT���"g�LV�@���s�@P�ړ/8��P8�M�J��N��g4���t��q��e����&�K.�I��O|����Uӈ���I���u��Ń��~!���������G��S���3�to�S]��v����i`gs�j�Pz]�� պ��|�p�jj`T-���5�:efr􍴫�73� MA&�.mJR��I?���,ҳ~W�U�"B����-)���S���-/��~��\@^���U�	R�l�����ܽ{v@�s��i~:_�o_���~r 6^��u��Zg,�v<�������Ԏ!�f�Dp���?B(�)P9Z�� u(F*�P��R�-�`~��+�}��j��Ƅ�0
ߜ��#��A�T�B��M���TS�����R�����b�W5�Q�je��A�B���ջfȃ0666�.�t�' ��8@�o� ��5V�PZ��px�h���#��g�G$�Y��̖��F	���@��_�j���C���wK��L��[��<�J�9���M�Ulz��ǑU[עGc���B=�8z����(\�ԕ���qH�N�����6����D(N=�����&�MD]Н�'�^eǭ�K_zU޻΂�	˔�].X��2_[s1���1�nQ���;ݓo�luxfH��/M�V	
8	3��83_�،��qb�����+%wR3c�晕��YZ��sIy.{4N�q�M�����?����b
�<�t��O��4\q�<�7�D�R�o�r��b��.�w/83����=*Jr��K���։�HĀqL�F�W��vNa�}���EF0���N���I�� E��K���� _�-1�ڤ��&<�ۂ��`�0Rq�d��B
0�M�+��JȂP�)D"��D�����o�T�eLa�h�aR;����b�_�T��}5��z���4t^j��d*�z�$/���^��]4^2�b�
��=Y0>�9u��`e'����F�"����f�@3�:Njf����������i���\z&�$O;�\O��"��#���#ȏ
��2=��!��Gy�4�<���|�0rf��>�u&���%`f��K�~�	&�9�@��2�OZ��G�e��D�:3$2� ��L]�!��U��y} �_����sҰ��M�P���r[#��������,S�0�2�+����F�Q��<2�u�/��H�)����<-��V��>��|Ej0�*����=,�������F4<��v���Ef'Y���1��E^�S;sR�*B�e��(��ǸCDJ!�ÒNF�fP@�t�L�k��	����XJJJ٧᥌�Mh-:���o��)����$P>�d��K���d��ԕw�(l��v��d���+�	ħ����/�$\��Z��2)5�?�$�f�u3o��dC�E1���D/�Qr���/���z�Xȸb���'=���p�&�Fx�1�L��R���sC*����>�I�L���rD4W�O��O�nl��<�?�?Ę������79}��O�����~����)N��Cl	~R�|ry���]��ք3��NcLk�U}�n0�܍|�D�Fz»�����3���ӏ�:�|S�ŧ�O�^���A�x��q9�D_)��I���e�jaГ��/zn�7�K���߿��o��S�w�i3��:k�дtrZ��
\
�j�Kg<�^���M�&��p������^�����zv60BҨǼOm���[Qm�ں�e�:4k�nH�:c�ϸ2D Q�#	����^�
�&2��H�ple�'q5$���HCK��*�p�n	�=�Xp�� �>�I7��y:��>��Od��q��"����fr#|���uK@\�ĪA��Hzj������2�Z�%�xt@��"S�$ۣ1l�ɫ��h��m��Ò)e�r~�i~� ��P���t��-Rf� �J�HH�!Xw�<ʻyә���6�'͖�z@<w�s-�L3��<�H�ְ��1�-��(� [Y$Um8{��hD��L����4���
�OJ8*O�w��"��x�z�圧���r��p�a��Д#C�����|?)����Qt��%,ٽ��EN�I=��8�9�~���D�:T�]�Ek �C?�%= �H
�fT�ڦ�z$�AU��u=t %�Ia*��i�F�5���Hԧ3�T�57Zs��wK�$��wֶ��爯���	����ռ-��j�eFw3cF����V�C����;9բ���7O����� ��`��D���l���X�\�ǏCV��BD�s�']���tɭ��p�cq��YhY�nԭִ@�z��jW3��Jq�x��(\������p����k�6�i��'_�v�sz�./�I�P7��yi�"�!�0���'+N҅�7�t$�U ���Գ^��ê��E�2d�>3�)�R�� !."٣b��H����Ͼ~�g&D��)4m.�ς6����Y���@ڬʵS�	R*�ֶ������}G�q�5��Y��{h�����ai����a�Zb�k�|��a�w�kq����4��g�oޡ�,y"0^J�3]J *w��|�F=���O;7 c_%��,�,��]���o7?R��A����ՄҮ��*,�Ō�+�x��U��;�1��07*]D�@_@U���
ns�4�B�΀�_UU��`-uu��Çİ;��LNu#�[��L7���u��� �'y�0<PC+/�(%�pC��U��)��%Qn�c��7җҽ�X�Х+�^�Z�ڶ�ڎ\]w�n�n?��6q����(�5G���x�sW��+��BMqNRn <�Ň64��[�B����^���qE��(���j3�K�O�f�K�V�����d/�P��_}}M����;����N�o5��%����:�9X"���Q�k��q�R�u��$C������fv2_�z�&���Z�!Jۂ��l�F��$)S�����pm�����������d��u=����5�#L:��[�M�\��W���.u���~��3�/?I�+R�}�'ېG7�C_gF����v����t˧	o��'��$�jҞ���g�&�?!�{��-=U'�!�|�ĭ4$e�� +I��[��J��]���6Bi3D�D��7W�%f[�:a�T!^V1j���0�L�W�`e���o�^m��X��a�/�|:���P0_,���_^f��ʓց6���kb�i�U�A�.���X�i��6�\���$�H���o��� �'�����zUK�t7�o�xj���~��w_�+����R�cD�2XD�N�24�dpq	*�O7�����o!
�%a�>�d��w���aJ���9��ʢ�f1v�,K�}q��iM�nw����:F�a?d�iM�'|��ޱYS��z�����������^�0�BsV��ۚ�m"��tÙ���k���!��]��b�h�����������dz
.@t�MJ�֫s93�i�c�7,�[Ӂ;0,r~t�O�t�.]�˗t��H�p�+`;j@z��ZY��Iw��߈��1_�f�@�� 3[�����:��:�FPAr�b�#��u�|��d�}�f�'��!w��a��.��QD|K��;0�=�(#H��L�d����U���R����ģ%;[���?�����|V��Ь�A��ߒe�+0��ʐ�?sʂ�!!�GD����aN...W �	m���G��1H�	Nl��f���D���_5t�#\�9��R)+�'T���7��[��T��z����L�7����]���� 1a,(���Z>Ő���H��lKݖ�9YdC�� oy:@����{ҷ����wvuI��k-.�'m���ie��իr�~�%��|N�u��2�Y-��vO�5� �Ġ�o��a4¸(	x<���
߮��7U*����r���I)9�y����8����6~C)�D1Gh^N�ԑ�Ƙ���j�_&iA��*T�%	N��q����2�(�0q�{Q[�(����NP���^Ө%!PL��އ��S�llV�^����Ĵ����ٹr��{:��A��Mڠ�CI 3?�i�t�eanR{fA��.XZߢ:��\�E���hu��j~�YX	�B.�8P��Q|3z=���������5/k�ϕ�|���$F�m[����8�z0���0��n<�oA�<�/ET2 �y^�rZ �v}����w�@k�w�9��9><)�{ʇbcc�&�ħ_��\*��333 ȁ	��K����[�	���f� VVs�}i\`3�3�ϟ?0X,W�4�-����7�Ԧ
S���R�p��5rQ�[��#3Ԩ�ݒL�'y֎�=�����)|A�a���O�ME-�D>�'�:��"K|e�<��e��0��O�+�s�>!26�[���X��'��󦨥h1�F�.�䋮!�VHƹv���Kp�qs�e*:��Q�R�>�ʊ�ђ8=�T�#	�ZN��P���G���ܭ�B��ӝ|�T�sg�o��e�K�F��_/��̗=�T'7�U>�%V�7�=�@��w݃1\%�ռ3�-�Hk��=���d����J��n$�Gc���_��|��6��2����O�������s��������*M�q�VVV坈{pp�0&��ӻv�m�����϶U~����Y��� <�w�BFZ��b˃2����V]q@ 0�x��:͔rg�����ay|��A�{󤢴500H204���8�Y�������ĭ�3ߛE�[x��UƎ�qJو��4�P��ж��cʘ|��e�q��}rqRzZ�OD���3��Zs��5g6s��١�K����m7��y���p��BCP�=8o�(fη~��e�/�M��>x�?k�����{CCz�qs{�K�y|��^>��Q����h�	
���A�3�uuq����j���(��e����7�9z��~�\Q�^�^QvD��o�����85���fYK��Ȧ�y Ȁ-�jo�-�@�H7O��3�)5z0��꽼i�4ж��Ҵ8t\~m�[��������91�y��W����qͻϤ��hkU���rr���~���6�j�t!f�u"���ҒH5nHB����4;W����z;�q�O^�pR��J����������FL��u
�'�ARy��~��e�kjč������k�3�R_6d�x����ʨ��7=�Ф��PKd7�+gu�G��|_A1�N�z(�@na�`��[��ވyY�!h�CgB�����!��+ܸ!G� ݞ��Z��Q��W�ـs�:i�����
nV�GKz�σ��&]X�k��ɝ�����\�z�<����H*�\.�D2��	~D3�qB����|�����b��Z��H��Ơj|=���l�O��x�%�R�����b.#SӠj�- �%�z�uѨ����W\�J{��7MK:졀�,UF�R�����Cٶ��QC��X7,�o���+���,Y��99`�~��߯T�E*�.�����t����Xc���-�*�i$�_�!�7��Ꝼr��=�q�Ɯ�d�8 ;��m��wu�d��GpT������׉���������K���􋇙Ib���������$+����Lv���v1�7.M�l��n�QX��;Z��y�R���~�y�5�~���b�˯R�0��b�7!��@��y�R5:��H��;i/�*Bʲ������e�8NYgKKK�V��,����6Z�&����|��u��{s~��GIi�r�+��.b���ɍA1�YINr�h������.���3��q�>�������}��o�qZPLQ�B�9�	��J��ߦ���ؐM�y�%Z3fX���\Y�m�l�t�u%�4��5�1lh4�\��|���p�L�N�i��,����E�i/��$eӑ���3$��c���������4���;R]�Ժh�:9��&D��p� �ݻw���g��S_g���eL]r.�nD�3
���`�L �����O����9'�pG0�x�Z���A�m��f.������YXX�SSR���~�9ZeW�����6
�J�5Q��i�) �0_�'Mtvv�XXXP%q���I���ޞ�
�T���|k�O?��E-a�/�9�br��f/P�	��tf#�Ҽ��vU�.bnQ�cz����5��(J����J��z����ǐ��z�,�����c/����6��f^�p'�e���S'􂀑�u��vz�#�����F����J�1VCS�VZ�r��;���ctQ�h�B�!w��$7�LB������w��A0V^#� �_i��B�G�N�v��C�qn�6���#^'�[u��oz�E�N���D�?�8{���@J���i�a�����1��!�kA;��_G�������2�ohUU4���F/��	8_)tgxv�i	��{n�}�o�U�?�̡�D�[1\(���A�x��2(�Ͳ�Bʚ?�T�w[������`��t�+�8lxnĨ�6b��瘉i�ҥ�E`�3f��8��t��냰[W�/�����%u
�%�{y���q�3��iwo�B��.��O��%=vT0�w� �8�B����%P�L��AGmoo�
��*O��"!��N@���E$��{fbɘ �/cBv�	!榱�˼/Rt�H�,����3��2�8zS\Nc��p����g�fqfr@�,�6�V�^K��4R��z��|�/��yS
��� 9ǧ���ć�״�Sp��k+}#a�D�ɾd�~w���'v
��Eȸ�f�K��^}Y�c�n����{�4��{�B��}�}!� ef��IT�U�{�`G�y}�y�+�����c�)S�ԩ�T��?��!����������},����H;Ïk�=-���i$������󙳗��0���dٗ�de!�d[���o�\�Ʀ���M��ܢ�>��16Ԉ~�Cl�>|_��۬�VNBb��e�i�Ʈ?�)pZ��iw9��ݷk:��L�F5��u��:ۥ�cu���dpa]���2���\:����I��'�`�@����C�,�	��`�OXI��x�G�_b���N?�L�V�%i��R�R�"�
L�IcV;nj����f��q����v�t]��4�c���������Q�����:%�Ry� P�=F��\�cp3F�D�e\7k��� ��Եˢ���;eܒ.��RTk�����Y����X���������e �j����������,U�Q1�>%�6b�0�#��%�\�%H◝T���vz�S���c�׏��W�ɏ�{'�uuu�A����ɹ�����2]R�!�:| p�@�pCﮈ�e
�b��	���ߓ����lc-(/j�W�v������-�۪E,ҾjU>	�����\����Y3)�����ek9��-g�>ѿ��=^���[��O������jy7N��j\������TL��o�T���궭� $�k.q���ifʤ q''���&�M^T��.mm&/����N.�e�Z}2R�&��#���V@"��*��gI�ɤGV�2�W�D���}�~��o3]����?Q#w�ȟ�ш�ē"�Ԛ��AWc��
�M^S_�:8=�o�k	9�Atq� �Nv���Ҳ��iii=�����
�J���:���]qE��|+{�C�,��WH���O�������N0�����Ɩ�����>Y=S:�$�����_&~-�K�>��>�<��y�IR�1��&����͡�Jtr���Z��!�i�*_�e�eMx�͟h�HZ���]�	7�p� T@�pXS"�[������g�.��SB�aޓ6�����/�����h׌olƳ��9��̝��h����Ɏ<֥�k���Ǚ��G�n�v�hj#ߵ0��^&����H�T�}�i�)b���N�ᲈ���;%�Ӻ_л��/E�E
Rm�m/Q"n� ��2��҄<U�gх��e��Rf��V��y��9��Gѹ��e��$��Q-�-�r���%�s�����u��{�+p_o�L�ϡI
Ó�݂���]��H�Fϕ�˃y)BuQD?�86^j߆V%�l������D�~����x�o�̍�Q%s�H���+��:��hY�������&#s:�TR.���9��%����p�e�#�x��v|��zSẄ g5i�s�W��fS����F���6	k�Z���ڭ������y����C��Y�?LV��Ψ��oET�����Ng�j�l���ȳ��|����KY!g�m,̈́W��=p��,���Fcp�	g,������5F�	 ���z��gɐ%�%��۞��"=�ds���
Vx�o]U�&s �o��ːey��i�������C�ZA�h-�S���T����8������?��w&�ej£Hh� 3�b�JR|�v�W�1���hO�)�˻|؋�����xk ����=p�K��tˈ��{&֢�e��]���I����I���l�%�[��N���O�dmR��X^�i�w���y+�5o'<z���w�PpS/B���-���ِ�_�� ��5�������za`V�4Y���R�]�k1�o�oL�H�R�/����A���'�����w�3��K�ztz]������P!I:`��N�u��=3�����h��[�D�aP4�&�V+�/�+U��'=b�w���)�D����F> �\��ϙ��*�|3x��|���U��y��?h�#ć����}�����bD0�1R��h/*���R��?soI�}T��+��9�?\�����
aM��/�!�ɜ�0��B�Nz�{��"�
Z��/�����:=�p�b���bM�(Q�Q�ὂk]�˷Fc/3S�H�
ZUݱh�h ��2i��%�s"��1�Ԯ3�g�A���X����#�G�r��lјYmƑ��GՐ~��c��Q�t6F�c�w��̖nS���w}��#�+��5ٶ��(M��ӄ��#CH�i)� ���T	���96�k�2}�|A��~�#�+**BG��O�w��G���nu 7�`v�?����xD�4�ņe�ZMf�z@��n5���!nЂ��@o�f �j������ba��9�p�Tۆ
h�J>QG�`��xWWW�ֻ;��xٽ������b߃��!X���ς!fe��f��2��n�b}jO7a�՚�̈��]��Q�vwO.�N*�E�ϰ����$��B��oƟ}Ԓ�s���H���
I���y��Yl&�J���~n�����Uu��j rN���>N��:�W����� ].=��a㳠af��$�,�$�\�F�?P��;��W���1�t�x~C@����#}=���K�*��0�Z�����66uA�4�����;�Utq�{,�n��6��.Ck�{�t��1���$5�k��xxؖ�KCahoO\�+��pCm��e��8����\�l0(����}ɦ�H��J-����g]_#�]u����cs8���S�!��eDY(Es��d�{ܵ�tz鷣 ѓ�˴�"�z�N� H�B�o�s�?�eL�"�J�,��-��Ic�w�)�=,��� �A���p�{��SYz�LM=:t=Lr=�zG���U�C��6�&����ǿ�j�d$�����vC���4aRxX�w]UKąTb�}dC���̀��Y�?.�~s ���AM/8���*X^�TK���s4-�Ή�}��q�����M��tY��q�:��24퐓.h��<�0��G�2����2�u/�<�RNd�+/�la�LO����Ă��1���U)M�!���>�e�tE��*Fջ1CCC��$�8%��4'�}+m�$i��߯�p�Y�t[P8�8;�n7N�F� L��I}UjP,������w����EM����[W#�+�4�t� �����]����^��8��0��S��t��bP�\(�·t1��C����#�;��݈m�������r���@N麜�н>�i&e�f�����:N OR���x�3N_���~�.
�*99��~���O���%}}}.���e�;@g� g�Z+�U_ral��^n�MZ� �������ޱ'3(�Jkc(����'���! }�����Lf�J B���M����T��^��h�>�Ӱ��ݣo���� ���V0o�GT3��'/<�#�K(㡪�͸��Ե�BNLZ�&�3'''ό�ΐx�MSb��2�ϖ�H�ˇ�\:�@ �%�X�Ƞ֬�
2n����!�S-њԩ�C��[
/U�_��&b�s��C;�D����;&7;�sZ;�W2�ш���P�5&���!�ӽ(/g�@���e�B��W���⢭3"x�W�������W��4�#�z�rol��[��`�ꐠ�fթ/�%�S32NG���VrRf�Q�!���O3]�A
��L!���@d?���B�3� O@���xb���ƿ)�W�͜��D�S5��`�Ҿ�]/�j���M�x�*%Dy�n��`P�}��J�^��1��@Z��@��Z���(�f�PYF���p#�C�jd|d� �k1HNm�1���m�xc;�)&�e���_y&��"Ǉ6��p
3R���N������dᱶ��g����"$��T'��n�����#u��ی��t��1���U�.��p��uW��a�P�|�cݯ�q�%6��gCg�Q�&��߇��<�Yo]4��8RY���kh�|��L�dP�<�I�N��Ӆ� �K`�ɋ�.�_1�eѭ�"�D�]=��Ş��4���RI+=&�d	�b��}D�]=$)��ļ5���q�~��m�a�)#-}�
�5���d꘺o*F�o�! ҔDx�(��j���C��GiW7�ԗ��8��R7����7�J�y"���K�/���R�.Y[Os���Z��GY���=ZtS�Ĕ����/8e�Ҵ�7=!�؇��h2i3c�϶aB4@gr�Mn�=�^A�c�ŷ��ʧ�p�MvTH��W}���*��R��M��p8Dطf**;S���N�W�� �KRL�RRR䉭���\�6��F�$n�RG�)�]GB@�h��������_I1�E�uh�<��񪕷�j�aۛ�Oj�l�a���&]$�j�P3�	�	��9�vX��V���)	��e�C"9���B�%Na
�3���F#0�vZ�S�%SlK�d�/t��_\\|}�r�r����{1�]�t%�0�x��v������Q�m�_�J��JR�������ч�ȹg[��e�#T�ިq��y5O_2-��q�zjԥ��+�WEG��A��J䕼BA����J$�y~OkDk�ء��0ڤ]�|�
�>�/W��܏Οh�tT9yPt% G���U�sL�UN1�]}
>�b����@��Ņ3���8�Y�4P�A�6��L�L�����$amȅ*<�"&,�*B�$�@�	wQ�!�>��c_
Mj�`�i���w��s2%��M����~?+j�����Jv2�C�Ix���c���)�"�=?�iN鼤�m�s�87+�&�{z}�"}8�b\��.C�շ�
̕%�o�&DDb�� ���z�� ��*�#����(��?�"[�B�;~�K~�1�Cvת_w�@�jK���Z��`���@�"hb�2?���`�j������i��lc�P�k��{�m�=E�+�o�����d%.p�F�Iy,�j8N]�I�H�d�e��x���1)��1y���w��[]��K��H�z�嵡�OB<U���� ��Ϋ��۟�B���<j�r��T�ҽ���]~�����j���8y��Of}}����X6v��?�0`KL(dF��	���JDs�F#�v��5�QO>�+X���`+y<�y���ݏ2$Q������
�HM���#'��:�3\I�knSg3��o}���}4ڏ��rD���}~����E����r�A������G����o��J(�\��F%�{�/���K��S��S�ԣD1w#���Ѱ��k��4fƜ�F`�����Ғkfٺ�Y��7��sE��LB츮(-���&�1%����&sz�$O����syI ��[��N	�᠆��>V�����9�5kkk-5�"�]K9.��xb���5���9壮pkW3�DI �W����2F�-zyL�Ze�����mK����<��J�L��m"d�sD"�u+YY*B�|� ���n����Q|F����j��(j�����*��"���E�24H���Q���h'��_�\������a��?K��s�?���[��	+Xp!�:@Jt	<n5:O�Z���,w�0H༛u�zWr�!�<��!�P?}'	������a��6,lVBl���	kFHͿ�0��PM�O���LfpYa��̙U�D�͌����y?���ֶ��T�"u���'"j�b��.�	 ?ɛ�Km��Ǳv�Wڴ2֨k혗&0����?��[�S}�T���u6���;Z�'3]�k*�/63�84-�Q��d�.0ήi�����UO��շ��OO�4��=����u���,-��<�y�N��SB!��>��5S)�;���&|�+[�GrXgV�7�����n��/1S�l������[E�2	(�a��{���T iT�*���m��c�3a���yMǡ��u2t���������'*������uU6���t+��Jd~�!a����˷���i��N�{�l�h����f1~��f�HI1%zΎ����^��מO���K|���F�-!'k9]��s�`�� �H���G�+�t����FZZ�<��S� %]�k�c��򣫅LsZuw�:B�Y���i72�GT0��B�9b#1��u_^��2��d�.�O0��i!NVnB9 �I2A�e��T�NN�\�'c�Xl���ux�'�u��<��h%^�\�ЌvD����;^��`��I��F�џo�󔢀/�[�fN��*�\O5hF��L�YV�����ڈ|�4�)?�ށ�,
K�S�������I!�Z�Z�Y�T��D�����
�'VJP~҇Wz NW;
������,�b4za����W����gɸ]�s�r��ǟ��Z���.�U�������?��\�/�(������Š�W����x���|0#�s��4��
9���*E��L{�p�����\O�#A�ת 7�NSة�mߞ98�e���B��r��;n���h(��Dek���ʕ��&�����K���M��7]�U��57���-�>�o!����c��U(���K��`-��:�[q�4�����[�v�����ӴO1���ߖ]��Vj��g��T�]�����\��}�N��*΃w�Jli�d,]�@>d����D�x��O�/O����	�NF�ag�8+���Q�/�$ߑj+R�%Ow��H��ao'+�;R�]5�`�Kj X��� ��JSڷ�x�2ӥ�<�¤�����iLs�с�sʝ'T,#��M���v�8��n��Y�M�K�ǜ�e�o�U.L}p,�#�/)�s���/��(�l�SO���s�E^&���\&`omA�t�O�~H�`�s�[�PU���K�Q����=���E�	%��;�@T���I�h��kT����Ӽb/�R�������-_�كz��]� ����C��ׄ8��\��=&(��(y�P�15+Y2�
�+�G�|��9L�h*��� 鴢�c3a���!���񝝑_�w��䅇"��R'�[wu��om��J�,#�p-Mͳ�(N�岻�¦Ml^��'�$4�����_�y������9e[�7��[�G`�7EY_�	൤8��^���D�Z,͗$�P�&��'���aZ�n��"�h�U��_6Z��SyA�Q�q�%����#+�|qoQ~������y�)�% ��$�,������J�؂��p�\�`�G(F���b��a~�T�KD'��\5��·���<��Y�yw�f��O�΀���*�%!�b�z���5f�4���⢸�0�&\9�Z-���-᳉��,5#�@t��(}
�9��Նй�Ff�R�I�P�+~�*Z ���9}|<�T�>��c�-��0x�QʷQ)�� ��16�r�QRa��؄��2,���zf��A�nT��K@�HJ�H+C�H(�%�]�t�C�C7������vκ��k�}��*FA(�ɩu	Y�|i;"'���t�� ���X��>rIs.�����5���k.�xK))�2����&:�⼸fI$��B��H��vF@\:��wo9�P�����O)Z��)���D��8�G�~�E��8(�ه�aĆ��4��E&t�3��7��F��a�W�P�����V2�0� �ۼd�<�1I�u�i�jm����>�rҠ#�fxd�vx��GR?�n�h6��D�����Ⓙ���)C��K�u��+�yZz���L������M_�{�m<׃Z*��<��������ߞ�k�,s���k��a��
��W�CC���(�����VDv.sA5��7��S����I�u��Lfa�������z2
8'p��N�P꿖^��4�ng�֍�I��i��h��è�xyH6���_R��7��ٵ�I��IK��q.C���fN�S�d 6�A#�W;��[�d� �n<	��v��]� �FSPR��c?
\���n�7�r��Ve�� ��z��|}�x	% ����g�&דK��BDĝO��n�48��T�D�NwQj��� X�B�6�z ��@n�\�'_=�vj�\Co~��R/���-_�W���� �������t��Ĉ +e�kJ),��)KA�A隣Ex�e��s����5Z�����������r��@�o���eM l���{���7�ܚ�]��:�����8�����b��«���C�n��-�60�����V��054��/ż�t��E��GtTk�S���x��)��%��n��+�q��Y��FPu��^̧�Q

`F�tpP�)R(��P�Wq��Υ�ģ����xo���W�����>���UcI��!�P�f���m�m�ʣ��M+Na��7������������*Ȋ��SB�,��D�Lx֫#O+*���2ci�H?;�4�j����HS�a�8J���7�B�2i��W��w�_�*c�舋�zc������i&����1���t�3�Ri���;��\gѧ>F-�;j� w\�[[s�1��b/�7m7<�Y`�4��r\�#�6٪ji��G�O�i���qϼ����T3|v
�u|�%7�+⬫y��so�oJ�����S�/Q#me�q"�OWv��i?`M������~s�4� :�p�im�G[��� �/TnR����P�_"5X
��\-�XK�z50����aБ#�ǰO�o_S{����`3��ҫ��5��A��(}��w�F|�i��P�3� ��P����g�j���r7kqZwm:��᥾��&
�sԼ�<PB��_?�����Gz�kj�mة�oAyw���`�/G�����J�Ȼ�$-?X�-�%������)hK�Gq-p���-5���#3��6�x�A�W��h�@@����V�hEt�#j�ɮa�0a"F۸��z\��Ռ��@i,�w6E�Lo=��^�E�0t� �N����YDS߸E��6������� �R���dC��eܼ$W�f:]X ʃb,Z�,P�^����}��#�,BQm�K����-�z2����A��(!|�{9�c�Y�B����B�~���bE����{~�OKN���w����*�!q���,�D¾�:�\�2ص�:�C��]X�������z��QS�`s�s�i9��H0Q`L��M8S9���%nZ�hBN&�Q�3&�|�Na����cb��]p�R�����uu=�|�)�߷�Ĩ�p~�'s��׺�~v�ib�օl��rģa
���vN�l7r��C�z便�E�/���-���3�(�L���&��~���s)��W\���I� ��ډ���W���,%�+���+��h�a��q�����?�х6� �g	�Zo+��ؚ�ɱ� ���N�cQ^�7"�fċA͌K�a>��NM����&+B��$�����{m5���:�1d�|���N��#余�����D

����%���	F����p�`2D���)����⟤lSX*�A߬Z���<���yY�<P�����¼�݂<�)�Oz�
��葚���PJp4�ڃ�W/��U�ǊV�0b�� &F��j޺ۜ2N�Ѕ�3A��w�u��s�-N��3�Ny;Rd��Uo�2F{K�EU�O��bxV��1��!a�Gu��r�C�cn�Fi���_�Oɍ\6>���IB6�.|;�������{w�,�}�/��<��͒B5�Z��>{�Z�m��4w�.d���x���v�K�
�^+l�r�n��\u����⬓n��Mxz��W���U�`�6�����G������mV�Z$���s����@T��FI��<km���@%��g{�E1���7��W���3Ǻ�i
��ʺ�?x0�Jz_����
޳t6/�4cO��[�)�%o���9.���b�0t%�G�¥�wƏ���=��$�u\�W(��,fC�]$J@�3��"�q�!��Xm��G�����:S�B�Î��N{���	�K�����{b{��g���P�:�h�L��|C1��d-�J��n�p�s�� n[H+�F�{��O����F����{^T�Jh=l߬{�"��5=�`�����3�_�0��s@��!<gq�<9I�gZ��\P������9P�9���5+�T�Ɔ)B��z�pJ3���߰����1��/�=gg�Y��~h��9�]���/��l˵KN�
7-�K�x�=e�*��'�za]�Z�����=q�d��55SuX�=�'�(�t�b愙�/;�;~��ƽ�SO��f$���Q;X �d7�&|��À	�ӈ.鍉~��&1¾����^b��A�*B�(���EM�p>��@C�^�
�����?m�^�ګ�k�ú0��Ғ	�S:$�Z�����\��?����<���}�/,'���r��"{�_j0��{Yx͎Ã053�Y���u6��a.��4'>�}{?a4ӏ�VR����"�ay)x�. ��a��4˿YdEOzP�u4�sR����.��$&�ɱ։Tՙ��!\��7���;zC��toy������X�q�y��+ϡ��[,������[k��fi�)/X��g�u7�{���h���F��H	qg��0��«Q��p����Pk9��*c��Y�J�!W�f�UσU@73�?���+��uiq �)�A�&�M����Z6�@��T����g��t1ٶef�Z/^�Ƚ�l֩V�Ϊ��Oͱ�aCq�E<��{h���8]���əJ��}�:�T&�>Y�d�̽���S9l&[w�ɩ�ӱ`ou���07�)
�{����-S�z�6q_�W1T�5�Qr閥r��a���_�|ǹ��#>�cz.fBmP���gi>-w�1�rwJl��^�����P����z�NN�l���<L}��M_�Ĵ�t���k_;q��"M�a!��@y�}���xnׅۨ$��G_�'�J�����2:��Q���Tn������F�ȣ�
�����;�����:Y�YO�J^q!�0[�J���$Ϫj(6��T9	���E� �rE �Τn��G��f�Psr�R㳺{�g��n���塳��_�hFd"�H�)��:t~0/���/z�^����gh���֭q�N�w(�H^p�����a��>ZK9o��;��G����`"KII�\s��3�u��p�������q��-��+�CԬ{}mp��h��;��������y���*C	�Ӵ�i��V����mtr����������g{��\�f�U�%N$��K�KK�_����K�	Ȩ���]�<�+!��uE׵���7h���C���޻N�ت���$��:-��f�J�:���nM�]J���y���h��R(�S���ۂڐ�fx���1>��m������ǉ�����?KT�uq��u��R!��co���po^`u���L�|h���������*��D��`�� �c�"=&�o��(M�ԖW��+�023O�|����}>�Q�Z5'��?#-m��¾��A����v���{Ε@���dՎ�ůP���,��ό��b��U�%#�0����mq�Zi}ցCb]z��5�c�%ֹ������S�?���@��P7.� �{�O�xܳ������1��T{0�Gn4q���bb��<m��Ga�(|)ԯQ�.�d>]��C�i7]Q^�y�Wr�>'[���R�#���ax�Z��H.m�i:::�㌗����;�3�-.b#-�8'�,�9��:U±K]���R��0J=[�ɱb}��G�j����S�J�`���)����^�FL1���� k"&�re��s�IF��0I�j�����7��"H�^���s�'�=La"lM�l�忓��~��-Ғ��,X�>,��wC	��7����%��T+j�*�+�
���g������.���߇���Jb����������seqV���d��qZ�	`P��� =m�����≫��;���II���6�w�xt����OUs{�1:�'''����p���#�'5蔃�H�Vߋ>â+���}�����k�̝~���L�E���]N���9�u�.���T�s���6��9o�23��\��sfY�2$RS-��/�:�L���s����V�O��cĄ#��y��P߈�Nf`��\����Ir��r�R-W�d��
!���!S�ۅ+r�(��G�/����6��c(���"�wv
D�R���8[`�����n� ���t+��J9m�CORSGˠ�^؛gO)ڣw%e�d���wħ��P>N�8�Z�Rq>�5���Ƭ����cX���q�@n�X�����d1�ݔf~��+�λ�}��]�gRT{��-q�0a*��$=#L 	۞��9�re��b!ߢP\�VV�j���]���z����;fBt��o��9�5r�˷ߢU�b�u\&�)>��w�1��/�lkƗ�i3<����z�]�f�>�Qł	f�ӧuG�$�@�ؾ=�H�׻�q;:�H��p�*,�9����������5�Cn����o�	��+��#����=�fkK�6"�� ���-5�є�����T�]ƅ]�xY��En�7O�k�P�<����T\\�\}M�I��Ɔ��cʾ�8֙�395t���Z����wtr���O>-h���o�j��+�@�����;Ȩv���gT4��� �����p��e�{�HTQ�������俜�jB��������������z0ʪ�,6��)�ȴ贮u�|{)�(��J���Ԕ�.�\mF��"I(�t�%gp�,��3�E�»��o%&ROU��'�X�+X��v_%z��b#�#׎��v�R���-����h��M��=@�$��U6��Dclю��F�Ĝq��֬�]��r>9F I�B4�<68�S+�(A�$�Pd[O��P����]��������:�/���J�Q�t~^��p�I�5Yz^;�w���`a� �v7>���{�`�CDE˦���-�!�e"\�؆\Di����EO
�~����ݐ߶����W쒮�'
ӂl��1�NNe'[��˝�����3����6?
z�؄�U�j�X��2��cjV$oV
j�F�
�ogh�u��}6�"��.0�?����_���6��-��d�t�~� ���۵�-3�ӷ�7ز;�[�Ʈ��@�x	�/�l��υoI�jq���Q	��W��3�*&m�-�}b����W��<�M
�=��w_7
e�B�>�.���OJ��Y��l֮�>>W|t�~���N���"�
g ��������:z�szm``��偗���5𙱓Os��Ҍ�'��띗�������S�0�z7twjY�}��b}�O=,���;�S��a��d�?�'SX�*�$j[���פ�aPY�R�U� j)'F6y!XY3�ݮ}��m��ޖ07%��p_�>&�{�D�sk1'�������g�0fݭ���'�ؿ�Æ~���?�R^��g_G���tq��)�)�Xo�x֋�}����h��hKH���d�\ ے���Ս��Z2����+Vei��{��#�4fחot�$�d����ew;��YCS�wT��M��q׍qw�E7�zH��2󶻓���{��<n���Ou�����>��h�� i�91�j?�|4��]Dv.��kT����Q���P�<�'c�.JiX�@�5�§�`uf���v4�s)�"�X!�8Q���M��D|��7�p���"[�������x��4�p�_�9��t�+xv��w�<�i�}}��槌A���Y@{��=��m�z97oX�T������|{�+OY�1a醷���e�P���`��/����'�K>��w���f���K�s����>qqq�>�a���d�����6I��\�}:ܕ�,{�m�����<�|�<�S;�wc��.�����\T�muI���(��1���l/�̬��̤�[2m('J�9� zJP�=��`Z���Et�ǂL|U*X���K?��O��:)ʛ�=ɍ'�V�D�=� Pp7�n�/4��Iz��s��]r0�h7<�c���Z���T����d8\K��r�� @�[7�$�E`<��{c���[Cw� ʭ����M�_���l`�zg3F���!����W��y�c�4�� �SG�c�Ul����W���mq;�X�7Op�������ry6���-�xJa�����65�R���~�o���ah�М2?x���X6�@���8>D�fP�4�q4���9iH����8�o�r/�-�t�G��4�����`k�;-���w�_6+?�({m�9�-��D�5���"P��t��'��A)���p��I���B���զ$�����*��7�%��@�üK7��#�#ނr�i�-��g�WeTz�:հ���Xyp[�N�Vҫ~��7R_6��z1H���@}v8�.ƿ10j��5��-0ְ�[�� ��JC��f��������|����}��o��>¼!�vV���Tn"��g�?�c��h2�����c�g����d�X�'���֥�iP��=����^�^���s-���U�/���;���e��2i��ǞQ�ŉ*^����fH���}�.����0���5�w7�S�� ���edZ^�';1��g��v^*�~���d���^��ؾ�$6U�>h��+��6m(حYs�"��m�~q��в��I"�ĸ*tV��Y����X��FX�j,�2�UZ��:'j�B�L:=f#Nd/��I��8=�G�E�n�<����{����|��"����ȋ*s��c���.s�l��s�ؾ�`�9^�?�΁�V�1��N>P��CGHR�Z�"�t��f]&|��/���5��β F@���ty��Z�t����kS<���86�CY3"��P4�mM!���ˉU��k�^y�1F����u���Z�O}�N�A�++]��rՖ<�;B�d%$�Sm����da��﨧��eѷM.w�q�$���Q�'/;����Վ���[\��0��ԏtt�Ԁ�����v�<��} ����A�o��_������ f��GҎd"ut���)���V�U��`�2痒���:�H����ɑ�)�}7O ��(�XUo<n�~=����-�?e�H'����
��W&	]�L�P�;���)�S��		Ҿ��AP^�㈋�z���˿/����<�g�U5�`IC��JC�NB�����.�;SĪ]1o�\<T�訤������O���ޙ�����N5���'�Dh�(-Ym�R/'8��?�<���������6��Y�ߧ,����g4Y˒D��X��-���~p -�^�лu�u���$9��p�G�R�<�����l�^�ei����"��`u!�Q�)gv>���W7���ED�&tb�E����p6ã�9���gZ�9����0]�?��	��t6�&]ER81T���]��Ҥ����6o	��,l�/�,8��!؍� ֚N�(��m�fg`�����=n�Jꝿ��|�Q1ޅ�v9�D�U���r�9��J^�v��
�Pdـ����u��6��[���xn�w�G�H*��B�ެ��~<V��v˹���h����u�o���/!�-g�ݏ��t6۫L1q�m��F�� y�
��˟IyJ��)a8��|���k�9x���hB�k�>�r�dd7\�(< Y�v�w�wy^3Z�Z�x���'��m��z���J���q#Ɏ��}�1�C
��>TIS�Ї�t��!+�GK��-vT���vU��T{�a�ImNT�`�4W���d��}�b�t|��ѕ�Xr���p։�vp�.GCoޞQ���Wy����`_��!ŕ�y�1VB�6+�b�)�ź�6�|,	 bwb\��H\�р 6��'Mq�>���;ژ^�O��m�M�fѧ��0-��eA"_����"�%��~J���h����"R|1�[��C�	k��Б�l���p]s�eA|t�r1#-!����_E���ǜ	�gU�� m[�����Q��7��
,�~o�	��b�c �a(�p;.����F��U�@��~n:�F�%�	��5�v�Ӆ�p�t�Czt�i}�fZS��m�E��AV���t*fLV�1�6��̶WT`S;D��aL�C��9�%3��I�ӽX8����h��/y'�[��kY�����]ՒAq�^R���ɶ]�
�&�S����������D��	X���J�.ң	�����s����榜�C��?A�&�ʉ"�龏&yhB�N�Q��O��^k�7))�L�v�� bʔ���p�<+�����P@� 9F�O�4�S=�W!��ÈBeQ��1*�V�HD�<��OI+n/��.u��i���/&�m=���$��Dm�	@�N�ch�-�O��:1HQѭl6���ϻ`�固g��ӻ�_Io}E�Û�D\���w�G�j��#�F�®u�qP1��d� x۹}��'Q���*����/�[�����,Nne9�Nd|X����[s�����)�1�1&Ya˺��3�����ÄW%�UC��!E����liI��y��v(�≫��h���?̾b}��1V� �E.�z:x�;�rvtL�C����ERڛ�%V�@�3"uSh��ӆ�<�l/B�U���̍w�6RYY	=�=��r��_7s���,i�
B����Ɓ�|�����8HڗزCN!Q9@���U�e9�R��=ᦤ�^���A�ⅬLO-sn@��8R�c�5Z��(���*� ��E,f�df���U�2��m��l��W���a̓�+=[������Z͋�l�2�i�B�S����o��KSH�3��W)U0��m=�fM�;&F7�w�׷
��R߭�F��j�&����N���� U��3Fo�|��lb�O��$#����"-������?��#onn�|����Ԡbǧ���U�,��x"����"#�4��孴0I�S�O�D��v�Ńn6V��f��h�[oL\8��s8��A���W�6���K�Ll��J�~pBQ�Ay��Bmܕ�@E�c��lj�����D�b�:�zk�5y��Exg �����~�<b1.���,���}�a.@G��!A��j7�<���;8F��Al����C��N]�J�"7nG�@u�꬐	n�K�_�,��X����7���Ɣ�@��X�6��C�z9\ޣm|�ꨁ�\i�g|x�gX+�* ��tq+=�e7���j��H�^ ����)�g�����~M@�"�����Z��������Ս���?������ў�E-��3�����R�Y��"8*���w�U�'�Sf]�f	�'�c��}m3� ���JvGB�)�,eAd�y�ڞ>?�$�]�~��<3��7�h�#X��y��x�%T��%r[������%.���ͿNOHII)��Zmv�܏MP�� ��1���8�hbx���B@��דQ���؜��!�qX5���~�@�5�	�0�T���r�,Ar0y�z�{�c������SoK�]¢��)��J�b@�U ��3�3�k������8l³KcMo���5<�4t��-oW�AǨx�Q'W�~������'b���C�5�(<�&�&��A����[.V" �+TȌ��K�m��F���vrR�[5(�=�,乴P|(M*���&t�}p����賜�4cf}����d���sܵ����ꟲ7-ꂑN�By����ɧ<����8�hm%<���Vg���bT.?|9����#�y���}vC��t��� ���X�zv��됛lpON�&�`6�c� j�l��Ad���X��q�"v�W��33�L��6���6¶�����o6�8���:���\�3m	S�] 1X��Rۨ��H%���m(�'��v�\�l�(��w/��$��H��9M;i�]�'>ݮttt���M�_1�q.,�}�����;�W N�<Qs��\�u�N
l߲�g�|�w�]HOHH�^����������X��wmW�-�2�[`���0!A��0'����U�q6��-.SL+8~%�Q��i�z�v1G?�X�\]mɺ�C0D���	]��6���l��\�?�	���n	d�z����&.��n��$�3����h���բV��m��:�4�88D[Xj���9�?���H$��pg�)t~�-�Y��2U�����iP�4��b)�^�P���6`�*�_ͧ��t�D�]���������ꦨ�� ���rRrr��&�\� ��i��B�y����$'�����%�z�0���F���p� x�J��nƀ����^C�H"ݒ�O����Lp#�w�t�I(*��@��<�&�rK��i����yz¶�?6�# �Y�|�}&�Xɣ��2P���uQ�@��B&����`�R:��[ҜE��@��� ������J 	��iE�I�w�x�����]T;n��G�q$�����|���Vŧ����m�ϻ�J�
�b%��D9�<�%O1[�jJ������%	�bH�Ч���*Q"]�����43��{�{ƈ
�[�n�r�O�o:+��~`I�~�g�m�J�6c������_�T{7�������0{*�������w��_���VU1f $[Or��/&�����&Mm��p���=!㤂�U����ʭn��"���v�����p���J�\�V����拵���D>���'���K�JUQ������ô~�/{�h+�򡸎'�2�J}w
�$9�:�Wä4Wi�y�?_�\��0Z���&׀c@�?m&2�/S���oL�����X��[����q�#C�ɫ���;GȺO�E�v��*~%� �E��*>���C������+���=\`z���V�zn/�Mw�;7�0���z�^��X������'''�12>��%Z�i�2@���{��`ce�j�a�q�)dO��B�	ӂ#�M�� bp`ޭ��ڨ�݆�d��~����*�#/"a�VE|;�!�K���"#�LF�-d\31V)��Y��J��?�=�$ou�΍��g��
��� b���ֵ���$˔����d�(�����K��Yce,l��=h�N�J{��m8l�?�ȯc;~4�����A7����R�j��*,������N��|�XB�Uϝ���<��a�p���;�,NtpLT���8��%������"}���)�1z��ߐ�0E~M�2V�&��N��8����P��������]��}j�3��a�����|S��릲��/f)��9�"�V��2�����B�p'a{��>���՚_��x-#�P)�߅��q?�Kb��
���ֳ�ܨr�d�+7�yͥ�w�� |�_=��`���%����ӎ� �S�\h�Uw���̜��0���"��5Y�t��A�O�@�2ŕf�^?�e߽<KhX�������H����j;&���4P�����VD��t,����/����/"@��1L�S)I�D���W�K�d��5!_0ry���z,d�����XX%�o��|�3�EM����P����q:�V6z5@����^X�C^X1v�|(I�]�� ���=-�w=EQ`͏�.�����΍�o'9��\����59�,p���~�^4�Wq)�i;�����^��+��w�G����Ļ���M�!WA5��<�.E�9��pfgA��{5ǯ��K"��g����s����L���y�9�V����A��X�?#����JuH�%�T?���A����E���]�[}�݊��>�V!�6b���Sl���U�����>{/�&�_O}^�d���u�-����o����U�#���ޯ������z�� �UXŮD��*Of0s��UY�w��:,J�|�J�;�/_�V�;��M�����wW�|��bv���\�qP��s����N�_If,E��|��.ݸ��F^n�� �yǞh��&���;��gZ]��D
j�9�qr�91���9��E��DDD��D��W���MM�����o#�r�L�~D�;.XL@���JR�8�4���gJ��7�������K���ˣo�۹r�W%}������I�(��ߑa�>G,Ǿ��]W��O�?ۅ��;��X;�k�&}Hm���ԛ�͍��gW�4�����X\��I��L1h����*0&t"
ȉ~�:������~�?�W͵n���D��V�#����nFS�*��A����x�ިho������]�xR��N�2�~��Z�����rl�e7��Y�^�i6��O*��9�Z��kV���'E
�嗢q���9DV}a��dI[9@p����Y|������A_�
���b,j�-���HmYE��Nb#9�q�:�XK��/�����}r��b��Qbx������Y\e�}�V�XH�g���d�<�.�P��Cr��M:���۰0�n�Uj��=��$�-7�k��q�w|Ko1��-��	np������$�Y��J23��v���g=ož@��5Y���U]��3�oL���(`��d�cC����G�7�ȓ#'2�ͼ����^u��<�<BE�4 �6C�`���QL��MGl$f�:��ڥq�+]
�e�B����N���ܞ�!��Q�V����ǩJ�e�Q�M��E����3U��2 ��!��%2��[��50ǹ:wD��3�M2���Y�N��������aG&�-�Q2�]����\E��&>�Q���	>"O&@W���)�!��=⩋���YA�w��
��N2^���B=����r����"��n��b���<���l�^7�SzA�I�{�d��\l�Cy��?����t4 ��k�M-���4�N��\��@��S��tı��3M�%���Ѯ:P_O>�p'�ų�F-.��q�V�?�@�2V�^i�w���++��I-��?������Pk�%4Up��z�1}I�su���<}k��C�k�#f ���9�K�[��i3�������õ0R���"̮�oh������P�dU�{��F8�����˼N_b�+�RF~��(�Jڙ]��p7�ׂ�.:����D8��P'�hH�n�b���	Y��|O���;��$vZ��)w9��v�im��M��M���\�K��o�L�h
�����毐;S>#��N�9_f���֩�F���W2r�Щg��i����vv8���#܆N3����w��iq���Q���y��W�3kg���6�����25#�tK��0�g
�w��v�R6%���j�)�W��_�i���u� [����_Z��ezVVV�#p;[ �Չ��$�j�Oq�N���b}��/���~�rEs0Ic���G�"�Mz1��'C��n���>�!�9�qn�4]��M��G�W�
�օ��VqQ@�2M��jU�H^�
�nz�D~��Ue�W���ma�턋?�OdV���G���96�_&5��N�4cb
i���RW��XJO���8�)]f���6_߂�X����Jb��9X���x��h�L��#JQ��zQ���Fb1rQz��ӫf&�5�QX���-���z^H�WWYYi��Sȸ�&鹰���$�!9Qe��6uNW����ՖN�tkΆv4`�NZ�+��i">b������D��#A�U��S0���qj���iB�Iڽ�S��>��6��{1޾����#��n�J{��Y,�7���[v���x&eӽ��"��vK���W"/��noޔ���xM�mH��8�?�m���XL0;Pm�I�\5[9 �T;���+�����8ٳ��Y�j�)4Ր��>�cw�R;�y<�}ڂ���iim[%�Մ��\��-��\Tw�Bs�zY��.�]��.�1bQT!y�N��M�Ķ���>͒1�l�X"##��1m:��O��Jj�
���a|P&su�s����Mm���0�c�Wx�B|n9�?
��N����[�yyG58�8��� ش<m�6���I!�޳ev^�+/�p�e��o�+�d��2��f�O:����10�T�3�[��V���f��z�����Sߑ1�1ABN��ռ0i�͔ZF�Wa�l}a���cé�	�K��ō�Pφ�)a��z*����l[�E����n��W��t��˷����\\��3��N�~o�A��v�C�~�uئ��#�A�?ܑ�����͉�Ѱ�=�>ؒi���i�����@,��]��\���g���-g|��$!*��/8G
�n���O��n4Y�������ows���[��p�I��_��RE�U8�;���⣓	>�4mv�t� ���ST�8�H��,�%'w2F��73bu����2��-U�YWQ��nS ��rd]x7g�Q� .W��@e �剞�-]*VϬ徸���ξ����.Bmx��E�{	.p�/M�C��p'�Ҁ�敩�Y�>���l�Z����/�졑�ML�`)T�=h�!��E��#��Յϐw���lonx��u�\]]]Z����:�i�$��E�9װ���'�y��+��C̥�a2cجps~[7�gR����.���r-�)��P�z%9��t�Emʞ7N0xKw{��[MFf�T��Ѿ���8q���{��Gџ��=�<�6a�����?:�ީ�/7b��G}Ywpv<@�*���?��%�wyA����Iy���焥 2��N֩:�K��E�$;%Ħ ���]yS>X#�(�5�w���e��_v�=;tެ��C���%{�6�)��;��O!"	��\�޳q��X��>����������3��bp#�5��2!���|���{t��v�%�5?��k���󼎃���E
�u[ɴ}c��s3Ѧ���e�.S�>�d�,J��w t�*/SF����̯t�3���Љ�l�2	O��6�&Eow7�DN0�S��l,����nEO�l��f�������,Ũ̌�ʇA\���[slFd��ݾK����]?\h,�9�ue�_����4���=��
��)��:��>l�DHr����'��0���?�1FU�HMJ<DL���f�NQ���)SO��Y����3���zFr���5P�S��#{o���������n�\ �S[��酟�������o!����U�O[3���_ÌD�Hc�	��H&j�f�7�Z~v���K��dW�����u�-��u�9�?�7��!r�N��䖜}q ��O�c���c��Eؒ}P /Ru	�ڄ��o������V�A
�0����K�r�>���I
[����~��9fQ7�-�H���6 �]�D�wD����Kz��J��0���M"BBz��8�]6�J��ᶎ5H��d�Kg�ye���?��G��.�!�. �3Ŵ��SX��@�a��Q]U]�-.i�������_�)��w�9�_�2 2��?k��;���$�n�6(�xW��9�7K�Wex�D�� ��b�쾺��.9K܎�"xo�lZ�@^[�0��g_�	�v
��y��;s�x�T��BŢ��=n�7�5�A1�(D���=���%�=�_���W��"mX��c�80���2��9�)��M��� 8��y7e�f��a5����q�}�Ԁ��FU'��k�h���p��T���9��[5Pt��	8��tC���G��Ch~j!����z����뵆;��5'�l�R�wf����}϶�H�ߥ��i��~��k�q�|��b_�C[	����&\�Q��hHO�e���/9*��gةݿ�ث�Kj�l��dd�jXI��c��akW���`U��k��77T�`�ΗM�Xm\^�"��K�E���?W�R���v%����&~9f�o���� ����j�{�Ipi���xq�+VA�-�_q)���(P X�P�h����+�!���3���Cf��g�=gw��`w�"2�:Oj��a��W^a#�|����������dLRn_ B`6��1��>�vs�n<|oy�f�-����.��[u%�9:=�����H*������x򴙯�"�]���ǆ�:S�;���4J��`<)�?�Y!�hh�/�`���r��]|#�E�0�4=7�M���Σ-��Ct[�O��%�L�W�%���b��e�~._�H���e�;X+4���	���:���0h<}T���Bw����&��a�ހ��4TD���1����&���T��Vfnb�����}�g�%�*�e��R��F�伱@�C����A7r��!��R>q�Z��M_�uc���:1 ~�)�����ހY��֌�������;ҽK�~�	�������e�	���3�p�gZ�|Ew�S���ɺ;E�8������g�ߍ�4ծ~�w��P`t�ж;��`)���7���2턗�}4���� #9���BI1���	���^ǹ��\>Y���m��1Ԇ���tO��:HL8,���|&�������.Y�!�e�uק��U����5O�uR���M6����Vd�j
����C!�U Y��"�����H�0+!��%У�8f����ń�q��"�Yz����R6�#�l�`�z�D^�x��\��ֆs_���"x_���Vn�jջ��rZ]�A��8��V溈]��]�,m���8h�@z3*
-�W��=��:?-��W��#���{�&n�d]���M�i�� yM%��K=L*;��wY����(2����?MhA8X�5�w�  ��n��g�F���\`7G�z=M{1gG$�������M�3��qp����DЉ$=���J����گ���*�ċr�ﵓ��j�)e���t��NW�/}���k��!�O>kl�#C��yk�a�1���Kڪ4Bj�s�甏�(���d?�P ���af��}��\u�A�h�h�:��s �%Fkv��!ڤ���v�O���x��hZ��r�H&)---/#s�D�o�X���'�^�P���pqs���8�=�轝)�=؈U�y���yI�h��o����w|���n�?��{��%u隈hfz��:��oF_�XsS�H�����x^<�=���?)���^��iť�W\����v��od����>�n��A��f��-l?$�ؽO��5������"-���Wj?����U�6xL��pCP.v*�!3_�:a�ƨ�s���J�L�O����W	����3�w[\���k���F�䈰 Fe��H�����傲���>^2��M�q H�g�n(��24�ۜ�Szw���9�&�M��0GKf���Ŋ����C�|{_���t��( �J9��᫵��!�7q�C�O뜏��~R�ګ$�|�f^w���%�Ć��@��v�'��Co &�uߩ��>�Á��
�<1vd#������qzuZH$���a��
�p������zzx����4�ߔ�����9{���г�R���]��������W����;����d�P>!�C���#�N��Z��0��n끌m�4�ΰ�f��x�H�Gk[	A��H��L��شb��l�f
�Q�L$c��8���5�7[�P:���3][��WvA?ӟF�U0)��<���D)��_4�:%H|:%��]l��G��G:��g�$z����t:���H��f�Y��H���b���e��0W]Xk�V�4���|`_���}f�fnhd�rOXOS�:����7B�"�
��
׋/�8�1�h�T_{J�d�Ͽ�
����E��p�rͤ�v"�ޞl�,�SjI��F64ҕ� K�I9�gt`�Gp�p`>t�^:�x�Y���g�����6�zD��є	�~�C`���h_�М�#I���*
t^�ػHG1h����4pp7�o����E�d� B|>-��<��q$?&M��t��Q�a�H�֨�6�%e�[�Xm�?����`o X�6��.]3P��;�oF�^5��|�W�����?�>�-]�䛥�N]E���^�q�w�3|�e89GE/�4�̋���X�����k���uF�]i0փ�0u�[�m�by���l�$��[�Zߍ��a�u��ɨ �;ᚦ������3)Cl�M�OU��`�X�`�ߥ�\�����v��r�����!�h��7�]3� �F��z�>�_��_�5��
O�1����
�I���ͥ=H :284~W����(�>��G4r8�=���*����6�}ҟ�þ#}��D���s�\9pיּv�k4���ߓ��9m���Z��[�8�
~,&=}?����_*]���!�TW��+��W���2�����1�Sf_���̾�����7��=�-�W���+�MV<_�D�6��Ϳ�����l�^�N�#�C�L�����K��(�npM[+�?�3#��k}���8��O��>�،�s���/��'�:���~g;�蝆1Y�A��G�:Xo�0�jJf���^��8�h�E�W�{{�N4}�䛏H����;��^�?'�'٫�I�-|F��x��ψ�L�m{wd(p��Ń�N��%�ù!oe�����^|��U��h7��/�xr&���ͼw˴wx����ޣ�Bw��?�_'��⩘������~&� M �rΨ}K������b�w�H��3Ņ�*� [�αo�3@���"0�P�فӰ�V'`\�NВ;;� �=�V�J��N���H8O����/�}؛��~S���[���!f�t�Y�Ys9��<zDɫ&\�a)7�tCXF�AOj�'H�sS�'��D�=wJ�6��\T8#ND�벸���JS�l��cM��պ�����ީ�XO�?��\�V&�E�[�,\@�/�:CT�[����jЪ/.��Q�]#�$���*��G�[kɫ��G t���E�������/R��-@y-zia�͟" m�X�[o�n�z�,O�/H��ru	���1,�^`�\6�1��wD�
�����JMb,\����/�G!u��M??��;u��M�7Q�����������~�P[��U�
�Q!�kBO��:��ݺ<s���g�q��ٻ�Ǝ\�A⛲�����b�*-���=�|F�fg�֋�`�qx���N��^.���������P�H��6�L*��6�J��Z��:ͮC=l����@�ǳ
}�{����u2��*wN��G,YiɈ�E���[?!�2��l�ʮ_V:��K��Vh��+Y���
�|ּ�l]m;���#�n�|g�Wf����̡�FәޮL.��ޔ!���Ө�Jg=)!�ֻo_��jm�����x*���l	�c�yD��i��&��-i��!��}߂h���Q�dGg_.`��v�hE
��('$�=�%y	Kt ���a�?��h�$ڨ����trP�؉����<>�Ο�Z888&�����^���t���z�/`u�냣�Xӣ�V����oH��!#ݦ����ΎIƈ\s!�}��̂n�x?_l�t�!f�c�c�-R�������������̖��"��-�}��k��ݟ$t3���/5<�|ݘL(��%�w�j�Z1�)��Øs̆�&��a�K��j�rV��&�]);��tl����#%jf�/�A�2R�B�2��֏��-ّ��zkE�.3'�>
��(6���xKڿD�жl�Ϸr,�wUh�vx"Mt��ӂϚOwg��no�#�SK�����I�8�p�	�q�(r�ԆW�C�-1 �u>[{8�;�i��)�����{}�a����D˧�~��q�4������T�w���+V+ad����t,�/�dXӟ��hJ�9��+M�c'p<�Q���Â��߰bf��Ԫ���Z������o����Nu$������9�dL�$Kq7�a�g�r���2�Cǒw:s "��DuA3�V�����L�-�Mc
�@pg�����j��	?�L��9�=lw\nf+�ǁ�?�~�=����c��.����y������hl��3h���Q�5�5�_�;�Ʌ��菔��,��p�^������X�[?���vw�I~�,x��FL��9�z������H�L¥lA	Tᾗ��G{�(�a�Qq���"��+�ޝ��\�Y��ņ�'�R7ǣE@8�'� �ֶգ�9`ff���R���oɷ��Ez��� ��w�gC�ӓ-���������������#H"���Ljh?��=iaJ�n�q}��)�U�X���Z�7,���b蓼c���3c���b��W��~�JE\��f�A"��^��J���v'����F�U�Z�~��Nq��r5�5sj�<��s�����3�m��o2 ߄��`��\���,����F${��1�.�� 0K��6�TcM�H����|���Ȼ_���ڢ����<ؙ�@kUj\��7����s�h0��g�6��r��y���q�c�Η���8=Y�R�*�^�r���C���0���V� H�Ӻ�Yeee����'���I	����1h�r��ɲ_��Wط�WR���W�U%�0���hf�.�r���G�Nl~,i�I�7>�������َE8Kz���p;)�qbU�p�5�e^;��}���������C�� ��}�ː}�v���\[x�;���t���ǈ#�����������]��C̼0#�©���h�і-<�5E���t�j��N���wg��R+϶��5�P�N�4<�����M����!��}���]]:@�����7��z�' )�C"�Tׅ#�p�2{9^v�}��(����f�מ4��ts���B�l/��|��)9v�u�K��R�$dZ�~����hG�d��
 UNT�uܦ�� ��e��(��u��G�<+�A���9'��6_h���C��W����X^��UJ��th�[�L�b��oOֺ�ɼV��q`-=?�"f̌�H]�Ow���G P]�^�؆��e���/�"��� �,��<��^�`_./�8�����g��@x��C��@���r��/ǯ�|ej����
��s�$}#��m�%$'_��l�`��[�C���{������c���^�3ً�ZX�#ϔp�C߷���\��=�>\1�PCI�"�����k�i�ƅ������eucJ�����ce�{D��C8
t��׭��I�{��ӷ��*�I�Fvv�ѯ��Z�*�f%-�A�0:G]nKWY(� �����i)�� ��(�lf��tcS��p�q�XRւ�|����?I��[#���R���Gρ��#c�niv�
���L�� m"yg0��D�w̾�P�0���� Z��)���4ΰ��5�����I�z� 	�<��j�xP_�%��x�g<���iB���儻�J>=�JKOt�}zuy����A�9��Թ=��#�o=Q)��+�$����kp�����/11�Y7�8�c��=�>����Y�78�� �w����� '����Pd��*��KPQ U! 9��{���k��u���* �m�+S��NħfGh;ք�wRf\�k�!��w�W�C��$x_/����--��~u��zS��*�G��q�m��K^W���D��M�,����k���YE�6���>�
��}1�h��l������e���f������rA9���
��M0�R�,��0��t�W��|[�N�<�������?W>E����̬,����֠�ۛ+!74�M8S!��_�w�K��[�4��aɖ�8�<��u�}� ̈ Y�V�G���T��~s���?zw��	�{GC�_,�hB10&u$�RE�
�,���AR��3-B�ht�����SI���J�{h�oݴD�簦�4Jw�$I�ab|^Fc��c��=b[�O�E�.�������&9Kx�LVgO���SC|�"�V�Y��Ӡr#�Hr�I0��
��wZ��t�4ǅѓ�ɜ��h˟^z��JZo<v�^4��ׄ���Ue-�� rJ�@��d�A���Z�v��rsq=��MTw�EC��a�:�n�|Z��p_��iܭ��o��%I�\~�p#�Fz�(b%%̊z��-�]B�js�m=��q�/Ъo�m	YW�ұ'�ix�qr���/��E9�����ʆż�� 4%B��Y�]���1��y,w,9��!� f(.t01�D~fؖkwh�yy��߉�8����SY��'w�:|�<l�(��jQ��Y�"ZK���WH�AvХ�O�:֣5,�	�̼�X�A�>s�A�����
2Y�-Y�]�o$�֮�n�P�x~�W`W�d�;㋿3=�U8��z�������b���6-:��Ț��{��j�~�;/�� �A����ذR߯9茹�&�!���#���U7�w��x�?߼�?��=�d34kH�7�)�44|������ƽx/q�#�	�gM��`��)�����C#���x+\�u�����DUjOZq;=������3�5[�=�=|L���jM��P���z�����&�D/o�S��]a`�~��;���_�N��C"_���p=����8�澫��w�2��$-���|6n=�odE�/6�9.+e��}m#��O�|Ϡ ����"�|���-t Uo~�_�%�Mqm�3vp��}�x�W̙M��|��D�-N��b�"���/W�6�� �0�bY���d�D���_Fd�^�����I�w}��/�;;;�9_}A��Cj6�KQ�0#f�� �,�黿\�v�{�\�(v ,,X��E��R�{�pݓ@zs�pw3�p���ŸS_g8Ц3̎�_/,	�{����6��I�꒚:��ƹW϶����T���T�D���� b��;�v
ku]2��i [�� ���)Um��z�I��/����j�h�)�{�0`;fl=`L��=��H&0Z?�Һ�c�qn5�=���S�,nXk��W��z����t�1�m�ɪK��0����/B�X̳/b��M�&����AM��HSϤ�S��	�Nr�����斁�-5�wl9��O�j���A�<WI�����sQY����W�/?�&ڔ�;�[�S�h�7��"�?!�jo�Y:*�Zsj�&�sn�H\S�N�E�d�=m�������>=L����Ω�U�j���wLw\��jM:���)�&���fY�<���m�?Ue����ش�/��a�@���, �:��xf�y�I�?��$�	�&����@��
wl�s�W�����^���o,&��X�E�|����� u����gڗ�4�.{z/���~�?[���� ��٫�ra]�c�$h:��2%��JO�͸"w�r���"��RO�%Y[��"�)v\����(�t4/;�_�oe��jUE2+U�
�ȫ-�	�s��+b1yHœ�z�����c���7�h�SN�3��ۭ��F)g��_���GG�Ո��9�i=�IxSwSԬI�Dn'(�&���N�{ڼ�)�Q2�F�~H������(��"��ԓKi�]��A��D�����JU*����Qc@Ȗ�U�w*���Z4*Zޮ�%�_:��@������&	��A#�y.�5�͜ɞ�=����@w�'|xBih�kj*�Z�:M�j�_�ܗ^��7��.kT�G�A�yą�i�K *� �����dQ� AB������_���N��.1��=53.�rQ�Vv�j�=�I�7H�׷�.�O�0�c���2��m0��Cư���� Q��ۃ���
 ��������GI���&G}6o�r�t�bD\���'#��N�H4NJх����c�,J������l�������^$|���.�?t|�����]�u��AUjA���PZ���L�s��`"�x��(�����a��ik�ĵ�ιj�)�8<v��w��;ŁM�8�ă"wR[�.��܇"q��J��mZ;Q?�C;MQ����z?��AA��jȘ!T=r�w���7Q�W���N��:�8Ex�Kt7��V�cEP����CT�!0T+#q;X�X��C�>&8M���*4*>!���r��=���.�W�o��*@" �{�����@���\1o�7"���,�W�g��;e0X���n�k��6�ӓP��Y!j��ݦ�Q�&490�f�ʝϬvd4? �}�,qA�9���3yjL�9*bj�O�hBJWA=�����=;���1���5.�� �n���a�*���&���X���k-p�eӝ�kܝ�	�%��x��������pVd�"gW2��{�o�	S��~��\|d6O-�5Q`�ek�eι
���Y���vY/��z�G
w��?g����/�$���?X�񶪒y]�w'r#��qh+M$�x�^��&���1p?�OS.������ߨ�Qer)��O�|.��ނb<�]V�����G\������L�BR�L���y���}=���� �Lv�"��Ľ�:���u	��i��p~�#��v��%�z�ga���zu���n��F�V	�Z^MO�}B:$S�B����E�qVϊ�1G�HIhH�'j�!B �6�JRã����~�7��uch�X�u��wn ��W�5��%/�:�ϝ�G�M���Ћi3P�jK�N�/�>�M�%�!�6ɂ�v�c]Z�N�\�[�%*gx���z��Ή4�I3�o#�.�O�=*nփoV�:2�ɓ�ע�O+,T>T���ؙ�Xx��!�2�����FE� ,��<�����5p���32�.VJ^��$��.X�O��?�"�C)O"e�y�)�����q�:��=�Ƨ�^f��~;P	�iF��>� A�J�z�T�bc�	���x�fׯ{�]���_���q�Ӓ�t�a�����km��I@�^	�v�?uffo��W�'�'|~���5(14���z�L+~.�N�N {�4[�~���,�"��0ԍ�eEv$��r�飕���=#7H_�b�WD��!���V(>n��u�@�������O��E���R�}덡Pr_�Uhl�$@�w�K��ŕRZ�e��G��xV8�؄��8��I���R�K�H�<�
W�L*~����V1ys]�`����~� ��2V�eU�oyp��ܛ���,���x6-�}y��G�5l:�&Vb�{���F��Z���(V��ef��]�B�~�_����A
�y���<�u�Yd�"��&���f��u� N�KĹfAŁw6�>P��p����Bp�6)Q�=cX]�[�r��?{��AfY?Gt]V�ǲ�����=3���F�'��Cy*��EN
,k��O���1���e���o؅Or���J=�V���8F�o�=2�	���U�����;,����7V7-����8�L��ʜR��K���&�r�k~�y���=]������6j���1�"�h*�#\���k!�Y�1߅�}�k���|�='�ѧU���G�<��NIm|:��rjm��
rŌa�G���lL����W�Sn����m���p$C�GI�5#{�޾ߙ"g�>��v�-�}�Q�?2���/7�����i!��y����Ͽ/�	���'{���͊g~���k��/��-��O�s�#I�;rƔ����Y�I%Q�og��Dk,����x?wk��}Zq�"[������qj0���� �p2����!�"q���.��Qg<������~�'��ņ+�޿Θ,�).��*� K|���!;���U���ª1�G7A+2[�����lt)��2�kާG��t��nk|�YH,�I��BHI'�~�*;��AЙ�Q�>��~��A��j_��E�߉���߶Q��H������u�|���;�٧W���=<�=�h(��k��LQ��[F>7��Ṗ�4:l��ݰ�'��Ƨ].�M���{4/��)���Nyo[Q�����n#���/��z����������'��I-���q�R�M�	|�l�LPԈ>�Il-a]�� �g�ΈϿH>=f��C�@���C�M�7�i隸�[V��_������j���v�Dp	��}���>�Les7�/.��Y�J�z-ўy?��$�J|�����]u5#�P�M� �,w ��woD�p�3�a���5D����<�J';�!���؀������/G�|֯t���H�_�+�ق�d�A��3]�p5pr国t�	O��q��{�u����	��A|���N]ߊ;��GL�'����8�lЮ�_�@o�N���?sY|��إ�_�Z��J�����9#���u�.�V�r����/��L��3�1�;:V� H������#3s3�KBTX2����{�� y@S_$�)�:����?�ce��U��o�k��C���y)��G�Ҷ'��R�zūS�h>�<'������Op��I5:&�>k��ɳ�=DN)�4�!�[���/1����|ŎZ�2��f���k� ��A	 9p�t���-� ��퇠1MQgvM��Y���J�F-���
�l����wc�	T�W��|���/(+��n'�.-�%�~<��!���v���zۘLk�]xݩ9��VV�טY����e�Q6��<io�?�������c� ���Vn�Hݗ_X����M�{� ��z>G���&�G���>�3P]�z#%��'+^�i<"H	)RR�
-�Uzm���#T��x��ު�0ԢN�P�x孨I.T1F�OT�ОXD}�z9������Ԅ|�h}Q��9�W�5�d8��q�d3*�?ip�<L�r��,�Uy&������W��"�h�,��#H��|��U<�@PK��ݫ_���3.���4K���9�'�r�<|�� 2堃.Z��댝�
��(/���wP�z�>� |�Ђv~T�~�=8wR�D��&��Q=�C�QF$���O���S�nwdŅ�<kh�BK�A�,��DE�6���H�n!ſb�&l(*���{^f}��-*����N4݄�Ur�mQ�۴O� ��:(�yNp��{��M��U���p�r^�EF�3O�I^#c�J�M�ز�S��Z���}�g������r<C��Īlsxn\�=7ޏ@��Z� "z�qѕv�"�"�5��� '��`���B�1��
{�<Xr<��[3.r�l�oA�t�I���z�.�x��|b�����F'��B���nM�?��*����<�h�xh�N8\�=k��g�����e�[8�J��²"Q6�vl�S��eD����N:����Ɂf�kc����K,O���3���,d��3u��uؘ�и/���b��x�Ņ�qa��l��T��w����\�2�����ğY��¿�c5I�f%��MMwI�Gvf���6�T��uР_)�xƶ��������9�T7C�BC	���x��P�9�EnI�r�2���ːo�v,��ͼsGO�]�>�\�.�-oƷ��6=O��\��m������S3r�]2������MH�V �3�i��Oؗ��'�g?�'���F����Y���p�߮p+4���\��*jf߭�]��_��X���"<U�w6�A�v '�D��XnB�=G)mp-q�Y�'Ӆ�'��@�G�鿚���-����Ci����a2��� ���-<�e��3��-e�A9T�a�mN�$s�n�b�/�k����C�C��nG���^�7�zG�HU��.�Tt��l9k���������_�hVCVz]B������@��&�N�̪����˓�#e���'w����r��Ż�	�n�[o�C�gj��7�A��R��I�����g-u��maE��J�ް�+�GjR�K_?ַ�,<�Ħ�A4�X)���#��=�ϾMC�|D�_��/q��x�C���RB7wP��N�M�����3<9 �щ��BQ�*�������|��#~��Ҁ�eF8]���֤�)�z+o����x��I#}��[��$dI^x��N��@��E5\������Õ�&�lY�bn�r�_	-�A[EA?����|`�-\��(��̈́���r�*�g���=_�q���nO�ghh��BYg�(�5��+!^��ɸW����Q)�z-7�yn��A�EM�o%^5�TI(܊�qjH1�<^;Kb}�`�+�ƅ�7��43�vBa�`�\Q=X�B����V����U�tU'o0��؅��Q�>��7I�[%!-������:�lNAd
/�}���Ʈ���Q@-�Y��S*�r�����K\�9��G��{sW�Ti�:t$�]Oa�p��6�"���԰�8����p�ÑH��e���8�g�SE���G�.%�)c8�L�h,>;-)1�W�۞y���e�T�3��ku �-��O.���v���-��w�	��\L}�d��#��e��U�B35�C�W��B��)�/i�́ŉſ�|�"w�a�=؅��.��cX�Y��%EdC��� �\v�a�CКCaML�����>��g�=ɠH��yG�fܿ����r��=7���i�=�血}f ������[�j����7s�oVs�d�{h�����_1it3�K�Q�[��}�B���9�PO��]`�������k�"�t�<�b�ĵS�Q��r��cJٱ�Z�¬B��<��� 	�y��i��mr�q��x#���~�>f���(ϧՖ#�>����!8ݙk:;MJJ�,59��w�X������d������~����|�*�r��g��÷HaG(��J�`��(�a-�+�$���,&�y*���E!�t��I,օ�H���#�%?�T�z�ц
��ٔ�����ò�'�6�%AœI	5咼���Z�$__q ��|>l]h�+�3׷����!�,ua�H����f�H�����b^�c�����"���Ӷw���'�I�z`t��L�ۣ�G.��¼$��"܂h�=���x��E(�a���jF똬���d��h���M�D�β>X�
�=~A7��
�KΩ4�(�@�M��t:2�J��k�H3�8���D�T�i�ԅB�Ө��f�5僟��~��e�����ω�w�g�_�|͗�!h �kMdy�ޅ����ډ��1D����|��˪"ᰔkS����9��}��t��ob�T�ݽ/�$(ݟ�>��0�<�3�pt�*MPn���l�5���c��</�d�@ɹ��5�Rn�Ӳ�L��gS��ջ89��Uch��T�H=��/�+y/vq���5⮾�|����t�0���+(u��L9'99��h'����OLZڷK�$�}f�-M+��Z�O��N�2���9�����_�d��l�A�}�����
�}9@R��GF��l*}���!I D,	±��hS���<�1�O��홷D)܍�>�d����QS�9֮؍�|��1���=!khuO�TOgF�'Y��-8/�;��|.N�`��p�=������25���/�/�9t�*r.wE�d%��/=�� <������H%���n�2���_VO%���]O�o��o��G������Ƽ8~��h�d��L���9P�� ��/Y��C�����?{`��cy��Ǐ�Q�:')O�y�9��!�}K����B�|��צ���ƺK�9�����<tI*����Bnm	j�d�r�t� �:��_?,���,=~!��Kt����ח�	��O�+�X��F��Z$ B�9fZ���kJ ���Hj�r��;8o#h�à���|׳'������0{X�x�7k��E�T1T���YWXxyy��
`�͕����C22�,Pdܧ;����_��H���7Q�f��"�܌���cw�Ɵ��Za�Ph=�}S~(��������\�pcz�e�nr}��w��~�t��r�h��C�G�F�!FM�u��侻eyccCN.�0�F�E�`����Q�}�ո��|�H��]��U�F���J82უ�	�;����j��;��"�h���i6���~��q�&��O��wpc�|:Vj�B�nk��hC0��g�j�����ը�]��b=�U�7	l$=]5D��r5Ab{)l��e��f�.�a����� L��G�.#�u˨��f�!wp���O� ��P��" ۛ���9�l��V.|k9wݪ�ʉk6d�¹uLB��o�҇%�|�8��*���ѓXV<��(��v�G�~��F�i��6Ur�I ���u[Fp"3W���󹁎�?����-�/o��jЦ.���I�5w����F۩��N����a�<#����0Q���q`���<�n*�t&�0���%��kW4z1���ޣ���z���W�]��'����czڜ����9:::R�� �ќ�/����w��_���WS���>�ltvv����U��,���M�����4_��#�Ӟ���bbf���t�Ĭg;U����q$����b��{r K]1%��E�%,ĝ��7}p��aR���8��_�u�Kk��-��{Rd�׊ii?�<'$*8��!�@��?�C��xuч2����<]�V	���B�;`�6����f�4�S{:��d�ӰP��w��s��v1��};M������e�V�ܬ��t�[I�T�l\���s�Ny�B�R����y,#7J��KD�Y����g?�% �D�?�R�� ���+��������g/ ��b��0�;i�q���K���ƯR��U( ��]�<����,:��ج��S��s�/�^� �[2s�4�ϟ������!�#C�����B��i[t䴥ǈ���g�����Fsn��4������ʮ�tz�b~p�s{�߾a$f�����%%�MH�d��j8���)W��zStg��'ؾ;8���(��Y�Tb,��8�C�ՅlWj�h��Q ���`���2>6�% �Gz+�*��n02��47f�L����!�����\�t������Fui>�0�����AuuѬ�V�3m���3��#�g��-(j6D���	ZKa�@��c��c��	#U��U�T#99��t��9s�u0œN���;�Ľ���x�|K���p�����w�6Xq��g��YD?qc���gܝ����O#�u���psS��Qs�#`�rX�y��r�'�'m#�s͚�
8��aA䈜o��oެ�s�&((�,����$�\O�qЋO,��G-0�-�7�5��C-�7B�C���ӱ� �ܯ�A�%}��� Q����H���	�	�`���W�_?0�g� 2�O$A5�P�JE���H��o�n(�� U�!�F��ƼR��g|3������5����=x���|F��\�~ ���W�%�M~�N�W����}9��?*�+2��>�B	;28��Uz r?��}�O����\�(F�P	��j�q;tw�Pd4ܭJSFީ�:�
����b~�d�S�4��,ѷ�DjÔL�4����]�m|5�وM^=�>���L�uS�f�a�A�����G2��}���?JDqU3B�ckE�M;Sz�b(d��f��K��K�u �H�?	
�J�Y��"O��s����=d&lp�G�nL�L�d)��Fk&N�+�a9c�q��2K�}��Ů0�q�\�ГϹ�� �ܺ�P1 l����]X�	�~0�ƚp����X�&�����x���!W��s�;��eP�-{�{�NV��n�(�����V*S��1(+���%�a��ܺ���`ni����[C$������G���T�����?�Y�*@��Pc��'�`��RԀ �`���}�9�ݒ��ק�e�ٱ�c�M�X�ysD �		������ϙPj��?c�]ZnP�-�[
��g	�¿�����G���;�y��䠡���l��{M s%�&�gV�"��d5�"��5�H�@?��ĳ���q��t��:�x4��3�柇�20�մf�Ff5k)������ �B�偸�$��&�@�q�D�{6J؏d�[��i���F� l��ؠ Wɤ�v��}��:����ge�1d(�l��L[|2����}��b!?��S��$��ϕdM�40278�8����D=��~BJV�'q����j��!�u�(U��4huH⠗�T���8A>�&3D<t��e���eN;y��^7��~���q�Lv��[�k��o{Se��pJ:i���ɔ:B$�j�9x��^Q��#4W=��Fw�Ɯ��0������y��o2A�}�k���e�q翳р�b���p����0�ۢѩI�=�-t_��������'�<�Ű�K��D��I�O���{��g����5a�@NXW�S�yρ�pp+�p@�ٰAb ���q�� ��G���9� [��R'3��Oc��8�������j�lrK;�Ph�D�ڎ�����I7�R�?Ȇ���sEޙ����w���#�n:`���'�- 0��`�b�c�*5�Y+`�
�2��@^a�d�������9�x���h�ʀ(�`��ei��	�Υ�K锖���TR�X���a���n��;��?���\s��3א
��T�m��-a�H������`%S��a���iɩ3�;9�lR_����Wj\_;��p9?�.G/�T^�[��؝�l�����)W�e���\l�*}�V�u��S�S��m�}��G�k�Ǫ�`N��J�5����O�Ur�j�I���|����V��B9��7��0�gY��ú	�| �0T��2\���r�ų�c'�6��k�5:q*.ֈL1����~�Yv����Z��C�2y�Q�����x�68ù/�d���P�/TO0��Ǩ�Y�A���%Z���C.G ��L�67p�l`?��;�|�^�����=/8e'41 �첡;�`:j�b�H��]�zJ�{�>lC� G�
p�K���')�:��!_iEú�b��� ��Ʒ�I*�b����Ͱ.S�_�J���&:��y��ֲ�ln�L %\�dK;팠xTe,���w��G�	�5���^MJ�MY�H��yZ��nU����l�n����|�(xTUNR!Νv��G�,x�A�;�}��zT�Y���D�(��;T����
Y�5�`���)6�6��lh��tlSg�!®�؆'�x��ú��I��Lk;�M�����
�U
̐&� m�?���J_T�����Eڙ������)^�ǘh�Y��_�Pߓ1�]�|{.�(^���C?|��a}C���4�[$/�'t�4��ləv���mũ�	=%r�`a`�PHt�����yG�F�!�^nnd��&S��!~*!�z�X����sԐ�T��C�8/?�i(u�~㱢k�G+^�.�z��,oP������ ����qQ�eCϲ�\�D��`�y�����c��3��ϗW�$��`2Yc~���x�B�)G^�.�7$)L�SnxZyX�ۄK�B{���o�DB!@�,x���.��a��ყ)�-�.z��%�;�.���f`m���=�	�m�f�=�����Y�˙�E�:�3�`�2N	�>6hK�~��kP7��\y�[v�u��oe�Ŝ�P�r�֟+|���,�b�C81|��l�h$��kή���ߏ���UJ�ɟ��g+~�$ٓ�����q���D�	�S�?-)��_A-�ǫ�

�����	!U�"�T�Mn��U�o�Q_���_|E��N�f�a�)�s ��(���Cޢ��b',a���ѓ'Q��Ě�S��	0��$Vs�^d��fS��[ ��Q����~���3���y�q��`���ɼ_��JCO��h����e5^9���j��\詻ı�xi������u��yB92S}[��:�.������I~�w6��ӎh8M��e1���:���q����9D�$�Á�Р�0r�)*e-*6ÇEd`����ww�)��<���.��%סHa�U\:�J{�l-L#���5��0�4��%>��\0*O1\�ZC!cr{F�)��\�~+���L�Άg)��d�eA��1�Ⱂ`�m�ݨ��X��g�� Ӹ�;�C��� O�?!d�܆u{�ޗ�o֎?�.
Bm��Yyր���,5J9L��EGG���Y�,c� �k��kٲ07��|��͆���&!~�T�u��Y૆��/k��$X�Hΐ]֩M�!��O���0p��k�ьoxk��¦nr�����i^cH�;zoh�����������y�+�9�pW�ݺORr�N���ц���l3���g��Ț��mWq�"�	�c�}���nc���V���'��QE�ܴN��Ó�&_@�8��_�ы$TL$�b�K�/��W_Q�Q��S�2	��T<�A� �����%K(��k��YGȓ��`�|�X����K��q��m���oT�G3l6g�z'�T�^�xHT�o.{G �g�G��`���3 _
�$����R�l�3���{�9_�D��;��t�SW�V�6��OtT��M��{�ޡ�࡫k$�����ߑ-�����C�a���I񠸫W��T ?��:� O �x��8��K���5��`�;��PR8�p⬩SN�&wTY�M�۳�nCu
��H ls�݅�W������&��4�s�4Y�2�F(��������Ɔ���9S��G4��� $�R��7�ͱ�!s��$q�}S���,��+�Q��h%���q�vtm��;�������%��P.P�b��B��uK�h���(t�m�'������y�{qd�V\>��o�����n+IŶ�>�����7�'�)��Ck���:}DY�m�%�P\x��?ၓq�w���1�&�pNremm��~Ɨ��g�|\��.��>Քr�;k�Sv&�i^]�����I�(πRek��sƄ�ʠ���s���f36hž(�j2�]���5��	"��}pO� ��s�f�E��?}'''�DASr-9���MQP�Fx��y7�	X�-����'��S�'�2?��\2��I޺�͸���Z�9�����d���w@h�Q��4CՑX*��-��ݦ�8�Av�5�s��"*�"�9�]�(X�=�G��{����8�̓�@,��:���v3<����x8����{%f.LV���x�����8Y]�QRs�{0��^uz��ӁЌe����@��/��F5��d�G2�
�3���ń���V�͏��{ߥ̌7�߲E:�kՅ�7C�&��oX��
>'����ߝ����3!����")���x��W1z�<�:�0�"o���L5��FO�J%��$A#�{LZ��e�_��u���'�~��|(⶙��z�F�h۸�ѠsZ���:�Ig�?��p)�*�.CȔN�t�����ȗ.z"b�%��&�<Hy��Ж� ���$b�ړ�����8=��<'T�����71����{�i}J^F!��K���0|e����S���@�0�(�gN��p�fG�2���Q�@dC,g��A>�Y�}Y�0�N�63�v[H<|砍��*J��C� ��8M�%~n�b�d�Be\�9؀��� �_R��d� &a|�N#��\7a��̴�s�E����voz�(���e��!o�pk�~F�jS~���x��Hw1ߋ�4��p)���V���$���3�fq�=Q�N��S�	�"�X�p��9��c{=͌,�[5*-5t��ACD'4�ו1f%AO���h���c\�O�¸�>Kg�B3�k������n�ʢ{����6x"m&�h������j�o�ԭ��~ �|��@�H�c�� �8X|ʓ��B�}RQ~�F�1v�A�5K�}tqX=�����呪��Uy%�7Sn��m#2�;�m_�Tx"���f�Ӓ�Q0��3�0W���x�jq��a��#�f�_D���1����l��m�nI3��z1�������1D�r�|���0��_��0�����+����0��kL���"v�'86�G�m�K�{7G��N���&]�vA�2��k!��j� �%������|��[_���9����V�T�-��	�S�M���RZ�����f/_��mti��X�8Q���x95�s�)�������P��$����J����EM8?��^t������x����]o��'<�6%H��tUI��,�������ϭ�lΌ���QjR���A�*GUM7�+LBH�9��4�2�^������g��H�C�p��T��`h�naSN���H ����5�@k����ˇ���{�������,�O���&%*��	<XH�=jC��)n݃�h
$KKu��O��LcD6��:{72��Ge�u��ɲm<�bC��w`�rߔD�C8joA�hi�x�Ac�q���a���Ǌ����*��ʳ9��P)���ɀU㯉
��T�u@JN�P�x�� %q&��Jk��{��&�t{��kN�Zsc��|1c�쓯��~�:^f�~W��cs6S�]�(Xr���gL�q\�ٶvZ��}��i��G�76'�<���-�G	���
��C��+C������64��~%9;Wf
��M�����E_|���o�J���ʮf�۷y�ZF�����#M�%{�>r��P:����WMd\T?1F���>Y�_��w���j�7���0��r��p^8���=poB�@4����ꡊ��Q����ff:�w�څ����fzQ1�����1��=ק�?1�Yj�^����XWW����m��f����k����s����ִ���/�Qb���p�>��gƄ=x\�$� A��ʪ�=<7f�&ݺU}vqf-�-��쇸e�J��Գ���������9OP����uy���]U��a�ƌ��c�]5"""��v�k�DH�󣔜K�y:{h9� �^�
�L��2�f�U��[P��"!�r��x?�m����xm�ȺB�;�m��,��_X�A63:l�<�(5�ɂU.����{��R��ݭ������?\U�!e�����@m��Sl�$�C6w��j@~�_|�l0��;E��(���}â��L�J;��7t?�$F8�T��6Eǧ��G!��=�1i��V�/
32���.U�����d`4�߷d���P���]�8�|P�V1T|�[c�R� �������s��T��~v����?P�;���Lv>.����� �,�w��!

��	�U�&���$o��T���K�%��� �7+�6�����=�߲n�8�����f��ј��o�e�A}DO��!a6�
�|(m#�WvGF��Mے��۷�	6D�=��q揔�����.���"���@�Ǜ����\) ��"�'yd�[����{����*��膷�����'Yy����/�+ǁץm�Г�� ;Й�Q����xZ:�b՟�7��YO"�~E�h�$U���p��S���݋��R&(��n��寲N-�G*V;�'A`R2�
k�p�4��M�,ն��"� �v�#�O:.5��a)��&5% u@�&�W�ɩ��0J!���V��y5��[gL��'�C���(�LÏ�bl�^�f:&6��~#.����Ӎ�m���[	̐��@�d�Q��DCʄ=7��
/�v����Ӊ��6��F?����Ջ�a�e��}�7��E�l�+!�s�� ��<s b�w��I�d��M��H{��r�.CP;D&��O����0�ő���iW,hg���|�nI�GN�Ӯ���/�}��$�j��.F���T��ӫ����S��X,P6,�^�P�L����4�#=4�����ė���b�?�a:\o�΀�K�t��:�$��ݷ�x��_4.DF��e<N���8˰؛�n���%�I�u聨g	�X٬���1�8���i����a���rƈ:N^�}s���u�w���j��x�,=����===����C�u�6"�+&/�Qc^��V��Loo*�wbh�w���yf\|���+�Ά~��p4��?bO&�R�9���n"a���M�4�8���I�p�<�D�-P�㖅gZ�6�cz*�Q���a�8��l��x��{nE�>�mHHX�RU�K�G5�Y�Tv�1}bߓD�)���o"��׫�B�����3��u;��F�ݤMD/K�1:��[�	ޮ~M����%H�,U��4qV�পLm�� �}]J1���$�`P���kHj����lZ��W�P��	`�Uy�=�����D�6�. ��7�P�o5D��~C{�v��P�'�xs6I~�4�W�_b�W	��̾d�֚�&����Q�`�mm�>/��Bw�":(��'a�Z�`K,�LܒKg@���J�Ü��lЖZ�����%�!)��G)j������b��η���h��)ؽ3�	����E�p��F;��+���&V�XM��>�-����+\�To� �;����}x�X��AQ��˖���'�ξ��٧�>��F�v(��=^2:}�z95�~$Q%}L���G)��g/G/�9��]�Ыï�^4�(hr�?A�P��5'�������\[�X-�Kr&0swb��a����\�����zoZ�a�"��i	���Y�,VqD��]�կ %�a[4W��_�t֒)&�n+��$�)�L�E�<S�Z͇��[g�2� l�zXjE:Q���>Y�n�{����2.���B�؀�e����<��Cz���T�u�+7�f�}r�]͂nH虡2z���Ҭ��|��p���ouu�}�'��gYL��!�p�ٽ�R�L�1�.����&�%�t5�u ���b���0;�w�;���`s��uOU|�/߿?�6�b�j���}��h�� 9�8m9w���hz������`��ɾ�b6�ۈ�wyx;h��8U/GsS��2ӤvxcK�����&��N�h�,��mq;��EtPc�Ȁ&�JO������)�Ȳ�3n�iKv��7�\<vs����]��p`:��7J�߃�0��E_�E)_+^7�y܍� ̈́�o��|:�;������O�]�T���2���a��V��S�����h�]|�f����@.�'&&��׏h�����MZ�4 PW�`�B/�I�d����'��:w��2�k]�|����Ʀ�a�d����0����4�ƻo�2�=��w�$����^W_k�#���n,`���~$@O�H �ӧ:�����J��6k���d��^6'ԃ��*&�ϼ�}b��t��lJL�4X%
�t��e=7b�����(�u;ؾ�G*K�+?|�K�.YK̗r��� �X��q�!�ߔ|�}Z���)�#���,o��!��cRܱ���03!K�(����@CN�]$~�_
�V�4�S
~�SA�Mq�M���m�Xő�ց�Z���b�E�G�4+��mz�&҃��3%����4���/ڦn~>>e���m����t�(=}�&����}Ч�[3~��6�l�����.���8��7qdr��b��	G��&��~�;]�E�
-�V�Gӌ��S��U�46N�H������'Z���Ɣ_�T),,`+,��n�ڥ��ȪW��М�֒�yc�Ճ����ьc�i��q�TS��)��:P�!�P��*���mi��ܓ;�l7o�����9�,lQ�Wdz-!pSzI�zB(�t@F ���״��T9�X����:4I�v�lb�J)�����{�W���+��|p5�+���o?��aS���>3�O�2��A	
�z��/��ؼoe�{FY����ѲNټ���58�/�@l��mT]<H&K����y����vbl�A����|z-�c�յ�m�9���?ٖ�~�?�L�+�G�&�����1���@���������ì�[�T^��������^���N��ů�n�i�<����4m*���b��,��;�W���G%h�6��a��V����'��ڈ��Mޫ(Q����Fe�+��V�<ҏ#�'��Cvt����9��6,�\�V�զ���ܪ2͝��)%0+4c,��K#���;�x��)��Lk��R1:�o]\��d�opss~����_���3��VE3�!�o/�o�-5�=<,()���;�ӕ�A��}��?�+�O4�����W�ν��T��L���A|�}O맖��U�w���ZTt���g]��wW��x�<:X�� ��'b�{�t1��v�q�~�zss323�!nz���V-�w�>ɦ)�9J���%&��aB��o��X>��i]��n�G�I2��/)�	�Y:�0�A^�A�1���6�I�۝+߯�7�z���Ɋ�>��)��c��1���N�Ev�;���>r;����^�/.�	p�v��FỼI+�'��u�d������4<�3����F�&�DJ�t�� �u�){���t�}킼���p�y��ѐ�T��{�c�R��n|�����N�q�&( ��lEx�����ZE�>�85�vX�3�����i�y(�F�b�F�R��j�2./�\K�����_��N>ԙ8�n�˯�܊�	�G���>�$r5�3A�(l��z��4^/w��`�����=f�RL�V����~1�jb��Cx4���� &7���MZ7Vi��^
�Ԥ���l��N� ��/L�ʑ��<��U���m��	.NN�.D�f�y��TM�	r�hI��
�gư��"`�+
ҜЏ�^Be� (��K���۟��\��<���N��ֈ��9��/�v۝�����.��C*ਓ���v%����lj[8	ϒ�0 ��Y�gQ�G��� ���
 ��o�(mˤ����%r��}H���iS�"�q�J��GZ��G�(���O�.[���z��W�Z;�
�,��Ŀ�MF�J�/�{�;j�I��vY�#�����Rc�abl�U��r�00�x;��n��m�~H�Rj#ܭlI�\�?U�:��a,M���Ԣ0�
�CE~���eCHs�Ѓ]�s�\��u{(9�@b�@����N�o���R��^a�b>��܄��ځ�	����k�����������������
����.$Q�M��3e��X0"�I������c�ϛ�&�Q� C��|O��)��>s;������9�l/���6�л�9}s�#�o�����Jā|[?�Pl�t��
��.%Z�R��i	��Bj����_�+H�7ŀ"��[N�L�o�B�s�f:#���Z[��8�X4+'� ̭ޖ���w�v��H$��Im�Nw$Y�uܓ%�"� x�W"�
���T<�[�3���W>���K�L*�m6��u�6:�Ę�K@��.�l��b��ׂ��}�wۦI��KG<�\���<_�m��p�s�.e�B�WE9�v��d�O�a�'��M� ��%q���>�*�k���i���9�������02�1��k睡l L����Zd��Q��٤	����WȭF��`����6��D>�&�5}���%�iL�oqʯ:��<\���lY�e��e�a>+�M����2��yϾ�5[������A��g�d�]�5��İct�ｚgYg�9Aw�[D��Ɣ�~�1liO��F3��%����1���3��̄;��@aK�K�����){Ơ6�"S�{:����6��jN��룕�����e����/��ȷ��Tt(��w�]Vx����qY~�JW@0��KF�Q�GL��Qk��n��T���t� �{	�������-�$E��s\0�/��p����^�o��C9+������,����Z�;��ASIQ�|��0L�P�����L%Q���uov�����^n$׏�O��o���.2�!d#2�=��^:Rx�#��үǈ{���BQ�K�'�X�է9+{p�0���_s���M`�\4Y3��}�شb�)�1����9�?�%[7��Q��䗚�]�9��+-h��-�-�vB���0���s��~��9n~'p��Ize\|�.�~�85+�:�]��󢯧�繌��m���(��+ 1ĨG��c������c����+�Ŧ�@8Z��=���V�~Ω�Aw�e8�!��g�m|�)g��涁� �O�*�F6� +��Ɨ�\{�]�\�� )P¹������91��dL�O|+D�#z��Ʒc����R�_�w>K�G<��>6��(�Kx��}��UJ�2������W^�U���J|:��T'��	ײ�}��u���	�;��Dݥ���w�ϻ��/\'B�w�xA-8��A�1������Vg����K�[��T{I�w%j�:Ao��
U �)^������耡��,~j�5�2w�E B����g�W���P�︻�����6�]M�������/qX'�A�ذ�^���2��-�����cEq�i*����rI�����L�Y��Q^ĉʪ��>�Qi��(��v�˲B���A6���2�3�Խ���vd1����'��dl;(\B�br��@�eNC��`�6�K0=���4�����V7X��˯l��-ڿx)e����k�Ӯ�q <P���yGL�C�Yy��"3����8ҿ�!d��M���1�G},W���zB��O�k���e"ˑ��`	=��C�P�8x���>Qї����o "�1!�׋��Sk������b=A�[� W��+V��dI��r���=���C��p#5o7;pH�p/���U��UVW�����'�oқ���8K��b;�׈N&䠥{T-�V�*�[_�؉6�P���������0nPa���4:��:HIdfN	��c�Ng�E6���?,	a�2eR��DG<1���-+�.����6㱇���
i��ܯx^��+Ҧu~��6xYj�^�ϱ�/��'�X����H@*�1&B�-�[8�,>����2���Su�ũ��y.Y����XX�*���!����Ra�e%��fp��44�ɜ:u��\Cq8�"�Mh�YߛΨ��XH|���$ غ�"�;�E���@���|q2H���1q�_��Mt�*X���0�G��iP^ݜɨ��Ϙ�
x:.~:���N^� ����E9r�-��v������"	�y���8�;C�G%�\ )�:��2X
X.�*��w�Er;��ߗ�+-K�.;��R�Ң�ik��#�����kܠ1�e*7,]����qea�k�w���+{p;S��!q93rP��0�<�u}�0-�B�I���w�����=Q�'�����l�u"���*W&4��Y��_z{�o13��Y��-��^�1{��4�n&XȮcf�Q��D]�uO����ÎV�TP��n7�+��_E��W�>�e|*Ia)�#�W��7 0Q��]�b�lݸ0|iR��&�c�y�p���lsW�6�$��Ȁx3'՝�,��Hutq����?��Hɩ!�m�.E����KS3�$0�'g홋�,�+���vi�2F�s�p�hW@��4�g5>Y�-"�]0X��W��>N{���"��[h����	������e�H�Q?G�D:���a���C�M��{�����M�)�Lo�/-�����>no/�������WVs��\VS�asKK��d���ע���0p�����wZ�+y��;��+�� ˣY�5�������/�%$��&��b�}�u7!c~��ns�G)�E���Y�&���q)w�D�A>��7�(*�G�N3�� ��4�	�"�Z���:�K���՛(Jӫ��h��|�oۤ9ư�|�o�u������[��ٲb��1��-xƊ��>2	�ܥ
�5#~���\��n0�%ꜰ��_��|�}��۾!��Mv/,�>^��e������x���2a�Gƚ4Nف�:����%�%̒鸑���˱3dF�n2w�"��=��d���I�߳�6�NO���,�����f}����w����6��x���U�~Fd��'[�j����*�@����6���&"Y�'"��zK�U����$�W����k�.� ���"M��x�Z�&���T��n~:v��,U2�U�����BBrp���X���Ng��5�f�~�j�ܿI	�%���k.ʄe|�]���h�p���&���{�[�O$������S?'��~�O���r'�垮�S����� ��KG��0��ny64�.}�'2
��'���۶�]u�oY����&��˃��ݞ.��[���O��+�Ɂ���Г$=KAN7�h㌻D��j���~�
�V��	����u{UY����I��DD> �v����e7Gw�x���jL�:aB	/�`��X��*�������9�$����9P�����y��\��� �_>��e�8prrr���m�|_^֙


�q�-�ٮ�5�]�	�t�mo�0LrOg�jo	�đ�T�����cY��t��(�}���ϷVJ������d�C?T�p>�'a8l�[G�cBob��k\^{+hZROh����`8S�N��O󁿃�Q��M��R1s�c����E0�Be�ޝ|w�-,_�e�+dmR�5/�'$�j[�H��S��������ni�)�%�Z�8�!L��j���.�N�; 2;�,��^w�ӖB�a�	������]M��\�<g~�^^�J�+���5�Ђo��n5����o%hp��%c@]1��DҘ[E�[�k��l�bb-nNB��tX�D<��̭a��e�I�O���K|YK���{�
�������$�[���;vrR\{4h�M%�z�K1�(�N�"?׏�J�1 �%��д���Pk�Ңc�1����ő�5�UE��� ]#��q�_�G��\��������a�R��)���߰��tvW���,2��S�� �Ж�l"�c���~f��ܨK*�G	���&m��1=!�EI_L�z2I���e���u��C�D �F�l��M��#���yV���LmL�	���&�{>�bb������fs�r���	E L<���%g�'�A2'q6��5"��!l�'qA���3D� �*k"n�O6�l
bjQmm�&��;s��f�1�G&�v�ȸ�ȼ,!�8��NBAr���|6?3�Bj���|�{���?˽�� wK���SG$;	�i�B��+L����C��ӇC�w���a���u�F�=I%T>�|)�uCO�A9��YR6+��J|���ؽ�^&$lq�2�J9n.�	���w��������o2{��~�ڍ��ú��5�u���/֯p_�������������Ln���L���u��R����z�#�}��]�,��[����e�w�o#�&&����zT�*E�O_-0+�@�W}vs�L}�]��S�0����?Ѹ�B"HIU9���| (� �2H"ʂ���:�D��D_*�^IfPIE}�&��,����2tٷ��DjiED.�i�"�=��E��"C0/5��_�& #��ڼ�]ȡ2�;FBK�),C?GG_M&2v��h���O'9�n.=l���$ߛ�{ҝ�?&�}{.�x8i��D���^@5�į����S!�~ߕ�;ޜ^x3c���9��59�*�Q��+)�&עu��M�����[�g�k�]�Î���Ms)
V^<=U���?�:o���*��5ݗ6�l�7Z� K퀣�G����7Ŏ�?[������\@\<W�Z[Ź[>����0��y���J�0��=�N1�k]�w�g�]|��S)���%[A�h7���� �	NFm�P��yQq���E�+(�>՛�O\�r�/h�ɂ�p�ֆ�{����S����#���2������T�9�S��v������c*��ҋ��_g����r�OiX��`'or x�?#rRmX�����t9�95r���BR�:C�#�Y�w�j�$ܝ�sv7��Qj۾�mH����Q��[lu��!@��V� ^�;��#�խ �w݌�@�e��H�j�/4����'�xž�&+�n�e�]4giS愥�vB*,��,�{���oD�}�#!����h���-��� hH�jI��U�����=�]���:4�\͒g%s>��u��n�{��ѿI���݈Wr �Qu��l��̶�H���y/J* �+� /)"����z҂�u�d������ձ*	�����}'��WJ����}���*j�V��+ קu�m�hW�-�ay7��@u*��ڎ�X�!��	�q5)�7�S�M|�@�H~L��ʅbU��	�9].�EH^0��e��_�)#,U	�Q�Wu��ơK�!/0߻���ғ�f%��xN����>�M���-[��K(��� ާ��A�{�U<�<��e�}�ױ=~8�-����D���hr�o�����w,C}��LI^A$���Ԣ)I��]Y�ڄ`q�̕�Z�����؇���@�x��mc���ǭ��NI˾(3�9�dx����]_��V9Jb�r���w돡����hQ�E$(s���
ې�`�#6�3iþ��K�2�p�B�t��* ��xq�9��zc�h�_��c�r��!��~نo��y���Sck��&�0\��k�7w�Uta����_�q2#,�#�L���V�R�#s����Z��o&6�
��[��# ��)����᪘��8��(X�Ld�-
��E�	n���
T�֜	�(G��� C�p7�/�{;����z~�,��tG;��ua|�֤U*�:���_
�6�X*:7�&޳���H��vM�zd��z���_AM|��QU;��~�~μ/+A�w�{���+1ړ�������iX�7X�W�_~A�l�� ���$���'�s/����N��|�O�*l4���\_���I���b�8�� ��W�R��7	h��'u�/Rp^!^�aSV_���v}�Q���C3�P��rD��<o�A���z�m�[ޘ��½�8U�B�&��2�P?���^���:d��+
����rUe�����.������;���G��n���eOYڤ��!�9����	�gu����`�A���R�"̘�5�?�n��	��(�n+�)�z5��©O�産sJk��id���߸w��kC�G�g�a\z�T�y¹"�_��E�c��<G�bt$c�������+Y�bA[?�0)/�����#�2��fuYz�,�l�P��f��dn���˃9:v�$r�±R:��zM����� �����%3򔜙ױ��t~6im�������6�i��7d�CtS�^p@a� �ٓ���*y������H��JoV��z_z�������[
 ��©1ZKv@��s%�@
�}����R!u��0a�
�N_���;j�q���B�&6�A��S9�)w�S6�&��x�����T��Yl��
�ӗH��֧�<H�SJ��[��蚂<���l���pl����ώ������q߃E��pf
u��F1�)U}> ������2���jc� G���6[��IKJ������#�f��^�Gϭ��Y�K�e��`f��N��۳c��� ���ˈNL̨�����y��)"2~�
{���3��X	�� ��S��趤�M*O��NCʁ��qU;�'8��6�Ѱp��hw�My��2�A��J-[��o�{Eή:�DS�L�ҟ�0�e$M<���<�n Z���K�OＥ�m;c7�:5�Z�q�$\�����xv����Wru�l��L��݌���<�Y6���77�xS�����dZ�B����1���Q~��d/�X�[Y����d`ն�{C>x�/䶀�3c ��كb� /�2�J-�&�nJ|�?��(s�nP�K�5oqp�Y�a��0�-�*�~�%�co;�,p�O�/�3�٭1��ʌ�W��P�g'��a�V��2U @�?PL�&�rK6E��y�tCЧ����y�i��Ȝ��/d�Cnj��D�8��Ud�6�Q���ZU]c�����FZI�E<�j`���O"�����/�'&�����=��|���ك�����*����J	��r���Y��?-�+
�6�F؆r�TB���(��SW��||�h��P�T���l� ���#0�p�opv��T}�-@�+x��aЧ����l�G�f��qUwE����'�K���c\�.$<4Il���n�H�=�'R<Z����42Z����}�;h)8X�;0UI��)ǈ��>%+*G�G�P�8.'���~k8MUcJݼ� 8i"cѼ����e�ʪjU���&�18��"�w\��Nh��܏����"֣	��DK-�)�a �_�L�H-m�Xp�}w�W��I�隷�d����Ыj5��с.C��D�mF����m��Ƅ��S*��R+�;��!��;Cy���D�o?�j��p_�BT㣟�����Rrl_�&�~��̩Xޔ����D'����$)syX��q|��n]��X�8����,��>�`Ԑ���JD �hr��v�c��M��������u�:��.�ֻ�a�5n�;w��:=�[�#xr�l$�b��tޯ���z���J�P<�d{E��p��:i�S�)C��0)I����2��W�����n���֯�^!�-2�7Ȯߘ��}���.CW���������hz�9��6Y�%��*	���{W
,�6�s��>2��j����S,}}0MԆ�#D�+���{D �i���|��N�ݯJ�ʮz哔Y ��YˡNB���Iި?�e���A �o��Up�u����4���YŚ}��UNN��Y&�֚�*Y������J�9r5؟�2��+(��Wi-��T�f�?k!����.d	�p���5��E~�h4	�ԕ�����`iVO8���cZ�o�2�w�db��bTc���?���IF�����b�����_W���=��e�c�l<�j<��mk�o!�x�c�� 7�g.-VA3��I���Zc�]%b�2��Ehm� Č�̥ �5v�5�9�
r�G^\_+�F��#�����{�줚�!�1X��v�]��"d��w�&�`���S�C�W�5���oc���FZZj��tw�H�HG����Ѡ�޴2J�1)�������^�`׳sǹ��9Ǚ�x�S�Z4�'�������N�߬�H��埃4�f�%ؼ�v�O�/���G^Q��V��A�"fo<uҞ�UQ�[�g�

 ֑.�[2㿂���z�!�頴6�-�iWy��I,Vi(�0e������6��|��e-G-��J��I�E��S��hD8�y?�pm?��1�{�X��dg��z��vPp�Gƺ��5@ O� �/�_�w^v�w��q'%#����ʀ���
J!ze���# �O�	%���Px��V, J�[���,rN�=jMC<+O8ŶJ���D��hE�9-�.����2sZ�y�6��E����Di���ӘG�~ ���*J���i�(<�����` ȘD���d>C<�2�i0�=�]3�H�s�b�<�a�7j�b�����tP�T�&L<������N�jb���@����Vf,�6���S�5�[�h�ۢ	+�}|$�nF������',�F`��.�0U�'�-�!�U2�q���Z��&'�q���Ϊ�:���~#rX��_����ٽ;�m_������1�0r�@�G$�kM(*3ⷯS�s�-�����ǟ�p���!�y
B[3����x�~�g'0�Z�<@���>��}�I\D�e���s��#J��d��P���^��!�����x0�<O����9+�w"]�'}�0nSm�{E�p#�'��P�K0ӆ}�_Oa
Dk:4$Vr�SLrE��{
���G]u�8�U�ѰO�
(�L�*����#~'�5*ֹ�\%�SF�z�X$Q��˸��p���]'�k�@�^������ъ5�^},L�L�n]^�<�Wð����ڜ+[���)nOU���Ub1sr�><�o�p���X�p��]�L�H#�DmP�/^�r�8Lϩ���h����O׬�İx�N��QI�O���$����Q��{ҿa6@I'���4Ƀw�µ�$!3��Z=�X-�"�f������o2q"�����=w����&G<��~tIM���5��:��f���y��C��|:�F���-�������ћ��?�@SJ�r�uϏ���O��O�DX��뺳j�(7lO<yQ��v�=B�|��C��K�z�Q)G�<��
h���g~FYtL��T��w��%ֳ33�~PΟ� vU�q�k�B#fH�����&�Ju�/&�m��H�ɒBȌ�������Q<޽�1\<ӭ�4>=�������X��Y��r�@�O��ħ�� ���5`�}���V����s�,i7�tf�{x���F��рFaw�[�+��f���Gho�n���1,p�'�)[��a%DE�	��C8�pF�%�p�v�w��Wl*Y��_�eE���~�=�U5}��,�i���D��!'}���ha��T��w���&��86l0�m8⯦0��r�}�B]����׺<�e{>�#������Ê>�uuu=��e��[[[����#j��[8B���v�;��,������_tد ���fj k���|$&=� �M_wl�4_O����.iZ�t���-���H�gzx|���xʶx}��7�pR([��?�Gb�.}�J�)T�\��ݬ[=Yv�c��A����#*�豙�� k��{�=� {��� &^=H���"�t���V�h��H�T�Li�k��
w����<>:�7�D�����'>	A}���������j���9����Eq�<�&�-�	<� h
���7�<Q#�(��k�As��ب����7*��s�?���w$�@���<,������LXu}>�)�4]i�j�h�\�YF�#x��iJ �CT�D�C/*�8��F��[TἩZ���s�/�y$���s��f~�F��(x��ycZ9���Ȱ3�b2J��#����9_1/ש����z���ų2��3�]��r���:�r^��;K���E�~��Ocj��󍢄���tI�¢6�$eWfS���� ����T����`-]rg�}9��ͷt|���5��)$߯���*�Of��o�����+6\@b0���c�;�ҥ�}H/i��C,z�P�N�6If>vpSE�˸q{T�/|o��|������;��8i�E�� y�/!��xQ��cZy�ɦ!�W�F@��ٗ�L�!����Io"�mU���ힶO��̑||�.?5U1�5pʴ}��~��y�Iay��2Q���I3�4��$cPVG!������zB�U��{h0��9�)蠗6�u#RՊ+fR�𐡸������#���h.2\����� D���N�$'�E���)tTQ�#�`�L{��V�H����i����<v,ǯ�[�!�ސ%��z.�ݷ��oc��&�m���HG��nt��[6D��h{�s�ϯyI�}x-��v�[�޽��gv��j.�� Ǳg��2���,��/�e̉�z�0ȇ���@���6yJ���=�W��['��AG�+ŀ�LR� E�\YֽBUS}��ŬMan�|��wx8���hI�\FF��@�мEN��ʂ��=,=M�B�'�NRi���=���sYTtg� ۥ�1C�4°j�&�����rC�n�!`�w.uV��Q�n;=��r&��
��ך�f�5	�i_����~��%O+�OG�:�[�����ߠ��~���%��#R$2��o�Ϸ���<����-~I(T������۲܋�.�V\��dN����G=9lI���D��&����!�DbdђzA���@2���~�Sf�'v�A���mn��-����Ͼ����`n���/��Л�%�;iI�P~�ʮU�'<�S��a� ��Ƹ]���� &��&��<B 0���)Q8�"M�cg����63�YDBzR�����4����#�J���\��o��&uA�>�w�n��
G)]���
�"�$��Ae�
���+o�$��+'|.�k>�党�Ä@P��jj;I�2�]&����Y�Ǎ�=ۉ���� �`Y���,�<�{( -�@B���=<(��Zep�ˌ�p~�j�]��܋�u
�;��|,�=v��`x�^�a<GTWL!�PC]�'�k�8�|�3�P�����4���l�y�y�) qJ�"h���Ap����V��8O��ET��O}ʷ�Z�@ �1��2�` (o�﵂�������r��r9��l�#��U(S�A��F����~�jHW�Ӭ�'3�T �KY��҆zjP���D��_��4Z :�b}x�i�֞q��;����TA�4�����}��q��%!�$�U������j�욛m_��fū�)	((g�*�g��r�_Vfrb��,?x'�=x1Ng{5���E��#~�,�أ��]Y�g<4���_j��?�8�������F��?�[�>N���'d�a*�n)��̫��/3��`���p#����~���"_�z�m*U�7����{Q`A��/�-dĨ{r/��n�j��H��k~¥rЦUo��`���˞R-�+��&��Hn��/�;+ ��p3�1�r���D�e��qSg{�x�a���;���?��jp��_7�B�6�^Rn���|��g$��b���3���;�<"۴B�����%�ym�4�"�Q�3 w�O��,d1̨ɑ�غ��b|`$��Ye�l�a�
k�Z��]wZ��onч@�[�M���E��y��4
t�X1��d��v|&#���^y��H2�(7r~γh��䉛W�0;-�q=�tq6�IW�辂$s�k4���B�j}���'�9Ԍ�Q���gΦn�u"1s.#��D�1#8��EfG��9;�C �婿+I��RJ`[λ�ޥ*���y�Ȕ@V| � ,Vvd!���3��we%aP��b�F_'�F&��>� V͋$��1����&�eGL�����X�m6����^#�xѿ�<��Ҹs���?#9gr1l���3�o�� ��w��y9�v���=�Uz4����@���p�Ze��:5�V���i�ID:��_�|8��ޫ%I�}^��mG�U�ci���hR�D�@���0 �.�oq�|��x1�dj$>}�ʾŏx����9�(�n:�!Z��7Ϊ��3�uз2�{0�K�ݴZTJ� B�pw���$�R���:3Z�͊�?�r[�.�G�aNW�u��S�]�=�B0��S�A���D������:���
`�X�%T9&�Y:>>.��|}���g����ΰ�KU����'W�g�7�y�a��&�\�^M*�@�%?�����1D2@bP���1E{҇�Q`j�̅�����N��|�V�x䢇�脃c:���0����s�qb|��4�N�����P	G�'��:���}�����$)��Hm/�ȝ�����x�[��>$?x�@��"ur����pB�Y��:ޒ�0�D��e}À��ΦԶ������?���U�N:B����	y���A�T��z��Q���������SG�#�Z���y��F��mĿ���"�OI_Y�v��hw�9��� �AU=k���وse��y��t��Z,i��y��N��@��{r����(<>Q�8}��zw|�'�%�\��|~�R
?*�^���D���!�⡞ڎ��v�Y���l6W�$���H�ϖݧT�E�����i
t����u{�j����ކ���6�(7�:'�l:Bn��P\��7ޔ/�\cz��[Q�ƚ���-)&���1*[u}��3��I5Þ2� m�K��$�C�
�$�S�H�<��b� em�v�@֊b�G��g{�����Ed�R}or�u���F�Q��:���N��{�m�dlTr�������Q\o�&R\c^ܒt��F2'�	=��aoU�������Y��#�?_ruk"͙{d�< v/{��r��
)�;���>_�!k}��?2H�+sX��ɝ8�g'iIH�d���"��I!j�s����\����	m
v���#�wÞ�`�{�iboA��ƅ�f<8׸�9 ��X��qj���*W�nLs���]�?�l+~��� QČگ]����zhͷM��^=�/�Cx�^�i!�.�}��!�pj�&�U�iɢT�%��"��lAϜ�Q�c�	���2�W���L����MG��k��0O��c,�f���]�O?0$&~����h��2a��'O��DGAj^A�ޔ�����S <\Թ�JZ҇���n�<�^S+3��K?yN@�:%B�rK'��7h�B/�M"�髛�]�;�_{����q�:���e��z):��؋a˧8&^'Mu�H�MN�=A��j�ݣƝz��ݏ�=BZ���4<��X�naHGnծ_�ց�=�I%@=V���%��9� 1l\��Mo��	��_��Q|�U�uSZd����:l��o���^�dҨq ���%t�����;%�4��N���NH�.�+���O�+ZYn�oam�y�����5R�B!V>�8Z ��P��<�G�3�,����}�^�]�M[��� 's���/=�{:NQ�W�_+8#�� �6��d�.15�͠�@��L�ܕ���x1��ޞ�r��nk���!�}C��A�n�D���1]�d$��k�#�1�G�23�U�h�n��+7�:���Q%�Wh�Qi۟�2Y-0&���7�vs��u��PB��ٕP��l���] %u��ͧ9�3M�z����/�{���R	_+��|F�C��q+%�!SQ��;��{�w�m�w;o�O��V�L7,���B�+)`���K�/��?�(ng
�m�ۉ�<����D�zU-Cc��߬�*\(�(b^��&Bn�S������H]�[�yoQ7pnӠt�!�Uij��>�Aa=)i+��)��Y�'uU$��s�۷��<�ml�u���y�~�Ǎ����/��������A%�O�/�ⷙ�sY��7�/���� C��~�����gʌ@�lV�������﹊�eT��s՞r�9��Y���=��)���x�����bڷ,d$�p���-9� ��T�֕��~�e�ɽ9�վkT�t[vC�;B�e���=w�Aܡ���z)*���'�x[�t_�!sL&�v�<$D��+M ��l��HI��iD+B ���!3����?Ɇ#���h0c���O|�����_�JD�r�e�||�9�R�CNػ���^X��R��9e����``�B_�:#���c�
 X���`��\7�{G+ht3�K<�h�m6��7�qM�D�����?��,M𛃾���ਐ���*���_KXGv6�T��2xI��&|]�I��鍃q���z�K���ͷ�����h��ِ���*��i��\�H~�:��e.�+t��¤� 5�y�7�_;ʰ���%�	<$n0��a�x�k�[�Mf:��JSu�L8���!u7�3��Vв�vM[~d��8O��Z֓۰H�K���\�31�C^�f��&���F�Nqs<���D�]0���i�@�bO�=�WV�,��%�羓@����.�MB)�;pz<!��>���wF m����m	�&�o�"�%2��!��a�7�b�9*T����.D���52��Օ��-��H20q_|Z��f��w'O�nWٺ�-��&���D 8��r�C����AĄ(>ۢ�̘r�Q�N2$Q���@,T�/�'�P渫*�Z����O�SY~9���Ў�@�X�=s3q��o�|��^~s;�����UA�YK; ��u��ʿ��ھZR�E��Zǘ��-�����L���|e�V�*X�Wd��B6[qr} Ŕ4�,}T��fO�ּ��5 ��A�R�Q���y�k*�G��T��� p��ٜ��uRP,�L��#9��8 �u���g������T����ͳ��㱷��I������EG�����������N�Cx�
����TTre wq�M�B�^B�B�ѝ@�@L?�u3+�L-a$Q���5�Vc�3��;�(���){1;-�X����|l��e]=� �$�;*����ISl�a[�%@{_��`V��t�+xl��a>���_�o�d\_�}����6iMf��:�� �b�?�)a4�J�e.74=x�(�r�hN8x�"|]$rs=Q�A�jQ�����b���q[U/d�Mu�J���o�_D@C&���4�I���
���\���/���2���ʸ��f�	[��;�& 3�h�E)q�D�[��|�<�#���0YF �Z�Y�2���e��anf9Dy5���X�p�X�����<�$2��Z�|n��B}��{�;��b܋�s܋T�>�f9~fD�B�Rt4Ԋu��R])'&7Ps5�&
�"����T�,3.-"O��4��{���6P0j�v8v����ڤ#���liPz��&<_;['�z>,~�����������v�=�����; �Y ��֞�"���iS����ףa�b��c�@�
zM�"���+2)Ӽ*�s)�F����W]�}�����y"�}e��.��S9M�e��?̡eN|�LjV�v[֯��w���W��G�j��ͺ'�ɩ���tbb�F��H2l5��!�ӧM����>�eq:�B�<
������|R�h�����G��G� -ވ���pc�-Ai�b8>��C�+lk�5�pV��Cץ�6���s�K�ø��,;]��� j>?2B �����sm��D��M�BVb�xo���\������l�R}��p�ū� s��4�ͣ��YV][��	���34[a[�!�M��;<������i�������vx&�vx]��c����,�Z�L~V�qwѬ��J�wG�W��lsv���������s0���� �.܃��9�bb�=��T̳!�nI����z:q'�+�'�=�~%��5��������gB�Q���:8��V�/KI�=��Ǌ���I�a*���$����S𘛥�?�wr�F���J���搇hn0�|O��xfx����"椛D� c�p��Ʃ���cz�@\���ǵߜ��7T��m�ve:h���Gq��t�aR�V�w�t����nt��(��e�5���8ñ�G��$�knf����ZPQ���?%��`�ʁ��zl�#=�~[w�Q>,�KQ�cy�g�JX�S̘#Oc��x�S�m����ތ~���#!.4��1�}�3�b��u�
�õ}�祆q�Tu����UIo6���~z��$�c�ǣ4�X,bT�Z!�b��	?jb�p��wJ�Û6��>�@�h��J?�+x���B�̆�_�R�x�]xP���""<�K�v������?OF����/��N�	����+f�'u�x!�ʻÍ��n�������mee�?'��7�U����֕��Za��+��U2�8�S4��� ��B)f���kL����чq�N&,ll�os��E��iY��Y��w'�a��S�#��-��Z����\�.��.|r��1�cLY�ҍ�gXÅ���%�H�0RvMu��
X�-#F�s?TGd7�����n�l=���{ J����f'��C��jf�B+V���!*��u�.��\�Ҫ�*�축�H�~pHeZVL��c�hP�*;��E)�j��XѢy�]UԱ صէ�O��x����mR����w���Fj�XV�����沰��7�_���l8�ʑ{w��=Jk���U�7�]_t�\T�7c.e�/�v,ɣ"���>��e�d���z��4�f r �@qI�|+!�_*і�Z�Q�h�����b�:z�q�#3"�>���v �~h�1�>dm��' ������s_Y�0�"l�I�{èǝ��������~i����I�?)�4b��f�m�-D�Wy���z�B�.�c����9�KMT�p�1>���%��|}��qy=r��YNxR�KR�qusX�����[�7�	�!����ZT �
×cEl�����~������\�����l4��>E̭����8�`\�����t�!
��gw�{��Խ�>vH�"]zN��Vu\��Ƒј�N�	`2������|1S�m��%�8�&���[��Z>Q���3.R�wJ.T7�w#�q���0�G�rM�SP��g���=Q�6�ƸEn^tn���X��W�lB'����[�9��<~�#l��pW����|!�{kG �i����4a�� ��~I���b�j���Q�y�P�#��&ϩ�Ɇc�e����XJ��tқD�mq�'7���@��m޷�C�|��w�Q'��{���+�~��t�`l47vq�~/�ʝdxwZȐ�ʛw��w[�+�mnoo�	�$J�!�_�.q��̏F���@@2�}�|�l��/	�a��{���c{�x����f܂�ۂf�J,ż
ҧ��t-k����X��Z��6�b�v-��f�F&�˼�M�b ��� ��G�z���D��^+���P�	a��c��,��T�lJ�P��H�AB�TtҒ��hwLf��z��� ���Ez�݇#QwVA�iU�P�̍�`��9%J/�
�:hQQ�[�kۻ��A��J�|�}� ����~(%^HH�}8M���/.�w-�,��&��g�S���\�����ҒG�6�A ӥ(߫�~Hj(�F�Ƒ�t���8x�V��
 d%����kZ��6�*�E�5ֿĭ�Ԃ>,�i΅��Oq�4|��z(g��L�&9�V̞@oԞ���b�P�[�ǘ0:�\>6�������,往V���5^9�9��?Bن�c���{���⛙v���gS
��1V�
`=O��&���A�x���]K� ��F���=\/��hQ�鈈F9)IA�r-q���1����p�LՄ{�?���'��? �)aس9L�nIrr2a��%ɊlGZZ}����z7��rp9���#�Q�N�=+3����Y�řG>{tO�b�g �����iZ<�IBi1x[X�`u���QzO�U�S�	��G�Q�s�v�@�)v�䪩�|Z����0�$s]�{�N�n��a��m� �����[��?�`��2:b�8\��y�c�����U�%����F�P�[|d�u�^�d � ����E������d�+#0AZH�e&��ĳPV�
;ROڄ���=�%T]v�[��L��
g�?�.�YRa�䇯�$=*^e��.3
�#�葝�b����>Ka�}�nϭՎ�T)rA� 	,au�gBS%t�|�|�-�9�Y�I"�Θ��Ud�k�#z�"R��)D[xk��EsT��f��F������Y>]C^=}�T<�T��3o�m4^��r8&�df^�E�飼��z-p�f�D�-�$e#�#u�A4׿�j�A���vl&I����C��ۓ�҄�q��dN�s���Xۮ��m\< �\�d�����B%�W��)�8�:�u(>���B�~h'�����7����9�^�sO�XG�80c�|s�G���Ir��"Ϟ<���Oz99o/hZj���/�M�e^�$��SQ�Ip|h�����F��i���ؾ-fD$bp 1@�,�!^ ��8ԾBÈ�<V"��%__���D�_R+��[֕k�QB>�� H����1?j���"�Dy5�
�f'|�4O�2�K��U 7	JF]�ƨ?vBB����>�Yȇ_��3E���������J�)"G8S)ڇc�(��dۋ,z�(���t� ³mQc�@��R A��=*bXd� 砯�~-������bLr������;�����ģ�:�y;������n� Iz���Yμ�~P���÷��{W���T�O6cXڿQk;����}��\iĨ�5�����.�b�N����ةr��D%%�	���x�/z�	��Diaԟ�M�̲@6���Oc ��ʩm<tu*���� ��)����%�%8E�5���>0�f�R����Z+DM
)���m�Z�(e*�U�Qh�W��^�a[��k�e����Tr�۷-���7��я�JZ2��⟄j�7�k#\f��p?����n�K\}���~�=��L�{1TIG����i�c<x⸹���!��?:V����u#�<��a'T��n�������}�һIϫ�߅���sgg�NMo�<hj#�(,��L�<ڪ��)[�^�x'���(L�^]��q��U6��E�䕜=E��v�	�C=�J���8!	.1.x���-o��:���t�+h�_L�K��0Wv�Ũ�d$L�jT#ƪ��P(��@O�	���",b�٤�4�ی���6�m�]����_�;`/h����S�r��!���osO�jث3X2/�K+��FP�Ֆ�+Tj�ȵ(�GJ �L�+�����W
/
���ǋ2���Hg��+>���н%�')0V�让V�����.y"���D!ןMMڟ��Ky����;�k�d�����@��@�U���*��.�P\�{��߰����)����yQ^�q�f��T1����N�X�5Ԇ�@޴�5Ξkx�(��gE�s�F����;�7�Uw ��1�`C�����:�[�ԃvҡ	Ä�t�q�G
��⛧�N���$�y�#�1��ռL�ͧ0�$z�np�X�I?��-������E�¡	*�]� &�-�U\�M?ar�(� 3�.�2�G~�����,�y�����)��V�|qt�\'K��K?o�;|����������߳������9�&s5u5���'��ž��Q�IK�ű��ku�0m�ޣ��ݞC���'{y'�E��+�@I�����S�q7��L�H~I��pTeϲ��X>{��'��vTS��봃��O�VHr�tډ\�;N���	��!~e*:i����2� ��"��`��|࿡٨�m��7�f�*ڬ�9�:LJw��[�c�b�I�@ME������D��|�̪���<vxr۹Z�}�j���&�7�5�uQ�8�X��R��JIt�wP4�1���{�?|^�����v�Z/a��օ������7?6����yG���MAt8�����X��^ۿ���@�'�>�9��7��t�ױَ�9xa+aߩvUZ~eD�U�#��ΤR7:� Ҕ��U�8*<N�[�*�S�C�Qj��NvDF㽅{��,�Ƈ���XΚW�*��ΓPϮ���b�d��\�t��K;�����$�Yl�.�S���Y^�˺�.wM.ڸ��w+�^v�Y>�?�h��8��m�Ӡ�p�b�������>�y�W�����u�L���!���2�~.���s!�W:҅@��
+�1̧�cY?R��+�j��-	�g_	������)�%��c�G	)>mxs��{Z2A����]�@���S�}7�X$ĩ��m	���� �4�����5L�ۤJj�۔[c��	S+.(4��Zi�Gʤ90�:��D���2_Бl���.	�Ҟ�AB���}$��O�
����a��ŖQ�2�<�V���h����E^䕲i^B[v�l4F��>�qu�h�Z�]��$�XuO9UE�A���J2�'|�l�$��6���^����=�z9%�=rW�h1�Bx�c��������=�2�g��x ���������Y��**�,�??F�l�e�����{�n�j�8�ߝ� E�u���ݫ�RRR�d����,��R7���f�D/럫z�
���w,l�"}=8�oĈ�U���U?�6m������N��"=�㐋H,�C�Lc��R��.NU��ʲ�X�{Lu��w�X��J�F�i���c-%��OY^��V��+�̺�V%@m����௕�flYje,:(��w�X�c��>$�J�}:��:PV}� R�t�_{Uױj�Ndx�q?`��z:��r�i�ۻ��	:��l�ϯ��r^w��5csw�\�;V��۾���
����{~�䭸T�f�-)��g�s�?�\���]3  �}�ڦx��@*��8;
�O}�1���+�%��eDN��ٴӯ��?���X���L�^��徺p�ɂ�^l�	x(+��@�-E���jy1�X;R�=>0�JsCm���'��x� :[�Y��tm��e��������]ɽ!�����4���,��o�+�\��ʼk�bd:?���3� V"M�/��T��ۤ��v쑥@���n�{���!�;-�uo��9��/j�^��@�ɷ����}����Ncz��D�������/Ʃ�i$�㷗��I��00+�����-���d����䬮!oe,�N8y���h�?�[VSJ����>�tV��L��h6J8[kW�� ��\��UL�d.O�ݜ����8��1�}��W��o�t������F���
�*v��
�����u�|:u�Y0��ʚ{��\� �h��Ԥ�8��}�@�u-����3#+3�k�����˼|J�[���	��	tt�W��l��	�p�����n�z��w�ɦ��}��A�����.}m��C�a4�� ��!jQ��8mEH\[���5��$<�kt3D7���K� ���a�j7EU�*�ymi`=�wz�Բ�2B^H�2���si��s����=
��;S�S�����y��=\�*|1Mbs%�c*�'�c/�r^�zG|`��E1�j��I);��?�4�^o�YJ�³b|���)���k�va�d���t&�' ��>}+z4AZ ��4?�6qU:�'�m�m'�?��il�{�{��U�-���F|�5����m��b��9�:�[����f�[C������{b������mA�y���=t�Q.օ����ћ�"T�/6xa  su����8t:t-#��>5}W�V=`]�D"��˕��;��'vI�	�<g��_��[�%�\�U�L�WI/y��Q`���iYGn3n�~w�˱�诱nO/'�n��A�޳N;]Y
�����IZ�1�
�#�`�9��F6�[C�^�%�i� �ⲐJ�[�$��׼Z��qݷ��(y2Z��z���/���ׯ&��nр«�j���\��t�%�y�Z�t��ko�#$�p9ڈ�ՠ�Ј��t����P�nasB���6̉���K���H�=¼O��9�-!����� @Vv#M���ڦ=P����^��Z<[I��euU�����c 2����#��C�?��%Ӛ� D��a�"h#n0L�#��@��aT���_�J��j场b�p^n��Y��Ú�Y#O�>@���c��`>xלzƬ^��D�ص�\�~���ssvz��G�	��F�A֏��\{�)
y��N{N�|&4o:�&J$5� J+�&$�a�S�B�f� R�m�e���l��(�2���K=���z����2���{�R��p��S���n��(�I���P[-+�5u)�i���&����\^$�%��v�>٫
�4���Wi�e��1��������ku�!�d8�$zs���J��d%��y(�������ں9��𹀳Q��^|MG�n�?��WsO�Z���_j)��"��������ٿ�����k�p�Ng�UG�S�5��.��/+sv56��ꍥ�h�4��c�j����q�Y�*;ηؠ7���N��'y/)5�YXa~�k��_i�U!�p���i���p��<C~�y>,���˅z�r��lG��d��Ԇ��2�(���
9᎕����vL=rߪNۃ)�̮���M"������@̣�1�ο�E�����~:M�jO� �)PXD� �\�����]],��U�)�r��`���(Sb�o�?$k�/�]bw�$�:��ΪX�Tdltt4�0���L��k���?5o#
�ko�8���&x�F��M]7`+��`��۸*=�/m��l}1��tr���aQEP�*c���Q��E5�#It����=��v5 R��@���:aiRfk	4#��a̧���S�a5�������7����5׭B.�F�N<��v�sigg'�g9���"��]z�2$u4
*.�oѶN��A_�3����BP���화v�#�fI���:��n�2;H��l��f6q����B��0T�����*h�'����&���s���]m��֮p�����q棍����y����0��KK�h���e�����*6VV�ы��Z0�`��60�yy��	NUB��k�L	p��3�Ls�+ʹOu�Tq��5ǔS��-�pa�R�ļ���E��ok����
�5ZǢ�I��³��]t�m��ϒ�K�%v��&C�JiN�6x�Ewɏ�@m�{��/��EӢ���
��Q�����UAX����1�~.[��\��ˮ����ij��z58g��;;��̜�ll�t�Ϗ	��-�W�}��>T����m�����Tc���((�����z�F�I������tk��,�=�e��/s���Y��Gg�����͍	c�I����0,`���&��k��buy����WF��ђ�"�a3+�>Yy�C�hM�ΰ$���S�%�pk�e�ìW�����I�LSM�4��l���i��N�=��i�8�jnC�ө�#�8�� ���a�ac��iLk�DB��L��~6v���nn��BR��y��Qջ�;�v����� (�؆�j���"U���+p��*=���iv,^d�6��XQr����iZ5��lŽq��ڸ��3�C1~Z�ʴ��ڧ�d�'�i�~N�i)FZ�@�6%r��$��sh�$�6��I��3��_���ʫ_�V]H����N\F�2H4Rb����|~j�Sl��ZU���?�m���*��}B�^*�U��|�@W+�Cd�i�Ӹ)��{�ґ�
�R���_��,�.���Bxv�:;'^��D!h��cW8Y��xw-�u[p�\W���zU�LJ����#_B E���^f6X�����6���\*�u�����?Ʃze5���ޮh#D���J��M�x
7._���j���g��o*-��ij�
��s��&'i0�=�.mhٲ� �H�JA2L��0N_~�
�ŉ��q��N�/�*;}@��X�m_�&�d����O���1|&h�
��6i�������9Y�Ŷ�iߺچ_.w]���-�(�"�Ά{в��((n|������ X��1�$�\?˭�ה�S5|�E�/Í��9�&ME�O���aN��D�k�aM�m#��
A�����kF��ƭ�J��Z�Ce?s5�&����	C'E�UA���o���iB탪=��(�j�!-�v��T�ZӌG���ߠq%��x�8�f�L��m�O�������I�+X/�����1��5�q��uWfÎG���Շ[,�I���C�ʽӮ@�
�s��~I<@��(�-��7S��y[�&l�>6;�zE(C��	�<��W˯יf�k�_S_�V� Xi	V�X[�xq���N���Ń{���x).�]���������~orNι{�w���>����]Z�*S��B/�3�W��k��S�x�6�����E�#o~Jk2��K�z�2�����JK��$x�h�X�{S�B��� �vh���d��ɰ���J�"�rj;DЊQ���l�9� ߡ�,c���u��V3[���w[t�/��Z^�u!@e��2��]!
au��}݇Ws�L�K�7Z"^6
��=��	�	R�̀:�C��ԑ���N�<t�=��ř�ȧ-T�o���Ɩ�/��%�ԏCb�kvsR�xL�7[��30��=]7V��FrZ����+�!Ic1�!)*���](zĚ�7u[-���~��+]묓��Xt�N$����nnS`��v�sbmY@��M����5"�r�g�d��"ԧޖl夨��=0q��G�F]�� �gSJ��a��{��p��2ЕZ�`4%f�w�;��a�Lv�����S���&x���4�����2�a�p��,"�[ˁ�����oHBb�S��n<����p��Li�.��iӴ�6�mt@p㸴1��K�C᪡5�1�9�/F����R.:ȋ�Օt�QQ?�[��hn17�_�&�u:/�.���<��<�P��)[����r����6�N�H�1"�B��'����
�.��S���?�r���d�ڥ����P�U��?�q�F�ʘZ���R�nm?�u��]!�y*Z�6���P(���n3l�6{"�9�ꯧ��w����;��u3������zݑt� [�E6"d� �1g\�CɛZX5Ԑ�VN��� ��'�����#�Ac�8y�܁ ��e�8@Z�4![�x�mQ.�t�G�s����9Z��wa�>���X�і�E����J��ǚ&0���s׋���e�j�Vc�bo�����)���UT����Oq�i��8_=-�����>�Y�nM=NӚꋋ_�VZ&'}�F��@�A�_m^�ZP���-*�������FR�?A�<�{7���S+0ǽ�r�q� i�?���q;�$�� ���J�ά��!,��|�@�WU�Nu��v��Q��ј֍��C;���9b��s�-���x�fR[G'����1���.�����z�`�R�%���nV×I���L7_'��`k�82OUH��=il��iV��Fn�G��ê��y3(��ns����H��V:�d�	N}!��w� 5'gϺy�����X�#�q���;�T'i>�����|��E)`#q�[�����L��e} o��Q�[~�
C���/��D`yo����w�n��"�\�moo��&-^�R�����8�������f*��jg&�8�����-�/w���t�Og���{�O���gx|*�<���D�{�Q�ّZ�����n���W�����׾��AمQ{�|����sM�g=�mi�2�R"1Lkj���[���vK��K~�}�K[96��f�C����*k����k�F1ci�?��e|+�+ǁ�@'��a�?�=v�����/^�����(�bn~�+�Xf�B�� hE�SHqQdX�:k��?�ַ�O�����u��(*J(�j�H� �A�al?������q���hz9V6/ǻ;>+��i����B0��7k�J\�{k~���Y�f����I㌏��e�^�H��'G֐��X�a`��z��O8�xz�yђM�/:ԁm��U��;�t�H�R���m���}K'��k'���`|}��y��6�޿�2�p�Hc=����}�돞С+����z�$�9D�L��Z���Y��MV*�\�#zO������kb�֜����,��`;�\�滫y�Bk�&�.̧��͘�"�6�	�� �/��iLB������{UP�׍��dgt��OS��Ze�
���fg	��s��K����+|�����Oqr�a�Tmo�V=}��*���HII���{��n�M7C`v���<v9��m�&a������Oɟ.�inO�-��j��NȤ8��b�'pK'A��u��qD�*��9ŉ�R2&" �C��Vvz�	Vs�c��".uW� @�o�W��ʰ/3~�J�svy������S���Y�q��k�r4�����p��Y1z���>�nlbM��S��<=LN�%��f�f�q����u�z�R͈:?�k��2xw,��G�UY�Nx�n���%
�1�(�<��(��gwR-|��;Dj��֖C�MZ�-2��+���x�)Q�&�ᑪSY`��^F��y�;kQ��?��zA�|w���e�b��G�E{F؟����*uuӺVm�Ei�qBc�͢PA����~�۶b�ȶX��K>��u�����o�544<&����^���?!���_DG̀���\y0���~b��o����- ��"Bd�E+|w,$G��м����®ˍ�}��s8���2 �F�o�(���Ι6��nT '�$�#)�<��/,����=����G�����z�3�e�>�=8 2�{�54{n�A-�y-�������bz�o$��qq�9r��չ���+���������C|�� �Y��ʍpj�hu}��tt�/ooo!�q���3������4�z��h�vys�J�MU���c0���@^G�v�j)�4�*+73�����b�iL;�L}�F\c�n�d�c����8���:3���
��	R�"#��~��s�V�Jf�<��6�>�r^Pc�f�5����O�-ᨬ\3ns�A��K�\Jy-�x�|f&�苵��� �������,�� 1�p��� ��?�I沕�zyq!����=�S��E+�`ꔇ��d��v��z^��tmϵ�b���8;�\���Y�v_����L��(77�RR�D3�$T��4Ui��|�%ϰ��k�˄m�b���!�.s�X�N���6V�V��5)������l��Q>SAOy]y��0�Ֆ����STz̢�"ݦ��ﯬ�&���r-窏hݪ����DK��VlL1П��A#W0�9�h��a	k�u��l��!�/��;d��Lݷ	�����loo�!�1��uջ 0Eft���/�}9�^m�V�>j��ү��ʥD
��Y�5n����/e1;�t7�lbD�&ǂ�z����J��y*;�D������w���ʏS��zY�vʙ�j��]��fJ��d����b�ړ�v�NՋg�]��\��#�4���#�`5��EK!#>ب^�a���V���ɝ��mP�B��?\�oܫ�M7�[0���Q[\���!����!�!���6��H��+�ƦO�!)��h.�w����<�v�� i1�V��Pl��Y��`A�]+�n|�~�S��녦����^��7�2؆�����ʱqz�ι����v�Z.G���%���|��Y��{����ivܺ��s��(@�m1�QsCx�9*�\{)ng��*��q)��{�Ep
*��X���
��W-U_����4�SM���b^���������&��=g� �~�ad���� ����x��p��.�]�� ��K/���h�jYҰ�搑W
����_�ya����X��b��"���x���^[�EҤƀ�28ۣXE���~0mfF� i���i:��_�X�1���Q��⼐�C�{�V�6݌���ȹ��� �1D%->���K�#"~��=��)ݡ�Ɩ7/�v�S4��C��g�P�c����
Z|��/����ݽ��,�u_��GtLv�����1Y���d�Z��A$�[
Ƨ8.c5cX�6��I��7ڿm�N�[)v��k=�X���`�j�VG?D���kr�
��_]Zi�^�[=�iN�Jb4��L1p��]N7��[5�O�2�ne������0Q�ڐ�Pv���!]uTI�fGOl��K�D���w��=|�\���Å�"ϳ)A	��� M�U��ړ|
- @խ�{�	�&���?5�2��pϱ��O�;�17�=���:�J\�Pm-Yn5x�|��m���9o�A"���(�k�V��~q������ݔp�㸸Xl<Z|�_,��\p�m�b# nƴ�X��僌��s�o���̃�H�*�|a̶��s��p.h��3X}z����)�3ٮ�K5R9�s�BL=��HFs��3l���zϯ��-_����U1s���)�����������/r��xJ�����&%��0W�����Y�h��Y���W�	=��W����Rϧ����?�	����v���w@��������b���ȭP<�<��bx'4A��ױ���댫a[V��v�8�����l7,�mH�qJ�t)qI.�<�8��'L�+��b@pV�Q�����W���`��.�C��*�8b//.>{spp�/��~�֎7����Ư���	)pަ*�d=Wms�0�턍Cq8WSN�OV�%����t��E���lif�P�C�Km1ɘl,E�kW�V�����o�] Z���cy�  �N,�z�l���!6�-��fǆ��ѡ�۩1q���M^@яBN>�����e4�����S��1���h\V2�W�.�J-`v]ފcd�ǃ坹�rg箌��N+�� 2!�p-z��x�`���\i9;�o|��~��sw�����i��^L|x܅�U!�!c�s��� ���>]�Y�I��@��FZe��
��ш.�4�s+ @�����@p�|FI�r}٦4��V��1�$��@��ȁwi"i��[��M69��?@~��]~2zZ�[˧=Iz���\��f�y�|Kl���Xi��cg�Xf���o�79���\M	�,��B�&��p~�	1��4wG|��+�VC������/��KnZp�Wo�X�m��Go~�#@lvv��e�C�*����Ψn!��]����<�DͤqA�+Y>G�U�h0�����l� ���TV��]/aJ쩥K����}qq�Y�b�؉�{���T�d�GN��p��j�ň����I`��|��C�':0��{����wEW���sax� @�i�eI�3?r�/B�z�ff�%�b���)����&���+v�j�S�����U�B`��Jcd�����,7����#J�.����;�E���ح�i�쳹#��N�E�,��>���
ͯh��1�=�]����A���+����G��"�C0�: d�A�V��
S�bQ��E�O?o�\>���9(��V��'���R���>����9�d8a5��.U��>���sj:��-����-���t�~�[�+�c�d��4+"��_��1)�g_.�T���Gy6Z$�_o��T07��p��~�(4v��w�N:�=%|�|�C�1]t���
�o��iR��FM^�w̌`�	9�6�uI=�q��%f  �|��QZ���h4����3B�`\�1��qm��|�����#?;#{{�R5�]������Ĳt��M@�jf�����o������B�۟�Psd��'4�����݀ ���C/2<

P�:��_�˗�[Hd��I����I@�B�K8��hHxk��K^7�b\��l�������Pl�c�%��
�G�������+FS��x�Sf#�8 ��0Ԅ�h8âcQj5�'$ԛ�
���s���F�u��f�n]�k"�#a���t�w;aaa����p�8i�5l_M1���gz��)QI� _�|4G��ro��$�k��!����K�;�j@?�t���
�3���_HA;h�Y�p �7���w�f�Lo��:D�qk��Z3�9��R��,�^�u*3A�KH����$�cK��g4�v���R�ҙ����4��3;Db�����F��[���[I_pF���g{)�2]HIu�c��Զ��q���/��`O��n�����t}M'�˰����:�ȲOO��O�eD��N�f	��ʯӶ[a�|W�i�w��T���5v���$6~v^� ���"���h����h���|����N��z�x��6/?f�3�X0�VU2a�:S+JdA�q�=7�"d�f�B���������|�f(5GX���\h���9ᖿ��,G��k��h2C���l`�*�r������N׍�k��a��^�9>��+e���"�������fJ���a���)�o�<j6�=G���=k�7��=V�h������ !P	�W���e��@l�� X��ԥe���~{f.O�)�����R@�M�,����A��gD2$%
M5-H���:�g��y���up�U�'J'Ph���Jё��B��^�]�l�����<_"M��<<u�?(�a�˦���t�h돡211��ׯ�gn���?a#Ƥ��)�x��h�[D�i8�=�}�Y��B�/5�j�_^�����=�O=dj�ɋ?K	��7K��7S���lG�����Zѥ6V�s�yC j����o�M�B�^li�<��d ���v�6K���T��O5�ŀ�)_|afk�^��A~.���l������R�~�� ���CRL�j�o���UR�5��Ȓ������ Ъ|������5����pvN�B+�o�]8�!';���Q\|�����/7K�1K7#.�`=M|dff��/
Z�[�n��9И�N^."��pj�;��{�Ȉ�a�1�5w]�j,�-ĊK$ht�f���2U+�h��]ez�>�7Y�0"��j�9~Wũ-y"12ە7�k�v��NЃ�[����p lrq���me�����Hi�<��u��?9��I졌]7.r����$���%XC(ǎ��Do7*+�J���ڬ@�Ԩ���hV 
��J�=u>n�$8~~���O�YLr.:-�[��� .�Q���2>��Aqb�z��ō�MF�%P��Q��Я����E˕;`��I���~���Od]�<v�]a�ܒ�#�t����d��3/�G>K�d��7�Gů+DzS�*гC���.��R�oS7T���X$,W�8��WyN�n֡J��jo��֘G=���<ޘ�z_zJ֮��j�٘�(ߋS:��;l�H���4D
�<�[�~����|^��ٲ�p��{@��̈Lx�M�R��q�)�3l+^F�v����7�Ӟ\����LF�J�E��t��W+�X�I
���k��������[��F�sM��ҫ)����'z�Ҽ�J'����M�R^=����N�(OCI	��Ŵ�CբGr�p?�E���sM��A�f�a%��(�g8\u����/��N_�5O�#����g����c�~U�w�NpcqWUv�|��?k��YS%�������K ���_��U֋=垐;��P����(�ٌ&2�x�/���0)�㭥p?���ڄ��ɤDY�ct����i���r_���L3>��q�g���C�gm=�؇�ݜ1{���Y���]6�� �z��0 ���v���Џ��Jyg�������M��~�ww���t
�Χ&�N(ݙ�D1G~_#C�(0n���$A�ۙ�ף;D�(g<緙JTA��z�@�\	��R�e���Q��(�k����i��#�;�i��GĒ$9���$����ݔ �æ�s����4�4�#Z��p��G^!�]i�Ϩ�uONC��T��s=�DJ�A��P�ymN�Z��s1��6z[lbb"����;*~�4p�ϓʛ�dl���$��z����!��ƝۇwRy]\����g�W+����Ad9�^?��z�GdIK���GqHy�F��F ޅ�1F	G	&9"wM�Hd�藈o�p��e�*H2J���Hݎ�3�w�1&�|����sw�srB����"������E��Z	�=:=R	\-��\)d��	{���:��q��U�NT�~��5�\��������.�F����6m��!��r��$#�.TT��uR�ի�Y�%\�2^�`D��vfF�(���7/���Yzi�7�S�������ӕ�4�(F >�ufH`d5�
����eߟ@�� ���4���TO�g�/i��p
�ACq�8\R�'yi��ũZ�u��7���yUH ��ML�Unpd�RK�ǽ�7,�>���.�xɽ��uu�H3����A\w�g�>�]�AZ:
y��Q����/;���C��̏�x������r�E�+1��27�ٞFWx���ιl�j�B�PP5��O�7l&Þ���Ԕ��V�ǻՇ��p�Z��Pw�f�B_�L܉>�_cqO	�ڒ��e���Bs�s(�f[_���rx{�s�I�b�֌��	��4���$Yl�>k;&-t)�HL�v��۞�p�x[t��	z�����}0NJ˳���9��j!]E8M�@�0S���]rR�KQv+CuO*�J�P\e��}���>�.\¿��	�e���H�/\���\yeGM����,^�)J�ZV͆�/��>>>P�6���ͼ���H��!�,�%J��l���2�x,�,1'��m���d��.��F3A)�N�=?���S����[� A��ӳ�������h��/� �&� `x\hyt�zּ	���c�W�5[1kN0NgB*��g%ø����{��m���붧��NԲk��X.�� P�(ly��Pynn���L,6��n{-/�U_ ��6���aU�Ј�*F����Ĵ�0"ҍ�b!dt��_0�?\,��A&�]�ʩ��f��Ѹ
={���v;��<ۢri�k�qj��|�vM�sC:��,��y	(#��!k�=�$Y�~a�B�F��;���Lg ]M{)$5�J~!��@9��D��rX�-~�uJF��*z�V��b��?�!P�`�Mԛ��>5������|iI�AvTYLly�e�D-��PY�9��LC6c�G@���zf�����&2 `�N�f���h����ƗBQ��ϝB�F{��L|@	���5N!�繇��5d��M���oSJ<D���S"��]���q��t0�Ԇy�߫�VI���z�7-mNƖ2�#�JdhtN���%�OaW�|-�a.�hLڵ��������6�?���?Ov%�o�m:���(�Գn��*�����Fl�7�E�-�e5@2	�P�{�왔�%�:-ܾ��T���C&�m�^(�Ic���GQ���k�f�3u�퓟�rp^�.6�}��q�ߢl�S��}�;� �q  �t5\ߺ��"u�')�N:���|hK�d��^fr��e��J�E�0jS�&��(�~�y@$[I�l͇�C]||���p\��4����
|ݐ���l�e�9��91λ}�@4x
u�vb����?��z�P�_][��s��&���8X���j��������k�+���W,AJ�"4��qQ,Q�u�D�ǾgS�Kne&�z:7{�5�Q|�����~������s%V'&&���D��c��7S�D ��5�{�}G�!y�q��d�V����4�Iɚ-�Վ�&-�x'jjb;;��Q���������3أ����Ԥ�BjR���<��-r���w�t�}�I9o�M�����@T�!b�8�M����;D~P�Ɯ	��vf�V|}ѐ�E�1�B,<I�sev4�'����2Nu���Rz3"���a�u���0L8�t�O��BW����u�_��7t�d�-C���C��Q�%>(=��X�
���+w.�X�qg�����Sż����Pǿ�2��(Yhېl���\��B7��S����?2�u�	*5���Rb� ]���������{����1q$��)�Zh��ݗ����1���7�z�)����*��i��������o)
?l'�?~�ð �|ʵ���v"���([S��{�)Ƙ�9�&�eP���ʁD7���w�[7^*{��uxh��`��"x�	ߊ���$�:��rBCC��f��?Dq�&�M����!�־ [K�q�XU���k��2�Y��>�ZQ�۟�"����6z�-������|]{�%�+�훎�Ǚ�A�T�w�g��ذ)�~���ٻl,^ʰ+�I���d�æ�F����a�=�rL��&�*�}\
O��;lV)p6�U���PÙ����J��!.�"޸��G_O����1��k'a���0�P�����kÂ$�zȦs�H�z���d�	�x�Y�P,Rf���ӂ hqb"����Ha���K_�
GV�Fp��௯?�pd5E��P�yn�ƊR��Au~�Wsd��B�a|	:#P�Ӻ�F7����䶗����>���t:���Bg3�Qc�]�\�t~��ٞ���99�!�:�+wJ�|�Af�G��a�,}��>i��m��A���(�z�0����R�z6��G4�H�0����pss+~�ݵ�-�"H�$�eJ��6�QD�e��LL�Uep�T��V=�C8������L�+���:��(Ȳ?A��`Z�ݱ�!Ak�W��6$��Ef����
��|llJmFm��m�ԗr>�h��WJi��^5�_\����
�~̊Yo��ҽn7	��ʭ\�+�.�����'W�N;h|tL~TE8�+�;v�IK�X7/R7�-�ʙ��3e�n�;�(��;����B���&x�J�Wxo�������e�r�/_�lV�SRΤ��Z/�o���L�:����jjj&KF1<�QZ����e��M.ڝ�O�u0e{���pI�7����^�������Y�B�B�2����M�U):JW��$���5{�v�b�"><�C#�:fu.g���4f��	Q"�(y�HI�es�����eN�'�|�/r%�6iCB�����AG��\���������a3v��:i�噵����h����/��Ǜ����~�"��Fq,5iUU.�*q6�~N�^�+���]Z~L�)�|�]�$Afqd�C�v`"�1�?�u{�⹏P��k�i�-B �W����n�}ǺI3��I��H`jii�e�Kjbb˝���$c��~s�Bu$]0prR�LK2x�r�N���3@�����kk�#��a�����
���}�*>n�[�HPV? ��,[��'��{D�]�E�I��e,W>���V������_��Ьoe�ݕ��������W�������ڬ4�s�ϳ�?=��g���V���?���.1���]~u�C�]��a��/��/���k>�)����5�\=��m4��W�����O!��f.B�����C�W6�z��B_l��W!�������^���ǫ���<�DgХ��m$4a]135�h����I1�E"z>�PK   Ŧ�XʀjV{ �  /   images/d1dcf8a6-8c27-42be-bb16-bda153483d9a.pngd�ste�5z�tl��q�۶ٱ��c�N:���mv��z�����7�g�3��{���kV�Zk�)ȉ#���  DI	%  ����9b�z��ysRTM $ IAw���/�K@���Ɋ��.�M���fsɯ�u��tcu��Zl�J�ˤՍ���,��iLCב�Mfg��.�,ٗ��8g��H��#�_~K����A
�q�����N&�x\�>��F�T rE��U�D��5�4}�|?��Ф�� Ѿ��I��J������5��^���cd`� �:����/���D�ר��}����'�B��N�:"��~ɥ����&��%�<�l�R��7zN��P���6�3�ԕ�B@�4a��&S/U�LAA�w��%���2u���U����h�U!/�ܝ5���4)�&:�.9%�][W�0HΞh�yM0FZ��]TU�;P�u���8n���:��d��m��>��ؐӽ�dBסͼ�QM�T�)W��l���򝘷�ܭ:���C��f��˫�8����C��6Kn�&�٬�%���ڞW�X���7�.�˖�x�d���� ����Ea�V&���:�kU�k�X��m�w߀�t#Nd�?}n�L^����@�Ko�.���}�ӋT������Z}#S�byY�\�%_�يu�E� ���k�D�׍wNҘ	?�Œ՝�k42VȻWM������ɉ���L��IkV��ijf6�}����Ye����C���Y���n�ɞ�&{� ٜKVZ�$�^�ጛd|��[j�q�be��Ru�QZF�ܑLR��������0rggv���Ck����і�xׅU
�.�+Wb������7���߲u����'m���y��_:�� Ư�w/��
������UhNo�XXv�<��ޏ�����_�C�#����iZ����5Tjk<�W3�2}�I��A@1�����u��@T�����b��%�&t��c��Nn��嵫�c�J��wt�s}Z�h�տhD<���7����21�S�_���BV鶫Y7�����zڬ�̸_uD�ʘ���H���q�5��W�M�F���fĜ ;|u|7�z��Y����;�>:v�i��`�I�nےtH���[{��JNgQ�'��R#��*>77W��i�o��a"��^{V�����f�n:)��Vz$��IaA���h]���2i�@�m��A������nǈ/�m�X?g���󚤔��뙬��׈7!Ŕï7l�ʕ�su��w���@w��k���$9��c�Ҧ���ߴ��u��0,?�JE+�-t,�+VC����%��ꧢ[@�"U(���j�����֣�����Z�Eϝ{�==k�4]��3m��;�5���ac�&�I�J\z6� xW����K�KҤ����󥥥��@m<B��z�-���'>X��#g����f�uͰ�aŊ-s��^R�t��j�
M�X� 	/ǰ̺a�o���iLɃV�A�"���p�^��J�J�\+�Q�?:*�5c��܉}��oHBO:����kቶ�����l�L�kZS	������fQ���9�!��}��+����޺~E��QV^>����p�BsT�p��
��Ę6� �C���j>�/��$��8g��9��E��~>H4���Es�`�Ȩ[���G~S�A��Yc���mӎ,qt�xt�Ҥ�l �`m -�)�f� ��*}�f�up&m�t��������S3�c���e��H�NJsAJ�b���@"�*e--Slz��7�sκ��-پ��$f��QI!5��.4��)����%t�/:�3-�
�����0���2�P[��L�̟��HSPYQɞ�.��F}ṟ�h7�v��&�"-��u;������z6���5A�u�˛�eY�ب��OF=j��2�`�T˭'���095m��꤃�C�����M���vfRˇ����5�1\L�x�kU���w5u�|�b LT�H1HEO6�G�K�� �)=�N��a���Y��Ѫ�*W+�61�z۶�5Ȟ�G��l\��p	i��6�MC��XN �#���غ�rс��Ï���O�0;���* .��Z��u����s�������������5��٘�icx�!�A��U��ê��Yo(Ƥ��JU�5V��%J������E�iG�;�9Y&�NN:4�-[�͸\a���&��&�l��=���$�xx�m�����pN �?ӜN�!y�,ͻY�La������>_���A"��]��x������5�� (�K'w޳Mg��0it���s����"S��������2g�M�u��a�1�����]���)�LKJN�(X0�޽�iK�7OD_B@�:�`NC�������v�$�RV��~H����Ʉ�5~;ާ��+Q�D%�[�=�c�^��l��(�q+_}d����Oh��m:��� �e�VB��!�f2�"�M�-^BN�j#�d<2A�ݎ��4��M�GO%#1N�"K���8E��k�}�X�����/&��2�`��� c���)k��X7D��F+u�\i�Cl�hhW9�1^g0��1�n�j�K�I'���Ǎ�C�v_���P����9�S����3�@	?66O!$��_?�
n��1խЉ%.=D�q{��Ⱥ'�LG�b�.
�L�r6�;6Z���V/�~V.��	rg��}�vxOL"�'ت�� ����B:TSM������vU`��q?��-�B�H2�#p۟5�_Զ"j�kx��s�K�zC�����%�e����<'�o�U�B�����)K|hԺG�1���X�(;�%��0rd��P�s��֚�$Q�O�P���ߊ��~�+_<�?�����8]�$�n�����gWƥ`��� ��`���t�����!?l�l�CI���bi@��
#.Pr��m;������t���}#��O{'��K}W��Y-�K�x���$���(!���0�Vb������D�P*��O:��{��ᨉ��×��$�p���K�A����WG�?\RdMR�보�P�b
���/2�l�]m��x,1��F=��TɌvv��y��6�⶷S�Ń?�.^(����:�b�S�έ�����������+j�?͛���'�+�nrS�#�f̺t��Y�}i���	��@,��M�;
�C�s������>���L%����$x����9	ܼe>�ò�y#�<�F�MU)M�4l����yi�@��������WHT�b>@��PHs�p������}�����g__@� ���	���d�Lڿ,ܰ��'���QGgg���N8�X�r*&������BJ3� �1��̝��z��B�7�H�[WX���у�!��c ��/d��q6'$�D��Lp�i����wc��{�ɗ���y���%�u�Չr�Ʌ��w��6~�~ �Agh�����d�iZ,���j����cl|�<���rP?�G�{�P��?��אɛ�d��~��$��Qa
���2�Kq�	2M�+��a<92~rZ3�`�ۆ��B�' ��~�)ԡR��~6�2��.e���'#-�`l-h���Ƿ����z,�|�+vpaF[�W-g�1�/ �
�'/��[s�:��ڿ�l2��g����U�H�;��u���	lU��w#�]�i�G���B�߭�i�A��Cl�m���;�l������۷5(o�?�KF39���L��8@F5G���s"�GՉ�?S�.x�!�A\���6F�y��!��_|�۟�Z�\E���=����ڏu�Z
ᆊ�����¦^o�ld3�Z�A�������m��:SC�G�߅t�IS��N�����iJ_��;�R!��cB��:.���.t:$���
x�8�|���߷��n��/������_h6����V-�h�PZ�B�J&�C�(���b#DY�mJ*+W�av˰,���e407��e�zZ8�y�\}������G�Z9�p_�pXj�6���6�M4Ȳ�Bq��l�4U��8���nP{Sę�9E�!�/��>z�P"���}ey��7�$6�s��+8�����j�c��5M\]E��H?1ջ]�۩���fBG3-�����T���z�X�ք\6��m��ipg��5�d22(��7A.�x.�5�!M
�^q���D��ll�DA\qu��.h�0D����H�_�F�|N{���	���{���N��JϜ�!�ȱ?��k<�3��viO��Wcz���q�	��	��e�s�O�A:��Җ��!!�ٲ��X�yZ9��SP�_��i���|��������<^���V'�զ�&;�F��ɾ"�3FY#��c����V�����T�-Ā��X�a�]�H�uB���3 ����>#5��#����dUý��fUT��ū��'�`���m�Ȅ6&kV�~DO��j��O��7��9�ֆ֙g+�����/[y�AzY�c\�`ӼC&eE�B�nx��S�N�C�>ݟ���/�a�Ϩ�:���G G������h"^K�������v�M_Յ�d[v���9�c�y�J�?S1w���ǯp���ޗ.�]���l��L�<g�f��%��?TJzљ�L)f�t	������V�øC(]�#�����y��L~�h'aؾ�H�̑����jo���7|Tc�唧*�z�����g�~enw؅�R�%/��p���~Ef��|}��Z����R�(���s�J�/���z;�Wl�AF�֫���}`����HndɘB4�_ɴH�x�ƥ]Z���^�U��^��*�O��TSӟ����u�!zȳف^�%��h/ꄋ��k�i���
�S}-j�1�+F.(���bcv	��.O߉���q�P�H���Q�z(�к&��6W�Gw�����b���|1ˡXp��������Ӕ�F�#_69��b�H)���FOrk�ֈs�FKΪl��#����8 <?:�({r���w>f1��28��Vd,W�J�64�]P�%/:ϫ�^Ū\H�k�%4�k�4X�gKS1�?D�xiΰeG�]���Ie	�z7��\�LF��j����ws;�O[��sin�c��V@oݥ������tf��U��x��yS�#<�~k���۝HН�������e7��b��quՑ���c�z�wNy2�8@|c(sʘW2����?�f���Z���O x���ƷtE��i���W�V����I�1Q�b����5L��pX�C���o���;)A���*7�|,�� ftP����y�i��w�p��(ޝ�����R���7C��: .X؊n"���>s!�1ߋ���`g�H>��t�{[��jS�z�[��Hj�@����!�ʢ��>�Ҝ��1�,2������<H�`��2�/</ح��'�� {WM�T�E��I�w����SYŉ�4��ue�ɓEkr�Py2M5?�o��q�=I��2ڊ�\wIg���F��sG<%ã
�u�E&��9�P����"q_B����*�H]�w��!��t29'�o.I)#��S+5>[�ш�k�E��{I�\�+�R>2���Ը�����
y�&>ܞ�����j�˧��Ftȳ���.��1��P�GxΖ+.�9a���!�Y���[)�����!��C�����AV��^8�gڛϋl��6�:�>^�{�5&�{d��N��I�����U5Vv*U9NNb���8.�(�J�Ԭ㩶�T3�.B��{K�y::"-U˰l�X͌�i�?z�&��^r�e�/0���-�*���)��P)ٽؒ�A�  �Ԛ�u Q�s���p�6!���c+fr
�@��'��F�ڔe�4�#��s�� qk�n,�}�-�u�נ�1�n�&����'@��M�mM�n� �?D`3(b�E��ؐ�?N^N_�������v�~��g���|{,��g��N�x�t��%���kb��Lo�h~ם������'��D��+�>��9�պ�d�t����n[�(M�I ���b��X�b����W�͠�xa�/ �����ֻg,�x$fQ)�k6��Aё�t2�d��/��9$*M�,��)�5h�tm����V*{����� ���4��Fְ1y���B�����Q���oH���MT@'lg@p#nD���<�꙱=#_��2���U6;C|v��p^\�[y��R9�~H�s����%��)zd�0� Q��'�{;�w��ӝ�A)�_Q�,W���Le�X_]��ni"�v�Ft���ns���6���<�Ɓ9򯇒�l&�F�)ֻ6[�.]G^���	�d�L��E|��bYez�p%\"�*�.M��`�= (/.zWƕ�lɉ��7��J�U��keY]��|��cL���I��r;�O�R��W;����zI�`�w�CULpg�����8Z8��Vzb_��2Qڥ?�i�j�K�	�ɕ�6��-�k��3�A������0�j�mFj�V��������[	y=�@���楩�����9�v��(�(<��z<I���}��LO��S>J^g�*���Pi���ܷ�ؘy���D]��,��	�a����2	����g�g�T�4�֥
-����V��l�oy���y&S��p���(��ur��>�.g�LlF�b�-��-`��nōeW
OS�ʀ��t�Q�
L�/�N�����:�_2-|���"jߩ�@ 3㠶� 7����Ŋ��A��:V�����Bw]�x<B�׊;c5t	|TU�߶JycM9��I@�y���422�A&�τ�7��.��Y���[j����`�u'iWE��z������j��^��u�A�G��5I�����^SƆx������X����h��{��H��J��/V``�#_C����������{��a�T@�'�@��IE��MN ��f�
���:�l��d����r&d
�H;��:O8d�K�8� �<g���qO"�I���w�ܙ���5� _{v�ԯ�BSv��©֝���j�y}������w�ʹ|C{��c`&:������P�����{k��.���X*�������W��Cov����v�'T8�G��o|�r��sE�����%�H7�AK�b��� �:#>>L�Wm���l�(%,���-""�{�!ߋ��.���`���=������:��y���r�Y�G���b��w���::8�I����GE�Pa,g�zjr%��G4�N�@!e�a[v�(����ѓ܇!S���?AG���偟��~ ��I���Y�b}\uB[G��1az��4-��$�ꅠq8�6�	�;Rp���Ϲ޷gw��/c����̍���]�Yk�x��F�s�y9���� ���G��:\�h�W�/T�&:�<�ֽJ���"`�<(b���7rSz%7Ӱ�L:o����o�Qb{d�D�?2&�D�cJY�hh.P'�i�!r�#DMAkB��|��-�vD�4�F|����K#
B��u���|��e����L ��>U�uƯ]{���LLL~����'I�5�Ӧ������U�S�z�����P�rO��~�DZ����� #+ˬ,����Oȫ�U8�g�:�A�z�(��Y�Np�,�� ��j��+mEG�T�����\TիK�<$���Һ��p�>U0-��i��"�S�^���$ (���.T7�3�6��˅I��nn�s���I
��b��r5�g��A���Ż/�;�`���%J���D��80�C�l�lo�r�n�da�jJ�Ϥ��w��tT� �?�� �������~����u9��CB�Y��;�s���n���)�Y��I��4٬�5�-�!�PG���v������.��pðm��ʐ���~��n]|Dt#߷RyoKފQ��>e-���(;/��u[;MMͧR��+d���J�����05Fּ�(tY�
�ݹ�A���.���޸�5+�P��4I�60�AA���ԙ?gp��ׂݞN�;�Cg1�͚TS��
"=7��m�h��R�d*�t�f�C^��(����z��ЂewwWZ��N�	1��5ȅ�_�X��f����H��S����1mM.M���ٞ"gL2��kG9_`}+#^C�M@_�05 ��B-/��b���Tz�%;%��K�fh���+�B簠g:`�}�W�Uh�ɇ�R��T?���YE�(�\��A]l�6�q�k�I�F�*po�	?[��&�VU���� �\��=p	
z;��&�b=�oF(�����ʹt����=���������pE4��Y�������1�w|�o��3_��h_gC}t���i�+i���9�2�L��Y�qnT��/|R&&�ψ�-�Q�q�B!x���	du �+Tm\�����k^�=��~3Wl�8�{y$���k'�θx+�'���uh�!ue��K�ϊ�?�`J�R���<�kH���;fz���"�-����sW���|�}Τu\m�FG�.X=�.�i`�
�B�U*�2l!���3x%;G9�n� n^)t^��g�����=�+���B k���"�;�h�d��ݗ1��P��G`�"<�y�6�׾��y� ΠP/����ui?�t-���P.�9&�r�7�Y�.s�̮�xwb;o��n��U8iἋ���K��Y���h� �^����b��P�(�q�)u����Xw/�c��^�k��>��|B�ЧB��Ǫ�ޘdĤ��ܗ������|�vʆ�&���H�V J 2W$d��XB�W�(�+;vd�莓4�+�[�mHk���b���uQW+�\O׍��17��FM+kk�Yrx7���5q�dѕ'�p��M�������]�"�]3���'d�bP�.����u����t	@��p��Y�i�2�B b�b�t�l�M6�(`P.o��O��2�Z"�)T�}��]uot?�e��q���`OG<�	�#���z@ȸg��a屴�$Z����~��z��"��%ꓻ���ӍN��v�|�'�꘵l�N�7��XR1�-�W7woqbL��M�B�� g �ߧ;�d���(��k5�B�ٴʊk��A ]�8���3h�q�������"��&sL2`��r���������n�[��˙u:s鲩�pfIm�c˰�����(�[�:֯�H�x�T� WM�8�,V�?)YH[8\	�5�/^e�UX��+��*��I�����;c
��u�tҬB��8K�Z�' �J���dsSè�;���s�ic�������j꧘�6�-Q'Q�j �s'r����n\Q�f�<��bx�}
_y	r��� ��`��˛�(�Ԟp`��o4��r.p6U>�g`��;��{�m.m�6 B���d,{1�H�0�p��E)G����y۳�6^,]8�2�_YubZ��'�[�Ij�8��XZ;�'�3��釨߆����a�Y�e�a��ur�!)h��7��Y��Ö��;�"���[�k&<d�!��çw��s����UkP�8>yqf1���0�ۥ����.h�l2�6EI=���sȢ��ᛱ����R3ck]�p���tD�w����*��7\�*�=�6��=���{�9�E�x��)n7�T����2�q�nG^�@�u�l`yier�L�G��4'EP�'�� �A�ۃ�O����Z�$z�w9Q���M�P=;�""6���o|<�/f�M6�A!8��@����r��ݼF]��aOJ�}������c��X������M�~@���u������Ԕw�R)A��}��j�\�4��^c����� ��t����}��l���I֘����{	m:-��M�bZ�����	Z{��,��D4uWn���2$ş�L�v0��}V!)Irڌ�Aֶ�	r��md#���K����w��:5��y5r�$2����K;�z�Z�r���|��l����6�a29�Qzd�hL#7TP��p�Vz���4nˍ�)�~+FT��U�>a�[?�mHH(ŕ:��x35^,�HK���u�W�)�y���qa@��(�B7z������ӡ��z7V�6����T�TS���$�7M*�DLK���Lxh�h		Ja�E�=�8����V�@?1!3����y!�o����ގOM0пZ7��u�90$��I-±pu�DܧM��m���.*��a�7��(��jc86�"���B�)F�G���"T¡�q޾�5�+�c��?\~�p�}'�,u�:�B��!���Z��P��qb��0��$����竨�j��޵�S"��[�Mi��������J�+����:�/���d�Y��8=S��9�&��VW�&cm�9e��u/3��*c�ZpU���>�̱̳�X���j9��;6
اb�����Ѐߊ�v'��w}Y>��:��5���\%^��A�X��� �c�8B�/�h�8b������!��Jl!I�@3���C{�T��# �Fup��߻�m�"�v��q�dܴ�������}M�~��x�`�@��n����/����JA�h�I���柱l,�R�b�JL�"C�f�`?̻XI��خ �qr�\?���$c,�L�L|�O���E�C\�!���̢R�?�$N��D4�A�l` l|��AWQduQ�i�fB��)�۷c���5��!8Z,h��zM=/�bRiGم��*+�W�,���|�QS��$B�͇����o~��+tEsGaj�w������D��9���T�Rx��a����q&H�<B�a��.�Ǳ�y����i�s@����ۤ�gZ�����H
䋬!������R�dt^��b�Z��0���8�:n~��$�:�)7�����H��v�=k�<v ľ��hӗ�-!�&���������_!A���$x�CH�
�bD:�y���>��-Qܰ��ztXݍ�����ש��6�q�뎓Qy�G��ḯe/�XXE��,�/G����s��T23�a�n���!�x{`˗�Wn5���3��J���O<�
HoQ���p���3�p��R�>��I�3���䉹����ny�X�t��QA�0D��h�,���CN7�DRׁ�B=;X/�u� V�c(�cQ+���e��E'�β�9R&r����-�S'���3�@�k-t4��	���B���g
��a*�\[,M+�K.�pu�|5U��z[�FȀ�Zv)��l��{D�k��_ڄCa��3M�k\��U�f����N�P��8(����AZ�o�#���/
1��z~w^� ̄��_'!����5o�v���eb��茉�;�O(C�t�I��T���も>�@t]U�y0P~/��()6���`��MԴqff�����m�=���$�3�����w�V�~ߕ��Ə�F�3�ÃϪ�E�o����(B��.j����H�pvN�1����Ǩ|2��+Q��>���d�<3/����I�W��9W�U�Ѓ����ܢ�1���m��w��_!�]X2������P��dC�B��k�@Ļf]�����a�u�d��y`#CI���ڣ�>�2V��ҳ���g=��=/���|�
�B�5�f����!xw�]gI�&4YM�]�N�Pk_�_���N��O�ܗ���ʓ9�V�oY��S%�y���D_ �k�,&D�'Q8�䨯Ѷ����"�}	Cw->r�#�h�烰�����H���Eͨ߾����B�<}�D��SF�]@�p��N]�o'�����y���0լ{�]�S�:���a.��S.�Fe�Y��YYٿ~���x��}?]W_��Av�xE�W���#R��p?���.1��tvP$u��1 ?*���d����"�ch� ..�v@�#�������9ʢ�?!�*[K�gfǥ���H���k�+h���W�G�|^�4Ћ)�f�B��zx�6�:��� �:��r
��e��͚��cdQYُq%6oA�=|jڻ���6�� |�R��z�1��E]��Tތ��=�E�Բ`Z�wՅ�K�d�!�3p�G!�*���H�qh�@z�5N�ƪ��Xł�lz��#?�k�3=��Ӓ
9�c������Ғ1r���6�E���R2ﭟb�a���R��o�	dt{	"�|Y�[�F3o�xY�4�|)�1�Eu}	�T��p�֕�{�ld�3�`z������[ךf�z�'���=�L�W�8u�nY��2�Z`F��M{���	�Ȣ[zM���H���xr�(}�pb���Q�����������m��������V������ߋ	Ț0�������pp!*��p��Nu
c�T��җ��)�Q
�ؚ���p��XR ���=.vC=��3�Kf�<�����l�W�uB�UC�D�<�R�%`/\�GM2"�+�.�Hǜk�J//+s�e�:��������@�y6x2b������u��Kr�x5����TU���˘��ػ)��w�F�6j��E� ���*�;&��k�y���S�3�y�E'���Ḙ(@j�(6��`^") �qE��a�Jr��,�����?��8���\�39Sn5�@-&�<��SCd�WFZG�Z̩���׉�6I��Ozx�$Z1�2�}xZ[��t?0TE̔���v�����z�6\��ξV'����hh�,!2��1�(Z�b�3�uH���lPa�
vqW�v�#�u�$����C��Ι��2y��;�2d�;:al��Fa��0�4�ܨxnK�P[��I�I/�j�����u�uݩy&y��n~�8 ����t����0�<��jEa�r8N���x�`�]=(ml������j�`�U�D͗���I6��.Is��J�v��%��GA�W�R5���a��H�6�	�)��_ �B׳�B+�:zd�:���o���)J�<��.�q6!A�7������5�Y�bP��"��� ����-��@�n6�A&<J��uC38,����O=� k����0oO���-���k�θ���(p5�ö���s����'�{�H���w���ZV>�B��A͡�1S�kù���m�etߔp�N"����m��۽������2v�� �=A*??�p�����9	�	?N?/c�������l�Pb;^fS]�z×�o��ֿl6:�:��ܞ�t҅7�~�Ӝ�	8ma���O��t0P!�n�~��uN�����&��:E1�<��$�B���[3�=Q<�)��ڶ2�G���%`.����)Ś�&IU����R���l3�(xF�x��.6f=,�Z�_��M4�lV3�W�[,��*�d���Y���0gQTl��@ ���m�A���|�T��� G������K�jR?�G_�2A(��d"�C?��dz�/=��j��~��x�0��^v�9_CQ�|y���1����Z�"�ޯ��()���e�<��)�c��H�5j���������k���\�i�����q�����
\�`w�[;זƀ��;X���v���ݽ���i��׭VY�;���^��zs���/!�Z���~!t�g��������=7�,<��l�����T�2���@����'崋�<?麳��`P�
��]f���9�db�5��9����d%�0:�<Է/a�T�&-��xa�3�����m��䘨��L��7Z�q�q��e߀��6�~�ǥVq��m�(��v�Q^�/J甆�����a� �5�$�����A�*E�{`[�VF<Cw"0��|��$Ė!+��I���X [�u�a�j˅P�T;f��v�����xE�{^��+�'] �B���O���!���9G�jN#nu�����ɒ �cA�Ƞ�|w<�jq�Ҳ�mE��u��~v��[i��Q��"X��sU�����Xr�S�pܯ<�o�ޗP�\��?x�x��ϲ����R�3���or���	�}	�.��!fK�ޝ<��[|�|�\����j���U��T���vlO$�~̉��ހ-lz�\�V�[�-Ƙ����Z��~��%|��5K%��ҏ Y9�ܲ��Rj6.���N�̬�G$�=�_�$����&�X��%�j�������ع΂����e�p�l�1!�\�le�L�@���C1����1Q�a뿾F[�ܙ�o�Kd��q������ڏ�#���S����N�=�v����\�K��y!�|^A��CH�G�Ln���~z�Yz`�(������*^�2�v���t�YẼ�dќQ�fS�$�zE3�+�J��K�m��q�3��B�w�������IN�Y�+_���G0�A���'~=(���G�Vev��/��B�g�c�l�G�ˠ������$>��`�D��=Ǻ�#/�W^K����G��*����5)�At/�C|���+�����[��υp���	���J��|�~�����U/��t�`Tx%���g���{�d���u���u�noo�ggǇ�6[�7���x8�0����pQ߼��A�jFj��O�G` �����q�v��A��D�5wWu�py~�c�R��yN�~�X=����dTJu�&�w�̥�
i�"��a׏�wێծ�	u�R�h�F��Ȓ^�j\j���/�(8D���h�z�����^{>"q�^3��ԉ$�����8�U'�s�f\�/b�Nj�*\I,F87�����c6��n�x�
����}�����>��ADձ��F����(*T�T?	�)���Fy�ʶ�Zi���)��dh�~��	�X2�%P���$:열���`�j�!�4> �zs=��O.�|��up�s�߶#J�L�n'��W��p�I�p�'�g������H<�(��]7�/��a��?c��y��.�wZ.P�
K���fnD����<�h,I��F.*�Xލ�Q땰m�ZO�[�a����k3T
�l\��}66[�<'˕�ѻ+-v��o�3���/1�ď�[iS�tD�YOwJ�#ũ�Y &MৌlA��+gf��C�D�B��`���sh�fDd�܏�pK����65ʶ�g�X6�I���i�������C�L���4�6\1i���b*8P6��s�3<Gx��������#��J`h�e�i�6��P��$��v�s����pk��pE�Ǭ>i#�|Pg�ծ�;�7)��,{Mg���DD"#�nsa�~�c��;��5�^?���~6�1�;�r|gT��H�'�0Ȩ�����p点Z��*$*��`}�\�ȗҍ�u.x�4�x�:w�.I�Lw�x.�S�˵(�v��*�"N�Nd�ƀ�Gt�O�����U�����uz2��t�	\(ʻ^[�5g|�N��rV�&��e���{�X0�@ʶl��
&l��H�xȡ0]�V������C�R���:�؞�����������Ђݺ\�nL��H`jm��4=ۻ�[_W�X3S�IC7l  ����K����ݮ�SH��"$5p�+��9Of�@���w4	� �d��|�|�#fR�'�Whᬅ�-���}*���6�,�!�6�֞X1����V���R�a���]��wJ��#�:�rXt>?٭�T�R|u�g��1��p��v�ַ�Sa+�`MUU�䤓�U����)D�}���ҁ��M��q\]����f7��Ib�ȳDc` �$Dd-F�{ l(���{ź�h�aM�ض�� r@f��=u�
�^t�F�)7�+R���3kǾ�b�|"Fߟ���x/��<nW��ם�k L[AG�ޞ�/�.P�2� <0���Ճ�!)�y���#�]�L��1����I��%�ibS%7ߵ�j(s�#��Y����#>v���OS��ZA��b��$�d�>��/w�_�t���t?�,CN_<��#W�^�Lt]xY8��[6����ۨ�����o�ju:��Ka�oM��օva�:.mgͱR�`��M���C9�ާ�g�ͽԒ�B�%��5>�]O� �u��0��5h�� �0:&����犢x��,�G�L���gw�;�ҟ"+"/_����{������W"��8G<O�߸�K���ϒ�z��������C��m�+��=��8�:5�đF��I�+�ͣ��a"����wԶ���F�����r��N�}Ze�73}�icZ�T�0:�N:�Y���
�gEoO���X��U�#�Ug�[m�
����o� c�`C�Ho@�c(������y�Ȫ��Ng��_�Ԇ�"T�O/�b���P� oqA�1�T�'0����,�f��MFCH��3��júI7��f�0~H�o��))i�w �0��Ә>�Q��M�Kn���Oz���Z�3׷�.r�Z��j��>���B{53Va�r��y �R:��<BQk�jt�.j�m��l�RT� �@~�D�
�o۱���X��0	���{�#D���s�e7�o�:����AQP?�GP=,Z�D/���\~XtT��3�C/z��nȝ�t��8X�=�H����t��� z���S�A0�;�,�����;�+�Kgp���JUQ�%YV��zV3�㪬�mYꜪ���44��ŋ���ʀ�7�g�,�?�i�MզY���!��'��Q�܈����mnn�---�.�_T���A
/�S��^���5
>�Hbt���Ui��#��7��X���fe�Rb�o�`���qjQ�j�W�n�I�����z��Lp���}���Wav��F���g!� <t��#�}Æ�qx����4�;:ȰN�q����j�Z�̫��&''��_��_���h���*	��7r��g9r���[�n}��i<��������v�<E��[����o�,Qlx ���0� �"� ���P�P�s��P��?B��IW;�/�
mւ\:~��w���\�c��ϱ2f�graȝ
�B��^��xQ�� / �60'�K�L��D5s������GT�r�e|�;�LQ �qA
�ҹ��/��*�V��89ETC�\� ������DƲN�1'IR�駟���kN�8���y?�x�Mv�~�ݶ3tu�$�Ò�@Ūb�-�
~�h�d�G���aT�j�� '��ރ� qad	 �	5�%�2�\�`��W�&.�h�_w��N��������v���~a�~�u.��z�N#z/Gg&t�?.3������B� ��ٯ����;�b��ٳ�=��#�&@'}�'���4E$�]�z��u�M΂)+XC3����ƍS���~v�*�wy��ߥ�����KG����[o}���������M�61�2��
C ��!r�T�LGC�{lx�`h`
y$�_�q��I"τ�3�Q�«�{�w�M2�m; ��v�z�A��j�̰�T�*{T���>�W8�	���h����G�2Y���pǗ�;�"d��{�4u����9IQ{N��u+�#�K�\j���a,�9A�K�6A��xT9w�yT�KLS9#�(�����тw.1����IQN��R:�����KO?����---�*�ŉ�����ޯ(�^�0�ꆾAQ�"c^
9M�Ë��  ��\�@-&����N�s��a�Vk5�9�ي�t2"�٣Z\D�Dx=j@�C�lB �&��2[ų�z�Q��m��U"DH爰}O�w�(�J� z��ƺ�1F����5�����?�?W�8�����c��|�c�>LiC :�g<n�D=t谓Q�@���chK-��׳i�ٶm�_~�S�Z\K:�n�� ��$�F�0�����}ǎ��.]�t��nmںm3��W��Pdo��: �C�a�C��;,Y�lE���A�"I�a��E:�-�|��-T��͂�T�������(N(Tt�ܳ�-�J�������ݢ�VЅ�Q6�{����r�z��v8��� {<�B=&�Zݮl��$ ]pIG���81�U�_���^K��E�>�E-@�w����? �7�x�8�i�U泲���xMՔ��ŷ���̓�1���-�N�Z���fm��돨��C��)��Al�u]W�6� 7�\�Bn0�R	o|nn���p<i@�:7;M�+�.�Ճ��Ԅ����V�SD$0��qƣb}�*f�5��
��÷���-�.��#��~`*V����}�1��x�A��z�w�ۺA��{�q0�+f ��ncs��M��O���@G ���U �ߟ�:���vϟ�5�����ʥB.��{���?�R��^�(�{��<����϶}�{���.\�)��LSg���$+5�N������>G�G;ٞ��(4P�"����NU[�;<ux� �A�;�A(Yk�Z����H�t�Iᚻx/{���j�F9t�4�]s`S��k�r�T���b��q���#
G(����ݦ���G��8#SE�y���e��`���g��A�b��a�ч���� ������s�,�N��+�T�ao�飯qJ���'?���@�����]��\n�0�m��>b��㲢lM�S���e=ϣ�6�z�	\#���gx���1��u�b�� n^��A�n5B @D�\wPw�������n���]��Ez�V~n��-L��l��ޖ�0#�^{��]�WEy�<��� x��#�%^���ď��8�E�V�� ő�7o$g�� @'�6ȡc�#�������T5�82n\�F��^���m��͘8>>��~����dw����$ ��~��O���K��h4���+�m����R�'X��>�C���B�����n4̏��\(JT
�#B� 2<6J�<��>����&p��6P6�! ����0` �;�0�_X @o�-tU��=1���e�V�>�&tѶ�~�<�����'�a!y
�����;yK� �":!���p�M�d�2���8�(�C
F�i����+�B�a���u�ԴW5M�Se�СCb�����ȑ#&�8�3$I�FM�K�R���QU�	I�
�ĲP��y;/��9���N.+-���Q�.�E��0l�mγV�賏�l<����X���ܩʝ� �j�6~n0�E������)�xaHƍ�^�QPeC���{ tZK1���.��+.ql�������; :��m��y���#IO	9t�S��m��F��7�`�3Ӥ'W�Km�m���fo��m�:t�'�X'���Ƀ�������L|���ǧN��U�A��r�o���W�^a7op�6��8��`iRYP�s���^�R�;��MNn �FhOx�8>�$��<l��7C�-��oMO�;�K�.�
���jP���D<���.ږr甏�ikq��~@GQ(�ųJQ� $��	���u�C�>G$"�+ �{�C3�}�o�_�>O@g+<z��{����7��ea�U2�쭔a�Ue�ah/�>~y�X+�ͺ���r.��=�3[�V��m��&˲�ɲ���H[eY�dL�K���]�5` b��G�Y:����Hޕ2
�x��G�B��(��2�htDӉgt�>2$@P�:�`tjx��L���&� p� ����9{s�^0�$�a��Ѓ�F�~��{46G=f(��
��X����|�����x�
���~����9�}1�����a�ڵ����� ��N'0d#:� ��+Ԡ�m��:����}�3�M۶_�j>�~����w)�Y[ � ��z�t7_��׷���7/^��z���kA断�hsߺu��J�r,v��\��0����
�6���M�(�*ux8�R��C���d)R�;EY^Z���>2<6�._�¾������C'e����s�Q��kd���}�*�!���,�8���C�z��b���38�� ho�y����'����n�л����.���Aѿc� s*��zig�ǎ�A���L&SI�Ƃ���TEyU��z�X�}�wm[�t:�����4m��(���
�"��UU/�$ ��3N�����X�0�z�Ty�x����),�袀�d�&�?^0>SD$p]!��y�W�H|��"9�~�ܯ��g��Z���QO\�G�޵�םHć������]n������ �9���;��h�A�}Q�����{?n؄����{�^B�����?�w7�;���Ӌx�^���J�V�;v�5�5�k��ߨu:�wF����/}��=)�5tP�k�a��|�k_{����˗/����"=CMS��P1�/ˬ���K.���X�T��u��i�V�M��b<*��))i�*h���R*WI���B�L-p���j���ŋ쥗�2��	СtEȝưDV�PH�QB�8�����lx�!.q]�2J��OY������>Lq��#�6�#��܍�& �c]�Q��
80��i,���ca�����Q� 4B�|��s�,˪Z�VƐY�� �r;6��|*�*�V��Ke�Y�V���I�����J��u�a�"@0Q�&��
�Ӳi=	�Q�OA���G�v�U�[��$wz��@0B~�vF2 �a�]��F� �-�Rū0{����{/ޭ\�oH�@�Y#}���ю֕Iod@�'��D���o�}���ЭVB�5\9��TR�}�OƷ��?����؁���?�v��8.��c/�tE�)(��Vo��_~�9>����ke����X��/}�W��=�{�丵#��}�kO>��sr���'�������L&�R2+渇Ľ9�������G�nؼ��T0��l��f�q��������S���r��t&,�C�^�R���D����\a��A�T�@
�k�!�pi�۝`& ��
�z�7��oS}<|R�^L��j�. C(�n������x]�+ZM- �kbr�O��P :U ���y�g�ǹ �)C�stnO�R�����(�aJ�T� �	f��u"����=��+�x:���L�P���^��âb��x�=Qx@�A�= t��)�.<�(������`�a�-��o�{�n�z�9�b�j��Vt�ѵ$<���D<�8Ȓ��o7V��Ǎ����� ��'�cVtԅ<��A�m[7�;�#>���'����(n�RgǏG��֍���$���b�Ϟy��kG��۝$�~orZ3G}��_W~�����.]�� +���k��ar�i�ʬ��:m�-ޯ�����iӠ����[ɻ_^)S�:���!n+�矋|;���M��H[)�H t���y�T� ��_!@��
!�w����AJ,��&���sJ�+x�a�=��I<~@�+�a�t�@$�n���nU��p��)�C��h�>j"!d�Dc�)�.���� ]��&�R(b�����Is��@��f�<t�smjP��H����h�p�U�x���
��E%ZE8�h;�N�#�#�p�vYt8���3�!"7+r�q'\ :��@���Ud�\��������DZ�蹋z��ND���ܥ�눾�m��Q4�'���z�H����!fD'�x�1�M��"Cn�w=t��:_�>[.U�(&�����\����Å��_��Q��x#	�ߣ���a�p��c?s��˿w���mb��v��mlӆ�S��j��z� 0�A�j�J��l�D
/ �R����6<2�[�$���B^��a���� @��Ekw��-��B���W�3�0X&���7Ecס0|�3"�,��Z����g���Ѓ�^��}Zw��Uh  uci�P%�n�x����V���z�{�h���XTى�{��)�"�łn������eL,s��Fn���4���'�	�c���58޴�0/��Sk��.�ɍIQl	2!Q����u�k/yRX�5���f���g�醟-hg�z�}�m���"�}��	ɒ� ݔQ�3�G@���(�w����ta����N�=��$��.:���x�?2��w��Vq��:�?z�+��w���C��G��Sy�=��4B����h[����D0�@tا� �i�^�p���,s���W��i��+�u��p�/��b�����_:��[�tnnn�Q�
���m۶R��H1^���9��@�.//R�|���b�L�A��������-(�����R��C/ �h��ls�6	�ֹbE�5B� �Б�;��k�������!b��q�4p�����XǨ7J����_.�ຫY�}�x�" �?;�	j�p�i-(^e�㭑9ϱָ����B|�h�6�%!E��ŭ�r	KĹ�^�u	x=��y�%�� �0��@�:
�oW�Lw������Ks�7�K�������FA�J,��k4�t}���wUE��#{1������J�f�m5���� �"c�<�ۈ�"o2��ֶ��C�5z��톈e�ԅ!���֔U�<�7��<�Q|�S=�H��[����r�M9D��'��F�RZ`��;��P�CDY���n��,��r�I�u{����3a�޸y�Z����m���_XW-k�\���-	9��{�~����~nnn�Qk��"��MIC����5@�,��Ûk5lV���-��.�V��<[�N��乩����,��؉�_cgϞcF:�
����	<I��1G�UX�����.�RX@�
�a��88D����n�͕��R t��4�8X���.�.�hў%欋a00�����ϟ�,���W��iq�.,�C�Re�f��T�d��p$�xݢM(e0�	o[�U<�;��T�S�G���3���^Ş����hD�����1r#q@�����}�s��!S��i���xu�X���"$K�_Ȉ'��c�:�B���E�3�_V{J`�D[�G?�;x� *rK���ʁG�p��f����M�-6tZ�R�^�z��h������_��_V���;��=n�u�y>�7��o{����Go�>�����a��e�P)�7l�����a�l~a�r���޹s;yl |RY^,�F��T]'��O�R=~^(k��,����@&(|�[x��V� �w��I����ԙ�폎+�Q+]x��ӌ�'��W�TzH��V�Ɓ��z\	��{�T�Q@'E�!a4b�5}P5X"�/%<m<1uOp��Y�	� a� ЩB=�@�T���h���2��㔿��%��g ѫ"��pY����"�K�����P�f���=k�;���9�"r������w���)�(�u���������W����n����(�-�Q�nJ��Ŝ��B����g��<�e��f�_�O|��۷/,�e.��������]� ݸz��={���R��^z����g�9ǟ}��^V�{^S�������+�[5��w_�ͷN���ss�E *�#,�]�v�\.�s�KK�X�P)%Z��������͓��(,�����B~[̌���"�}Ŧ��U�nw�6��Q@�՛��s��rY���C�^}J!�U�s�)FFY�w1�,� �� ��<�nȝ_El�~�[U)��U���b(Q%>S�B�&d�t�>��rPT��{�C�y�"�y�ybj���X�$�Jy%�bV����� ��h|�+�"y�\��� �5�������߭���f���~7@�Fw��ҫR�/���!�F�5�n�����W�(��g :EQ�|x?CX z���d�Ċ���ط�S!\�aQ�*�v���O��{�R䐮Ԏ�Z1A �����s��\ R���оp��wdY���/���?����oJ �>?�w{���������o�=������u�<g��,Uо"���׎V6(pA��~`A���b~����\���c�BӾ���Pn@� :�`�J�F�~��g�M�䨮�����fF�hG	�¾l�!�'|Yl�'��?�����9_'|�cb�l��!�1A�ٱٵ�ІB��Kh׌f����sOթ�U]=Zg���f����֭{�{޳n�d*kkLee���%L*Õ�8�&j�"�N��5����f�0P���͵b�G��]��
�<��b���D��e�������]v��zV
tL%�.? �J�5�A��vؓ�    IDAT����p`��`-�NΖ�y�x6R��Xw���͏�w���(`Ԥ�9)p�*�ߋL/��G�F+����4.C�>�q�Є�� ��u�n�X��hS���`��S��~37��0n������_�G���ұed�ۜy�x��O~���K�{������ Ѝ1�׬��, =۷oo]�r�+%�%��/���T6�����7<��ᱧ������j���߿�BL�0��;�tuu`��#(�����!��J��c,t�� ֥�R�͔���\VF�A�U���I�qll@`�3H1B�13tt��1�}����-[����ZS^VmP��v�Fb=�Q��Ѐ../�
� N�D���@���w�>�|�앮�S�q�̡fra���t� �$E�����Pv^�L��Q`ۑ�܎�����v���u��sd;٧����qn��`]�U#@������y�������%&w��{�X"������X����V"%O?Jq��]�INGt�P�����=�{K�%�F� ��"
*�<���E���	�ǌC�+���j���-��C5�a͊�0��iӦ�+W�~������ǿ_���k��^�(��c�=4f֜���Y��3�*�ve�Y�*vEE9	d���)R��$Z__�#Q��#�L9���aZ��uJ�6� d�Y�遀,�[QQI
Ŏ�����ر���0e�Udr����&Q�+�ıR�܋>�t�����3RB��������?�b.���WH~4Khf��cP"熒K��*���]���5 �M5��pK�Np�v�m1�u�c=+g	�� �Q�y~.h�}7-,*x��ݑT��:�>�<�	i^�`���+��k��
`ؼ�`���iP�����=P���8��O!�Q3�0�����0��J�UW]E�ZG�c�I�& �-@~%yՇ�I���r���֮Y�TYY�����o�Ѯ�S��~@?���~䑟��9{�֯����Ù�vnZ1z�h�����|��e$���ށ6��R�5��� ���q"��{6mF�L nM������׀�y�6�����z��A�$SF���p:������<�5�
����\�C�
Q=��k��{�=�]��RH`&,���q�zF�\��Wл;:m#�.2��܎�H(F Ӄ��իW��Q"���P��@�N��	�YT޲�戹S������le�=TȊ�?��?>&�0�};��y#v}�.��f�ϥ\�"a����P�]�'�ә*x��_d�T��*vA�l�J�"���/{�UV��D�A���O}��pa��S3Q/��,�S�����% }ݺu{�oX�hUE��������z�!����I�=��}��}�G�6o����9��50*h���DP4�E���t���43:^��$�(�'�`Ӻ��N�,��T-5;�����(l&����7�6[�n'�����MU� t���À�[	��nOa�����cAar�bb��Z('m�ha �S��Q>ܔ�@$��1a�����l������~�Ȓ��QW�..,�/ lF���1Q�!�?.���K��3���	�� k%�mZ��q����/�4lψ�v΀��`	�[/&:���Xc5e��
���$ύkqL���d�\z���W|�HM:͖?\W��P��vz�����׭ZM&w��Z�jצ�8�����ۿ�^�#�u������衇~6q��Ywoܼ骖��d�;G 
�5y�dSYYAt����/��b
���#=I"�)�-S�1,,pzb�v�i�y�g-������h��߰�z��6S]_G
����b�"���֩s��8T8:�<t��ى:�����=��{�*`�^r|!@�襥
��Ѓ5Bn���r3k�,��s�Pv�� ��L�t4&�`�1Ak���>�cz���=t}F���#�+z6�<n��8��?V8��G��kQ	(��Ďz���5�R
�M�v<��$2�v���T���+/ro&P=m.��rs��.�fP��}��Dh,�CBq]�r��"�hժU[w����!���_��"Y�:��{���/�ˉ���{6�_աC�������TX�`�Cׯ_O x��?F�� 0��0���@Гk�����s�Q�`�N��F2c�\��,y�i=�ij�t��dU󇬭E�b�&vU�bm�jJ���8 z���yi=!����Yk!�Ъ@�!]�å`�;���Ǎ5���Q��40Ƈ �C����̝;�>��u�J[�Y�Mr���O\�����Jw���YX4h���9�� �"0����"ꤱ9Ct�{�k@֧��U���:,�Z���]#l�� 9��-�e�a��( ��gonYj���K/��46"����|s������m�	�)�J�A«V��p��������[n�su�i��f������~�Ȥ����woذ�J0�6n���5�m��
@6��4Q�,rEE��!�9�}�~�&ߛf��f�MA������8W�klD�p�����>4�흦U�� t�.�k���j��*R�����<}���~�;6���ps�]@]�R�2�Ed����G�@�+С��w��4�����h�|���O��c$�d&C>t|���C+ݫ�K!@�`Oҗ ��q�E�0����u�b�{|�=r={%��v���z��A
w��u�|v�jpJ3��'"��<��Ț����O_c.��b�k�$w����Ǝ��,/��������L@rV�X�����GC�4<y�M7�+F���c���=����{��͘9�G;vl����[�	Б���
�&Q�0�"�����r���{���Z�ަT �����z�`Z�^ƌpР!���ּ�l��p�J���e*k�L2���5 :�5�O�НJT��bV%.�tA�) F��vM�QAq:J_�6��}��ܞ�vzc�cp^��[�:�_�PG�%l���֌�d�z�u��SO��F��Bك��+ąK��|�
U�k@�(�@�)����O6�z��]��>~]�a�d���Kj�a�ޝO��(��������\���Z"�6�u$��5�{�!��R�9	<�D�44Ԛn����IQM$2�̻��*�i�Tֺ�������7�7m�:8�X����\���C�����}�@������Џ|���|��;w��u ���o�Y���U*m�$3.upbaa\�͏V�ٺݎ����n�v@G�	��9�sȐ��]�x�Y�j���ʚ��Z�R��*ѯ�S��;~ls��>8t�o&�TAT^wج��C:���Ezx����r���p��t���!)����8x���C�9sg�K� \z�gm���h��(@�2�dp�+M�8�ڌ��9��gK��L�>��Eҽ�����Vt��,������
O�t ]Ʃ=L�����/N= �u�z������{2g�7��7���=�d\*���N�ET��\J�	ݿg�ٹc��hoo�^����D�uu�o|�_�s��hn�q7��$��=��y�ٳ�ڶm�䟷n�44D��_{{�WP��?�����B%�OnO<��v��YP#��WS�0b���]hV�YG�=�M �䁊�F @(�N�_[)N�}M�,��  |%��&4�X�~���H������|-���Y߷^R�P��n�P Ⴁ:�Æ�:�X�������l޼���t裂A	�A��(ؘ	�����b����2�TD��� ��.�N���(���gT�!_I*W,����m���u����c��z㗎9��E�ݴ�D��Ța����3e�Tۉ������u1P�]��!�0���h����G��[ZZږ/_>'�H�pԨaso��F���q�}n�Ѐs�\⮻n�n���?ؾ}��(Չ�2��"()I"�!ĩ��-�38��jnc���. ��[X:UTJ0��^~OR�p8Aq�ֱi �Јg�yǬ[������5>��+	��M���䃧����L'�	�o�O((+�2�wӨ�侧M�aK�"J���j�N�	0uz�,x_ ]-QP��Y�8@��w�P����Hk,�������kj�ͪ�+���'jX{ŅP��օ��r���K� �F.��3��8<k�)r�.i��-O��=�zbk$����g��{�Xz�|�]ֵ;F<�0e�=��\mP�
����u>O1H�D�� �օ�K�Pm�:7_�c;�93z�p��7�ΙLk)���=E�N.�D� /�#�H���}{�R�fsssˇ�>|=�H�1t���7�t�����=��f^~��?�1k�w�Z��)�'��Hې|r�ҥz�/����#�B���Ƒ"!)ʓ��HV q�pw�������B�9|���EK͚��MIY�I�T�]g) ���EC���jD���)��r��%e�ݿ��g�c�����5�#����]_`]�kA j������s�~�A_�/18�ܡN^�ۦ*��L[�=
8b��v�" 	�sl���������T]YeΞt	���<5�	R��+o(C��!�ºǱɗc4":��=?��[�a�5���1�-
���X�b��y�]ˍk��q+�U6b�� p�����p�L��=����q���ɼt�`WE:g2�)� ��`�P�T	�訤+2c�9�)˘�g�n>}ݵ\�`C�Θ��N2�����ܓ��%%�\X&g��vQA%T�ܾ}��5k־R^Qv��-[��Nk��~@?^;�$�gÆe�?��?~��7�����7�v�9�PZ�h��4���I
�lPt4��j`��:o4^*胵�6Gb����i�����������,L�Z���(&R��^���*-h��!E>� (@˃l�B�L�t����,��Y@���w��ک�A`�?h���
StA��!gV��0���P�Q[[M�Ǎg���g~�!3��wh�󁇕��,Xh]8R��W:E�W0�(b�O�.�O���+
�}ޮ�]��}^/]�Rϩ~/K֖l^\��s�gX�СT�{a"��>��{�Lg�&k7'�C�R]��X&��3�{�<CD��뮥5�I�d5[�:۳�c؇.�J�� �-[6��ܺu�5��<_Y]y�_}�+KO�8?!���2�'�s�̩~��4s��o677����T"E��L��ne�8�L]@w��~��ϳ~��=����FU��Z�yc�?f�X���ɽ��¤2�F �$Kб95Ct���v!@��!h� ּ_���t<���	��ﻀ���T�ߕ~�컓�> � zX�0D\v�H�=a��s��Z(�G�@���P��-[fz�A�q�Fb>��}skR��Sj\@�R|���}�^�P��f:�O���+����L�G�1��(q�j�6K���&�<��@a#�a��$�ɏߖ�5��Z���0��ӳ� Y��A�0��,x9�`!�M܇X��H�T��ܻ��טQ#G��oC����m��	@n�L�W0ar߱c��q��=k׭�^WY�_���+�ǳ?���S1�Gy��_�ᥗ����޽���u8E��u����s�%_�0ht�0��/����g���8N:3M�j���wv����n���N��R&ǭVmd:L�؈s�~�lܰٔUT����P����@)踶tM�*q�0�gV 	K���RzRϓ'̔�W����|��
Cg+D�L�.��N�����rٖ䁳�=�@n[@����c�ԩt�3f�_��G��W����`%�@��C��cZ)�-Ѕ�G*q1k�hr?ʭ�}-N!��\�>6���%L9�&3x4C�t���{~1�k@/�����[��`��LH�I������N����4eUe��/0����4U��dY��`��t��	��ܑDVxԻw�6���!��ڵkw�[���A�����7���,B��uM��$��K/M��o}s�{K���|x�Š9�G�T�0eS���tn坓�3��f�V�1�'�.�W�m-������\�!E)QH��}��a�>���-���������U�H#/`r�`%y�to6�=�8�2�Sg�I�gBQW�APG�ƈ�ͥ�Z�>����z�4;
�����&~< :�Ժ�:��C�۾}�y��g���?�B�t��Z����,��y�Nt�X���1���!O#.H.PO�֍�~���c� 9�	�V!��KǠ�q�������1�c.�yV1'�#&������t(�PP�T��.��\���Mc}��l(댙x���p0q�~	@o>x�d�ʕ+��Y����}��_�|��ŉ:?C?Q3{���ӿ�����q���ɡCP�p֐>t)�@6?a�Q� :5�~X���X���v�`3@�QF� )����Qۑv�0#G�0GZ�̌Y�̶�;Lum�ɔ�Sa�ߐ���M�l�gp�K�.\1��+\xt��m��d��s����zသB��5a�8t�t�+p@�ϝ>���t�^ؒ��X�AE4J3T�����6Λ7�L�>�̝;�����Z�'�h��h@�q��w�ۋr9�s��=ND��tz
;�gꮀBocP��خB ��u��Q��6����3u
��Hw��ɝ�yRpi�-��.�&C���4�H��슏�+������L�*������T�C ]���͇��-۲f��:������m�{n���~@�O&d\�<2m����j���9�R��' �S�l�B�F�J��5���.�Ŵͬ��;6L��o�48�$%S��0����2+��G�:���Ϛ5�l߶���0�����Щզ�5�@�0��7��4y&�(�#@S�kAF�T�΂�g��H�`/���������)l���P`�&�9""�ܚ�)��X�!��l�c�ujH��V�P J�>���7/�D��5�6ȉ��6(�>c��I
����{����(h��;/�����Q��ǐ���X�w�b���]`�Ɲ �B���Nk�~�ݭ3�}��]9�	�ν��Ӿ	s�4�m]��`�>���
/^L6P��L�#Fg@��JS^^���f�d��\���4�Ұ�� �Ȯ]�L���oK�.ݸzժ���{����7���~@�O&d\<��i3g����k��p�HK��MҜy��c�I)�P� 6w��ߔj���M�$	l���Y�3p���K+DK) �8nĈQf��}������;LMu�I��P�8�<Ora0}w�k!+������fh7�<_�^�e,��2�<Ɠ�"`�'w�e袜ty�ڷ��F�1t�&�2�L�U�4oM��P���iӦ��������c�6m��l@w���h@�{�0��q��j@w��wTR,���~�p��w���;�W���lg��K,����Z�u%�6ݶ:��,�8��۟��imm1�Tʌ7�\v�e�+?aJK��:��w]��L��JL�yЗ,Y�v��U?6��ѯ��}�1�W³��C����Ǽ��ooߺm۵--͕�,��!�.q�(vm��<O��0�ZǶ�1���[[��!�Х�%�ɛ�$��ѧTX&�m��&��2�7o1.�&%�
SR^F5�y��5�����u�b�!-(�
/qJ����ʧ-ց(��
�e����Fȟ���ф�xLǉR�S��s&�D���
�t��r�_=z�HZ'K�[l��>�z�J:���rOi�@��K��5�f���0����UB��@�����t�+Zas)�|��g򏻷8�Û��ֿ�X+��!�G?ﬂ��Xć�?���6WR��B�|�a��0�MJ=1���>����9������A2d��s�E�\L�Se\�d��UJ�,0v�0��P/����?�i��2�Y �hѢ�6l�wx��'��o�fo�s뭟�zo}2!�����9���^�}��-�9�R�����L��fp,�Z��T{��� t,|,n(
R�M����~=�@
ՠ�L�Y1��WWך�C��-[����#���lNL�a%>����    IDAT%�JP\��#J�*��1���t� 5WH�2��v��0.�s�I E�d�; t��UV���}�9���?����<`���˅7ʐ���^��6p��&��B̪|^��j��zDz����b��'"��z!e����{�Ŋ�}�R�&r�
�g%�ܤ	��:�C�/�����谮#���K/�֩4���_��C�<@�&�G��f�����*,X���-[�4h�3��Ɨ�dc�o=Y��Ǟ��6�'g���o�ڴe�m�G� Ε�Ԕ�.]��R��q8m�eK'�P�b�Ng�`��`�����@�u8D�XM�,XD���0p�3��O���q����MA�8]�Ư-����a� "��Sί������ڇ��>B7�(�������
�T����*��$���]J�L�eTT_��g�����AP��n���khi�C`h���A�F�s ������Y��p����Y���}]��ｷ�sGO��zK��eϿ�Pq%�~�M@�Q`JKq������^�M���|1������	�M��wק)nџq����k�nrєS�VO����_�!��۰�֬,f\�2����x�:����&���h�	���A�U�NjL�*��X +��Kק��mƗ,���8M��ִ9w�g�^>�K��[Ӻ�sO@��w�@�Z�ْ���+\���^.�|�Y�Z8��+}$[��bb�N�����N1Mb�.Q7���?��G|�~�B����(��غi��@ڝh4�L�f�J�??��uJ^}��Q�	h�I���Z�?b���5rs��9�cI�7��D����/j�b1�����R�*WRV��i�9���9��ǫ��˕��i�w���`��	�`�Xr��l`�G�����@�Q�<���S2�G���3���;��:��@���p��I�3�/��y�-q��c[��pd�υ]ۆL�@���)Y�Is�abb�4r7�`��$�W��K���z��/aЀ����'p���']�q�k�N���g����tT�}�K�j�L���r���}'�Zl�dvt��`���&�x���yd1)��eL���j�_�guSNַ����q�p_ԓlF�X}�0�K|:��T5�1cV�j�p��N�3�\���X�V����<*��=��/��i��
��Xݬ���Y���#�
���D�����`x0��������{{Jh�zoJ�2-0���uM|z���CSS;��3�:�҆�+'-#�}*����a������T�k�w���������4�t9��_�����P�q�A���^r_��B'����E��+�
,^Z{ $�B�:S��.l������� 0�2UO�[������^��le���U�R�̥�{C3�e�abc�m�<�ߎv�c}g�k�0t?����|�7��P��tU�/uO�Ba�E7��Oё��v������,B����BiO�js��Ն3΋���z�l�Z�V�o���g����~�� �h������|my,�O0��%��ة0Z����z��o�+
��P�9��JGmd��f^ ����������t8L�*C���<���4! ��-���&U�M���0 <��ho��e+�L�QG�lS�d���3�t�2!����� ���֝4�Y�N�f�`_JXdp����8�L�������|s<7ُ�H�,�|����MN������$|W)�^$ �E��{�@$5 k�)�%M�����#��ؒн&Xe}���֕�kYe�5�B������a�p�x��
��G"	i���EǞ���~��˛w<�Xw�]���%�L�m=�	z�M���ڟ9�����T�{�L�����Uv��f��kˇc9K&���1�#
Q���hU�j���@�)CqW��8>aƔ48�9ͷ�Á��:���&��|SW����l	���$[
u"0n��oJ.y^�G�=BzH�hc<��ҵ8R�/�c�ϴ8l8`�3�FB38����}� �~ILLWː���K� ���z�� �=r�M��m	���)���A��g`ܘ�lc��<W��0�DX�kpA�K.5F��C��|�a����d���� ZF6��Ct�R�(t�W�߸]�(ˉ�p6Wt �1��{=�[�����D��������F����]��%Z��&IJ���^<zիq*,���H��������V=�����궖�n�񂽬��� F�_b�e��(t�c&(�Z	@��Rl`h�>͕�S��宨-e��-�x\J|�]�����SI#4~�&x�&m4K>2k
</i7��7��W#�%�t�(��ё��c.�!�=I��?�%)���p�*���*(�;(�"b�J�Ƿ�^�ByX��=|`��Y���/��TG�ġ4���ʊ|JL��
j�/���u�7����I���s҃\!q�;�z�}E����EyJ�J۱d"�W��JLќb�$��D��
� #?�k�.s��Ʊ {�}�`H��O:b�l,�g=�N�r�������ki�|�`��М�Ц�f+7Cz�] 05�����C�����g~��#�����U���^�����2]��ʈ,?���W4NTu<L�	Z�=�����������R.��b"��?a���f1)i� l�E�tW ��#�q\�!U@�k����y=� ~���xpc�v�Sc�ڑ��@4K��W�s��q�B1��R��w'^����aN��&�p>�˙��H	%�x�af���F$��^{�@x@�8�[�w��xqG�&�����|z�1#̼K��@똫�eL����(�����%\�U���]hrap�j/����*�q|?$x,'n�u���9��}�������U[
��9�����嚂�U�)=gOG\K�Կ�z��=���e�ؕ/W�k�0:�Z%f#��Ғ��H��ϲJ��/�
w�Lv���]���g�*�aa���F��4AUg5�5�ʩ�PRP�o���٤{4G���S�ci�����5	�ޚ�\��+�|�:Z�Ɔ%��$��SSS���0��*o§^�Z٫�[<?W=ԣ�Ȧ���b��Q추/覹����Pd��xC�حEx�c1�(�@��w{���~���@C��3ֈ���@��L��=����������t�]��i��z �P��4D��&�S�ْ�S���$}����J�L"Y=�!�	��Ć�Ł�U��O(�1 A#iF�>�Q�zk*!�E�U��"s�e�v@��7�������;��P��~v�%�L��Sf�Lng!d�\�qQ��|Z7��4W����8��{��
�,�)wb�7
֏��5���Kp�������aӇ��<Gg�Jz�߆6�$gU���^Y��伻�cϚ|d��[��O�رs$W��b�6B`����`�9v��b|�nut�5�\-NH���\P��z�j�:X8���S���B�"|C�z���\�� ���'^��Y0vU=�g��
����*0��.f�u�o�����`��㍿tӮ�l뙞A��1t0G{v��0�F��{w��oUO�{JZ���i7X<sN��`��;?��V�1�Hѯ~i�������@+��������j��<�j��{���m� �v\��;�$�o���U�r�eqAT��v�}%���x�'�=lX�4�%tYo܈;.��p{�Y?�2���������ή<����Mgͭ���!hb����� �w~�Ӹ����L�0���W��s5��ί�4�P��u>Nپ�x���<%tߌ>q�'cIdٔ���k3�V�c�L�j웸UO�*:���a����/V�/��۰�=@�2�z>��C��܏aEWM�2���]�"0�v�i^�TQ�s�F�_����/u�u��_ȼ-:�����r����f���R*��x	�a������9Vxe�I߈�ܪp�}_�愪ͪ}�JNRqI,�K�$�[C�FC�7ע0!mX��m;�2HB����0��_d�_M#��d�Tܗ<�D��2U���
:�����/EZ"��1��9fU�z�<�61�yMZ����|80�ꦐ���o?1��?dR��9��������kZ�����^X0��틣R��M�5�n��C'���g��0%�	��;�ǒ��I��?�Ͱ��F���1���e|O%�!�b~XO�˓1�&!�1vg�az���<�D}���/�K�1�G�&�K�Y�U�_
͗1?���y1�~�3�aE�RI1�QsY(�/��;]εܳ�Sm��y��]brݠ���?Yw�J
]9�6^vVm�S"��7 烰3r�Qaߨ�\�[;������@�e"I�o�k@�t�oo���I,xe�,�,���7��Euc%��o�\��*�'#xsD�u����ļP"��]�x-Ϸ<q���x�ټ���r��k��'�־G�n}(L�Y8���m?_��qvrt�G�%���$����H����:��>��4k�ݼ�J[���x!���lCK���/�|�t��Z�e�3���f��=4��;\�xy�D�Dd����'6Yd~�,&�X�"c��R��{��Y�y��E	W �����h=b~�HБ���];���r���榞�t�[2R%��ɘ6�&p�
�7*ZAbS�*FWF�|�ߌIN�p�˛��-�j1E��w�T��K�p_�6fl�S�D]���� �q��ػ�-%<�~���=�z��hz;*����q۱���0Cs��czӇ#�����) ��Xσ��р�Li���%5?5�{�Ϋ�ʮ[��]n��] ��~�;_�E�"���,���c�=M�Ϳ ��J��'k���7[��,��$xR��� �P�v��y %%���I/m� <%������MZ$�y�J٠�o����ȽMO
%W��.2̋iR�u���s[��朞�wE�vƗ�ܚ�K�yW/��d�,���cq���v�܏��1dZ�b})���*��=^<�k�r�	){5&_!~u?o�T��0$�4�Ȝ��b�Y>3�F�\X�_�Sw=���!�4�]����9v2���ZrI Cn��<��>�9�=�ߨ�ח-��h��ɝ���{D�|��Ճ����7ש�ώ�D��R�{,��Aێ��8�r���
�� �d!���{�k&�9±5,Z��'3'X�����54ȼl7����z,�<���6�,��_��`-���_�5���t�H�I���\���Bf�UT%�1��hqC��Gk	�E�H�ش���&�{Y��y*oVt�Gr�q��P��X r����öT�Cf�|1BE��?<S�]퇩&�\"V��8{�Y�%�ץ�?�~��p�/%�_��,c����ZK�D��ҏR���c��
���漴N~qio���^�����to��0l�8N�|Ҳ���_##	�/:wd�+\�g�e�Ζ� Ss�uy9}�UKkX�F�3�����v�y�SI�
��6�謣�J�5��Yk��d�=�谣wwOmFq�-��b�w��f6.�nG[�����Ǡ&C,^�k ���7aDj!|2�-(�a��}\���N<����<ߒqޝu�<��R-���]���C1����a?�$E�o��3�ݸ�y��m�q(] ���FFӻ;Lp�n\ƞ��12�#�*jpP��ڢ���N-�4p��ՕsT�|>9ub�����p+���P��D��(֕�@����ʢn]�.?|����1��Q>����f&��k��[ڒ�ߛ�N�<��A7v�n�/FԂ�˺N���_�[��5��D�2$�/�h~\֙u�xTTTP	l~�v����;K�?ٹ�I6���MB��X�_��p�����ǐza�:�\Uh��;�D6!�$�'�H�2ϓ%ϖ��w�DA��*{��j�zbP��>�P�W&�,P$a��w���s ��W� ��z���:Z��!�_�\]�ό�aw�Mr���0oq]4��Àڟͩ����W�ml����ƺ��ٖF�*'�,��)��!�h�뎙��Hu��0&/�z�!S
L�9�T=0]���&=^,ښ� �!pnM�4E������׬�,X�[|��P����.[�.��)h�߸����5�߿�_�����w
ɔH,1���J>^����e{�o�f���̤�Җ�����2V,N6�x�/�ҙ
��Q������~2g�ڷ�Q:)���c\�����.3�����e����)#
����p�����D�xp�����+�_ �����Ŭ"�	 ףܔ�$�
�C�u�B�Y�A��'j�����vBa׎��{�ݻ뵯�g�����1 4�ɟl��+���ۀ�t��Nx���^y����6 c��¥W|A�i�Ic^�G3�ղ׺�(:��0�|�ϴ-&��Ьѥ��qBP�� ��X)�I*5T�9ZO��o���.��]�<!D����E���^��C���i|@�r�F�x��4���s �,~��v[}>n���0�����{Y��L(M7vpS��1	E��m����y_���7nRg��e��x`B~$ЗF��Q��Ĭ��o�k��?olq)�����Vލxk����9}�|��)�ʈ��m/��U1y�}�ݬB��0%%�d�݆���x8� ���Z�hZ\�@H��`ǨC�R�]=�NZ`j�t2�W��}	�������Zg{�H��vs$�Rh���:�9׼�����F��?]Pr��p���N:�����e���S����na�M��KJ����'��'_ߚol�5��:;�*+Q?�ۓ����o��������9�Q����c+�gk����"�*��|$C���O*��ݢm484k_�:$���~e��N�ȮN>�����`����GR��Ϝ	u���{���KM�����5@����\t.l���5Vtܟ=T:<7w��}��Y���� w�)���h��0�Gn�3�"Q���Z��&c�˅H�Ē� �'_M3Js}�3�wy�W�ފ<DxD�r�A�k�UY��H[K�I��f�,�_�@��g0i����k�W�_/�o==#'�]l<�.�fQo�n�
+m�e_��l��[cm RD���|q�n�Qz�@ưּ�пL"]��'�8^R��H"�������6逈�ݫ�Z���d�5Y���d�]���k�W�q�|@��=+$"�^���װ�r�'Ӌ� B����نR�;��4Ĭ��,^(����:��LE$�p�/�M�D\��*�\� %�/"�U)����[ҏx�����,���O� �tz��@��zmg�ux�7^Y��k��Z��1C�2��������ӫ�T	%f��"�J�IpR��;.�k?��, i�4@��d3c���UDeW���g�y[�6H�7����`�M��I�ڝ��̻�ݗ��w�I��8&�C
���������n/Y�І���)����6�'��%?�WU�yV�Ǵ���s���7.�e�L��2��m�L���<Q.>�����k���&�X�L~)��nE��������'%���_���<�}qÂUwg�����t����}.���0U��(�p �_Yt� �@c҂',�7�&��E`��w�p�y�pL�\�f���'Z�m���+-v%S���js���ܭ�揘�!y6j��q���<x��.`�+_���[�U}A�Tb�6�o����J	$���	��B��h���/O���7��Vީ��/�,?<��y��TVg���Y�K4Kp��͐RY�
�C�p'��'�����1>2��E'�?f�p���5��+�	26۹���t�Z�v�ٶk�������>�Q�V^�nooOb;n��G����Y�d 䗻��e�ԗߪP3�3�ps3U��rbi��i�1���௜��}�w���UP렾q��m���`��|{0k ���a��̧�� �{t6[Qݥߵ )�-�˨���F����UPhH��ay'��(���g#��Jo���(d�|��:[5��>��;,Dz��4����1���\XSZ�n*˭
re_���Z�ۛ.��30q�CGT0G�r�l��\;������ǐ�$E����ϗ�/����8���$��>:���6
 ���$�̎�%I��.͠v���,`gge鷧�"������C�H�B� ���;�A���O��7�SSS�;ΫB{��u��-X�r�2���zk���nk���ё�(9a�A ���\>NJ�rS�2)��c�N���=��h�h�4c���ڀ�Y�n=��j ��mˮ�c��ߗ\앜���I#�ԧ�a���Q<�]�K����R�6�]���f�OL��c/N7���R�d��15����/h�T�ä�f!��JL�k�fL����dgE/�!�+�Z�b�����}n�\W�$!�Xg�������mF3��s����n_BlȈlw��hq&���3Q��(klI�2;��G��oF�6�Y�y˃c�L�)`�p��|�ޏ"%�?/��_��}��������]�t�_��iE�l.�<��Br&A�X-%�_pa�ur�J	��w/M-97�	�:c��_���E>o1���!�s���D��c\�j�Ƀ��vS��[���4�u�X����~T$���Hg{u0��0����q�)2;�B���^�$�}��Taq����I	7Z�Q��o�5ߠ7��uQ~%"V�W3�$�=J��+fS��)�~A��1�;_����4 �m��`�G����}�����{ޗEub�'���`ڎ�U.*�En�h���ºo�l��~��wI��Q�)�� 9&"�����d����Ɣ�v���L	�;cz�Zv��f��]`V�1�}�4<�8ȏv��P���c������j~_6�s�BQdpq�A�1��}R��ʜ�ϠD��Y<�~�;�C��FG�g�*2��m,�����W����^�ø���Q� �#���d^�ߨ~��^��h�������D��g�k�:��G(��Bt{r����t�=IH�9���F~VĮ-QY����ܵG!a���?�+aY�EW���-9CJn�:+Eu��K�p��O�ge�������ع�;��y��w���/��BD�߃����p_��%�mᄙ-�K����%�	:`�YS@s��.�%q"@0{�ٯ�j��q)���ۜ_���da::>��b_O	kz��,քRJ�J�3�L�d��L&?o&��^�Ln��|�2ϴB��V���F꘰ۺU4-u�����R��T��_�3��!�0�~��u S�%�����bP�Uv�	Z$2�$����}��i�c ��J�̓�=X�5���6�B�V^B||��Wnf�($��Λ��c�m�~0��nB���g[���� ���o±�Q��E�7���{�X�`fM����ꋡp��.�u�ِYˍ�W�!?9��y }::ƪA�C�U��Fx�O��ܠr\���d���l_17���G|��}iM!�=�CX�����\�q���+Q�؜�uR,$��SD+͊�R17p��<�:n̎���`��@W�VF�/ޞr��|���',O9/���V������< ٮ��	�������`���}oj={���%��}sƯI��[��|.�[y����Q DTk�T�輚�k����9�I���JJM3���/��׎#""���M�d X�sDȀU���
�����BZ��2��T�V��#8�c'iؐy�w��x�.%�Ѓ�v�Ӓ�E!��/���8��/ #(ጩ���'��hy���ޞ�x�`�a��:zQ�b8��#ߏ��B�:r��|��,d���dG�k :(���W'��l'��s+,4��������}���8��5�ߎD����o�����*��O�摞9�mH}�hl:��2����t&��}�òV�wO�K�b��B�n$]p��\=`��g�HdܞP��5u'h�@n���Rx�73�������xE�p�$-������ܼ��  ��U���m��?��F����xq�k������v0�69�8y�۪� ��9D���W�'Yk5����AUPfq �,��a[1:�Z:N�$=��K8{�I�=��X���A�� �kP��vb�:8&�R�j����b��y�wYH[d���~���� �J�]�L���G��v�
c��]c�"'�9�)���9�ٷ�9�H!
����f�*�=\�����%�����?#\�9�6�f˧ ")�тy;��N˪��Ez�����.��E���K��U����]VEU��6;��(G��� �<�(���3��0���q����J�W����Z�N��ښ�YB�Y�4Cv��Ύ�^1�l99=&�N3���0yc����,�!�H���B	��;�Huu���mJ}B�Z�qi�d�/��5�H�39E�G�|���}`~~���Q�
O!J��@����<�^���O�Ԛ�Wk�)b��	���}����o^�>����w�R������q�ZT� �>!ح%�E�,�����B�CyX`�Y{�R)'�V`A RȘ:��iI�[E1�˹���!b�7}�ky�Dk����[���M|U����k��8��t��I���o��b~�_G��V8֫��J�,9j@����~�,L�u3�ns¿�e�8��s�ܽ�K�͏@�7F���C�����������f;�I.���S]���hC?�7�f���m��Ǥ��K�����KR���ۼ[e��@�*�"Qh�� E�K����R}d��u����b`�v/R��?���r�(N��\�p*N?s�g[_e{W%���!�sJ%{�vZ��-�^�lW��l�X�㗮��g��텅}�= }�}����B���m�4R�O>s�p���\�=����\R�R�c�H�R� �9M��բ�^�Eg�FgI!L>WszhF�bGX����"Q�◂�b��iC�����,�C�����k���N-�g�Uwە�٢���X8̵x���K�z"��4]��p�--��H� ��¼s���nܬ�~ş}Y��Ħͤ�&��=���n��V�	U��k+�����C�K�@g���Y�Ɠ@=�4'A�+OW��[�22�J�7�o���Dy�w��ٝ�����>;�Rҿ�`X�tf�_���8��;�ظ��w��s��|��o�{Yk����Ylx��{^���׼o=8��Zsi�%��~w}7[SRa��f�EV4��m��PbN�e�kT�/��&=r��M5�G�C�K9����O��G�K��������k5�{�](�C}'�m��W� ����ǅ_��X����*�?~�R;5�-���]
�-?�Zݣ�:$/�f��/�i%���ܶ�J�(&f�$��̣�G02 �^4L��$T	u��C�r7- ��Y$�� ���z��������P�#�	���Y�ҟCg�`��H�� ���ǡd�@;��c�
�N>�D�פ0�j˒�����,;f�X�EN�譶���é�c2������K���<9�9xvv��`\���k�2�(���������>�6�g��D���&�?h��_*l�TZ�B������Z�y��V�V�c�����O���l6uc�
�?�,�4��I�3�ȭ�?��M�j�lm�{�!�w��� ��<�˕Z|�Tſ{z�ӰF�֋i��܃=���p۽�x6/.5�WL���"����n���ʄ���4rN4�� 	��q���&��ԝ:��p/Nƒf��`1U:�ه�RA�)�?����=�[��X�bx�)ik}���h�s
���T�ࣿ�^�Ro�
��2�w�B�0�<%9>�n)�ua}l%�e��d���!�f��Rq�r/�V�|��8R��$G\_���5���o���p��]�W4�Dڀ}���B^���j}
P�� ,ǋ�?_2�*�)R`����a�~R�&q�	�~t�&{X<h��1�Y����i`t��kR�����!1���{E��l�e���y�f\���ޣ����'�L/沚4v�OÜz#uvl�E�K��jP���M��e�i�	a�Z�P}/+�!N0���4�D<��lO�5Tʠ�؆�h��K��#%��*��y,c�A2��_K�gPT�+6p��K�}M"6��G.��		3#��ԟ�WA?��X�q���X��9���
t�tXqr��~���`+enk�J�0�xo�����{�Ӄ�L�f�2h��$�� ,at��7~A��p��22��ݓۺ�^���7B�ޔ�U�X{�<��G�e.�F��R��D��P���ru�� �@)���\���=�O�I�������a�<mg3��m<�^i������p�SV�Ӝ����㷘�FCc�f�@t���W�����2��5�����pS�h���a��ą[���΄2�ާH���n�q��`#��
~s<����/�dU|94�~�.&��.�!=x�t��I�(��G��g=�:	h���r|�w��d��7+�z�x� K�Ls���T�z)-VH�d���W(���3e�X��d�>M�$��I����3�MCE��|@d-�k&�)�G��z��Pl�04�{�y(O���-�1���>���Ӱz!W�� ����0�@�~�폕Fm�����p���:�o�qCb��?$>\8wx���!��}x$��tLe;Ur$���%�=���Ȏ|ﲻ��V�	���Br�����u~=ض���Ԓh�[f:���FG�άŲ˒\֥TC=�eƜ�������o��+�m�6�������3�e�EV�n��^DhRʎ>�u�ouq��o��y"I�<��t�c+^�;-��Ny��JR���'ˡJ��z×J�3��#��װ���ܠ6�XS�����K�s�A�#�� �����;^T�T`Q����\�-Լ&CC֬��j��,W�Һ6�W�˪�"&�"	�׀��P\ -���Thmf�sz��^�qԗ�A��8���D��]Z���b.��W�&��<�d
n�Nd�� \�@��w�@u��Y#zG��V[}uZ���*_:@���7��yc��Rl����v��V;c9V���Ҁ����d�2�2��{�g/�c"_N�J�P 4oRC��1�	�i�����6�l�չ�<��z�
Q�-X���4�N�5��u4��!�q3]5O������x�oe�6)�e��xދ؝�?�H@�IL��jP���aM� �%Y���aK�clxKE�`���'@��j /_4�����4v_*}�"x����Y�N���4Ie���3������ ��ϭ_[��7�������,��"�a<��D=��|�}|Qj�`~����k�9LӴ*��0kIQ��B�a&�{�r��'+]Hʅ���͒� ��ZQ���Y��sY� .tp�y�i"g{�H��x�|�)f%�	��}�H.�񬄇lݨ��>v)|ĹQ^>���]�OW�*F�s�F��`���E����<~G�
n��m�UZF`F	5�%ǌ�Trߏy��w��f���fc�d���]Diz�Gv����'%xgx�"����g֞��mR|�	6�`�Ok]��XS$@��Λ?���*��9���1�\�y|�Oh2����k�@��>q��c�P�54}Ԙ�TQV�WF�H���Q'M��W��(>Z�gM��"m�:	����X���d���Em��0�(@���yޫ�Z#}v�l�wal���e�ch�Դ.B~i�<�p����bdYP���w��x�D2Fo����!{>sR�1W�gl��>�7���>�v�QH��KR�sI�7���X%��0���|w�EfQ\�(�`I����IF92�%`�ۈw�%z�ǲZ�<���q��*gy5B&K<#%���J��p��Hڊ�rK\�ڄ�tG�]�O��'��H�6��!�-��і<��%��㑰E�-}��#�<������t�\ӫ�S	,q�=ݫL�w��iLva��w�<y)s%�	)ׄh�Á޲o���+}jb]�.��%P��*�#����X� ���N~T=J�a��8n1���	�/���u�LZ`���7����'J%WW��n�[D�ͦ�vG�����+�%F<�MuqsE�v�]�TT���QY�(\l_�b1�BF����(!q��=����ss�8!͔�i:��*��v�#�}����T���&��À9x�i�%�G֛����3�4(�<(ax�^�;�G�d���q`���ک�.y�HBZ;r^�O�����}$�b[��~:�C2޻��-�}�Q��O��y�����z����nq2�>{�9��B�ZuBxF<Kb��A�O���sTb3U�($)�� s��1͝��9j��G_[wz�p1����7]�ͤ[_����t�9�^N<�6~����)T'�K�-=�_�=�>k�Xlr��������ȞTc���^�:�=fB$� �H��M�(����Js���će_�O�#���3h�q�CFbou�-5��� ���Z�wo�o�&:Ƒ�jh=#��#�^I��ŷ���ݣX��|
��`_ʌ��`'�1�1�1K� ��*� �Z�Z������l�c|b���`b���$��1N_2f' �n�����%b���N����kT���!��9��Ak�� !k	���~��"h�ۇx@_͐k|c.���(�Y�=���-n,�f��;pB�Ƀ���S`N޳�#�5����J፾8A����w��; �[GW@~�H�;�'��W`,e,��M�>��6����}%`������V��{�!4�3&�h&�^�;,�/(�Ԝ�^�C�\��u�Ȋ�yV���<� 0w�:��ϡ��6�Xn��t�藅����_�V�6#\I�Z�U3S	6|le�#Ϊ$�,�KY��J�!��%���k��cf�mW%Pz�����Kve����Px����M)&�Q���'cɧ�kj0`:�r��8�;�=�'�.u&��
W��+��5�6��[�/��=s����2�!������3�{�+��O>�nO���߂�f����ʃ��4�d׏0�z�E����M��n+G�y���s�=3��r%)��a�w�񁱮>�;��ſ�t��[�`I� ������\��m�o<����>TIz����W4����R�z�?�笄��DKA������۪ԕ{{{�I����";�~��U�f�����LV�4�5d#� �u�p㚒X�ޢ��)C���u��p|�`P�
pFV6��흛�3G��: �Ԃ�Y*��� ��wSG�'o�C��+%�$����P��E6o�5��3��}xi�;�X�[8Ŷ�Ǝg6�7��L�3RǿI�s�3�Oܞ�}Q�(`b>�5<	K3}�7��;���ܗ�����;s ���?C�eb
��*z�X㽙�K�3�1���k�8o��/����(a~y�Q`��'�SEa�˓�yz�>K]1�Hv8�������ͦ[֟:�(�M aJi�����t�d��Z$���:^�Ð���'7�pì�}1IJ-fHHR���p����ɕUU��U�[�ά���w���@��"B�~�m�w��2~�3�U6��U��ק4�Q!�C�%?ERZ�@T��q�� ���Q@8p����������Vg��O� �	!!���Z��|X��tW7l���p�q���&~�'��Q�s��El o�l;C.�$�����A�cn������9��f$B�*Y�,���MMZT�u.K����z���Z3�5SX�垺?)on���{�2/�P���/cϾC�a��OC۸���l�E��k�����j���8��aS��W5Q)�c�+6��|X8
(��s=DF$��
�$x	��_�\�4ؕ����G9#K�� L��&�?�� '�`����/+z���;����w8�}��9	�#�o�K�Ȝ��ܦ��;�h��H�6�[m��m�Z"����ѹ�.R0@ 1(��2쫼O����k��nK$�`�<���ԓW�(h] ���ɿ�\��_/�x�tgz-�H{�٬�z#����Xto�/d�f3�FzU#Q�o1�(�S��|��0����l���ũ���RT�.�{���w/l�{���
E�����j��	eъ��&b:��6gqL�U��f����C���M+��9�������>G�A?���g?N@�VYN�g���ǁ��k�8�����7�*�4	��<��s{ ��h �s�{/�ng�z��V���02��&���et��.�2��o�(ēVeҌ��ihhh���v0�qӡ�+�;nq���w4K1Z��/���6�LWZ�g㕵~|xC����K�j���K�ʲK���E��E�W�V\l�@ֿ]g�5���8�+�ee?$���u�!89�l��4P�� ���dd}��D��@�_��4MC� ��_�1?�U��r��פ���/��o��h�������k5Y��y���"�UK�n��ç�6nGN��2Up�d��fH����ZUw�V�� dV>�=#ǡ���;%���ϝ����Q�y��"(�,)V���o p���	�P�op�_��}dL��2�M�Y�λ���w�M�w�me�N�l�xoI���	����9��!��=���,=�.��?\��W^��g��A�����;��k$�����[:fh����k���O�g��9������p�8�3���w;�3c�9���#��>��u���gp`C{q�cS��T�uJ��t�]�7C�|�w��]~i�=��ynC�d4/)�h�. =N
 ���[����<���ޑ̱ ��yZO�Gg�#A,��i�w�a�y���O�����V@��T���f?+���4i1�XI�6��ai}��+�@^=Z�M&H�%�nRZ�-�t���?�fEj�Wd�RO��`�o��eRe"l�P䬕D2�N����O�\��{��F�t(����-��WPw\�����N-�A���Q�H���v_��<�CUB���k��yܛ�xւ�Լ_��-1õ��� 6�@Q��<8q8���� I�6J�Y���B�˗ ����K=E���9(������/�2���ɜ��Y֣)l�͢L.ViӖow�ZtPq��V���Q�rw����85��	�臮�c�[���SV�#=��Xrz�L��K�PG���p�g��P�����̦Q����f�� x�;��R�q�n���(��Z�����{�r�D�b�!�ݗx %�'6�K!���՗ֺ����{h�螺�L�<�!�U�����~�k��{�ذ�ji�R7������eU��7�¦��c�~p!z �_�!����װ������H�֖$n��s��܏��@bسC��������7+���R4Q�W,#b�f���O�	z�	_&,�nI�O9�G6��˵�y���t߈� _�ű#��T�����[.�,Ƣ�d�n�'��K�&���Q�u����2�q�Ûݔ>���6���#��t��+6  ���m���7��0�Ԝ�N�n��`-�&*e�pw�ʥm�'Ga��4û�3n��\qJj�� s��y�a��E�k��0 �P�-O;4�^s�.�ŉ�'���N�d�"̺'��-�|��9����eb���Ny�V<�	O{��#\`s��6
R��b�� �<��V��8^���If����ՌWEB��w��/��3�a��"�ͺ��c>�%D4�]��+��{	��I�1����*~�M��v��'�2!��ȵ�0e�+C"�:�Ei��ې$���l}}0�62�������mU��o'������m����j��3Hl�:�[r�r7p0��LE�m� K�>�%i�wc��V�~r'�89,�IAV���e-%1(_}#���S- ���?G+m����7(ى�#����t�wG����3�P��sa��"1C\�a�?�`����H��Q�ˌ61�j�r�(s7��rĬx8}�}g`����9�E�}ɩi2SC�s��SF��IL�����}��� �o�&:|�Ld�)� X�z���x�ߍ�z��.4
�eR��,��F�+"��
:P��~}��wj	�>�����=�Q��"t%k���fq]%�M���:���PE����ׄh�cj���HХ�i�ʤ+��r7�|k�upVǤ�,���R�>��Sh�RF�^��͚�ͪ�A���+`��&��j��\R2mr�4d=���lA�/���wa9�\{{q����~�>j��@�ite�5ٛ0ܘ�3x3@�^)�����j�2���3�y� �J��;xrѭ�����Z�vn�#n�qS5=S?�Eb2���O�Y�U���P�)��w��?�ͬICP�Cؾ��o�j�+��ƃI߿�Uv��g�C���c1Fu�ͽ��Nww����橚dk~���0��u?�t�!��4��>d��8�VC}w2����QS'G�z�&}Ò*5��'��WӃY��.rӋ�,��)��h@��c�g9̆��䈲��\�_��b��]�A_&	u��~9A�`�#0���L��*t]|�ٶN-(`0(6��1�/�K-_FU����8�4����r,6��sf�� ��3��4[��+*�}�٦q��_m�T�=�Sye(x��ͱ��I)x�E����Lj:;nJ���'�(İO4a��0w/�و�KٸR�>s���E���k]�?�z�й	�ډ�m����؋0��W���:BL?�[���=@�l�\v bk6�,HsIK��o�W��cp�?0��tT!~!�V����
��=@����P�}��E���c0�\�u�/_'�)vޛ�V���S?���&�֜
������h�[-`� �����W~��Sx+�îbA�3���z_"�R�^^4�ߥ�\<��QOjx\�f�:�g�t�$�G�f�Yʢ���p�Eư�Ef�k�4��͙G��"�$��b*@�S-��_�q8�\�ݿ�F�8�gh��<@�]�DDǘgT
�gWN������Z���i#8�I^̑T ����7�m{�%�@��Y :3�(61�l2���*����~�J1�.9�v�� �,Ci]I[�!{\Ć��/"ܠ�@Z��\3���8�x~���v��x�t�n$��������V��C�W�|�
�aj����^�F���eᕽ0A��hG�����ו*x�А����2 ���$���}^7m�Y�>2��k�+�,lM� �r��C����[�Ţ��~�X�0�f����Q����5��K	@�����=^j��ÊP�_�8:@kég��Q���i�9���z�X���5V����E�y<�qN�,^{�����[f%[ ����6���ۊ���߹}�0����F{��#� ����%<mؚ�(�4!����ofN;m��8,���-yÿ�J�1HjmT���� *�bI3䛼>��Ba$�:ݼ��8}3�LKPX��4�eg���ț�l�@�Gb| ����`��HI��o@yyꡝ�^�9I���.�琇�M�*��}�m�>HxԸ�\&�Y���]�Y�Q�c����R��J �>�.b+n�I�):��0N$^��_M��b�
K W�1.�#�,�>уx�Ct��r�ˡ-C*>��U�>�"�!N\X/���H�]��ΦK�$����w���G�a�r��X��_�r�-#�2	��Brz��ۮq�8�Zl���ʍ.���Q�,DL�tW���)��o�C����W�2�e��{I�����p�_�W;�ʐ"v��w�=fک�] W���.4,,��� �F2~�Ҧ.K�o�O=��w��U�9ޓm��p�䩣����O�͓-g5�u34Q�*4�U{Ҡ%��ҷ(�#�9�z��x@��͔���R��>�?����q�>�ho�O����6D!vr�k0Vo7=V�W�r�i���t-�Z8�D�:�4괶
2%S[�|��/,�$�9�u�i�T�?��dY�:a�"W����oT��(н�>�s�v�u��w�Nx�[Js�μ���wCP�AZ�4vC�G�e�ٓL�t�t�`y���2A�K�yd���r�x�,^d�@l���pP�����j�ݵf��ftG��]� qv(pdH(�+KL���+n��؍!U������Ndx��)���3��y��D�f��t�h*�w���ᵹ�,�(����i��J\[]�>M��2:���~m�5�ᆴ��y|��N�#�d�@{L�b���j�������?%n�pL�b}�c�wp�R��P��&WŚ5�[$��&2��g�ώ�%]|	0�N# ���{���$��'���K��V�F/R5�4�P@!u��¡!>���dC ���̙����:��C��K3�c��m�S��]@�1��-v&��[ě�
w�3=�fT�7u]�d֣[f�Z������7�kCVn�_���¾c�W;"�Z �随�f�lĵ(����4������YS��T���h�,��M�+[�5��q�+s-@4��\V�za�o@����G��`����݌��o!e*�N�*ʢ�W&�����	���8|+�|�Z�J5���&�5������5�wX�V��I���S&�z'�;N=n�0z�\g?�\�Ddx�Q��W#US�m[���:���H� ��l����!:��@?xZ^�9�q{��.J`���G�7q�?��� ���
&=N��v���P5��k���)bk�Q��ʟ��?VB�����#-j�B�Ō� w$�~�� 2��!����D�[���]��m�� ]�DZN#�����-P�)���C<s��|��
�DPo���خ��8�؛׸����T��}.�/�
>�W�jr��ל�&2��98��a(� ��V�mR(F��#^��t�k�[+�Tv�ݲ�G�?:d�����L=>�
n��9^�.��K)���t�V|�MK�!$���Z�G��(#7&	ţAB�#4ӭ�!���{d_���8`��1���Z[��=44v{�v��]t�_��\�٭ߙ6lb*�xf�e��	�����m�)��+����a���s�C�m0�� .�.5AW�.+������"^�6�~+����AU�Q��A�*K������&^�J9~7-6Ae�ε�`,���2�*����q������~b�����f3mH��>�ǫ�i� xuF�ke~���&�������O�R k�{@ع��	qO�B
��l\�.����ۋ��?�(
=��G�z����h�?c���v%� )��LTX+����i���b���(@�*�݊�~橷��O��#����'�Q����\]����o	m��W<Dք��X��� E>/�L�E�����6�E�l�T.	�r���؍�l������c0�<������g-�s�E1u3t�>�,� S&�c���ؕ�"�ɤ�0�� ɨ�1?8w���k��G����Md�Un�֥�o�0�?3���Z��vY���S-M�+{F<��D�4�?���-&��z����O��l\�����'����W>��R	���ڦqz���å�3���l�!�Z3�U�^I&��a��q�Y|�t�$姪qc�������� ��9<X������iPo)������ۺE�o�5�5�!b㔞G������ |ҺR`y�t3�7���K�߻�Q)��0{=��y�=;��5+m8�F�H��K�jŋhg\#@���?�I")����T�}Lb�I$\|�&�S�%���
�/v������2=���,�D���[�4�M15�CU��
��A~/(� .����x�8a
Fl\�E�u��}�8�:�K���c^p�;ox���B9n �O�]�		��'���4bϙ���lwn����W3]�h�V��P�D/��N*��<����+��?7���;Oҿ�ԏ���^��9�ޮ6��tI��d���&4�#E�h�j�-  �4�	�D�m�����;�Q��wJIDJ X�,I����|�0�9
�HE��y�!:[:J \��z`�E�W�"�ip�+��4s7��z��y��� �����7��C��oa�Ih�P>6����~�7���e���zS��f��0;�}{o������'B��C�a$���\z�"�?�l]��g��KR�
�̣B"hr2K���賻`�tE�Z�����y��1�(�� atSnD���}`�*HDb�=Y^P�)P��B��M���0��akdGz���`��hWt�����$M�hD��k3���L�Ӭ�B��Hd(��� Y�m�Ҭ�$bcc�b���ni�o��8�sA]N����1^���?:?mbr�WS�� 4�,��?����B8�۲��J�Mc�� .�f�tN��b�Ǉ�?�X]-�Gnz �� C������K�l��.��)�΋��'aĸr>S���*�+���ށ����Hv�����������3���U�1�K�#�Eٍ1h��8p<cx:��<:C?�� ��`Г���x�̷h�\3�9����i�Q-B�i��zY����O4�*
u�W�f�yF*	X���M���r��%�
��)$N4�{��S	"���5U������[��2�i������W�*���r������'W��	?{��).й�ތD��DbZ�=r `�~ۓn�~�/O�9�NN����i��PsV�c:������E���'L�tJ��n�"d�))U�V^n�;T���x5���Y�~;�d����������j͔�o�GV��� ��ȴI�w�r.q/T��䩾�y�R�E�aa���U1�� �g=J��b (0f\��3�D��:����W����@�ܮ��TAC�2�J�T�e�L֕k���?H�۴}�kz�\Q{BL�8oJ�v��̓�Q�rݛ��F�f7|��Q��~|��BC�!�� �o�?vv0�>%��̀	o� =T��v/�2w��I?��p�,9�'�a����|Ҿ/� ��4dkI�D���8�X�SD�#qH`(�8*�2G)����a�h�JǤ*���� �K-GC0o�憱��au�od���۷o*<�>�p�ֈ~�l��^���T4�mFF���$pY���i�=�����d�"(N����X3��ɷdDX�S�8�B�\W����=�P�t�Gj�V��Hۘ��+oHXN�N߽�5���(5i�;�XKf8����VU�-�x�/�p��ڇa�z~�V��A��ND��E�n�o�*�R�;����'�=KǕ7m�T�I�����Q��K�����&�$�_�v�\�
��Jwo륤�{e
�:����L�~*a�i����}�.f�'�9|㋗[㶀����8'�gV�Zf��T���ۻ�����Ilp��#
��y������Ì��_�O�E�˓��\�3#�LXt5���{���m�M�;��+'�Uz�F7+�y�("_p��#k���9"t�R����V�-ש�j�7���SRR6�.�X8z�����ٸ�,
u��*)+Ͻ�S�n�>�������i0+�����}�ܟ2c;�lЗR���@\�O:���u?��+����j�P�ɤ�
j��������VO~ꗷP/��mT����X�nX��f)1�aIcA�(�z�'vX�GlF�������#�iW��{>=�PN � _S�[,���ۈu�p`���Q��jx�E
 ��2�WȾ�-k��/̉X*j�h�=�K���1��8���rȽ�h�g��v��ǂ��v�G��ak���89l�G�al?��}ă��K�wo�#�3�n6��4�H�x�6&�H��ؐ�R\��/���~�[s<����c��¼5S�Iv�6�s���If��j�QIGun�W	��=k�+D�����Ak[G�s���������q$��P�8��T]e����o�����6�ӗQ��8��9_���F `{� ���NV�MD��L$ru~>�݉�����m���yU|<�P��qΠ�^F�l=��O�r{d��9�nK
�;�%^j��V$q����*��.y��f*��B摤�2�@�g-��E��=�np9OY��.؋�q7K��������]T˄�m�G`��vb�:��r��\eX�ni���S�b�z�t��4���w#�Oi|q�*�
vFnx1zCd�S"S�Vn��,�������XK�"���8��������^��<�>l�%H���D����T�R<��4$���� ��
���O�� ��ggL�b��Cx|>h��뀀��9ަ�GO�]=������B�{���M(	���Ș��q��Ìlkm=988xh{yy1q\���q9���@�P���yM��	�m�٢��d�(�����-M$��P<�n=��"�����C7_���du�����UJ���[�F�u�F����7�����렳Tҝ.p����q�tۂJ� |g�S��G��E��6T'������.��(K����2�]�<�4�ظ�����(0�����&D��}��ٚ�B���:l�9�hI��dD(�Wѧ�B
V�E�b�N'U$'u�S;����O\<�+��w���w$���&m�X�@aB[{��S�~�Ke!��Ef�v� »����/�bU»����l��o��Q�8n��V"�Y(�@�z��UmJ
��pW���w�<��m��d3cӣ�Ν��#��S���KD�B��k������S�$����xo/++�:�a����q피�.��Q�ǿ����~�����Y��{Х���E�����909?�:(��ܖ��Y!"Ƃ���iw?����t���$��~��GzJ!w:�F8��y$����ys��!�����7L�J�me�+P��U���s	i��f�R���2��G��u���D�$N�P�=�ƽ���4a.3b��@pWMp�Ӑ�-�ѲW���0������t:�_��-�-�o��a�^b�u;Aa٩i�V&Fx���[v�s�g�Ń�s�'�ni4���S�zd���Cd
k��J�l���j��ed>����n��
G�� 
�x���&<���K;tG��,UVTQ�	����N w`S����2 ���2������n�oi��\mo�|�jm8�m>Y�*uPKfn������X@�G�-��o�b�����BY���ħ|||���;]�̾���]�#GP��u�O���.�<��a��y
,�<�Hn�g��G
40(����h�PJtj2��@E_ۑ*�����vΩ�D��2Ł�E���d�4��4��{�K�
(���4	��O�T�[T Yɛ�F�$�p�+U��[�����kׅ2��Ð� ��ӯ�
��h�C�'����B[o{':8cIf��2.I�o�����b��d��aH��Ǹ"wm�%aĿ�,n9��;,��a��$+�?h8�m��I�~*���;l۹��Sf���"��SY';o�>^L�����J���G�TU��e%�K<�W��l�u��#R�����d}?��ٹ���[�Ղ�����@1>�3�}B�G�}"6
Ͻ�l��X��P�[��yqI��^��j�w. 8vI�!Zڎ�i5��ݫ��2A����������m�mn�����^
H�������|�jЬ���hu����:���n $���Ǉ.�a�.��Kz�Q�W���l�*���NF+6�;��/�����&Q��A�T+�B�*������VS"��Ѧ���4�u������g�d�q�[q
F>2�?+��+vH�<o�"��Hn@�ga���99]J%�Aq�g_��ij0���X�*��j�ΗmI����M���3v�ݣۋ��ǨҾdd��G̦Z��[����������r�X���	���90!haX`H� 6�cutR���GD�h }�KW��K?�� �v��X��e����H��Ri�\N[����ؿ�+5E�3��?��T����Y>�������Z8���V���l���ȅ{����嵺/�9��ҙ���W��_�Nk~-Ol�����g�U�<�,t��j3�eI� ���Ab�[�LZǮA�}R �P���6�*����*�Y6��4��m��z�����ȧCO���Ϲ�ws��+��mǞ���B�A�����Ȇ�Y��
��������3�i@����	�8Gx0�3/���+6B/J�Ja	���j/fS��|���in�_�f:�I.�@ԁ����0\Pyb�Q���ܳ�U���T �e3Ʊw���:
ֿET���7I�L��y:��CE��ne�������x��^����U D�V�Nؑ��oj�`N?r���9�j�#>�8���1?%l[��a_g�)xyK��ˤ��"��Q���U�֤s�[N^���ߤ�H���YV����#��׉_U3U��Zf[�YtZ+��
���ߑmWr��d���׷�O���)()�["����F^��D��##S����r�\^��㼄���">����\&�E^��9:w�^6`�ī��Ḕ����-�
�7;tU&m��u��2����΋�i�<��~�!�>٣kp��kK����%}�cD{��'��ULO�cƃ@�����ʎٓ���������-+"�QU�R�t@h����[r�O�N�!��E�d��d�/Ӛu�G,���˹�u��n�5%X�Y�v�Y[���Kb��t�T�4 &��)i�O�L��7)���7�
's.׿����2�9��(�_��m
�D�h$�	��X���'����j ���.�?˽!h	�Ӹ�l>�t�> 72�����E�����6*]LE���T����F��T��8\`z�Xey�+s/�}b�t�n���@��K�.A�F�I^U��H[����le��"�Kbv�_�����`�$�Z�Q����E���/ԮQw�A��\��|����;�M^���*��=�*P�����?�Iɍfo�ݿ�7y����8s�3A�U��Ń�V�Ȍ/vp<�v;jF�#�(Z�����.:k�Y�q��zc=����(�=�{e���G���c0W3�i���["w��U\̕�SaE[�B�������AhA��-�2~L��F@�|
�	;�k�t���@.�%�l�-ۉ`���F���r�}Y�*y���x���Q>U'�/�����ZS.�e�;�k�����i3S�*Ǒچ���5����֙-�7_��s[7eX�Яp��%��ʉ��C���%ˑ\��]��4�N��|������h��U�о+u�9�g�9ߟEb0�����wJ�
�l`��˘�S|�l���>�U�=&hŚ�1��IY�Z�j8RX=�x ���i]��lg�o������r^ǧ?�NK83�&.�{�e�������i������a�l̞Z�78�<���r�]aH���IE[���X����3��I����A?��&�4�ip�t8D�ur�n�a�z�GFP2cn�$k`�[����}�e��<a��g�D�~^-	-����9�ߖ&�"�~��L��NWv��"C��$Ś��8Ac�So6D�*[v�nC���Ne�䢆����%��*�����a%S��+���B޵���� +g�pL�<&\-F�F�'�-��ק�.R]�����
�$|��7_[~.��qvQg$cUڎ֑������w۶v��Q_f`ld"���1��-��I��
�v�e'��V�}\�B��VW_��3�O�l������<A_����M�����f�d�_�:��I��������rc���2��H��<�q�IɁ��9sn���4�}J�"v�Gjj����\q�F^�iu�(��:RJ��F�a6W���h��������Ƙ0�P"X>
��'�����J8�*�/EJ=���r��&��F�i�����[���W
q���I-s�c��σ�6>�J1�yy�QcV�&ź�M�ʠ%V_���n�y=���8D�h�wi��i����ѧL����B�M^Yհ\�2��h���Y�ڭ5�.zhb�P�y�[V��YD"[�`���%�Y4f��v�� ^&}�TP�B)H+$�#1��~�=����yΧ�\�|C�£�50X�422Z3j�|�_jt�f�>�@��]��%���>7�^N�WeG���� @8L:5�b���%�����jD"�g��e�����#�Y��N�ӧ�4�fT϶�5�Ë��F���pG|*�6��{��o[Y��}�r^$8!݈!����@�����ɷ�T�k>>z�8�.t��������v������[5
hP��N�����u+]���2�4���/�z1�pKF���a���=f�` c��<���+É�s���O�[�4M��������	U��*�9�C39��BH�m��m7�M�>	�f�n*���J�V�ɦK�׉D�!�hB���r�Rҵ��ȃ�{y?��'	��o����� a��קK#/���?�G�J�cl� G��o���-��pt����� &���,JT_����iҜ�z��_q^��|���y��yR�`b��!m�PD�h
�l7F�`O� 0G+C��7����*����+��+�S�cB=�*��Ȇs�9��0��B��� �M5cn0G�(��f��c��T��̈́G��+ď���
�O���A�F�y{���o���`6��b�h(D	�`�T/d-����$�'z?�R H��&�'Z�an�HDle��/G,��t'	XKVB���A���	,e�M��Br�Ҡ8b�6ݫ&���`c�����Z��	~yW{&��#�$-�����/�MB����E�{.��;���F���V���~��yw��xZn��K-�7W��]� �0A�x����|]@���I���T�r,՚	+�z�\P|4~�{�rrz�}�����g�����������?�V��h�0����٭bz)%ަ7. �6�4�ty��ԣ_�8�t{T$�$8�a;i~��r�����ѵy�"S��$Ƹ{S���gS��t��F��cqA�n��w�W���z���p"��T/Sm�����zk=<��i]#���`�d+~�}8�	ο��E
�KfG�2�0�/}����O��kS?����VMԖ�В��Ә� q[(k��qq�? D�)��ʟ֧��׺�_�2�^3U��J���X��I_�B^�o��c�6��,/c�#;������]�Ku��� ���<WT���l�vZm�����&ׯ����e������L��D��ׅ���\#�mj�ա��L�g9�M�n���680�-���{��{�B���PJ�@P �����N�>8n���>gX	.Z��)���e/�p���E�^����z���-楛�-�6Sh���h���6�=[�Z��}���}1[F���X�8LLy��w�8���\1�d2��P�vo��4ڝ $F�0�h�#SW0�EIZ>�nNݟL)p$�����ܢ�j��y�փ(�|���'Q�u���Z�����nW�ҥ�T��xM�|��U�X�U	4����ua�7�F�8_���!H���P�����8Ҍ�&\_��C�p�|s�o��::�w��A5��0LN���Z�5�?��܊��5;?+��~)��|�@��,�����}.����u����S̆o��~46:z/`c]���m���.�,�$%�o�gF���S�����О���x�.�M7������@R��
����=#/��L�8��uY7�[�U��b�Ə)�u�͘��Bڣ���2?��Y�P$k�� �/�Zo��wU�T^�u[H��@��X��=�qv�z�������DX�����,ǥ	�s޸�0sI�����R���G)�xO!��l����7�{6��a��G;�U~�Sc�������^������Wmn����v$��W�X�`k� �>q���>�x��3��ToT7ݲn?fx��A�?.�l"y�` ��$���ˊ�����E7U����aT|���3E���d�-'��%Q�ܦKs���2ţ���^a_�hg��R���틶��?Qlh�]����m��:@W���S�躷��?���z�Z��]i93�Z�eP�����]դ��f�:1($�il�k��� "R���e�ߩ;Àae��>��}O��_ҳ��k��Qn��ģ�V����TB�L15GØ���5��i�F�&M�|��6�4ˀ�9�x�﹗T�xm��-<����*q��
���&Vl'�>�%{V �;�S���J��� �|F{��<|�­�Va�D[�ף�S���6e�*,_o�6�����@0�u��@��W/٤p'��(+�9:��C�Q<2&Q����P�̬��'lع0&��|CCFF�����aI^]]}lk���.R��A�;��#^���U�_�<�w=̊�>��S3cB��)����%k����]\b�`߷�W�8&��$�T�f��g�����<+��A�D�)r�\�J��{0�[���O�����
l��X��o��0j��	�kI��ƃ?�R�rOFkBH��yp��/uNJ* 0b��Q���@@n��1�mZ�2� ��^�L�
�v��^��0W�̥"|^��w��+xe7#&d?�ݖĢ�į`�t}�]K2����6�Zܶ>�_���³3T��}�P�4���f�p��}���0,���۽d��w%s�)������k�h��%�\���g��H-�������q?�=c ���Z�K(���=�t㐽+F&���Rz���poj�8�ے���ttt�===�mm~�{���s�ni.!����Fx7��Nw��>?]oL��_�pFoY�{�0T�G˟�>I������������2!k4i;�\=Ƙ�1�vrz*ݍv.��Y��zjL�SI��9A��g\!ڜw�������tg,��C���� �H32Eu8� ��Z9��3$Hb���(��E�8z!�W9a��_}�L�Z��\��3�X��(-i��Gb��Q���㕎��� �l���5>�֯�h��hEs@aY*��,��S�[[�`� >Ζb�ͣ�X h��j�%x�j��0*����b��4 �r��	���ӡ[��iG�Ϋ/H`R�ҁ<��@���*hp��Ul1���l �V���N>���������#��|���~j���2/�Ԕ�ebdKpy������Nla��S
��ш�ُ!��X�$̖?��L}����F�"��'���1�NJ��$x�W r�+%hҵT����{3#���H�0�5��5t~֗Q.yE�<C�֊��iBd�e'Y$��B�l�,"�k�V�֜rZ�S�͔ӂe�l�)��" �ީ�����͜��)�ģ�9ؙ�'z���6��vs���2|�[�
��XK��5_��''��c�my���4�bW�ߋ?�Vb�XH3]� ��B�7�L-g����ɍ�Юx-����B�
�)g��;|�����
�I�3t 
XI����Lݲ�
�<���~��<��:�Gh��ȗn��Y����A,�FW��S����oǥ��z7�����X�������yxx���.,.^�/5�rb�[O��A�y�,��b�
"~���"W�;湲����� "6��=\�ܼu,��$�i4/"�{r��ڌ!(��^�:��{c�M@^�d�����O���}j����2"�k�o��B)=���Z�b�����<��;�$�7[c_���
(GC�(��~������rp���ʈ����p�:�HF0:�c0��9#�� ��$��>��5��E;����hk��B`nl��t��E��\8X��Oo�?��8Qm�{:�M��6��|/-=�8hp;[g'k>�Y�Sb�J�F��eh1*�ƺϧ�|Y1��n�����P�Ej��'��ZW�Fo|k��=�%qo����"��O�.'����wik��?���E�GL`w�W�#�!A$xo:����,,�s�p�XN��Av����b��$�rB׽M6�_�Dq�&n�YHO��ui|����� �#)>R_w�D��A��`5���E���]���������qLe�����w��I�-s��(�>��M\~�zA�J8'��-�ڛ��"���_/@�T���11וk�����,����k`�⾨N��	�/�W6#�W�����,lm�N����v�f��1��4ƐD�F�S�w�ܺO�3������iE���lA�bʂ��;���*H+id����h��=�>�S��/�IŢyޠ�-�{%�.��?�}O�K�lO�ƃIb�F`y1��<v"_�������?zz�`�*sJ���m�֝�9�I1ɝ��)k��f�X[Y�� no2*'���h{Y����}�!��ݰ?1���x���"7�[�����
�KKK^����,?�$Pǀ���k/7Mā�AC������ )�����z
��6�1+���]Sk>���P�����4RܗFh�iŇÇ�GjZ�N�2=
6��i׷�/'ܡ��ym��P�Gԫ2?��tf���Y3�:Z�&�=�[v!�F��̫�Nj�ϖ+�cD�2������<��C�R��A"�0���/�T�al�����f\4�l����pDK��.��۱�g��������$��:���a���_&�oL�f�L����Y��F'-�]�b�e��"�:|����Gp݄���!f����XĢ N\=�$Y� B��Ϸ��wYa�YL�og�
�p�H�0���yGȐ [���s{��F��HW����Wö5� �G�?�9�"��-�>�����L2D�^�GS���$��p�p`*>����9�>âF����q�^�SRm�͵E�[Y{
���[��~��I�;���n��]܊��� �Ci�B�ॸ���������7��?s���k��Y3��˘���W�xm�n����$DkQ������5s��	�ǘL��JY�i뽵Ƴ�`����qS~7`N�o,St%i\QO�ދ*��%ZI���m���/P���%�Wf���WT�EF�l��Ryj�M��������[�tQ����2x\��{��n�?$�ӹr�N{���?�e0��v~��P��B#kMf�e�,��s��6b�F�N�]�7/c�+)�䲋 d�A|��F�����ǡ��J�߱ۑ��+�ڇܤQ}a�S�\*<x^�\V �nl��j1���6#���P�>'��/�	�W�)s�ۚ��遄���"/P{�����E��$�t�m?L�3��Pgrq�n��sA�;�?��p~ �|P[�>Ye�16��L}x�4ir�z����]�����G�T��#���Q�������j���:�M�6��O�+�/B@t�20��2�[��� �Uj�)����,0�9�gM3܋6ht�Yjl�?n���!��@ U�K�,E�ß@?Ö��af�%��T?	�,�<����?���i���)p�k`��8a����k.��_���\�ߊ���q���E�K�V��>����$jL��Z4�� S��^��5Tſ���%ƛ�"����׾>�CMX�n���Y��ֱ�������!���0����0��yE����(A`�n7W���D:�FO����2f����.q��e$Ib�Q��hkQ�W��"F%�(�nX~=.��%� �B������I�ax�[^�������Z�;�����jP5��������u�o���8�����։�Y��;;��3�H�=\&��5a �5@��7
/Ν���H�& 1�5<�~�Ֆk���Wo.���+�p�A��B�ԉ�xڃ������Ƅ��	��H�;��������b�gg��3��舻�&(G\�����<��,�}��|��/�9u|�=��@'��a21<N��s�M��=*t����}p��Q
�n�JuΌ�b����cB6�Jl���a�9�Mr��S@�[Cv�O�@J�� ZX�DɟXv���*�Zz�x�v�g�B~_|o9�Wk�o�2���ru0��U�a�)j?�E�� 6P��Z�-�-�aɮ�\�'K�这��F�?7��ƣ��p:��g�����T|��i�����p��^��A,/)�II[�EK�cD{ر��~��������D�D$
S�9���S��#m33R�5�2
yj?-۾�e�X���  �;�B�U�R�K�m�|�+/�Z��c5�P��w��ѐX���)"��TŘ�
���nm���/@%�������"��1�%ą��(�z��}����"��\q��P�7�qO�%��B+����e9�%�Uo�W�jUqr�����D�Hh���EhAɀ�1��BhJ�9�2s�Ɓ�{�$��wkf(�^ph]ٚ��5���쩢#3�/��I����b3��.3�����1B'3T�*�������-��N��QK�N��	T�m����lj2���u�9obv��Gr���G�q�}����Y��=�AE�Ns0%咺�n����j*��WԻygGxl�N^K�Y��������r�O�ƭ�4ʝ֧@����ڼ氢���F<���/�Y=��,��(Ƭ�Be�<�v���o��H�ηdN
t��V���h4+�X_�\�?Id�	�V����|[���	/N�;��7���I���k���%�/�7�O8���ھƵ��t7�B������UC�B�}�,�%nR�q�T��%]��4EO ?4���##���z0"�z�i�X��=�5���'�����q�ąR3|�s��}�a!�ئҼj����MWߎu�y/��P��Y�7�`�����C����(ԺMK��w�Cf�ҵ��ޙ6VT�t��1�l��o�&i�4�o�/bV>_�J�^+K��Q����[�H���:�l�-��;88��3x?���wPQZ�E��.C����@p�/PDX"��4s"h˹ �Χ�et�( O9�ToM*������h� �=;�v�&�_��8H�)U�2z���|��E^�N'��;�}u�r:E�
���v���������klq�>�B��:��`��)�?��v��YƓ���C]ؤ���`�V0<��0�j�4�� �XÍ4��vl����e��9��L_LحKz!������m��\Y��M���E�#��P�3�Vi?*���yY��WCr�g3Nt���Q�C�C�c�D����Z}��՜	�y�kjz�C��������_�\�5m������U���l�ԡ�V�4�H��z��F��דE�C2u]@Ǆn��+�ߗ?BkOl1��_RO;���FF3"IN�z{]��f��8�d���wY����y���p���ẁ��؝�(.&�ȏ��M���V��}��U�7�h��T�w'�h�Q�0�m�'�_Yqf�,��`�X{8��h��G�,�=׷l3
�h:G(w"S�k�٬�:w郳!�[EHe��ה�xeH�D�	��w�I-rB̰�\j�d���~3!�엻��q�k���6/��M`��w�(�#?�(��pI�4m�K��t������>�hk{2�����P�g�A
�M֘k'���J��fD�!���+�d���Q&���}�T�����٘zl[{h�Y	����[�p7>��<v���
��%�	b�r����m� b�dd����6��d�����]S����� ��uR�J�� �'���"x;�LoL�{oX�r1�*�?8a�L�jg��{��4뢘���ִ]O��Ez������׈�ٷ�w���}�o8Y,�	���f���N����ʨy��1SjZ���J�2�)�[E��?�qw*���� ���?�R����:��UK�82��@C9�x�[�,cz?�e��r&���Hc���a@%�H��o�U�aq754x13��v��v�Io�_q�됞+p�-�LS]US����l�ppۇLlȅ��^@���z�]p���t��+"ьb�U��|}����+��E0#VB�TWA)�s}��ڋotg�:.���)�F�l�n�T|��b�=#q��4�1H���	�
�^����zZC�]vnRƝ��z���L-؄쇩��I|@VY�����1ZtM݂�&�oP$�uP�~����D��,����
�!9�8�[�n�����U�n��ta7�[-��Ԙ�1C�O�)A��!����^R9({N��^=����I�C�i}���8���(�TE�=A�n���h�m�.���BM�?w4*D)�rOv<`�/vw�	���J[��l���û�f�	_�B�l�VT�J^ʙ��n���zDA�tGJ,t;�}{"�i���o"䴃/FZ��\�м��6es�%�,:����}��{ͤ�������ˀ���Q�ô�l����}^�#�T�������ㅫԭ��a�$��М;�x�e���D�:��T���1�o�GLc�y��	e��
�HH��j*Vc���Piȭ��QlW�!]kc/�+��Cn'܎v�$I��r3���f�V&�=�"�L(U�'Ϩ�mZ�S����$����[M)/jp�� Ż5B�����/�:"05�.��\.��򰶣��e�<!�j$Ks�.#��̯>*�_D��v'(0�W�7��
qC��=q)�H��= ĕ�Q�.C�'�UA�;�����_J���A���^��8��r��b��l����>��ڴH���Ŕ:M�=�1FN���X)��}�)LL*;4���1g ��	$RsK�Hm��7+r�-����IpsG����j=k��p0����q��h��v�]�8_�f���VqU���~��9-ՋZLY/|,��S�mQ*��N(�R��ڐ��3�	 �&Z�ä�
�t1٥W�a�ᛡ��y(���,�	;9_���'�O����g�׬@B�R
��bΉjh���Hw�FB��k^C����!P��w@����Sw�-iNK�?��"�׿�}�$��;�����"j�f��rAj���u�{�k��?�	ճx�)��j��ٖ�:��k9��f$V	�Ǐ=�	��8������$�}�o�?��V.�
+��6����y:�A���n�M�`�IJ�������^��2��0\ӄ2���6Ӊwf=������7�������3x �f�/
�J��[�`���n���\k������EK/N�Y�<�R0���9�3
��^��]mx9,f̾�2�j4�6|0i`f,՚�Uz�Ip���m��7D2�
 M+[�G ���
9a�po�-�1�D'#�p^�*[���;�J]k�N�s���0h��������v
�n�=+�p�/B��s((�'OO���\����$�~���F_j�4y�s�P��a����ʰ����Tݖ�?�=�5�~����/ߤU���4>�G�<������)&�k4t��rԊ+��ʰ0�ϖ.���:va���hp�0'N	�RcI%���?a4���Ü�r�-���(i�:�yk^�Ӏ����&�O�_GK+�Z
�>�*�OU��J[600`EBBz��~�������}V��ct�a��P����2Z�4|�T�C�`f�fn�!�ũ�[i�q2�#���d�%2�OcQZ���9�y����j���x��9 )������ �2&o%�c�rX�Ɓ<ս��/:k�Zƀ�Sڅ����N;r�x�)�����J�G++!4Z���(96	��²(�.p���!0�k��� ��_��;@zC"�b�9���e�C�����)����V�-n�)�Bx27�5��j��zю�H�၉@��t���\����P�.���n7V^�y6 �����o�~B���}�x_qp�G?��땚S�=$�r�!4
Γ`��ʚ싸X�B�{`m� P�1k�K��x7��W���k״g���<��ِ�"�G�n'簆X����r�����՞�:֤�����Az��˶"G��s�K�u�����7F�� %���^��1J�{O� -��>F9�D �7j�M�S���I&���~��t\�4��#����z ��s����~�ɷrC�0Eڗ���|��_H%���Ŀ��z Z.m�.Y��U4�	}�e�ׂI1����M[�EK���!���� � �삎��wMĘ
�]ڮ��
9i��
hJY�o;��� W�W�O�@"��,�3�8�f/,u�i��m�˷�z���Bl��}�Mvv��d�8�%�/,��MΤ^j�e������4�G�������)�ՠ�<ܠ�,��K��ꜰ�Q{gl�#��(��O�ȇ��t��tV�'9��7�Rkk;�qYޫ��*/W�no����~��;[1����^/S/�,���sƻ)�F��A+���}}���V����2�Ѽ�V���Y���xlZ��������uU��8X�O.���CS���E��8���5[!piRr�^J+�)]�sp2�"/E��*��M�F*J�"�����h���ү~C��s���2��������&����a����Z_��?̐�{x��7�=���lἺ��@O��?��on�"�/��Y༴��|� 6� Yt��,J��Έ�q@��͊�h�ʝ��L)e����ad��RU�_���x���v'�=�hG�q���g���fM�}mM��=ށ�?���<&ev!z������������1�k�:Y�wZ��CV8y@��O.����od/N��v
5���m۽���\Y�w�\~��3$��J�77�C$E�$�J0K�c9 �����F��R?��zO�<�p7���4�T��H� �һ ŭ0u�o�Q�Ā��B�S�r���~t�豇S��݁`[���dO��ݡ/��"d��b��Jh1�G��Bs7�AMr��o������F%�离��tj�c��Nm�J[ͳB���ʳl�{���n���?s��-+c�@ ��q{tZ��Y���Sn�C}��ԝl�ת=����r"ʟ�prY9ᣧ�p�}���a��sC����xެ�7u$h-Bv����.�㍬n ��%��
G*\���`Q�Pφ.z�������4��Bj3��=[m��J�B�(b�'s�@A�����쮲{7X"a�\�~G���+���@H_���R�$��#�;*i�AyK�����m�;�����YV^�_&C��L�I�qλOX��j4p��D�v�A��`Ҹ�QƆ�������FJ�q7V6o||gȿFrJj�^��8�|��dy��m$�� D��^�'&%y����ܕ6��u��u�Cu��b�Ҫ���W�w?S/�)jl�>�Ŕ�m���R��l�@o���pđ1�ɲ%�1��%��M�E��m�$���"l$��WP(������Q�4}cF����Xw�_������&�)Ֆ��}�цƳ$���E�3\�'KW����Ǭ�r��A�r������`F�OQȃ��㉓�k�~���	�y#��<{��=;b"}
��2����Ŵ ��Ga1���*�2���f�1G6�Z���=�oп�I�vO�S�ly����;�t���2�y�c�P7;��i`^J�Q�ŵ��8F~��2�1�Y9��x�!�w���RL�D�\5_�1r9,i+��}�E�	����u-�!��4)��&�Dʾ�Ư	Q/'{/�E���o�[}/�V'&<7���-���x�|�z~"]���A&��*�P��<�7-�EIX ����W�ι\�r���gx:�s1M�ۀˢ�dY�`<���7u���x{?�
�d��r~c�0\��,��RYe<&�p�

��rzl��n����en�p�A-ki ��2�b{�)�R2�K  s؇Zim9�,CP@����@�]���V�۠p��|�cU���yS�	ϔ�`�Ұz�{v�JL+�͑O�Q�+� �3�Ŧ�`{�d�k���.&��g��` 6.�5a�M&���XLk!iDF ÷l`s%@�孵���4�^�U���L��Y�a�\7�!Q5[��(�������@��B9�QN���[�5��{KU������y+[�˟U����� <�*�a>�|���`�S�D��I���OmșqǇ�� A%�\B��� �[(�=h��<I/���� w9޷8��=��I���)�a��*1�5'K�t�sP�2X����*h�Fڍ��np�Ǩ�*�mLTo��=�h���7 ����t��Qf��q�����H5`e�f� ~՗�S1?DH\MkVGU��u q��b � l�Ab�aԹ8����7Da��4:?�vm"%�W�rs\hP`ƴԮ/ߘ�j��MllZ6�+Z� a����sntώ8�'6��4�WS��KY�O�X��f&�XPO%׫�M�1-k����}�Q��X���Y���7O3��"��_��j�*>��d��੡<���'��l�M����"Y��T���r`T��k��
�(�j"}�J���c�C�K޾�8$��@���'��C\L��C_9M������Ȥctc���D �� b�⬪:���l%on���F�o��6x��4(^t&6��X\�*��i��O�d�e{��9��N�aH0���FΎ�l���v+�O�!*��
�������uB���pKSr���b9*"A0B�ہ{T^����i�i�6И4~��ۍ��Y-�ڨ��J Gs�{��q3��FF���"�j�S��.��}*^Ə(>��>%)Z���2�ͯ�x
_e�������K)�ҡ@�ʿNLv�@k��mp�����s	��GH��k�n
ҷ�=viAUhz+�=p�e\ї����?)�`d��z /�����(����M���E!�!Ir�����,�~++��
�";�ޥ��	2D����a+t+���݃g�e껬��2��g;������:�ތZ��nt�}*E���۸j��R�I LH��)2�/��l��!/Ic1Uޞ�q�78�s++===�6�*�PG��l��/GO����w�� x�T��'6:���q�)v�C��xt�O�x�Z�w+U�-���Aە����GA�n�/=r�_�r��c�6?DP�D�"f)ąj�ҙ #Ꜥ�u��
�]�IȜV�d0Z�0jGd���#s2�9��Q	!\v#��w�(�����h<8�y��r��������ﮄ]�	����%�N�#��f�{�,�/��J�(Q�/vҙs�cj��q.�OЄf�?@I�_��b����c��ۉd���VX�|D�W�u�~����Q�)��k�b�9�A�E��cW�4;[X�T]�Ѯź^M���ÍJ��A�/��x��_�Ƭ�2�k�~��VS���AJއ�i��%��߽���LGpM�x>X7��UP<`J\��O6C!� K<���@�����Ւ�����m�Q����H^TD�?��	������n��˥b�����
�}
�McAQK������o�_�p����V���ؿ� ��,�w�m��76��-�s�r��+ū C�z��/4�s)ʿf�͒hx���5�����6�֤z�e�\�e� 8� 	@^��ʜ}��{a����0\�/�T7�6��ec����6�ڈsϾ��O�F�b�[%ź��&� J���S�F���k-�8Q�&�H���	`��0H�B��
�f
�L�ߞ�U����݁P���]S��]���=�	����Z�gT/;���ȭ��f�:4��_��X���!N��c����g�����ô���y��J]��o�h��-R�b$8��@��_��>/�+��z�"�,}���nǠ�,
ޑJ P�������2��;:j�.)y�|��j���Ӂ���>[�L}ۉ���v�zQ�'o��5N]P/)%"hV/c�[���:��;�\8G֊AA��i4����T(=3j�U�j�H�T�+2"��:�=�Ã]�Q@�;� �d,%j�����/y$���U1�D��h�+�T��M�����%���D�r�0�6"����ԺE�|�^:u������})1yJo�Iw���Mp	��g�� ����t��D�MB�8��.�����10�{�%��b��(���W%��N��Pv��X�����J>Q�EYϕex�	��x(N�;��BRi���e�8$@�w>��b�l�4.�,�|�v����%���w�v�Sg�R%�n$0����M�x,�W������wӐ1�?����o��Θl���[8r/^YU�>�"k����kne�J�_��
 ��2����R>p|����d��@�ww�c�ig�Z���=�Q��5���mF�\��v��l�;��FK~�]'����2A�$�(����G�n�ݿ�G��B(�w�u�}[M7}��9�޾���+��me�9�=($�5�FD�-�'�|OlIu��wKa��K{����E4U�cR\@.v��%�<�VCs�lMj�tzd��y�륙�S-�'����l�t<���էn��O�fI}n��
�ڽ�}�i�h�;T��n�Qz}����eR��V�z6w��T�9�7�P*n糽>(И�[��R�)�WzС�RC��cIz��jj�J<o5�;KtN��� <`�0K�������ij$�P��y�L�UxE�7���ۥ�\�"S��3{=]{��-�ny�Av���ˢ�y�x�1	�a�dOr7�b�N�|�N2D��[�a�q�I�g���HTE�L��VVT�Ĵ�=������[�2�^��a�����N�sv���I���b	n:� ������0�;��\���r����7R����΄���%�ˬx}�!��H���.�f�4u�f*���pn���BM߃&�X���f���x���^y�P�5���Z	�t�J���.a���9�ҏ�tV�L�ܐ솱��sm��$z���h"����a�j��hDT�FY��&ϲT���¶놽��}uXuxh���G��#��9��c>ng:���5���F��rh�d��i�nm1��;��
�����ͅzu�/+W�`	[Np�C,,107�H²g\[#�f�����O�����O6G��7�$��t&	 ����6{�q�*���'�{�a�Й��!��$վ��4}����>���y�7M�y�~���~�B{r��=�I|~�¿l	]MLy�䑬%����� �N�����7�d'f����&&&�EM}'����N����mHa&�Gu��W�5U����Ƣ��<f����Ke�9L؍��<4^�I[�џ$�v��4K��(p[�/>�̌PQT�c��?㚱#��� b�9SD���o~��c]g����0��RX��nHj����J[���nQ3�m�3����f�Ai�C��?�Y�0ˡRw{�,5�|\��q9�/���ߔm/��w$C
���2r*�͞����ǜإ���i�ht\B�Y��'siؒ|Y ��R�&ɐ�_f�o�Prj�)Z,Tj�U�W.��:�t�g�����P���8�녳�&tfcҘ�I
Qg�fUԣk��u y��v��M��@��F\���p�L5���Yh�iI�}�d�@����T�dZX�E��JE�(�������G�.��r��|�;mZ"�@r�d}o�#ب"Y�p�c��_�s{K������ܟ���L��6� ��}ъ����F��v�L��ŷ�`�4W�@���ҘW[���&C�7澻��#+�V���e��Br���pgA�7�[�R�=E�D�v��\&$"*X)ܮ��o�٩�=�N	?���)~ԕp�Hb��l&!|��}���}Z0�Qh���ӊ��_��Z�q�{���1ay'����KN�����%H���'3��3�K<r���<����l�DRɮ����QXµ��Iˈ�b��1IZ��wMN�ʙ�1/84������5����X��\>|�q�_h�;"R.1�g���f
���Q���9(`���2��ϫW(�lyĻ�������Pߊ@�=`�g_H�ِ ��v���^J���ղ�?{d敹%ۼ���Y"�WȠ*���a$��e:X���!���V�/oo�@M̓:V�R���]�ֱ����]ɗ�vr��	ꓵ����86�Nv"0��]������.�
�M��qV)�t�c/w�d�C�|�p��cF���������wf�y�Ry/��ƪ�2��>ϛ+�"�&��4�;��@ ���KX��70̀�!H]�}x�ԃF"&�+��6�C�>�a�\|]ϠWL��y�?�H�.��*Y���͋/UdZn� L����w�(�r�H#GB���C��������1�.���5}"���
s��L�H�>��[H;W_�ޱk�[�-jB�m�
�%�3��y���o>u6�=�VTq�Aіڋ�Go4� H(���� v�� 5�)?([�����p]�@H$��gq_0��"��ߪH�ߨL~��f^t�潋�E�x�
 e���? ����q��R@��\raj*x���;M�[�����3N��P�����jB�l6�S8F����&�w��*ř���*oL(I����a�Dx{���vrf�]�=8g����Β�-]�� r\&��|1[�w����>� ���K�o8�G��q�9�*�����T�SA�p%}vr��8���fr����w6�`x��~��h���K5֙�7���+>[q���H�j�_���G�_��z%����
ТWB;���ar�c8ό�o����S����/JPbC�o��Ƨ�e�����,�59��}�<l�ڻ�ˆ���<|�&V�g����l:+��<�>�y2��L�(�NX�����o>�Ԏ�~�*С�1��1��:������z�;��cA��?���
��ie�ط��>f���"㢇|p�%�[`xiER<� &5��r7�+�#l\z�
�~�3�؂�&�H��РX�����h��%>�8�Ԡ������=�_n��_F������O�ˏ�����у��#�#swTX6�8�ψ����c��<�� V���F"������kU�#灐/D�w�?�J~q�T�1�p��2C����(X���&h	�.ET�Z��{��#���\Ӌ��#n�����B)p*Hk��%Ն.�w��μ�
����nҮ���|Y$����IK�s�����DO�6�J	����֥�^��3T��N�"Ccq�JY�꪿̉3ќ��2�X�Pz�u�Tד�m?�{e3G�e`�����s������2�TQhu����������:���㙑�&ʻ�5��l�TB����QIu�J�����
 �,]�QBL̇'����+-(�Pd���ǌ�m��]s��>��K�o��	�0�!����#�Q��U����^;h����5;�^�p���I��}�#��e�؉�36!rc"�����\֒;D&� ��0HD��@�%�_>��������B+۩��g��I��
Te��iݭu�Z�,��Au|-��Q{�m�{�9�-ܗ� q:��	�w�5��5ޭ8����jh�ڮ���ۡ���%�R}@Z�+ ��-�I�Cn�C?6e�9�>B��Ȱ��42�䷄��f5D����\�W����fY��^��ι�
3��%���|����I�b�q�(T(5��
{�o��o�i^�NXV�����>�X�}��|��i+t�1��v�nη��@�V�X�j�����Mrc�s`B����ǪI��z�`�sA-!��Ip *��J�v�x���"��-F��B�����ȧÞ���/�p/*��N+(�C4���oy"v�eE=�K�T�H�\h|��4�潧���G�]#JJ'������PL>)����~���|>{i?�=~:y�>z�<�JR���#l�}#\<-,�����'�[8���4�����p�@���q�zs����P�E�~lo^��^N %Y4lߵ��C}=�'#"mj~$˱�,����ˇ7$̈́Y�Fi�O|R�蟕��*�M�Vp7@���=�^��u�=�<�H�ȗ��쿾 ��v�J�Cq�����_n�%S�+�b�,�<	���vrt�M0���̲\�Y��~�aF!����K�ҏ��+�&6Oe1dQ��8c�F5'���z�K>�� ���jggS���1��𓯒'�F�ꏧ[~%���=pGkP���Z�i)����z;}G��H �����H3c�`��2��QN�3+�H"�y(�Ϝ�q�HtNJ/��	�$Jӗ���*BQ��wa�K��&���t'�DQ(��e���-?L^���[��N$��½t0�m�!^ e������"z#�ʆ�Һ��"J��`��&b1���/v��Sk}q�c�i7f���
�+�<�Ti��I�0��,5��n�*������Rx�'Pz�Y�i��!���G�p���O����)q�Np�B�5�������w��S�Ѷ��&��p&��p��zةA���r��͟�]���κ�v	2+v��̿��y +r��Zho���T�6bV���|P>A��`�^�G)BE/|�&gY��Fp��NO+E���{	u�S�(��ا���.�3�|i,ĩ�T�C��;�V�[5T�Z��oe��O�����LA��9,��U�;�۽:��G���;[,��bI�o��z�.��/g�?Xq(�op?�]wiɽ�Ř�V�Tʆ�E�ac���t}�`��.�!J<
�-I����w�m�#����Ɣ��&��ַ�t��x��\��?!�e�5�	���/uӕ�c�#�?�{L4����\�e���n��,±�*����>9	��9����ZY����ٱ��D�Ң���PA�3��l��C�|-O����9n+���Y%���]�����!��j�˳�F���G���7E2��n/��_���).k{J  :bք
��W��Ǐ6|x�̩4�q���
�����	�p:��l&�L��a9�_ឤX��w��:��OS>|
��;���"鄇��zt)��Zn��&���ꤪ`��g������Z�h�t�gfh��6A!P�ͫ�s��(��%��JW9pX[qALDR�	%�[qV�lѴ.�r�~r��"y`zM��kJy�33��R�d���'��UJ��/�g���߷�zm,�ѪK_��z#�JH9�i�[������/�1'�:�?jǗ �T)F�x�2�^6��)��,%��@8�PR��0vo3�j�o*�`|2�|~�D]T����I�.P^,���*��<:9�_��d7�@� Y�Rٲ�[aԏ���-�-��92��� g�����ɉ��1'�>c|�E���?�7ZV�6Ϟ�,	х��&��D�\3�tQ�|k�!�CC`�JCx��_C���/�� \���r��!`�bŲ�UI�ۃꨉ�)3���F��		��z���N,1�i�+>h�>Eq�}G/�xY$I�!����x�S`u&�1���E�t�G#��{G:�SK�'BL��h�]��U�m��PB� �~y4vpΠ�����݇dqd����#�W�|�xrm�Oy0��Ti򆼉"���v,p��-0�j�9Y���J�g�&�7���ġ��R�Lȭ٬��CH]p���%��%��3�R��;@-�?��47
�lO�Cn)� Z\	4���Bo�'�v�>=���OH@���4}����w,��=��8��>"�z��.,%�yw�z��~(��x�#�dU;��`9�G�Pj��,���Γ.��Q�_���,T���%g��^T~w��Q�䉡��*yRMg���X i0��M7�n}#���'4�2'�È�Y�	z�'�P����xH��D��$D�J �>у�&��Ϣ#,k�X�>��}cdZ�~��������22��.��p)Ȫ�Q�Q�8V�oiR?��H���(�>�+�}�����Y��Qp��ƣC�@yՉ���'����oŝ� ��Eͪ���*��p�G�݋Wf~Y�Z��=���7�E�4t��zX�1�[{����yI뗭Z�T-4���u��h^�r�X�`�M;;S��5�3_]���+,
y���	zx�PŵD�S�U��A�P�E%�3��ގ�Hi���["�,uM��+y9ػ��3}w~n�~ؠe��ž�6��G�+��I^YY��00��[Kj�������>���ڜ3��.Q���sv��o���ƣ�_��i��U����f����...�Ѣ_��Tο(͏�HΝ�:�1�s���ã䣩�IF��Ok�%&�l���D�"�!�1?���)fse�'��{#��?����A������7����c�A(�Y��2��bL	��)d~�n*���},�o�Q�wr���:���:~�� ���:Z��N��ј�>W��7�v2%=c����T��	 �a�
��i��:ߛ�b&j'6]������`d:�*�غ�(D��C�����Q-������2�-��]Ͳ0uZY�j�:�_�1���R�w�4"w��r�5�Ch��ē�)�/��
�Fg�x�V�
�V��<�b� ��z3(��������m�]_��"�,����������z6����P�������J�8��㟨O�����
.��+���y�$xT��"_��?��H�/�D��h����g���NOL��V��҆~�kE�߭�::~�O���n��-��U&>N��n�?n�o���͓�����~f� Ξ����MG��`c7!c����C�D FR=H"�~x$�?���d�L�
��S�W��I�H�
�/�,s��R3uU�h�ߴޅE���F�E{�"G@�lj��?b�MN������h&5ޱ�U��:��x�ķ������s������M��`�[[���]�~޴��iP�mEF�:N8��Me�o��+ȿ4w1�W�4 �z��tW�!O�vz��Gx�㔞~T�������!�F�&y��nM�.2��u9������P��E�w�6�ܻ��.V�]]S�\�q	޺RS�K�Ú��2�)�8�W�pY?���f��X�P$Rj5�n�l'�<�(+�4����yv�C)���A��o-f��k��e"�8�`�ap�M]Zi�wX�33l�!�G�M����6D��`��j�98�6�tƘ���[1B�[@�-�Č0˵�JJ����,�Z <xd�Gh.��xw�ō�Uu)aE	[G[��)d���:˨�������*]J�"
�� ��(�H�� ���(5H�P�#�C����������������ιW���/x�$m?#���'�O�^�)E;|o���Jj�K=�Tƾ���tLY�BBW�n��fc� ?dPV 5_���S��6���n�q�7�C� �WUTu$N��(̯����M�*�ʃ����CC���zR��(�4d���������9�Av7��%����y�}���S�g��>32��?�(�3h�m-u~~�l�����o׾J�ܲ�zi$v�zy�xC�Ԇ�o�:��m)>7�iM��3"�@BФe�h��R�튅����ݞ��xBB��ï��	6����Z�Sk,j������I�\ ښ���N�b�*�����S�O��'r�J�%͋� o��CQ?t�����ܞ�[cꔁ|l�ʳ0�B�Y�Q�p��֕N<^~�Z47)�z�$�����C�T��Ծ���6���|_��4��̟���M�C1f��yX�qvx�$�w���3��D���Wױ7�[y��YC*!�j����R�S����(V�k6�u��+6F�\i�	9#�j���'���I�I�m�X����\����m�ճÛOU�9X��K�* ��o�|ҮdE܆j�w2b����1�<����Y��lJ�+d��0���J���� ��VT�ْ��앸Q�ͤɚ	?'����ŋZ�^��W�R����k�Q/WGz�s���	�>��[�_�߽���3|�BMڿ�V��{�Z�V�|}Eٟ�7���{��ICyk���]ή��Pq��A�Q.�M�լ��C���*t�ލLL��������gܣi522!n>������$r�u�n�'0��\��31�S���R��>�CVE�hFn�V����2�f^ߏwb�E��	�:��@��;��#!k�>-%�_jE(�������i3+��9j�q���'�Ev��y_��s�6��D!�u����tl����XRy����{���8�~�)��|�w9�\Oa��53?.�q���#\�(�}t��ƭ�k��_ L=�́����u��+��2Ƒ%��+�&$�#@�<Iwg����q,v޺,�^T��j��C����E4�5~Qƚ�����3YE��d���F���-���ߺht#�Y_r�l�zXzW{Wp�le����b�X�p5�u�c�gv������F����uP �Nz���5.�T``�g��~����F�:G���O&�����jW��V]7�vC������?�������sܛs�s�'�3�^*���y"�n,�%|���8.h�����E�Q����g��>ቩ^�0�enJ�C���"L=��;V�Kv򎼤Aa&g�B����k��5���`'�A�}��\+���w*�W��}��^0��J�C�E?̖1���3$3��]3؃���3�FB4�s�Mټ���?�R��WG�����e�
��&P56,��&I_��r�$��irB9��{)&�hY���ߴ�%2���5ǲ���?Y����L	�e��(��]��yyfV� �}�BVV�* ~���4��-V-���+t1��H���[�][#Ϥ+s*q�`�v�A\^��s�T�׭�R.3��K�Ag���
޼��lJ�Cj1�[�e�&o��H�
<�L$Vk`�}�ntK��΢��d��D�E��Y��Qq�-���M�y��y_TT]Q�Kl�Ӷ7XGZ���ݤ�x~LL��=����p���x���JIV�zc���ޔ�<h˸t^+z�.�f��k������8��jǽ�-������i�m��)�[ЀAc_Ax������G�������R��^'��:�����&��ۼ&p0zZҚi�6���&'{���J�9�AO���S���30p��fڢ�V�ğR<'�='�w���D�y�����i��-���������O����4�֮����@7��cp?'J�@��.�B�=FR�9V�*����sd�%��y�0��0��0�dp>�;� Xq� 5A�������A��X\�Zg:Kl
F�СO�9x�b��]�}�:uϠ�K�^<�-  ����7T�BLzCZ�
b��KY�����!�kK���Z��5>�YW�ï�p$ ����Z3� KԪ���k׾m���6Q\���k�����RT�!�D]O�@�m��o]��{�j�7O5v�*����/_�+�mV_�x���|mo�H���O�0��=c�;u��zj��f��Q�9�%�%V��$����w�ș��ېh��˒x�NK��������;C_��$q��г�lwɠ�Ow�s�����ݽ��פ`�=��F�Z��©�C+!�8ē8�t���6��Bv]��b���h�~:05v�%�r�~�u�U0��dF0�h� Q�ݶ�8��[��JJ��HM�|s74�\.0a��"��UW��:hzn�s�
����}gU8o�Z@�	[������g��7�A����bs*ۗ�Fܮ���H�iM� ��Fg.ڠҐ
Ԭ��1�rG��<�%zԍr����!@�����l�#V��{-w�%���.�t�����|�u��K�*�����ѳ��p*��$�.��/
�Ls��TsT�x㊕���I+��g�"zj��Y���C�)S�L[���� ���R\hQ����%I����Q�:Gz>i)1�����('���>w?[z�������ܣg�	�y��˥��`�;Q1ƶF{5iGe�I���y�6��ެ�sG��'�8�zu������H�\����ZE�u�]��x4ù؍�48@ʡ���N,�4����Ꮚe�E��
K'Sh��>bX��u=ݭֵ���5E2Ib�~h.T����g�!����)�?\�� ������9�O��%�R^Y�!͞����o�v0P����N���r�2<T�7-␨u,�Q�Aw ����KR1=�^�&(~
�����bK��r�${�p��]�A�oO
H��1�Ap��dKg�Ŝ̀.��E*�'�/��˧���0pjߖ�2��E�a�S�#�����Z��i��S嚋�~f�U5�-Rp�
qY��f�2K�֟����@��H��XQ��9�a��j�}2'R��v��{��Ѿ���ϝ��M�����/��.!$f׆:��ri�PƮ�Ҿ�','n7%Ȑ�\�y�%��eC��Ղ��=����&)��x[�I��+qө�665o����ɨ�#ގ5���M	5������62���t���eǊ�����QV$�c=��e�1�+vg�,��A�:�����>���I��Nz\D�m\�B׬��G����z���P�k��%6�*I糃�we�b��Ĭ�N����W��d����G��ʨ;�C;�雰�ز-._Hыݬ_�%!�*�����.v S/��t5v��B�2aE4}k%b|!�����6e�B�O��������~���*�|U��m["���mKF8aԺ��O^^}>UqR[��"P ����n%Γȹ�-&��XǀbH�x����%��ik��X�$u��	W��~�<�>����#�&\|�!�P�%�ZǳXo����� ʆ�B�.ͷ��6�[@�k!��_���yV�-/a����F͖�� �+	���t�'&ߝ�}�$u��]���c�v���<���Ar��bfPD7���	+e��*�=1���W��rgW����v
Ξ;;�(�ZU��ȵ�^ݳ�C�٥�����/���l~�d���*��<���pz�St�0��1���.���%�7Ej�-8����ek�#Z�3#qje�zOhj���!��`h�E�͔x�n^��Zб���/
N�R���|<��Ĺ�𐠱�\��5�hg�U-�G�ym�J��q+�J�݆�N�F��7p��	ҩ��@�&��|I��GE�=���6�+��y�M���˱Xus���jN�In]Wo)]|��c����y-}�Cw���ϵ(`���k����L���yY��}촼��H��؃��+G�i�n��B��/ u� �ML�ۏ�����|�u8�Ȁ��f��j�]��M�(�,/�t�� �D�yJ8��؋�=#�N�|�TȒ�ݘ���>��&�*��I�%G���P����2F�L�RU�%�g�h{v-�0r4YW���62[���d�1�\n�ϰv3Y+_J����Mv�4Oz:�����M��]��]hZ�$������|>���{4�����i3_�Wp�?=�g�98E��ھ:O-�T��!Pc����e<���d����~�R�8��EWD�45�"����Gtt��A��ey���%=ܙ���r�$Jj�k���S������Y�%�q�����j�t��A�!x����xxW6�Y*5$)&�鱆�m���V=���ʆ���t��]����;4ick臰�q��V$@�R]k����:aP"t�gA�Q)��R�� 鬖�������J���a�h�7�!�-w]f�<��sks�tD��1u��]��p9&�_?��Ŷf��č�b�����ؓ0���f!�- xT�P�k��
kr)W�q�NM�x�_�ǞO��0C,&�-n4W9��Gi���aυ-�m��h��"�G�a�E���=�{�5a���_-��{�:t��^K�5������`}o3I�����Iq��M�X7�R���>l>Uy�L�b���s�F�E�8�t"�^ح�M�K_{LT���u�j޷$�T�lQȥ�63 ��� �!��*���u�L��M�fz��z �5TW�fP7te
����i2����a��V��1qJ�~�8L8����d�7׃>��c�8�fG��᪣5%����m�y��<dZ��2g������9)�N���oɃ��STJ0�,_++O;5g��s�f�J��\U4�3sd��BQ�k�ëm���>g�#�`4�A�f��������rv��&����e��c����J�� ���<e��)ޢ:iϙ��H��Cb��sȅ���@@��\�+��r|<�,QU�V��3�M��Zc�bngU����A�IV�A�%�|���	js�Q�LHB��7�a�x��K�Ԩ�Ԩ��#�w|�m�<�2cQ�9���D���p��ѩ)�c��-���(S�Ǆ��yG`g�c�����;ݻw��>)
�%�	?&X+KU,��N4���0�a�tnɏ��G�r����(�̐���T�Sz��h5�.^q�|�K��.���������s��n4��`�B�$�թ���UD��`���\`��F�]���ڛ�T�/��ip ��tC���HTP��&�B����j�Ƌd�=�2��w�z|��Ԍ/m!�*UO���9u�y��N�J�
>��5����r�����<�S�2������k��i��i+��EZ�^����P��g��7�}ݧ�u����<�/Ut����xX�ڃ;*����f{{x�;��%dz���.�"�_ ���R�\(uq�?�[�e��V�i� �4�jV�h�rJ�J�*���AlN��h�F4����>���.�o��]�*�Ls\�|�5U�u �{���T�K���%:���d��l��CC�[b�В�J�D�せPԕH�������s�RjJ����1����M���C N��Ӧ��:��p�M��|�#k��A��q�c�����֯��r��d�@�Z"����]VDyN�38oF��3f$��a��Zoa�D��r��QK�y��YHI�Ջ!q�T�V�<9'��L[��B�{�E�P����k�8=,�%�� �-��Z��M#�g,)i��&ݚT��Àm�Jc|�R�=��Vi���r<�*Z���V�2ǽ'
�����d//��6�>��}���8�3�pTC��?��A�ţ_��j�<P�r��S���"՚�h���jrX��z��t"�v��\2���@���)�Q��ND��՜�'���g���%�T��㌓O-GA>6C�FT7ߵ�Z�2���Fl�d�>�Ǉ�hS�~Ɠ�]�a�.+�
�RO$gupT�V������ymc�S�.1ěa�0���,�xg4#ʯ� ���'���6m��\����Y��)^�md�9X�bۜ��F�	��=HO�C���J���B�&]�)~�X�9iVWfW�y`w��o�ş!�]σ�`B�х��
]����O��يS���@�.O��,�wW]�vH�����V]|uC��vS��Y'�s	II:�]j�1�`ff��h�k�
vG�oT�.��\R��U��,÷5�K�{k+��Q�~�\���T;_��*2W����M�b�I�ޑ���N>m��a'X�F�o'��\���p9���n�u�{h)-N:q'݂�G>���tJ�0�oqTu)R��B�&��1/
�[�|k�i�����L�i�Yԯ��fmϽg��r�����ͥUWHw陿r�]J	�wŔ&]�q��3l�x��(�U|}�x\�[��O��k�{�(a��2��ɹ�ۮ+῵��m�(Q��T��ֵ���T���_Y�N���]�bk����X���Խ!�����rm2��������Τ�=��v���M������u@�y��ڱ?�����[�S�N�=t.����p_�^�3������۾���˻�&�j|�<c>|d�߁P�����Y�v�/�{]6W,�\Z�Zo�7�C���s��L;���}�ԝ�V�X�"E(�1��K~Tj�G�Õ�R�(�>C|b�"���A!��75t��҃��� v�̮Q��e�$V�}E'ɿ�"uL�e[>ˊ�L�fx�u��T%���I�n�I��3C
F�E�=�jǖH��c�V+�@<�n3��`
	C��2�r�[ڟ���]�!�c>�燧_[�S:��������&�^W���h��aZ��8�t���O���G�=��>���{n�j0�_c��謅�!�jaսsA����T���gy�v.�}�K����VF����@�k�!��d���e�̠��� 鈔��sbS������'�;�r�>�3�|PU��@dS��G�A.�J	b�8~��	b�I��+�F�}�~��)o
͢mj���zo{�w��Kg���a+���vj!k~T�op7=���YF��?Xs"|╤,�����\{�
����U�aH�7�ߴ#�%��MY��V�bu)��D\�֣�Z]�Z�T(z#+c�N����Vp��ΏDA�Q��J�'�J���q�!5�R�	�P�$�ݬ����x�b��'(8Jo����ʠ�ӌ��|�)��1h���p�O��
m��{������Ƚ�X޽�����܏�[:�S��{�aA��◄��x0�Cj$�6�M'w̹��E��:���R)�%�S�\tH� �x/�{Z�ԑ`��~�f� I� m/�'� �P	��B;���q|�%L�d@8���#�hK�Z�E7��3��w�T�nJ\`�A%'r�[���6�����[�-���I�w�`�#W��b��6, e��lei����M4�mD�c�0뤸�n�D�[}fC��,�-�O\\�S�n�Z��@sX4�W��C^�Ξ9���ڈ�W��:&�ٿ�3�U����:״/���M�$JX/?�+x��}�cayl�r�6Ȱ*��7�	$�F3�[�v��������W��CO1V��ʁ�y$��*��d�Dȟ�ZLi��B��)����[���/{6V���[A;b#�퉹Y��<��3򦚌F�?�W.�]���S�ࣺI� ���/�,$&1�A��w C ���]�n��P����4~�#��m�`rL^	�
B��H)���P=�t��{�H
��������Fj�otv��<�U�YP����gg���l i:�g�'1oX�W���{T�7��,5�⏱@$7�5�2�]{[�P~ۀNLf������S#̋8������Z�Q��^o��b�)��I���"��u�aڦ�j���.	�M���Y���+�*�n|�:b�����y��E�����-�H֨\Γ�u��H���q�'�8Cjg���*+��N�6�ۚة5��@�E�X�z���L���f������ �[����I���2��fpc�޳��j)�h�,9p���b��L����l�Y��\�!�Ya�ɗ��HIV۴��]����ѧ%�9g%O��b��ŽJ�e���&���p5� U���B}�އ}��ߺM�k0��˛�Q��S���u���#�:�
�ִ�7��R��"o>���z{��ϒ�_-�����q\����˔��:PMxB��X�r D�*A ��q��F�W%��T#)��ͫ����b�����g��� 0;��kq�y�`�17�����&���Y����Mй��N@�^Q����-�����v��T��ō����&�[�0ylj�	�d���p!�~���b	C���wQ�����a���1/�/"���E٠x��fJTh�'5Q
�|9��J=\Kg�K.���;p��ݜ*>�a� ��lj�.��Z�w��ho.Q[����E��6[S�C�x�&"�W��E��Bջ6� U�'O�,���^\j��1 ����^n��[�s�xЈ�F9����0����R��$������*���õў[��)��S��۫���+^6 c�]�[~�g`dfV�.�����w��x>S;�̾L�-�gj/���j�0}^������ �9<1���I�rʔN@�'�ޔ(�|�9�g��;���_dG-�N&�-;ܷ+��]���nYn��j�W�D�d%���״�LR�U��)�d/���;>���:���?0���W;ˉ靗Mo�7�)��Y�#�@�!�o���9����]�[)
wI�:�ʃ��@j�)�SFK�?�u_���'�*�n�_~�#�޼Cw{;9mZ�>^�ʅ,X>�]2_3Y2M����5�,����~����5X�$:�i"t(�)v[#Աm�fN���8b��-\�]�gwa%������)�e�*�J� ��0A��|��j]�覄R�ťt~�pA�G��Jl�f�0C�]tbه̃wF�*�����"G���M��h��L�����?Q��o�
�  �-k�I+:;5�o�Pl�o�3����t�Az��}�t���Ȓ�[쟁ݯ"���m@�Ob9�I�~Oåm���&�n�h���[聐�E?�3�����֊��/���HY��=�W:3�&S!���F����Y���o�?�7��'}`�/��Q�?��n������&�h��� �m�ߨx��BR�8d�^?��]���
���N~M.X�I4I�3�_��$�0W����n���s��g�����	T�+��#zh��0}�hq���*i���Y�a�����6\F~��ob6%�]�,�N#�v�y�d��!�>�8��;6Z.�(��՛S�k'�y��D��T�_����m��� �H����7��iib��Aln�X���>��oH��py�`滟_w܃���p)�:�]��j�w&n�X�]���מP�Mwqrb��+��P��O$���S�a��+�#\h�	Jb�1��	0�k��P����:nP?3~��9�&���\�F1.-@��6����,��S�Q�B�^�b���g2�� � O>�&���T�����>B%���&�F���%��>��M�*&�)},ءJJ��i�-ZcJ.K�[�R�፴��u�~I���^<d����2خZ��ep�%�`ߋ�j���E�rlD��n�ڻ4����d���iα���0Y:���
@hc���U�+|�4����w���O����h��Eſ��p�����?C�?��4����_��	m��Δ9�o4�e�����¿�Y�
%m�E����$�ϰ8�L�:�>�@>����D��%���/%I@�0:�๐W�`�� ~
;����[��3_���j��"B�$�xA"���E9�U"�RO���X:��lG�6NM�xL��M;M�g���}�I:>G��n�3)�#Ks���8 ��	�s����EK#�N��s�'}�+V��hA$���$pݨ<cѝ�VJ��Q�%0��'=,$er('n�aW�pusp|�p�}��?��������~���H��oe��� 8Wv[�����n�a���=Έ��&luw�fɠ��[��/|JG����V*>�q���� �ew���H~ t�WM��N�}���)��ԥ�YO$x� �|*S�h�oTR⁴�c1�8"�R���V��"P.̨d"�菏c���
���'��|�3�!���M�.�����s��pԾ�oD��f C�\�|�KdґO�'h����b@�4">T�9킃ǺvDk��5��1�̜�����bFUho�e�g`���w��V���=����*T_��t K�\�z^�Q����i����Lm�U�ٕb����!�t�MT�0�=����ϊI�'Kc}�c�:m�T���]W���#ȔE?��x+cZ������N�IVFy��ʿ�N��qx|Q�?��1�l@p߃:\6M�{�r����� G���c����Ωr���4�kv��23�Π�����&a�|���j��	�X�!�ԍ.�.u�/���l�*�|>c�;#��Gq�(J.�%��f��l�)�Ǆɽ �o,�YDc���sq���q��iN���/k�c.��������M��PT�7I�	Ҡ�|ɒ����qo>/��Z8q�������H(�}�9.դ)n�̏���_�ت�l3�Gϲ�K�v��� :l��E'HZc���l��jd�rY�v#F:	�~�l�����\�I��Q�&��u�f`S�k�BK�!h�ק.&Ӌ�����CЂ�f�b>73���S6+�}c*�$U���f��V=87�^�Ҏ���C{�?��F܈�c��X=��.M��G���BfG��ǹ������PDm�c�L����?=��e�Mt]jږ�W��C�U�G%��ۡ����
j/~�`����̤�A�nY~�A��'&�W8���)Ƥ(�Q	�(��Xn��;3D`�SC��a��V�WkT=2Ӄ���߹d6%�-�O�����DO�,������4=w�k�=�?�2��p�L�����B�u>�6��;���^����%X1�7�����ʱ6���]=֞F`�-u�p^�����M r�GR���Џ�/4Ͱ8�j�}iQ��;:箮�<�#ۭ��t�&ү������-�����W��=����U��URC(��r����q�n�8j��+z;�>�fHD��E>�Ĭp6�9騅�+C/�ο���^8��(�S��F)*�b#%K��ڠOXY��qk0r!5�A����-k�_��}�1�A9� U�Q���R���J���
Ki�ar~��9حWxО�?}��3�t��υ������C4-\����X��%s��mK,����Q��h��]�D�5?�L��i�a3h�r�D�O?�v~?)))$���k5����;lm�>��2�}����x}���Nj=��镽;��/�� L�z	����,xq��W{S������Dl�I���4S2��rX<��\6���f�,��9 <aajD-��φa{޲�����?[��d��W�)FZ��j�t@�q�+N.����Aj�	"���Ʉ-N;X���=0�^�yIgࣷ�^��������qѰm��]V���J�2�`hA�����۵-�Ʉ!�O�+�4����p�%��V
8�|2���+�
���=v囃w��W<J,��a������:e��+�ӎט��w��RM-.�O��NaqJ)Fo�ٱ�Յ��٠�x�������>u��D�m���Oq|�Š�4a։R������?ȏ,�U��e���S���*eLx��%��$�5 �7�p6Z���R��N�O��nz��5}'ڒ��9i��J+��@-�6ݰ�^�|�I���9�c�s2�}����iQQ�T���;T��ϯ��^���9!���G�����5�#���E����b��a�Q1������.�i,z�^���}��)*����7�d���=�5F���c���|>MJN�V����tM�/�e�btF����)R����u��/=�o��$�\Bh��M�
i&]-w/�:#H�K��^�����^a��+��h(�|�݌��AN��+Y�X�C��= �G�� �{���;.�B�ޗ��иW�_4*��	[[���.�Lm3g{ڂPy�^[K�a�S)A����{������8�x��D?D�ߴ��1X12�#z<��k��X_�=Լʝ����8�V����h~�$_r�����A����:�9����3/��ƕ}|h̃a�;�\�����I �nv8� 06�_�םg����`7Y�]	�������ý4�e���o�km��G�C�c=<�����u*xM �"�������Px�Lv���JI�#M�x���~k��-���6�̰�О�n(����~~C��������U�����`��=aGw���|��
��a���v3����:�q�5�> tP���'�Ű��M4�Ɲ�O�}#��E��K�M�ˎ��!����UL�>T�P��fxվi���2��'�ن��}槀�M��#Zc��6}�栠O�G�������\t���i��Ȣ��ξ:�I���������5V�.��H�U�Bl0�ZYT̠�:ύs伤'(��K��}u�Ө/�$�/��~Qpz䎑���Kn�ѥ����JEv�y"�4rc��}��A��jZ���`X�{�9܈�/8��a��=�ê�ȫ
�ɗ7���Ke��	��}f�{χR�}�����v�0n{P�yk�� j�5B� +t4щ�R^�#�i�]�\_,9����I�>��;�p
�Y?���f�f�!��u�z���0 �p򵡂Nw��2�H��IƀHa��s��ǎ$��C]�~�UT�.c�ۀ�N���B%�S�:x��u���܇_5;�Z�w?b���pi��i�V���J�G$z(��Y�W��~����$#���FK����m�m>Ƌ�g�]-��s�	�d���[�k�>ǲ�;� �+n��F=�m�!��RQޣ?��|Y�ᛪ�xK�}��`"W�q�����������r������R��xu����!%�������5����U�'12�(-�-x������ʡ�v��t��)��'�g�ﱁa4���e!ou����s+ڸ(by�³�h+35�v��Iר„�*,���
��w&�`�9�O'z��-�7!ϳ;&�?���x(lΎ$'��g��0�_�@ZGx�m�<j��H�̊��!��ر���\ý� �e����H6:}:�{�\6[X<�5���Q׆0@f��k ��7�Ll4{�+�Qɘ��ӌ��V�CN�[>lĠv+��0�����I�QǾa���6Mb}p��e�Z�X��w�?������o�dAT?��Ϻ�-�&k#<��'֤<��e�����^��B�ǧ��lVi���1�O�5_VE?�LgMz,2��h���g<Sd���� �yP�Ⱦf�%V����eԐ�笘�`.��NM������&���Zt�����|�7�އ�����y�P3.�ɥ_���l���p6.�Qc�'�LG5P�o��h��ٽٴ�b��G�9;2���$��)ֹ�:S����!*�Y4eIL�7�\��%����|\�\)������� �$Z�'��:-��<}d�{~-�>�M�ݚ������̯�V{܎��4�V]V�т�2���&-�+��k]��Wg�G�Z��m�d2�>%	��z#Qa{77Q�QV��7�e�@�iEN��'�g�-%�v=~=��-Jn���@mG� �������:E|4у �^��=t�C�������Hn�@��l���_�H�+�� WZ��:V^1L�V�F�7�F�`tE��h.�����F��0���L�w��_'r�h���{�n�:������X����&\�h�l�tm�#"fճi�[�4q*�6h~Д,,�)}E�.���������ƹ��dg9�eB�qX�Q�����H½�Ʈ�F�.~G) d�Ӭ���t�H���D�+3���5Uw8�8s��sTʿ��?�{�������:BU�zqȫ�)kF@=Wf��D >f���Ԩ5�^_b�w�W��ˎI�>>�8qh�Je�tn���g�s�7#�/b���Š�K����ACHs��]P�f��i'�9?:���=�g�3��>O��X?o<��Z�
h�����-��0f��_6�#-�Պ(��υ�	rY�˜~���A��]>ո�\���Aӹ�֤�������X#ކPa�{�3&���q$�'x?�5L�u��Swov�$�*�G�'٪���Q�ʩa���6�d����3�+xv�&?�fW-�A�r��Y����.
��W��MZ\>�:�N$%�fu�6��ۃ�n�mZ�f][W����:���G���O�z�T����j�Ec~z�����a30wNt_���������Q"��hJ1`.г��#����^ޒH�� ������#"�3��6��a�dE*^�8 !k��,ۃx�ݥ�d��\h�`˙�5��פ3BƄTC;�����D3���||u[��ќ��Գ;���T"0�lw�4������Z��Lt���;5�Rb\;Dٌ�V��&�g��8@�Okȹ���?I��邈N	X��t{�N0�����h���܌�;�)4�'�$�P"�_�w.����E����t懋��A|�w��bn�k�J�f����y��9�nޞ#���c6���\MIR���c��\�@0�PV�A�x��m<[<�qvϷP����wJ���ÏC����e�Aj�O�9	'��e��H�?����$j�'�!�����;�������H%�TKh�Ii�[�\j$/�����?lSE��Pk��Ztm~��D��u�UD��4K�߇Z���=C�d�˕�?I^|e���$7�|��F%���Иp$�HI��YU��g�ύ�9f;<C0�0�Or���Sc!�kdۏ��`��޴�U�Bv�p�ti����+�o7i��q*/���o=��d8������%vV�nQ�$��፻�L�	�}��t��v�t5�/,� ��t.%�ff䍈���sc=;p�&������®�i�@����B+�)��WZkRuk��>�7|����l�cp��
��@O��5��J��t ���n�x�kTsm��0(����Q���M+����%J��Qx�/��@L'5w��`�EV����+t�Κ���Z>+ֻ"ļ�O����p���m?m�j��Jv�O�/]qͬ6i��M=�K����Y�jjJ
�CVȎ<��ׯ����E��Z���jv__�:�{�����ĜŢ\/b;�/�ζe��aB�L����i{���aee���=S��V��&��L�-E\��O��/���]}�����_�$��L�L���D}���4��:-튋N��K��J�D����PB�f������q���[��1�D��˕���b�����Q|M�&[:5�_׀?yg�ց�=a&��B_�FL��"�o���q��Q�H�Z���������Z��aG�>)����J�t*���V��,��tFˤ�T^'0F1$RM����j�%@���`㨺��yR�I��NZg�(�����7?���L2�l(�Eu��h
�.��M���y�c���w�]�L+k��
j�D�vbjb�>�g1�8\��΀���JJ���A�P5�j����{e~�D�/�Ϊ�0ຑ/��K�C_�x�kC��|(����'����AK�Hp��� �n�u�m{�I �Ī0_���S��vi�Np��S�$b���f�F�¯����8��c��M&T���|s��h���~�$e�U9֝⭴����<������'�8C�B/��XF��kb��XG�K�����"�bd�=%���m����AW�'H뤙�s@�	9���2s��֖��?��f���E��GI�w�^;F�̜�Ψ���ߗ��y��{���ۯ�q�Yy9�oY6�j�v�{�jk*%P%G�'�c@��<O�_�i������}yʏ6�lm�Fb�AK������/L-�v������q��εF�{�#��(t�P*���c��:�a�%L�RH���� �pq�"oN�[���K(�G$rJ�P
Q���j��r3PC��H1-�~�Co�6��+`�K�/̥�e�ku+��K^N`" ٺ�g{L;IQ�Iۇ8�쥥���4&�?�L�^�z@Z��(hu���O@��c`�b����w����e�y�z�Lg̃ͲR��+�  #��aK���<7�/��T��;@e��s��x��l+`��D�Ȃ0��m���r7ZJ��ZP,p̹��y�;�ܗ}��q,�-�%}Ce�L�IJ���YmQw.�;Jc%�@곗�2�TS)��� p��ݒ���0/΄-W���'��h�&�v ����u�61����hi�@�&������fd�j�m�j�n�l����"c0^���҄>T�f:��##�Q�V�J�^��&AP�b��q�5�C��B�+U�2���c�BJ%o�u�f��W�4Y��d��ݶ�8c�~�T�ڍ���C7u�^/7�|�����~oll�i���0B<p���F��~�T�\]v��ewՕ;���z��?����Ξ�!�MK�dh#Y�t�B�}4w�H)}�<��p�'y�!xۀNK��?�!�VϒH�F�M��*sk@��~1�٦��G�� B_����'`؊��.Ӎ�t9�AL��D�
 ��1���]G,f�S�.��������c�s�P��R�A?�ꆕP@ߒ!!�Z� E�J���
�`�1��q}��ˁ�x���~-��S�c�/��;�˾ c���iM�F#k� ��Ƶq?�^[�����B�6i���� f8`?=���p<AqT���a.��!�����ųa������Ra��g�י�� ���;M��hrL��]\���!ŏs �x�*�8�^I�ל�|�~VRX��� ZbV�{l�DEs��/�.���]��`D�\	L��}�1
���^�#
 ~�Q�"�uP�q]��y~?I�0���uݤ\*AH�XQ�i�$��F�R�����:��49_�c�N��+�O:��I���(�V*�F�$Q��r��(�T�����~)��f����0G�A�t �U	�i�𢡊o���Ien�Si4�(��q�Ƅ^E�2A���{�����&�8��nA4�O�ޤک{��}����|�c��u���7l*�cl@� �����}�V!�,0����o8F�Wݶ���v�OL�f��XX��YYiJ{�-^I�R��Y=��l+�m<;�xlCam[�%n�;��j-[���+��3z�>V����L��T�j��s�> � ��s�b���2�	�q�j��u|��`��D`
	>�$&�faႸJ&&�D C�H!�%`�� 1�ӦZ+�f<�1���fk�,.,��E�l���?R5#c�~�{؋��) �n�;�G�������Z�eQՒU��a5����]�8��U~�0sa��1�ᘣ�������F����,����K@�k�
]L��1��5׹���Q�"�8���Р;5�\ccu�K\��� 9�:�fz��l�&)� w��
��U���Nƿ,������Zg�Ts�CWߑv�1O1nT<�=ƎYh#��H�s��{�3ח�f���P�X\�,
�O.��5�1i�����&�ӏ��_.W{q��Yw}��x��1N���F��^�����q�
�pet�~v�����˥��.9A@�\��~�i����$M[	�p�ZͤС�j�Ϸ�8^N?ܴ)�o߾��O��j �k_�Zueeeb��2�raa����$I���pK�ߟ�(�+Q�_��z><���&��_P
B��E%�����o�i���Jed���������҆�񕩩����t�����7߬���������?�O�(�W��+:�IZ�X��j�B;�������	s��;�B��mk� ����39� ���G4722���R  g�,, H*�>��2(��-�P�zE;l��{0��p�7��RpK`W���� �kC)���%��%@{!�$:;�R�ʕ@'�'�A<RW�9�i�5(P���@�0����Q��݆r�`�:�e�i��b/0��A��#��he$r����� !��7�� � Rk@��o*�* X�v]d)����%���ō���E[�sM+�(t~�O:����_k�z��9)�_�@���3� }��ǜ�X���� ��џNW ]<��m�.W��[" ��%Nh�����pc\�جHƻ��)�\�9�=is��uτ��F�Db��oL����͗�J�ǼD1�1&sm�Zļ��B ��z@����~c��F#;�5��ş�\4�f��0�*���(s$K��ken&�]t���Պ�?��+��@F �.�Z���i�q�ľ�IF�^9N����M?��t]��~/uҎ�:�I�AP=W��S�I�@�~�x��L�x��K�ng���q.��w>I�s�^g����H�aj5DF�r�s�ȑ��^��%�/|��[9��xn��3g������ťk�+ӽ^�q�j�U]� t�c�$��D��Cx&�����$�`���cb'q�(I±zV��_^.U�ˣ������\�Z;U.��n�8u�^�/���7g��Ma��NZ�V��x�:������}?���}�}��+�KP\�>8҈\����A�LRʶ�1�BW���j�Ӫ'�0e aA#��H/�-�0q$�����~F\����{bJhO��4�ψhrZ�B�!!$!���� <�!��_#3\
�� ����S��pm���E�q<I�ZW�{B"��<�].~㬰+,��r5�Ծ��P¨�ྫྷ˯~מ� �v�;&3�������_3hձ�'�9�d_�u���K�^���"��*�T:��G� ���9�T��r���)ۃv�"�eu���YB����;��3^ s�`���ƨuZ�H��Me�����Bg�"��L%���O��e�������e��8 ����+��EQq5�Q����?���-=�m�6�`h�q?r�ٿ�� ���9%���3���m44���u{��m����a��̠XO�c@ �K�΁t�j J(�!���8�֜����^\S��=�䚃�%X�ڀ�A��s�Eڇ>F��D@ޱc[�q�F7SDS���g?>�U�Y��Z�R/+����3`��$m�q���Β��a�w:ݕR�?9:9r�M��n��rݰQ*�Yٱ���\a���˿$�����No��_�q�٧_5w�����7�:���8�r�\���m�eAe$�[Y�rQ���i�ssfye�,�ϛ��e)���%/ˣ��K4��������t����=�麦Y)+�Zeqbb�l�R=S	��Ng�ۍۛ6M{ӛ~�B�f���v[�J�g��}����>q����_�8N`��`�`�2���M0(+`lIQ�������"��k��	�<��1	-8\syIw��U!+BK���>�u���ׅ��Ҳ H���� 5	v�"�!�H��]P P:�E[Ha�Y�Щ��a���>Ľ��s^r�5�����v��
���O��{B��SV��4�g�3��tA�gAhL��aYC)% ����ǌ
�
�*u��i5���GTF0�tG<ms��3K+�`,�g�3�'���x�Ѣe{IQ�$��d�c�����umJ�;](x^  ��"�'����v�I�Y��0~����P��m��A���2d߇�sllB�9B��K�嘑>H�� �� Ee4����P-��`@��� Ʃ�e} �1g�O?v�\��4<��O�6𾲲$ diyy�Be0��w��+r�mbv J���G2���}��H����k������
K�����N�BTk�Q������5�v�5��Ÿ\��*j#�L��/k�n=\��0|.�4� s�� Y#AY �F��������b�v��u��iuZ����p�^=�m���l���v�8�gff�Q��%|}_���<s�̉]O?��m�N�z�ɓ��,-/o��x�V�9�S2aPqilr��رKdEh+T_RZ饶�>��#����L,X�Uj%d�A_76�`��ž�&��%���{�v�]���{w�}fll�a�-�����FG��FFjK�֞љ�O��O7^����?��{����a��"õ!����FD �})�uD}Pӛߦ݋:
&9-0�@X�_��<
\,,F�O���0�I:��3h
��`(Z�x�}p}ZN&8�
�1�9���!�%��}aF��'�N�0�@�0��X��($p( ?��v�X :~G�2����X����l���X�g)x�h;�>�
)�B�M�8A0������b�p�<�Iw�R�E+�V%��f�	��.�4�
,Z�08�F�l����{2{p�A�B*Xh�*AM���o���.�Ջ��d���*צIŖ:���E[�����fZ��e7S8�(q~���,���fܾ���gj(d�K�u�/V�JJ��:]\\�!5jl��Ν��z��g�����d.�J��ftT];\)�w���A��9;{F\/x1��o*;d>���U6�pm(�h,t�%f�~�̆�:b|���1��?uL�ޞ��L�R2�f��}p)��?u�i�f���Ă����0i&ƧĽ��E]�V���0����x�О�gϙ�{L>#}���=�^	����������fiiA�1*�E|�799�޶}��k�9���y��8}����Dmvii������}�/|��Ǐ��w����=u���.�l�ۛw��Y�`�p�ްQ����lӑ�X�n��JQ�u���u x����׿�����ĉSy:�X.`n�`�#>H�U���EQXm:���nw[�[j���n�^=7:2zvÆ�OT��'���m����w���{x�}��G?��������(,S���\��Z�X�Ќ�a��i��_��kЧm�S0��QA���{����RQ�^�5K
�c��@��w,x,.�Ɖ�,��c�>k�χE BצFNz�π��,h�oh�����D��̴,闷������mF?0��
�F{!��,@�W��!��5�g�Ԕ�#�[��u;[�R�t�8n��&7�_l>���w��>"eϠ&<K���)�xN�Px?�K�ioa�k��O�ϭ����d�Yu52 �����lq�XJYA�J )mZ֤VD��,��V<Q�Jıg{<�k��8�T7��OW	R��R)��� �ژo\c�h5�9�{P�c!�Xc,1W����'��ߠP2���㰆.�����Q��8c��GZ�f���sc��Q����9���= �# �j�u��7򒶸7z� ����m���++�T`M@A-�l'�b�J�;k���ӧΚ��?+�Ȩ{lP��h�
ǳ�т�l�����;w����+� �+���m�
�f<��c"S���ϛ��O�a��fb�.F�0���\���������5��r��{ve,��oݴyyrrr��j-�Ԝ���>����M��,
��q<�B�$ͣG��E��8�?���gϞ���S�~���So���{GFF6LOO���Ɯ�{�Ȃ�0J��Q�H���RU��H���Q�������@ �<y�<�����_�����G�x!BT�@Ԣ��� #��%��!��:���~$ ���#�8�$M���.�i��sێc3�6}i����<x��3�������/��:��O�='O�x]��\dJ�����g6n��\AJ)HF�*+1ؑ��|��A�3���5�}�}�vI!��
`C� �-!O%���ԏbB��Ap�׆� ��SH������m��8s�Q�Dh��Z�(0��L�F�z�R�`��v�;֭�JYy�0#��]�C�1�y�,����=9�h�R�����kj�����$�����)��1z���̙S��K3p�3J
X���n|V��$��(�T���=�� �42���B��j܇���T����<%@E�����|����KŎ�o��'x���%�PA xI��%������Lq��@�r0B� ����x(֌��qGd2(��:�T<_�R�9�ؓ�5�Q��YI3#%���Ҽ\x��3��v�e�A%W�i`n@P1��2��fJ��H�{Vi�
�K��F�P$���-�/'O��XX�`����a]�� ���oٲIb���,B� �S�)�w2�2��� �/}�yΉ�1�XZ4��7	bI<5 p?��HL��A��K�7��ᕙ+N�]�2��z�^��^�q\��;�vs�Z��q\�	�s��D��sq4G\�U���{��yQ㴮�#j}qqv�O<��Fs�m�f�R��iff��عs�LXD	c�%j2�c`}�~��_�I	`a��`a�� ?r�����K�_��y��_���@�Rp�@��G�o�\ ȟ}�Y�� ��JS �2��Fژ$�gܕR�t~jj��w|i��oپ���}Ͼ�����v�~�}���O�<��4u������i��a��~�ύ>Q�����l�����u�i50�9���uQ����+$X���!H$0���J%-lZd8�F���;��q=���w,�� 9�:-V]l��F����K���A�#�	l6��p
X��T�OaG+�ϋ9(��#U�˨N������h����~��Fs\����F��}�5U���)8h�}�d`(�q�0	�B����)Ɓ�F�+Z�2��i���gܮ��q܇~e\C�{�%���nb����R�8�v��� �g'��\n�N�
�=޼+݁��vd��J*��9�~��F��(=] �W����D�LO����p�)���`' ݹcW�e��i|�-�z��E�F�^W��N�-i��ܙ��`�>ØqΠt1q��^���|T@;{��`x�����7g���A�I"s�̬��p�,�/�r%0.�4�I�/��JM��u�f�^3�S2�n*c��j`dn2�"1Ƭ�9G�,���v���fnpaA
<��Fe<�����~8z�:yF(�׍6����� T�_�و���J�y��q.�A�����}vb�\��    IDAT��l�\?[.�����`��~���� ��>���K�74�������:::�w˖- P�����9Hg �:,a4��]�����`�f֘�
F���O�@-�Ţյ�<LON���5-�!�@-�D��JY0FWrC)q� ��8Ί�y�J������k����������7�����������;��o>�/�}�ٷ�a��3EQ��m�mۼY�W�a�Sxp,T����!�]K���4'�P3B�-�4� �9��,wNf,��aH����E�E��4Zm]@��ׄB ���kc���X��' h7�1F��;��w>p��Q���`��>Sxr�0��~B��~�s��$P�^f��@��û�~�JSf��/�����MAJ@dIYR�x6�fO;.Ħ�m�V�HC�Ye;^WJ�f4,�B�� De����jM�8�^��g�,C���¡9F��-��x����Ɛ��ZO���)7xZ���uC��Y��hd?r��Z[��p�v�c?���4ۤVF>:���\��������*N�g��A�����zܱ}g^L�B��c^i��9~�YctE�2��f��4�.{�@^R�a��2P�:P崾q<�,ޥ�ey.{�Q1���$�̭��j^�WP�:uR�c��;�1�Ɏ�l���8t����7��YA���C�K��P�0�]W�������"{hTປ�B�����3��l�1ű2��J�g�d�d�GZ�83vB�I���6c�K��>2�H�Z{���R�ΦA:[q*���ˍk���yڽ���O��Ξ�qiy�_9�����3[�A3��1�ywTi�]$b�-���6lKa[V�d��J�,G��U�0����#�����21�Y-�Җ�%T�b�:�"�0-
�V���Q��4Շ E�PР\��׫O<t��{v���m���7��M��w�1��C�8;{��F�u���o
�p,�j�R��8�͛7�����w��~��$��6Q����|��.@e@����J���C����hr��
w�� ��xvLtQ.�ZT���>�)3�=��%ү��&;#jq.��I�㞤ιs��\
�W��g1��g��V$,F��T'�� �k�����������A�ӌ�-�*d��e!8����U��@�)Kv���h����O�նF� �RU��x	�(ЮR�3�s,_�Y�z����d��YEF�g�p�;���?U��{ �
"Q���EA�ک �~~Qªvߓ��Ոq�"ǀ/��J��Q�L7���8�G��"-�c�gF�&�",fR��cz0&��IiUt>;��
��h^8��ğ]�M���a�@�%�%΅�RC�V-�7�5�V���~��ZP��&((`�Ȍ0 UY �Z@�p<>~g�:�R�"����n+��8�[�7p!�	��^O�?/���8x��];w�N}Z�_�?P6��Ϲss��y���\��z!���k��o�����S�5��Fv
�3�{��pO��޽�%@}$�/��=ͬE�5�e�}ݤT*5JA��J��r�\�Z{*��'=��c.\8{�E�^T@r�ɱ�l�����������{�T��u��A� ��x�]7IMbP!`�b #0Q;O-F���E��O�'[0��c��Lx��m��-4��AK�ha��	iz��PRg&� $�~̕�T�lG���8��n�����<��7�|�7�t��G��\���~p|q����bw�ӍFc'
�$IR�G��4N&gf64&�'��vc�Jc� �
���LE%h�5�|b��Ek�PJ+j`&>�óB�s���R�U+�W�-4E@q#�T�7�pXn6�^F�UD��u1��ac� �8T< _�^����3�Z�S�=�)Z26�>�2<_n�e�QxV�j̍Ż�UY�o��E��%���`���j#�=(��3���63������z�(� rW�=�/$=N3�F��p����R��SQ���Jvt<��P�?��:Z�� δC|f@�>��y�)�
V�d��� Ö:�k��,b�3�)�Hm0�qR�t<?�E�'�B�������䬍}�u
4� t,�}���2PW�L3�ۄ��gA�|~�W�n���,Ū��� �͸�VV�
W�-�ͱ6�l�wq��>�r�O&���me{�/�����������xN��p*"T��6�A�y  ��F�n�Q���;m�[����`sn�ܲy������/�ܦP���Q�׭����#�)יrz�k^mn���5�v8�N�!;����J���8x�9t�P�5�WU��:����/����wFGG#�ʢ�g\��j���4�ͧ/'j�E�c���к�����8�^E�4-b�(T�Q�������μ�x����8F�h��t2��L��9���������.t�W�s��"�IV��T�W�ۍ"eBw'��iE`  �?h#�65I�%+н���ى��'o�����z�뾸��c�}�k�,J����я~������FC��ո���0}~��᥅��5�+oX\\�7;;�	��������2G.tY�=����G��F8sq��IaB�3����({Z����V��l�,ew�F`��*PiE7(h���zX��	��%a �#������M�r��Z�C�Sk��u�=��=���Ĳp�\2W�Mpl ��&���X)�J%TüŵT ꪣ-��Q���������Lp��s>+�?�B�#�<�Mexo|fL�*�F�*�rM��u�{�-��ֵ*	
�4�B����,����Xext�Ri�cb��'CE�ö�U�r�qj|J���d����6R�	*4�`F�A���Q� �K6)j#*}�� =p�Thr-A��5�n��݈JG?"@��ET�>���e�2I��qa>�R�9����g��H��f��.CQ� s���x�ڈ�3��lǸO��I:+.r�p͉�gd�F{m���B�J#��9��^��pa;��0�}���:�P�M͉�Ϛ��=���ϯ=z�y�k_k�'�2|�ثl�}\��$�F
��8� l�TdG�@ow1_"���0���22ͱ��c��~�I��|�С3���!^@��'�ͥ��ϟ��V��� &i��E��XT��Q�%��l+�`fY2��� �	Nji	U�4P��)Lzl�ؒ򙤘%�[�tG�p̣���|�$Ǚ(�IJ�plq���S��2����0*4�ڧ���*,R��555u���_���_��{_���~�[n��� Ga�M���:��+�n�_>{�[{��ʩ3g��ذ�F� �F:�V:��
I	N��l	&.�������dV�,hl���S9�`�(�N
}#��
j��N����td�k���b� TX�,d��x�2�!��M����`!�p-�>kZ�,����t�u0:b�K,9�]�2��]��#90dm�E���'�P�M�OH���:� �`	���K�j�0�*Y
�|F
!Z��;�5�j\C,�D��&��2&�Cqõl@�{i=r������c>J;3&�P���f6l C{�A_�y1ol�K�'���F�	�/�
��4�-��#�+@��YP�I��˷X�@�W�'R�%������[vd�(���bna\U8�
Ҩ� � �xW]�WVE\�+���L��(��s}�e7�fS�1 >���������.�ϙV�m�����I�	�ؠ���ظ�Q��{���������3��t��L�|��;�k���"������ʳ3��Cרȷ�o&�����3�[���dGQi%��l�d�6U�%�1+=ej�P�%�=Tv��Nv�kZK0�n�J���\���]1i�7�ׯ�����e׸�s�ȑ�.���������?w���¯t�ݟJ�x��]J1��ж T a�F��(%?�j��dd�I��*U���F�N_&��ٳ����	�a�F��R�H:3�W#�&�qR�&�K	�Fd��k��gR��&���a�*C����ƓP���Az���� ��s{��}��_�����?��?��?y�������h���_<�3������O�܃��hI^-ry�m%@%�����(3X��4v�y�{��#��ʰ# ��=j�S��0� bZLD&h�"���<
�q(D�?��Ƽ�jН��QX�y��7�鴛�P�yfX�ض�B� �~d��2�>�n�}d%�zբ)k�$&,D���x�n_3Ȑ�-��S�;�YI������ҋ�Z�g2/<��ж�	��X��#x�*��В乶�@e�U���٦��46?G��ML�styQ 1��` �B9C�k�m!����8_�-6nn��| 9��e������c�B��1� <\�o�����������]�y�����{��5�U�A�(�"%�	=(E�Ev�0��$mF�p�m�v���6� �_����u�[��qG��x�HY�$R"Eq,V��Po��9�����s�=�zY�*���
��{ϸ���[㷰ƍt����	�5���V"�׀kC (�J�������*X�x��G��z���%|�ڔX���(�!9XE�;]/@d����d�_�6�v�s;����5��ge�^�y#,6�	�2o}��w��+blQ�&��jBN$߁�I��5I�.`���9;ʪK��Ξ9�[TL��UAh*������O��٠%-,t��/�uxN=����/x��h�l�q�c��S��&1c�Hy>{=�3��9�'��H(�]�.������W�����~� ��+�,˂O�����l�7�;;?=��9!Q��D!Z� �2�j��D)�H�KX2&Y�y�9���uq�_]�����=��� %�����W</�1������&��fC/ͺ�X����3<��h����z@Ek�}�ʢu��v�p�  �14�������yϻ��~�)���u�����]���'W׮���K����
��w̠Q��X�}X���K<����4�CY)����4ިnM���r�6� @s1. ߩE�R	��t/0V[�4���"�6��Y�s��Xu6њ�B%�M������5��X�d��б]�T01�P�dB���r9ម������,ڽ��}��u�"��
,��ٳ�Ş����ÂK�c��BF����ؠM��4�8'�{<��0p��>��	��1����O@�	;<�bL���^�Q�ޚ�=u�⼐;s1�\q����T��KYk���~�2��C��E�be�,���0�z��e�k��B-R�K[^�1#b�K(������3R�c�7\�l�"�_M�յGA,�^�Tn�z#^%q�6����h� دo�dKk�����IE��U�z`��c?�A`}���2��f�k.��YB�TN��O0��3�	���x	Ѥ�(s���o|�c��s�{��6ô�\�{�n� �կ~���~D��������1�s34��%�e��5�;N{G�����Q���V�L���P��+���4���5�]YY����~i�=���ϟ��Z���gO>w��?���w���f�B��4'�����&�]��t��5��!������}�ya��4���A�Y���
)�����,*Mъ}?�+�g:C�?@}�Ⱦ&-����2%C�X�ւb/L�����q9\�qsun[9���z��?��������K�d�is�œ;;?��z�C�^��յ�K`4��~�O��`�V6�qI�ứ]O��	t��$�+����S=)�L[�E�r�+喃�q�S�lt��.�0e���N*��5��;th�3�Cp��{&*����"�/,�����l���+G�o��x(��FZrF7��ye=�ľx�<��yXS�@)���O@�"�}񎶬7'$�GC���1j[�T6�g�9(�lb��.���m�q:vt�s����ϥ|�\���d�j�s�N������m��DL��4�AM�]������ljX�Z�����[�	@���Q�8�Q�j)kxmx_�C�h����{��K9,���DN��k2�Q-��%�,T 5�#�T�,�Ʀ3a�b�dM<����@�TA\�q�'Ҽb@��>x�X3�#2"�����p\�Y`�^�Tz�@B��\!O�'��T�qn*e8�n�z׻�2>�;X�,MĽ?��ޟ�ɟ�=���ŋ����M���Ƶׄ�v(��g&u��,���?'����������nX��H���T�:]t���c@�ǹ�\#Q�s0i�����z����������h��l��G�}���buu�_������}���H�-W{�� ���<@ ����b�1��h4&`!�q�u� .�lF;g�9�pl�& I�Q�{Y
�H�^:4MM��*��
� u��}		��\��Ե��ƒ��N����#F���.�P4@T�߱h���=��������~��x衇��ӳ,WW�]���^�����������1HE4fw�&���$!��m(^��N%(4�th�\3��1E���9	��{��>\�Ţ���m�+��s��:R�X����LdTYo����.���ݸke���6�H��mm[L��8��y�Ȳ�ߤ��Z1�vh��J]�a a�v>��F�m� _�� ��G�uP��"!^��f�2dBE�~/+c\t��~: g��z`ƙ	me��-5�o��V�x|۫�g�����-@<�p���r3Y�L�����7�h�,��$�*���a����BƋ	�БeOi�X�a�N%Q��Zf������:�1$��$	����a�@��8�)	�u4�ߡ?�����0*�rOw���/��[��M�� �m����d��Uq�s���2�cN�k��O�
�'ʀ�|�,�
�_� j�d<���2�4Qé_�r�z{�o :\Q����n|��ȟ����"
=A0���^���7�| ���To^�[^^��E\�5?H���%*¸w	�l_@Fȼ�2H�]%��5N]�r,(�����8���JX����_	Rn�zY�n2��x�_�����F�A��m�3)ƾ���,� �[�fx�FA��(I,����K)QQk�B�xO�tu�-�t%��+b�Р��/�4�������AjmY���I�[�;&1�X8���ҵ����?x��>�3?��ߧ| �O?����Z���~�_�F�waxz}}�x�G�p��t4KW�!�I����ZV\�Be��w(M����n[쐿 �a^�S�RᲷ����]�9}��ȪA��v9��D�	�)A�� mp�-L����_��˱������E94u�L|����.�l$�I�I��b������J؆�9�iYYZ�E��	[9�k�z.(c*`x���s���jlO�/{�QQb���r� �\Y��R�*�=1U؊�a�7 �k|��3�^��-A� \ *�P���O,8��^ܠ�?�*H���g��T�B�md�*`�B��P������a<�w���	�y�IC4�}��xL��b��xM�Z.�%�/o��)��wx�Z�9�Nr67e��k�a��$Q��˂w��Ùv[�ǚx���s�cs}/�z� 7}/�!/R-�z�Q4ŋ����],mZ��\Ƕx�|x#���/Hn ��R2ԇ3���c*#���Jӗ��%�8y�;w�|>���+p�{�/y��Rw�p�&#��=�)R=��!�'P���	���WB1lA �(�;�Ro���V��W���vu���e��?��Ï?��C��W?���O�#^�1�̓�H��A��#{��ӏ[��/�8�a0�C����Ky?^���˘[-
ֵ#j�nM߃{= Q��	�nu z�����������تq�*��-.N�Bb,
I��IB+0"��n�J�ȉc�;'N��;���������cǎ]o������V���}���9�#����< :&\qEV;4i�QI�mh�`E2�½.5R�    IDATn_ˑ�{a���$,HR$��
���+U�؀.�CdW :��HG�6���f!�3��<�45^�+}�j�ۯI�.���>?�"��
J>�j>��ҿZ��jz0���'��r��a�G���� d��w*(l0ì߅9M����-�������h?S[�x[њ�7�m?w^�����>�rP���Y}*��j�b����%�/��=�兌t�gzYh�bp������g�L~-j���4�}3�At#u����X$�ߺ�	�Y�,a����J����g(�Ϟ���򔘹i ��$��+kZI�Z�#1;;g,��(7?���y���ɓ�+��xͬB�Q�h���%��r�S�n��0� ǅ�+��j���f�����^1d��^�V]Y� k(k�J���F78' D1d������I��u���.J���%���������r�g�]�uW*]zv�I�d�n�'�7�C6i0���޺���������yblA�����O~�w<��ӿ��u>���Ղ��1K2 Bc����g��t5	�����<\I�W#<ؖ���X�<q��"��6$Ɖ]U	1t-�Q@�;@�q��Sw�,���^h�؉;�d�rq�-X�P8p��WA�R���,%a>������}��?����j���8�;;?s���4��<<������%Q��b�� ݱȺ��^h�C�r����([yO��H�����"A�-Y�$l�ox��X؋>m�df�ET�]�n\��s�eO�������B��{�!����	������*>8�(�P��R�p�Q��'�1��p,gõsQ�OB4E]-�Z6H�Wk_]x���ܰ�)�@0�<��:v>���t���2c�Vd�*�*ع@a�3ƣ�oMY1�ǂ1h93�'J�`�'E�����:B&zL]S
��+h��ɳ4�t����*����@�F�e5,�*��|�43�-Y�}^.�i9��K�� K�y�9Sb��Q<�!�~�� ��"����!7����_��$�.q^�I�4q~xV�r�>�3 ��c0���5��X�9�ַ����"� �92������k�y.>���$��}�I�3 D@����x I0��v��E�{ ��3?;'ָT4����>L���1U��
*�m�߰�e������ǎ���k�Xi�~�'?��|�3�ϟI��_������=�=�ؿ�<��~�[ec`�rǃ�KP
� t�M8�a�@;�u�6���0fk���1��(�
�2�J�ߒֿZ��\Μ��R�.w-cS0��`O�q�D@���ą`N�M�;��Oo�Z�������O?���w�Z�����ÕJ4����XP!G|���ف)c�LV���T� .1r����E�x$�1��}Z^���W�nE{��{-<ZqHʳ-:.�̎�-s�yIЩ�ٮv�;�>Cwj)_x�]�?��2e@��6��۸�y�|� Z�� ��BXQO�4٭�L��).xC���8.���.-xZZ�˒�2|�En\�,�G18�&Yݼ/[	���o�����<c�d=;[�8����C�`%Kڠ���M�|&ַɤ��H�� �S�I5D>Hj��ϕ<�9�j��"���P���h+�r�����,��� �-�׵� )9AV�zIP9�6�/�=�r�ϊ�o���ٚ1ϗDGJP�k����x�1�ֵ������#�iT��V�<��h��|��~�_4��9�l�+��zP��c��6�k>�$�QY��"�u�`��5H³szH�>�6�u��/��`�w����HȄ�F�;\d���s����ύzK�C�\*���k�砞K%���]�<ةtuS«����S&=&�b|BI�u4��j�����t�������F�,@�����w�m��ow:�{;��6.��J���W����
�^8�'�`�C���jؠ��ۋ��P�m��0F+�p=�腇f8LJ��T�S��b�põ��"����DLնU��5f�j׼&N\i�gJ,�?&�S�{�z�;�<�@�'~�'jˋ����z��X˘�"���ua�,I���jR�Ը`�^'���sl�z7z��!�kT�^"�F�3��	��pQGͅ�����K�ŵ���m�3G姼_.SI~�P	`�Aْ�y�$�p{Ѧ��
["��El�r�ϙ�jV�8���B�����3�=~���!^_Y!�g^��.���-:�%�n�iLH:�ym �L���	*c�lq���؞�#0HY�"���,b��: ��N�a�눝ͮ�Ͻ(Y�����-u�J����� Kn~�k8b��ڴτ��~�r�s��o��cB������'�E��O<C�����ˌiU셁UQ�o���P������{"i`g�1�������k[,	��G$�wX���^ d4>Q\��\;H0@������ޓO>���q�nw�?����g�j���3��Y谸�����P�g��ÆL�#*1xΒ���J��B��\ɤ'�򤪋aV��7�p��X�J����u�i�U+�7VV���3g��ȑ#�V?���e��?|������>�0��A��I��$�M(V�J� �w����p@8 ����F��(߄�>V�6G�9�b,�z�xx�XI@�*V��qF�F?�>l*��n�v���2�w�C@-]�>���K�p����}�{�${��>1�fS��5��y�H���3���k��mp��X�ia��Za<\ ��Iu�(j�w됉W*G����:���|N��=��m���u�㔠���"��BK�Ϛ�`�1!��|�S �l�I�@�� @��TX��B�=c��uԋ�%6���q5���Vh)Kޗ}T&���%�m�R�j��m@/+r�b}�� 'Z����-|��0��Y���2F���ҀmFH��ަ �8/�Qp=,Wb��XCV�9�F٨�a�<GS��e�j���Ow��d������q��Kl/+yE�������J�h� JYi��F��#�T�=�k  @LIX��/��.f�r�5 (^ ��~��R��DA ;ʻ�Y2ަ"π^)ܛ���@��p��D��?hqqL�S��B�d6ḏ+���9�&)	�ڊ�.�k��N���L���E¸�����Ѱ�����t�E.
��,��~��ju���_��Aq���7�U�����k���?~�߼��8�T͞}/�?������>�/_���{���Aw���Ւ$��,�P3�7�Q��Y���������٢z���M�=K����J%�\�D�T�B&�|&��ޒD�I��eC?e�*z�&A���$I*���O��YEa� ]<���?�� ��Ie2y	n�LNN��������y�}
|�(�Q$�dq�J�z��՟���?��?�SS��v�$�/g��C�"P;�I �2N^���M�����!ծ��Iқq�K^��L��CaB����.���N� �ʦ�Em�:+?+��m�.z�v����B:�i���� ƑAUZ�lk�v)���|3vό���A�4K�xt���}ـ^V(8&Oa�Ͼ����'�S���z�(%�wҺ�|ʞ7ۍo+�6��w�r�&����\��:��9�Q�k��e���E�ϑz��G����2����^? b�2��"�P�0���)� �(cu&�X�/I���z�@똣���RP�/<����Z�(�Ux��{ *��q������I����zv�-�	f_���`}��?~�|�b�r�PCP���z��#���E��a��8qB���[[]ג>4��Z�֌&�b��~��b/�����q*|0|d���r�GYK-/���)M8,x�)���.!��K�� |I�3Լ8/�Rq�L֋�p7I�G������O�\��~���?��/|��_?z���ӛ�Ƕ��������aeYZE�YFQ�e�4M�$IcL� R,4�H�EaVA��Ȣ(�5�h�U�y�L�e��D�+��$i�g��z���0!�R�"�Q?��NV�3�J��gY��IR��I���=܉�0�Ra▝(���O�,�pi�j�y���V��p=P��(H�4�}��0�� 
����j��?���7����Ο?�������w����<p:``Ra�u�Ԙ:���(��Z.�� ����=*�����1@��`d��M����4TpN0�鹋�)�.�nʪ��qlK��E�ی[�M-�cn�[a]�u�"��W �lf%Z�GŜ`���ۛ��̜
�GK�1ƛ[�P�ϵ��ϓ/���Z���_��m��P+���$e����	L��F��+쿂������-Y�t[6�wZp��}�E��z�4���(���?��ku)]�E8D�.�
���D�%�5�\���bN��s�`��2c{[�~�JiG�N�y~����X��[K���@B&��\��a_q��=
�>�|a�aQ�<1��j�����a���k�d��o�]����y�˅L!gX��~�s��~Pp@x��iΜ��Y�8;���P�(giI�����V%��DB2��(f]��/�ou���3x�T I�VH\�g�3����6L��o3͖������߫7����o��o�� J�W��t��߹�x��^u8�� 0��n�W�����
�(�|3 �@"nF�X�iE��3|wwWf�a��,��Y�2lk>�Y<�d^5��|����ԥyi�Z�������^�ղn�`N��|�l6qr��fS����T���[����>��~����#G�����؀U�}�?�}}��?���6���~��h���@���$@Y���`�B�Ny��9���+ȣ��=��^_�Sc�-tn��LS�}��5��uZ�t����͌�tx���s���d��"_jc\������KeiB?�X�T$v�� B	�y|:>�1�;���rв�z�9�Y�i��=��m�,i[�6h�oZ>���d C�+`��1����в;޶��}���K< TVs � �(��@�����P�-I����)ƣ�P�Yh�ki���6l<�� д
���$�r�
�6�������R�*�k��=vs��!��=���y�N�e�P�=�(v��̬�Ÿ/+��
%���T�0<�V!N-��i���M�0�Di8���/������'r9��3gNKY�;c*��j�̨����u��E1�4���2D�g���h	ȓ��|�"+�@��<"��zZ����,�^���<Q/	��%c���nZU����2=�nG�4�-M��*q��G���ݡCG�yo��b�uhҗ��J����w~�/��_����]�GW�f�%�@�⌄�`��$�bp��/�-
L.�j9k�Y�6��y�肀M@���l�`h��r<I�ݤ���8y��E<�~��8�����"6��a�f��H?�꘭$:�W�����|�`�d�u٥=	�'��YV���$@�~x~7zp���bb�t'����0��A���� ~�����뷷�++�u`�����:f�@�Yd;�ʟ��1X�g� �;K��u�2¡C�iuy ����5FsLZ�xШ*�(��l�IdLֲQ�H�Z��S岲 ]K��h�nw��8���`��|(G++�zk�Yv�N���CAK�D9���^�֐��]�!�y6���`^S.����8�ϋ���cn�������eX�؟���2�3mW�#9( �ĥ�۳�����v���b%�:r�Wh��%	勑�r���6V�Z
�a!r2�%l��EmVD��eF�2M�����ڧgg�~oi���<���/�L��v�l��t!��}�|����G��k3��gΜ>�|dQ%)���GR��.E��D����ԋM?v����Ž�{q��ze�v������B8���cJ���lH�`�lPbɛlz( rSW�=�by=CTHӛ���V
��$�a.G+��c�`,�b�S����mQۣ/�����$����*d�p� :,3��ַ���YԼw{�|�ؼ�FY��ao����P���/���d��

�C���-(�%?Sqa5B�(��p\�#p�@�� ��ܪ�+���.�|��*�v�fƸ%��zf���c^�A�#%)�t<G�.Kӻ���B-�L�|t�KS�i�]W=i؟.n\X�t.�v���$�rNH1�U��s�Yh(�
��<źn5�!k��c�ZO��,�h�O�ns :���}�� ٱZ ��FL���0��Z+V��3c�gx��yO�~��9 �LHñ14Fn<4&	���J�v����� ��1�{��)H�81s���h.r1^;1U�.����E�������ѕw������=��,7~� �@����?��_��#�P����s+�������]2q�lN��6H�<U�W��33�ۢ��E4��d.����֨@|����M�gz���ogͫ�^cM�;;��3OPg\^�(�ä���̊���a��3@���x,�.V�X�U)��$^
�x�^��@10Yn�=�	�g�Y�e���,���H,���Ur���$�����"��m&H�ϣ �I�T"w����xv��V lK|�2A ��C�~�2'P�_�*�XK!șJ#��TnC0����k�q,6ea%hz�0c�`��{�Ai�6MR����i���m��QJ�K��eqJ%׻֖w�JG���A�>[��B�y������	��&	xA�0S@�PE���+�� ��Dl{�ЂTA�0�8̻@�Ώ�+���s���#�/ֶ�o�/��Gs���K�=��3yS*"����ݖicL�ZÐ&�6G�֠�����*c�(�H�F�T�_���Y�4<8�l פ8�F`���'@{0���|�٨���[�z�/�G���A��F�;@%�{������G��C���ި�v��m3�N��GQT����7��'#y�J�AIjh��;٦xX�u�(\�ܦ�LR
C_���:qS�ֹj����bB`�@�u�&�-�cr���k��� ����B�rG�|�t�\�U�(���x�\�D'����g�Ks`+��� �)�q7�mu�L�)����~�mY�6e--Q<��$���]���V��]�P�`��]�ܟ�6��p��P��nz�%?&��0�ؚ�UX�v���~c�:`�t<�/���g8~��3�|C	,U;��	�I���XX�Fc��(*Z��d����r+���̒<Z��1gh���s(D�(�T	��8q\!��,�C��@Uۨb��uwy�5#�5P��Qo��=�n�����פ|�mP�Ԇ�t��g�s�!*�k�7��ZC�h�4�d�+�+�Bkd}4��4�y�-⹰m%�\	��e��2%�p�K�sxHL�<�3�ל�l~��W��@KE	�PO$�
�h�U�W��>ݞ��㳧�~������ RdW�T��`����������n��Z�r��ҡ�QX9��|h����L���0l4��j���M�w�*(��;I���}�ք�w�gP���1lU�����K[�rȉ���Eڳ��0%[^	l�@�1R F�coG�fQ��}Y�^t{�s�b�CaY��%��Y�΅y`����!큹�W���Xm�s)�����.q�d�;eoz�r='�3�P�й�=Dm�@�eb���7��3	�����)�E���W�my��W~v�#�S(�8�|0�r,�
�~�ﱤW�UP�c��A,#^.�t	�:��p/OY��N�{Ǎ��8K��dI��*<�xIP�w$�!��4\�zi Z��A+�]mT��!Af�G���2��d3:�4A���5�*�����@l�ĵ"�"!�n�R�j����W:�'X�ҟ����!8tz�6j�@1Q�^�B+�\��z���iz�Qo~�ڨ�_�z���>��{���Ls��|    IDAT#�q��
 �f���O|���c���z[G76���q�Ҭ��E��v�y�٪-7��f�Q��4[�z��� 9^QUKK �p�
#]� ��1�,ъ,d܆�ԃ�M	2
w���q�&2$ak��_ۈFlb� vu���|��u����"	������ՅZרks2O8�s�K`�s(/wa^�k�6|��T��,��I��{�,;�B�?<b���m8h��[�6���[�|����P^�ˀ�fF���z&�2ȗ?kv���r��
�PJo��Mh�s#@�{?��� OZv7|���]�Z��X��9 ��(�:���[~ޘ��6��u��y��h�C�&��I�HWLw4������f�EzHt:�f;U�d��2׀�/V-�XQqIW�^G�e�+ �R�"�!�F�17���h$�1���Z����*M�X��+�3A�z�
B ���\/+�S�p����Ź��}�^m<��W/-���ҡG��.\�0���
���+�4v����������K;;�;��~�h�,giv2��j�d��:ڬ�ەZ����W*��j���� W$b`̰@ �"w�I$�"����}����� 1N��5���ݮ��i�����Ρ 0�`LF;���
����@�����"3^��I��6�e�C?�˯H�* ���"5-+�`�����Fi�Q���ܬ�z%�(ܴ��,�V���M�D�1��e�V�� 2vo%�{Ҿ �2�h\���d�����VtU��e�`���\Q���x�<�(t%!� Pb0,:���1c�����r&�Lz����
�)��1`��6�PX�_���sd˄=D(���-�{G���4lk�#a2kC^%c�}�ݒ�8�18'�!9���D !����܆�G8��ܒ�8��dZU�49>���C&b�	o�g�/J�%�t&��(�SA/sza�;*
x_�ZT�p�Y�u�(�����>�n��t������u�1��͖�M>�'?�ɸR�m\���X[�4�}}��?8��ߔ���q%>��b��n:<_k������j,��J)� �A&Z)4� ���D���.��*�
��.�W(;GU'��n ���xZn|�Ѝ�
�[��6�s�c�ٮv�q�G2�)�#�S3G�]*(���m��P l��$ӊ��ܦX���W�,Q�G���$��e��`���7��z�Y�f�ʓ�ϿC��e����I�1	�o�d��3��R��h���I���_��'t�A)Y���A�Wh�#��g#Ǽ�G��T"p*L,��<�������!�rMX���(��p!C��^�]_����o�E[k6��,�פ���4� �v�3�k�������S˜�g���N��d+�Ύ̉b�Խ� %�gj�W�p���:�@��W�䉙�T�BGJ+�$�)��[yM�F�q5I����.,�}�ĉ�O�����52��d�p1��-�i���|t��ͧ����nn��l����93��N��[�Z;�h��f[����X�4b�.I[�(�LY�r��\պ]X�SwN�]&���ٞU]�⾷��#y��p�\g =gf2,W�f�.�|���k�M��iي�����l�v�>zt�����5vE�d!�^��Z����_�&W#��X�p��BC��cݲ��n��b/Ť��߸+_�+=M4�ʲ��!�O1(�|��q���@L��,�F
A�~��{?@��� �Y���<{\�^�\�A���J�	f�"6"�kF^��a�"��e��斗ڷ������E� �WPh��6�Z:�!�cL!AN��)�#.N@�����Ro�ݐh;hG3}�eA%1�/�k"��`�}5@�$L��nGNX)�g��cQ$in<���,��JeX�V�*��sQ}af����+'��.����?<ޜ�&���o�@_�����͋/6WW//mml���{=/8W	��s�s+��fk~~�63Ӯ�~S�ׁ֊�E�X��b���	���h��e���M���[�X�#6xI���Z�k\��`7��E��q�:�dҘ������3ꊥ Ox��&/J9K�@AV�7�58���|O�y��u��MM�F�����r��r��)�Z�\���@hZ��E (��D7�@�� z.��;�PB���4%{����b��)�<�r&��|y< 9fn�?C+��l�gV&&���h*�v���D�%���<c��SB-Kf_��2�i�e��vҀI��X&�q{\�����k�ԅN9���>�iS��X�����VDN��δ�/���8�������qP��n�/S.d;��ɔ�Ub�P%�v��s+x�U�+��dNX�p*�U*�-����Z���엛�Ɵ.Z~��酋7+�� |q�~��^c����A�ʕ�Z�z���k����ݡ�D��8����斖��p�gI��Pn�?/�su�聯���I�k��t��uNvfr�tF,qvk3mi}�M6=�M)�k5_����V0�m8�ӷ;��	t�2�Za*�2��G!_��������Y�V6��+d�Z�'ޕ](G�YX�;�A@��Sm?@��}��s �N�/�����C�"}@����>�1~�,�u���3��g[��~?@�(:��X2I��rKm�'Ş�=�C�Z�,�PCU� d*�[�1�����2��r�%�����T��0�>	�2O�j]#��!F?�\�x+d�w�{��/�����{(%f�����ȱ�u�^�?_��4�9�}�z���7����c��fea��?������ra��˕�k`���OT��Tf�|��/^=���J%~k��j4ZǗ�YZi>�І�	�(4�z]�#��CMɼ�h��a`G���(��Z��7��9�x�8c�^s-�LhZ�
�E� ;,��K^�W��Բ�g$�ـ��"�F�����EK�I��e@W���-�e���U�C�D�W��#���P,��~e}�<^�=_� \��N� �mc'�Ѣ�qM,�)�_a!���ur�A�1�b��|-7�`|l���ƀ^>~���Vx,G����+�]�8&�ʹT^��v<��U����ˊ�j�<���:��j/�iNb��C����d(ǘ;��5J8 ]�)[�w�^P�|!�1I�bL'�[ �s��^&ס���`���{C��lu�̱��^�J��A���x�+����F�������q�����?��[x����~�����J���+��kh_d�oll4�{��������</;�љ��Ӌ��/-n��z��I�w f�YP,ĒLf���إ��R_,w�#>���e�0���Z�j}�X�V�.�nx��X�c4�p雌x�1c���c;R>��^�X�B� E ִ���nw�u�����X��7�����2�ɢ�f�<c t ��A�~��ʅ�ם/�FA)U�ko��I�!ߕ��͜�ܠ7����;��aqx���&Z��8�jS=>�k�/)�����J�G�(n���*���}��)��5��1����B�{;���������Kꪳ$�v����R�W��R�|�Q��%�jՅ/�C�3�
�=VT�%�.Fxh��x }�ı.�Z���V�c!�b��
�~*̝Z٣dp�z���eٵ���Zs�ߨW�/,[y���cW��?��^19�+������û}oE	dم��~ov��|����#��[ww;�{/.�[Z:rzeey�՚mT�Q��P��[�����ժ�v$L��c�\d�`h�t��d'- ��
��lo����p�gZ.#�w,�X�A\��V��z{��}��݄�c砫��@���*W��2����e��hk[Y�0W�Y�'tis�$H�b[��/os��Kg������	��Y��R�o[��we0���loe��|tO���QP>����75�v��j&$E��X�1 ��Up�c�e�ϐ.t�:�-q�z������u�M���a��2�sgpMʫ�xQ���^J���5�u+��Ԇw���CY(ra,�Ws��ɋ�^(:�Q1#ꑹSN����X��qQj�!{ᾱ(w�0��x�F�O6��?�T�??y��g�m�}���)�0�у~w�~��� ��f����ٵ�+wlwv�F���ٙ���F�N�̷��f�Q�������B'�]��6�-]QȦࢅ$9}O�#��^1��:�S��!��cvE�բN��,LX0`��c� |�h�=�u�y��Xb��=_��u�CY�]pp; ��_��ahI� �ظ��[��o{�Qn�@���^p�~'���ͳ��ؐ���^�X��D�t�med�k���]�7QJ+Xy;�}�����d�\���,���IǶ��V�뗴,�]��!�7�Lm�̘)�:���ȸ���-]�*'(�L�'��a\����?T�����1��Jɀ7�9]��2�09�L2���z����%ϐ\򚴇�1����ӕ۾�<�!3��ކP��ON�mx!�"��� i�/]�V�m�k��^�=1�\mԾ|Ǳ۾�=\y衇ƻ#��9t3wq�~3��?V�e���+�Һ��>���9���N�^v�V��l4k���q/�ת�kՙ�L�h��%-o��/�4yx��*�5/ݛB�R+Ք�0p{Qȹ�M��Lh�l,x�e��t!�ߋ�x�TW��i�3 F;Z��2	cI��<8���8q���*ZPvnm�*&�0�Z��z�h��x[S{N�~�Ct?˚������e�w˥_t^�o�
/�o9��cM��>擦w��{�gm���{�W�������w:��V6]�:�4v,����o��ǟ��0�4�f1��/T�pZ�� o�( V[e����{�9�/�:ʿ�Qۂ�
6@b��¸�u)��S>�ǖ׸L=���Z1r}f�E.����E����Z�MnR��� ��0|>K��KK�=z�g��<o�f���L�p�~3��:;���ۿݼ8\ol]�׮_;��uO��w>�3a�r�^�nʹgۭ6\�h�c����m�O4]I�+4�<���%]t��1ղ��[� rC!���O+�qd��*X�&nn���=��NK\����27z~,��:W��S	�� �]��V	����ql@��p�J�ݦ��=<�>����9v~��ǳ��c�x��^�#�R }?��F�2�A�-mٌ�I�vś3�n+Wc20���6�yX��ha�ʶ�m߰<�k�BU�Gn%���b�h(K�$Л� ��`�3�5tL�t�u:����#�}*�e��5��ʍaJ��=2\*���RZ��~d݀��4����
־o(��X����
��~���� ��A�D����xhi���g�~��3���y�Ҷt�������F��[�վ|�rks���v��{G���J�r�Ѩ����sQ5�(h�aܠ6-`c�ʹ$�;R��F��݄:!u�d�ʁZ���0Et�\'�K�y��g��F$0aY�<�� tp�s������M�^nɘ��*��E~a_�q��@a��%���ڵ�{b����a(ߩ�����qp�=&Y�/w�g��3Ϲ��TA�/��+�5��$k����<�w�}��ǖe4)"a��F����`
,+3b1�E���� 8S�U�.s�:�/�1�Ͻ���<pZ��>�`/�~.�ѤUr_�0���q���'x�j���w;���5����r��1s��aN�*�d��г�m�}�Γ� �&�-�N7�Q��9W�rh�1�����T��j���`�����G��s�Z�ۋ�����n{��<{�7?�y���o4��4���%�Y�O5��;�������- �J-n�+ީjT�-����vj<Z2��0��J(��H�2 ��f���8����M<���
ds�ϙ�� ��Qߴy��Ak��d�����NyɚW���{�����౶���x������m+	ߡ\O�l�3�y�E�Q��� �֙�P�UO�s���%z�U��7��p5�9|����Ff2]�ǳ��sh<X��m��$�ݾ?zi��el[��L&;G�$O�ea���h��	\�>��C��*�t��xB}��70��\A5	>�"���}����3��/�:�~�c2�].!-�Z�aNc�aϻt�w��U�-J�̑KS���_�+U&8Q�ͅ����n�i�ُ�n�+��(s�?X�(_� 8>C>��x����5/��kߝ��������Gannn�6�4%~�;@�aJ�ut����߭]��D��g.�lm�.gY��y�[<ϻ3�;j�x��h�4k�F\�5k�X����RzI���DE��܆�X\�|$����Y"�ķ"i� ���2$��"�k����{^gg7��e�,
�T��'�<���R�3N�a������@o��X�\\�x�]�@��W�=�d�lơ�k�3�( m������r+Ԫ���^��W��p��p=�ܕ�N��r����$o��-8ʯ}��ÐYaQ
K�} '�/[q�PG���Po�}�*@�����3��h�,r)�;�h�DA�7�$�I�cS�V�^��^*/}I.�IL�|�EQ<�&o�Ϋ=�j�c��;(jP6���w�����+�����[uAI�I��[9���@i�*�����k�%R��R5|�����3&:���Hϫ�d�(������8���[��]����ٹϟ���o/-�6??��я���͵�� ��H��;QH���G?���67w緶6�vw�ǲlx�V����i�l4�G�8nG~�h��V�Å�V�����M]<LyZ��o�GH��;Z�ZV�mPe�2��p��2�u����������⊇�b�c��4�A�8C�c+ z��GA�Y�e��W�,pj��1��o��P(���}�M� �Bs��"�Q�� ��T*`q��g�]�Cˮv�>�I��J��I?��n����2䢩ؘ���I��I�Jr*'9�.��8j��1Z��f��3��s����X�%Cb	��Q*��
�VI6�!�s��x��qp=�Z���jx�^�[]]���|��mt�J�IdW��ۢ�<rn�Ĩ��:(
��\g����=��kՍ�=�u8%�׷v���T���gk��7Ϝ��so{�[^8{����zhg� {m~� ����^sW�/�Ň��>�kw:���`���=���\�_���j�j6[G��J��hT��f�Z�����=O �ώ�ApA��u!*�ɢb��VԍKb�����H@�E�%my	��}Q:����arGI����v�py|�Ʈa�<�����Nxҹ�$��y�ӞP�^��m������Am�J6�l���X �� Y��<e��v�[@��\�>Z �x�W\��#GT�`���+�b[�z�枘���
�E��X�VZ�?��)�R�E�,+8vH���i7C-�,�?�Ĥ�C��3,���an��l}}�K�b�z�Z�@��Z�N%M�7]ߌ���nh<=��&�qn#iP�ctmHFY6�vF��v�_���/5��o�<y�sǎ�o��#���A��������{_���Z�ۼr�߸����;�c�ۻwfAz��h�l�['+�x1g�JT�׫�f�]s���M]�X׆���.�E�U�;��cb�SI�Ӥ�:�e��k�DX��G�kv���#�βf�� L``�n�k��E?KPW����嘥_X��zcVWxLڳ���䔕���� �L ͸�˖�$@�]�6���E�|rlӃ� v#@7H��Vl*BkK�t^;����Ȕ������.�ܥn(k54�WQ%���M�ϟ�Jb,Wv;++��O���ov3"�4�a*|���HS���V�V�ArkKB<i	�a�T�t���:�M���N\]����@H@�و�"� ~29�4M��$Y���F��d��ս������ۮ��[����cm� � 	�ߧ.�.�n��Y[k_ڸ����q|�KN�Yr{�k�[�5��~�̈́a�
�*��aX�UbI������]��5���~��J�r�<F>�v%ƧpS>����W���J��ɜ�� �[����:e���.�"��:\�!���&9#�E�ʼE��  �IDATG۲C(�p��O�3֔�Vg�W��Aٲ/�{|iA�T�Nz��X���d������* ~o)�����X1t�"yO�3g�+�
v��##������ʋոD�v4^��g`�m���x�9$�^(Z�6��K�$����y��f50-�يIEY>�$g�C�ְÄ�P�Z����ښ���&ɂbM68(���g�]���k�������Z���71s(� �1�rYT	v���x^z}4J�z��t����'�t��W�g��C]��Lo���7ȃ~-�&-����hl^�6��s�h��_��D�gKY��7j+��ss~��Uk�F�֬Vkq=���(�)b~\ D�����_���q(A#��D6FMi��$=����sڣ[�9-��b)�K ]- .���%�\���hN$c���e�p����K���Ԣ }m��ֳ��Z��Fcg�����Yq9�G��pe۠T0� ���KYt�\�7 ��b袀��~����I����裼�V\�R�?Ȋ^��%u<'A��!�T
'�G�D�=P���`^S�.�%;-v(�c��,�R4�o�HB������317c蔯4q���!�����ް�A6:g��$I���j\�_���^^8<�7ˋG�v����'O�]��_��Jc�[a�u�~+<wJ�R����ָt�ٝ��R\�g�66�������Jx�Z�-�jq;���0j�J�F�<OJBҬ�1cq"{��NW�* �q���nO�LK�t,Ht�+p����<�IKƪ7�"�rtA6��%9<�	J`�Jǵ
�[�X\ԥ���Q�;\0�����5y�]ePpd�� �q9۠g�Ͳ�s����7S�|�V����.;�'n�K$�]�J�1�4eRl�J��m�I�2���ч�JV����ʐX��/%Zp���  ��2>���
�"^��:�EO*�����o6�"���q�c�Ű�M�\&��0���Q��LF)�@�����;A�U�Ջ�z�ɹ�ٿ��_���ʉ�7������qAܞW�����(��wvv�[[[��`��������s$��3/=��	�OVj��Jx3aXi�qT�c�˅u��p���`4I�<Y���2��Ŏ�q�
� �ɜ����~����,7��k8��LY�)O@���@�|�?��~쭪Jkkc��.j�hi}lm�Fb�5b�FQ��Ub���WQ�1j����~�������﹞��9���~_�yp�[���S�\�k-7���9F�!�aW#~|	�6�g�H��z�	��X��g���h4�7�t��\�Y���A��Ga3��n����$[d��Q����A�	I��w^
F/9�7�����1�e���g�;;�V�C�Ė�&*��f���\�g�Z��u�8�4��� �ӆ�{4gҮ\�W�n�uj�W��z�.Rj���R��F�f��������j
urZ��V=������؉Qѓܜ>��n�q�ٍ�r��{w���d�����uvWHRf���.K~V�!d�_`�Z��Ѻ��8��̩b6�����60b���Z���:�wd|��+&?}X�mU�y�c���_0���H雺�h�n���Si�2��4�K�oK�L�~���~m�'�D�iq^���V����A�<���}_	˴]���ǔ���L��Lx�9O�5ع�1.����ܩj���smK�4�� �!+�al�������tЉT�iNd<����(+��/6�h/����g�,��2-_�D�����`�$��ߋw��������k����u M
�>�<\���۹��y��iY�"r2�ܘL�&�HZ�]��(P���j�������-�qrqua疍X���z�:�"��������7W�w�3 ��e��/�@-V��9ă���L�mߖ�wM|U�ϊM���u��f3�k7�ν�bF��Z��1Wy��J~H+	�O�o�j�ֽ�5�!P�^mj��g@��;��(*��q��1����Ǳl[�v4��K�Y��|3a4�v�{ٲ�U5�f$H8�4ذ�YxV�"�[�9�&v�f'�1qJ���5(�6��m	��uL�]�>��\�a��nf�^r�z���ݗ�7,�*;���=Nܛ�"�ӻk���b�~5.�`��::�(��|A�C�	5�Ej���V�"|��S�S���ȑܣ�i���R�c���ޝ���P&O���3JT�*��J��r�{��f,�r_?���>�ǭ&��3����
:}͛�Y��6�4:˗�����P�h�O�z�|ǟ?��m8�b���$�&��5�TT0��P����&��cnN]1'ݞ2�|No���s�\N*:		�}Ĭv`�.-���~13���A�5
��Q��u�.��1Y�C����X�9�}��l�w�5'U�}UD������Tm�7�����$�X�JpY����G����f��4ƀ��Oscݢ�uP⟆�n�R��=q�ݣ�&_<��>��("B��ltŧq2�&����cBbc(6sO#�����ӆ�9��z��ZK
��BYJ�>Ȁ��[�ajF��(
ܠ-f����l�S��2wy�yCB�Ҡk�$�WriiIh?�����t8M��S�t���i�WN���	���������z�?tl�F:�07�"�ȹ|�L�)�m��g��o����s�B�-5�S����&?E��b�[Rt��S��T�n��o�4S���=jJӫk��	�T��)��O������2$磢5n;��M쮵�o�~�����ro�1����}��p�`e����TC*k�c��O,~��QoFcXg*��l���'Н���ڇ9a,6\���tD��M�$~q*y1��W��^�2��J�W⚶{{kK��ݳ��9Kr���H�>dj��=#8�*?E��Qω1� R=����i߂w �##�A��c�|�Zo�\��,��j�#��`6n�e��� �j���|�
���2|��������V�G�8�h��&BI�̴�H����� �����ղaAzW@ ��L��^����!��(���Brn��~����)��	���<�b��e�b<!��{M���sfZ�q��FTXw��i�X�mژ/�bj1:��ȡ�w\�����41�UxP�!�牺�L��A<��� _5����؈,m��X�a{��B�I' �r{�p��ԯZ���gY�2ԧ  ��8�ݔ��~E�i�s���'�����]X�Ѻ�J>b��c�s�����l�����q���ќ��}��C�������D��Ͽ���UW�l
���ustt$����KoO_����m�m�1c��s堬m�R)����c�E��	������oCp�����h����%z굻c��Q{���l��>�J\QGT�?��Ͽ{X�ޒ�7���xgWE���� 	u�f�J�y(/��wb�k^��#bI�6�i��^ІBY�Y��pD����j��� G�E�}]]7蝬�*����WE.7�
���첒*��>Y��hG�^QY�6U��;f�L_D�{�w�K��w>;IS3A1 u-t��k`�m�ǖ��/FP[�Y�T܂���;j���Z>;n�����:�I�Un���7u劥��UAH��1o|;��s[�[h��lq===�K��zx� {�by���x8�De�ǊR�x4�S�������Mei%�*[�P#����ʽ��/�ػ1�b�
�r�?����k���Sj7[�S�Ĵ\�q6���m�fs�ܑߖ|2R_�g���jG���@���q@�ec�6�)�j���m����T���ʔ�:��u{���˛�A��#L��?hA������>%�q(��W�}�	�:�OpS���
����$���)��T��;��g٣�1(�T��YY��h�~�I����;�uynm�}�blH餳*�ay�QN=�P�)f����d]eFG������.���ʯ��=W����؄�g1b!���԰.Xa˥����F�*'U�`��N�>�h�������W%y��O�Y1�x͑C�� ٭��������"ͫD#{ɝ�O����6A������h}��Q�#�?���Z�j@��i>���2C:<��F��؍�}�CA�G���7�������4��7����sm�O�]��`ݐ�[�5��Y�Xۮ�� �dc&�֙u���jO�=���&vv�T)^��+�[�T8
�_]iw����p��=��c�?��D6H��H��r���Y>�!��A��n��ζ1ow��͖\��k��ࡧ�o�W�f"��F�x)U" �F3)D��T�A�E?R+H�Y�K���ܔ��'/�^��ԅ�s\�Dr��]��Y�Gh���]->0@Ir�:�h�z6dpO���l�tg}��[���ǡ�k'Xw{�/��Y�����]ڌ*�������"���UՉ��xS{��t::����g�76�6�2��.�������'}���N})�pnK��h�a�cf�>s�j'��� �_�G(��#u�ϟ;����D||�3{�C~��w^��Qŝ�C�!���Z�TjނN�Lsb.5X���ɫ��/9�D5��B��Ჴ���m�WY\wܒ�5m��s�G����	�YLO�7xդ+R,��Y���>UJ�M�r���!��`�˾-o4#�`����X�i��s􌡦j�_��@��ެ���!�z'y�Q죋in,q����-1�'��T��]�q�IJ>��V2>��Jg�~ ��!7�ޡǵ>������)e %1��V�|p�a%�*/��.qJ�'d-��j�֖�r����\x�A���x?L=����Q��2d&��� o�B��A�%�|}'�,;��^�?�D �[b����-m��>�;;�o1/	�;EtE�'�Ь���?�i��D�-���_�����W_3e�R�f���`�L�2����_��r/�����~c	�wk��,�S���<M��2�}����̃���X}�8�-���0�����fL���qEhH��IBeBWݭwnN�l�/��@���Տ�E���/f7&޶\���W�ڒ�����s�O��`n�t��)O)�O���'.V%&&��\����l���X�C��q8Q�ȹX�2��5��R���
}{�j�}���pR�*��B��LX�4��Q����>�QǤN��>�!-��Nx0[�Q�����R������!̏,Ū����7'�䈶�p!*�v�i_�H����j��ìi�<�z�Ngp��$"�Θ"��"Aq�{:�޹+����̟зjՏ3�&�n�����+���[����h4�����ǽ�^\@i5���Ά�gM��LR���1��}(T���c�P<�����+���-���!L�س�Ȝ��\��
�}y�V��D��n��qp���Cz��%����C&t�N��tZ�q �?8k�K�����o��&�+��;��A)|@;Q���YF�@��K�~P���P"�k�z�V�� ,&��󍍚v�7���'g0��������<5��֑���Ksr���uhe�"ԁn�Ћ?ʥ�b�j����ߒ�DÒ�Zs\��=22�piM��#���珼Q�sCm�^��7X-��M�5�����;�������§�3C	��Y���v#j_�ކ�9����e��]�}�[;Q�<[\S(�IB�ooWeԁ|$;�E�J�����M�����ie*m�S�)�E����-�phw7����f�I/�挄nx�wy�/��K'(�Ao���QH� ���o%�7y-PJ�|��"
�A ���px@pp��v���p�1��2v�H���we��U$F��xL��S����ʋz�G���QBwy��9�5m
$���)�Ij�{쎀|�̎�d�n��?�n�'��n>�S��=P���b��^g���+a�wh�iN��&��{��u��n��3yL͞&"�ؿ�)�&��.�kŘ�3mE���:z�����#��	�1�A�.���aT���G~���;���)s��[k�D..��;7=���Y�O,����B aN�@��䓞��?�|�T�V�u4����a��/H ��gȫ�Ғ
e�|�!��Ah��I[��7�H��*��v��KR��e�I�3���J�o��ho�Y�W}p�����n�����Y���j�7b;׼ʊ)�o�ިV�N��ۻt�993p����eF��3��	�+4��<�+�m�����Z�f�������sY���l�ߨ�J�&�^J�E��A�^*(*����膲��I&���7�?�,�,��B c��{���њ���{u��cb�9�����OL8J�ρ��@]��z���1݂X�Tf���yi�/M�b7�"��\�K�@��� `A�C����W+�[Â���_C"ْu�Ř#S�[��Xtn�H��,�Z}de�:?ܿN:�c�7�(X��$~�+ʡ��kI��d����Q�	��4�)pY����૔ڦ� ���t�1��з6E�n0��{�zi^�e��1=���~��>�LRP�L�V⵳>�R�O	dp2�և��Դ(�9&ᨳ���j+������G�r��,�M�w���rJ�Kc؁�?5JR.�=�ht�Qr�39��~�`�1kݑ��� 
<9bY1�W�57N���ض���������V���£�'I���L*O�x�гk����j?GT�(J!�yO=�qtn9��"}I"�"w�ע��U�N�ĺ;%���Cۆ��%���\��OF��N$�Ʊ+yi�����[����%��}���f�*F�ّ�+)S���%�T`����BS���a��L���ԻMmH�/Й��Z�����_�l�{�=���zM��_�[S���I���^��U���xB{�p�/�C�4�;�7s��E���y�U�����ڿ4�ǲ��^��"��R�%�_r�%�_r���.�o^��5/\.]m���Z6�PK   Ŧ�X_��.
 �	 /   images/f557da7c-7f17-4077-a29c-07168c914697.png 4@˿�PNG

   IHDR  �  ^   sQ�   	pHYs  �  ��+  ��IDATx��	�d�uv�Z{�}�~��t��s�hH�R�DJ��HdX�"��$N�8��h'�b%NE��H��`D��(s�q.3=3=��{�~�������s��2e#i�E����n����?�w�ߗ7�7�7�7�7�7�7�����B/��ŋ�����o���)��d�����������2"�)��W�ċs�[��O�)S�s�Źν�Tǽ�V��{��b|�o����ܻg��w�+/������;��=��Zڽ��>�������]��}��1��W�d�c/�>��f��s�����IE�$v�B�I4�O^g��,O����{�����,s�<�u%��Hә䅓��Q�f�����ۻ�#gLw�����f;�4��Q�u��4ux��JPaG�H������;!������wj���	(.Kk��5ZA��;�������Z�pj�(:~�߉ާ�i��ӛ��Ⱥ�V~���c�8GI,�V(�,Qb�wfQ\HB�\7s�ɜ��
��@\��|/�@����"�}e<'t�s�(r��ƙ��L�i>�R���9��y�8�A�e���:�x�7Kr�����17a85��b,�[�|���V5���p�"���^�����p�t�YPk����+<�������IJ�H��	���ppX�8Ju������s�1%p� ��B�յ�2c��7/x�?g\,��_f��9΋���^��Y��}���t"<q�aڝ,���uC�S(����� �t�8~-t> ���3��$O�Z�����s=SZ
^%��H��n5�����/a�1�<w�8ﮮ�Wd1h��g��@�r�̜����p�s�	��7��A�N'g6M1�-|�Vo�3�Q�'(H��G��q�F�4C���C��NR'��4�w�%Ƭa\n��y�>��������a��
:��s���s������ ������`����u�@~�	�+O��s���LF�48�v�8<:
�Z����$i?�g���(��(��X�F�ǳ(��!x#ov:N���(�$������/�����?�����?,:�n��ð��9�!�P�(u$E�Y��yƏK^K�ÂF��K�.Ϋր�O���$�\�o����`4��������/����v����6'O'�Y����.ԟ���=Tւ�<���$@��!���{��̷'�� �"O1���_ĉyVk6�o���I ���>�܌���|<c�����`�o��O��M&�N��ΒXǆp��O_��y�7�����,J@&�S�W&Q{�U`qj�i8���gnel�Td���G�9y���A����>�����s�:i+hd�$-\Ld�]�_��?������5/T^��o>�΂���Z�z��~���?�������=r(����R����垜��K/��W���ʒVO��G3�]�b�s����F��q�u���ϳh�y\1,�����C��Y�a�Rh��(]�u��x�}�ђԈ8
�t��V<j��LDf���.&�Z�4+����A���G���(�3:����j��ˋI4�Q��n�i��q�,,�Į�`
���H��,���F�N�L&�����F�X��;�Ef���9�Z�M��D���/���\Ȁ����PNB1H!�N'x�M�V� ��@�� 2$���b<5 �+.^h_��5�y�L�%QQj4�� �1�cs
<�kzIa�뻼��.f����K�ە(��ݽ��tii��~`�X6,�>�K����Q��4�91֐k-� 5�Y~"���-�,#�9�r���:5���%w��l:�d�FB=��h<[X���fˋ�(#@�c�3���P-�f���~
�n�+�1�'�6�u��&H��B�Ҽ��U�q=]%������\R�
d��gT	E��vr�ρ �r�e�YNe��Y�%T�4 ��Y��Rh3*P�sf�@H XK}�S%B�F����� �!���>7��Ƹ�C��^�sN�LUFA�'J��.����JP��\�h�HNQ"�T���~� �a	!ˁ�Ʌ��e��B�����X���gY�����I��-��9�����[�t��j~���{�Ԧ���d6M��$j������������v+0@]�A�8݅���c���XXX̩&�{G>@{�D	�@�H����M�r�b.M{P��y�a�x޵z��S��I�5B�Ó!  3̒.'�8����J+.�9��"��h˨	�0���EqW�*aR�a�=��0��|�k��P��it;�D~u� �`8$�����o7�<������~��"]a�)�"p�,� ͆$�8�=��t����J��ci4F8���f�x5�ԜP\�Eg0�A�6��,��B] ����Z/�=���� j�� ��`D���R0�*�5�l�VL>�[_�w������[P}��B�����_}���/����i�o�GQ�I !�,Q�FhQjaC���\6��%��`��rb}%�aNv;MJ.��Q )h!�@�0GCwi�S�G#�.ᣌ�P\y�e��	a���r;�	�L�r��Ϋ����d4[�xaqY�h:����%�Э�~��kN�uQ�(��p֛���x��H��P5u��G��J���J���HjE%bS%0� Li�d���
���e���:i
�����'s;T9�TA�p��)���T8i��q:��)4.��$�(�����Ӽ]�>�A�@X�y�����3s��1%3�=D=�P�S���-��c>�q��Pz�z(���0&�v�72'����)Ȃz��^O��a� BО�Lr����<I�
���B`�G0��5A����P����(�Z������ۋ�k��xc6C�jfQa�2��Af��?�
���`�6��a�h$0f�V��9)S�[Bb�����3C� �+f-�RGA��d8�5$�Z-?&N�7���)��I�E�]U-p�O�KD3-��@��i ��-n�S�8����� ���F� �̼O�z����7ː���7�{5XU� �����:��vʅ��R��.wVA9cg� 4hj3U�������J.��x
���ST.�Ҁ��q_bdB5c@�x^�;`R��-����ΜZ{����I���t�^�ŋ�q1Gn��M�~A�n6�a8{)���aPX�J ��ѱ>�,I�ޘ��x�a=I/��U���GJ~U�E1��h�����L���0�d+έ�B�Vn��lR�f!�K�n��� 0!��2�wjE�r5q`d@�M��(�DF7=O=)|O�����Swiq) ����Jywq�9<9��=
�Ϣ�~�K��?�,g��~�J"	m!�bV6Ή��%�1�
FC��W���ũ�Y ?�h�H)m�� o�n�bʱ�YZL#�?�c���vS`:�~���àSo'��1�8�s0������g�ѝ������P��:�Ţ?��g�v���Ǔ�����A��ѩ���$���f�-�$���$��ޮ��x'O�ʓ�^hLGGd:�T2�T6W#]���n>��������O�w�?�O(� h����s�a��Ȍ$�K/~��T~�#�G{T�z����{�Z�(��Bw	߯A��dqy]�����ի���j/�z�T�f����N���1��@�P�O"	�M!�N��.M%Z�m7P3gjS��N�����i�9:��r
��c����<b~qe���N<갥�[��uX�X0c�1,4�R�������,=0X��0,"�t��iLW�3Qk,�z��p$ C�nueMT�r��0!�S�en`�8�|�ve�g�v�t������j����N�nh
�\?OאQ�KD�'A�~ =)t��CF��l2�������K����k�I��2�1r�uMp���'gΜ��h�5��{�a��󦳱ފW-�R����U���{����7��2�����
����a�W��x�R�O1W �@2�:�6���Ů�Z� ��T�4���=��1���hp���@ϫ�V�[T8x=L��#��%�_��X�5�zb�`����ʿ������%�|>3ʧ���9���Uo�������P���y=��.vkG���Y]ꀇ���PF�]���'��񁜃�988�ӧ����"Y[[��_>���e�'��k�����4G��d�ziB$�1:o�*��tbs�xM�K�X�+���)k���S�+�SO�l��1�2�s����=q�P��5:D$ŘS��wC�{�I#Ý6�NZ#ݧ>����K�=iB��#�
�I�)������L�YI��W��@(��+�A*�d�V?x*�Z�y���Q#�K�^̟����Ε��H�5�҃W V@��6f��O�0�����^k%�p��&�t��ww��kY�����'�^���q�s>�;�����L�erZBW���BGFN��=Yjvd���p$�I)���ăci�L޴�(�x����@��Z8J�T�|�`�������oޔw�㼜:uJ666UXo�8)����T�|�@�q�-f`����:sK2	��E0���"wH����0��D�`�m���̔��*XVR�`�H�X�Hs6��S\,M��p4������0�Al�z�<T���C�UAG���#ˡq?"�0�r��x�!}o��<RX-wۘ�t �J���`�!�=cë+#��EZ���b �[��Xvoߒ�Ŏ��T@޴x�S��P�y��&@��Mdt8�טV���Ǽ�BB�� �̘��Ŗ
�@���zC -0r���4AnB҅w���Rc�hh�pf!Uʘ����,.�`�d<ʩ�u�E�-o&��+�>��t8��L���
'^���Z��}`]�A�b�~<����O�C�t�R}�׷ytJ%�	,��)�1�z5�5����^Z��8+EV� � �u���^_?�p`�x�,Xw> u�ݖ)��ׅ�b��`ܗ��-���lt<�^��߫�5��{k�s0��~^��LaН�Ȓ~J\�J.tcn��EO�����R����;�'����$�!��2������}Q��_�{G�m�I�2�<�kक़�;پ�<�(��h�筬������Ғ���v:��zv��T��Y+ޯ�lm�BIֱ��7tqOi�z��S�S�tCoCa�'��9�2�Y��Fi�
Wi�w�Ь\�a�5ic�j^"A-��c�k@ᧉ^�kY�	דGѐ �J0v@M�"��`E0�ES�}��jK��aI�5<{�@��7��S_��F����gs�? !1�Ǉ2���,AcEˤ3��C	d_C�Wz��ɡݓ�G���wH��Z쐕�t��)<̩9�l:�;y�W~��3_��jQ|�M��y��N�{�V������cYA.uZ2�}M&��Ի�ȓo~P�;2��8qNKJ����ce���� � >�0�$��TaK�eO�!M'r�;�$���?���~�䪌���{�RLT���`����!�����{ 'W��3ix����`,u�k����J�C�D}�u�E9ؾ"^R&��M�8񀬮��7�h��W��̅�
��7v�dayh.��}9t�2�������� %q�ߧ������& �@�=H��[�����'~PNo�H���y&\`@�����˗��7d����A�4a^�����H����my����C�R��<y�,�*�)��0��aUX��p>TfQ���#�֠x�`j��D�}���o_����rt�&Q��En�37-�"S�%��[0Z��]97ADG�ǵy�;�)��[���kr	�s|���r��.G+�	�7K����VWW�گ>Eֱ��׮�3�Z-����{�^��3*y>6�<�͹If���稄�Z\��Ǻ�^��}��Hv�<�ߣ��,�յ� {�Q��*0L��pl�dq=�UE6C�����w���0�4�N�n�^,Oήm�>x�W�<*If��c/s)�k��7�|C��<�/*L@u��R&����%/sW������5�A-��+����<(��9�My_ (���FWNn.�3�}Q�Pj�t k�K2��8���d��!}) O
�Y�<�f�j�[�#y�Ժ>W��%�i^f ��?����_� Ҁi�k�l���͛�Rw5�`J�J��}�Y��mN�L��~��0D��.��6=6t׫r���Xg���`���Q�C�6��yF��a��:�Q_�5����m�/����wyqE��������O��t{tt����/^��7n(��Z�ܸ�|6��O|ʹs���]��׾�߭x�����o��$��<���0�$�fs2�gӕ+W$L�j/�gs�m��Jk[�vgA�!`��r��ډfI���|�������߿�/��+�����G��G^��}����A�.N������B�B��RX� ��:��,�:�P�,�i$�^~I�w��)��59���JT9��K�B �@O"E�5(���@b3������T��y��Med	�sͅMe�>�5'À� 06��L����'��\����*]��~O7�d��o�rQ��ڦ����o���\]�����=�z�ܸ~V�<���˧��3��uVN�?AS��K/�5�2��
�d�D?���B��an`�Aɮ����&�Jח[����&xϻa�v �D����!o��P���Uypk
��|��ɷ_|>�\q>��Tzrb�I_�L꙼��W%�f�@�5�i���M�$S��{�rcmE>���K/��!�K���xtP�i�lR����-z��ҏ���rɡ,Ξ8)�<�\�t��S(#�@_״��y�\=�����{�qQ�Roll��o}B^{�5�=S�������Z7<�{�7{:� ��9h�:֋J����q$X�˷^��Q�o�R��OS�P	��u�����{��N����Jo��)�H�����%��sU�T��}Y]Y��~O�t����Ĺc�� 0��W���M��I��2,��#=P/c	P����'�[�d�`40����D!Ja��|���={VN�<�s�;��J\N�5���\?*7&�Q��S��yR?�:����St��g�<� v8�2��^���0G#�7�q�٭�C)4��z���>�ߗ�7���rG�����.6d
:ܽ����ss�c��qj�X�$rԵ��z��'t�HG9�_[h鳾�·Tq%c�X��l$�L �MRy��<�r�
ρ!0�#UF��󉺣��
s��Z�z_�y���;sV>�����3gT��{x�����d:�z��#G�by7�'� qo>��|�_���%Jhf%J4������wn�h:�k�����W��ը/�m1*x��{]v�[���d��y�txSi`��ı�Gа�sA�����]��{�1��w!��s�q�Ϩ��,�@��H� ΅��2�OO�K/�h����8���V����x2~���/�G��_�'��K,��^��}����8uLN�K�d	mׂY숴�f��.���V�tzS���n�6aݖ���{�Tu�[�nG�e�0�D+��t���j ɪPL�h�nʘ,c�S���2~��P��5eC���נ ��1�m�+ׯ�&��@���� 7`���ч> ;�.����w�E<�!�x�|�S��o}�������?�C���!��7~K�PP	�%��\M)��"j��}0�!��P6 ���w��*�;-?����/��s[s���W���eL�e^�#�s,��b�a���-�◟U��wd���u�6k�p�����2<���	�?5e¸8ݦ !�t�n�* #�uy̵_L��WfS�b�Đu�ql�ž�VK0jS��]�1��x4W�\K��47��c=�i�Y��.J��� %T�m혞�� �ʧ�B`ԏdJ`�1�=���ЃbX���e� ޢ𠫑 ���8<Ig:ƹͺx�����X붜Xn����{Na���e)W^&=z�'���V�H��ٳ�C?,/����%�,ih Z�(��u}i�����u��߭-ɛNm��;�P�Zz2;��ڕ�I_��x6�B1wz形Ǭ���,�f�X���U��Y�#��͊;L�C3�P�!4rIR(�)l�u^Y]���F�2�c��@�罨@	ɿ��4��=�}�+�� )�˫r{gVYWN@Q,��h�B��`Eb�Ν9)K0+9�4�Y'��z�����N5�kI����E �Ul�>��	h��=Н�ӲV/�y�r���<X�nε���+~�g�¯��r-O��	�XW%0� P�����1��2����Z�1���L�)��'-aq}�EY m.u[��mK�*a����`ޘi��A�N�R2�'ׂ�e�p���N��3��W.OT�R��O���\"W�8�k4�ߛ�6�腦|��? _��3���*7omK�f<b�L�+��f'7O�s :���-����FCbK�����M��@�?`}Z�`�7�+���Z�#k�r��v�歽�V���������7n��vQ<w�q&ߋ���zB���@���%�P;��^�U>U�4%3�D�F�	a��z��K4b�(��-s��ɼ M��Z��D�o���0� �����K�� b˪6�UW`���q@u5A�@��+z�$s��I<f���r��)Y\Y���U���BPܝ�'+�<��{ǰ�nɻ��~��X�CX���`e&���8�,�i��&�Bb���:�y�������ໞ��FY�͊N(��IսX�����2���Y�|?����e�����}7��:P��H-g�-c��ο�,|����]((z^��+t�јA��L�V��qP�3,R0^�ysQŪ1PQ-ab�B�i��]�� �k�Z��+- ��/cΒX���}ta����x4]P�ZUo��V\�Z����)��Ռ^�?�����0��<\�-�9׋��s��zL�`O�Ź �o�N�̳ES�㾚/�0i�t��>U��0	�w�~-Ƣ�,�	c&�;�B���)�����<)Z��,�lm`c9�� ��W���͠�l���hG��Y�N�\�@55��a���N�.Nz�����L'��5K-TBŔ՛�r�bYl������3�qb�֤�YW����q��;�vv\�b� ��0��-G�7�^K�Xʘ����5t׺q����<s�D�S�w皚�V4e��I�a�����.,��,I��2ɵ	���ԩ�0�ϊWs^\��V���:T^Zm�߹�L.�K�4�c�:Yހ�jֿ.�UO�L�Zs^͈OUv������\R�Ur+( Q�@c��	@�����[FPA��[A;qn�<���[�7u��
dڭ�@3 	}\V��T�̱�2���h�������YfQ�����h�d���6�[�2lW#`�l�L����rx���*e9�n���(�>uⴼ�ꫠ�@���c ��͎!�,]���|\{�;���?-���ZkW����^���͵�7}�{���B�#���h��@��6� 91�\�$���%�A�:�֋*ҝ�9>:  hYK!U����!�"�v�Ք��ɾ�jkj񫐬b�d&FܘY�&��BhE�VK1���,���y�hŬ#U��D=�&�qrE�\�$;�=".\�8��kWe��o(���-���~�k��r�$�U|��G��}�sR�׈�M���s�tjw��<je�'�_����_>���d��rr+a���*ɠLHd�Z����Y�+�`��8+��.���g��Grvm���c�;~B����P5Y�Og�KJ�?J#�_�Y�Zn�Y�P��)a�ի�*��`���åۗ1c�5�C%�Ϯ�8�,��J��J���T��I�f��Ek�5�>Ž"Ƃ�n�)c}���@�"�ƯAy�N�f9� ��d��1���4J��|���D�q��ʵ!-rLR�4�-���b�vӔ$�-�!�bv�QA�|'�g��hޗ���e�+�*\��:&s���H�)�u�T�4d�e$��5)�qO�: �m��P׹�{��h�LT�	@3{�d�XX��5:�ߑ�co��N]��rkp�6P4�ܺ�z�R���3O]�L���f r�y2�:%�$\'���*�\��,�n}i�
%���%s/X���[�,Q���Ǚ �qLpm]�NK�Y�y�TM�*�s���k�қ����&}��F����`Iʾ/�ɯ���s�1ыV��t(�r�Yתi����ڴ,{GA_~�˛Ɣv�R/�T��q��~%]7|��z�XJ%�ǹ�Y�*�#?��e��#�Hf���<�� �94�d�4��T?�Ƿ�P~?;r��)9><³�C��,�Q�H�sp�4}�\�j�2Le4EO�%��8Y�j�h8��(\���[�����������=� �h9�#�CQ���錭���W�o�z�����^-���K��}��i{�qx@DD�t�Zd�\L�~g^��2��8	�uw[&����2>)�fQ�L\���s������Y��-~DB��y�D����؜���@��"u��R�|ӲE$�+KҰXo�ʑ*�e?�F@{CYXZ�AA]_�G�k/�	X�ׯ^�Ã�n(�?�O���9��]� �9K,&B}���*�,/�sApt�o�.����,7�Xn�_�?���wڗ,�D�@�6��Ia�T��F�d4k��.Z>�rŃ�x����˯�͗^�܃l8��2M��TMyi�T�Wh��V��0�UH-��)ˤ���s�U�eI�ֈ*�v� �Bfٯjm��A�74��D���F.3p���1�+]�E�B�(c�AS� ��X7>]���f��*�L��r5����z<r)�0�y�z��}o�[���!����Qn	МJ|�D�[Ě��Y�==��	�����:WeDړ�,#�:�T�w��IZa+2Xw�Z]�Ē>�d�9a̗VׄcȬdҮ���C��S��$��t��*���L��f]iy^fM5C$8��Ɔ���.e�t����j�j��uev�/]ΎV.`�`�֠����ο39ڿ�H�pW6a�y��g�
]�I�@���ge:8P��e�;�b��{�`eZB������ ޹KP�]�z岎�,=y�;ޢt�<U�@�9�Ω��Wc!Wo�S�e6��UVXWV-�c�g5�	|u��@��#̇4Ip��Q�V�� �r�]���HK��C/���Cnֱz$S �^-z�
����s-��$mz	��6�������њ%X�����yE�������7Z:�dWz��*�t��5��m5*�F]L����Ȩ�-v[��Z߅�fC�u�g�e����v󆜼����@@u�: Pm�����o}�X7�B�?��&�h�N�e5�H�����@���hx$�7��>qbS-�B�ΝmL�+b�I(*��Z��)��J=�m5��A��	�Y���جjQ@�Q�G��ebI2�@s�M\����J��+39&�i�V�B����+2��Ϟ;-���$�[�^�=[� �v��,}�z�5��ݑ�4�k�n�no"w��eeu]U���Z��œ��*�{B��K���\8с����V^2-}/P�2�����u�T���?��(y���"_��g�"@3I�xG�j�$�Y�B�����4�����#7&�a��.h߬�0V�C���>c��3��hR�P!P�xU�4���E�k�_��F�&N�,�M����@��Ks�2�Z�{��RD&��e��2����2�f.�t�^%x��K�E��@��nk���Y�w1>%�2�\r�\���^�י!���kuπ�v��4tS�,{��iv�cƲ_�}i8 ׮�Bu�3������*?Ԑ����|$%(�Qe![������ք���e�{ٷM�u�Y��fa���W����h��-=4l��͔�"?�J0f��M!Y�I�H�=wө*���/GG2<ܖ�3dp���U�Dg����]�Dk΁��T�r�\Km�ƙ[@ ��Y�ΠU;��n��e
|b�,}k(c��p�e�;h�s�9�)k���-Ti���&-y֫[R���
1>�H�Sw�)b�HJ��WIe��$:%�u��esZ�K)�<�
m��קȪ�p���ZU��h�n���LxR�	k�d�`ieXk�x2T�ǩӛ�g2/�������TXa ��]����f��=#�YZhk��?8���&S�`��阈�_���L������K�.>�V�֖%��5�k�Ӗ�þ���E@�� ����N������	!2aK4Sw8M�didY�X�i
k:ʫ�n�`�N,V����FwYˤ��%^YFS��Қ��pbXpU�����\�����.�*��ȭ&ݳ���	�^̘7��'�v���"��3
~�4`Q,�7�� ���m��:�u�8oo`�<��
4�4塇�G�|J���/>+�v�e��
;5�̹�ڭhM3�+dւ�28XVL��~@?oB��ϏG)t��+/-X��B$S�s���i��R�����!.��Y?�y�&��A��)�DѶYfj��L��$���V�]#i*���d����ךVeQ�NIݡ�"U�*]�Z����{�q_�o�
]-9��j`o� �,�rܓYZV�Q���_�1&G��
	�"W���%~��v�%Y�?��D��V^�^
�@��i0�۱��Gp1���@6��z����5,�3��� �Y�r5�`2���?R�$H����@L4"8u��w��lna��������~���А
A�,�J���D�*�?W�°FV����� �1�CN�K�R-J�*�	��Z����G~l�����,�����S����*:�[yUY��G@@����X��%`eBe^o+0|�W@��!�'Ù�R���7{
�ìJ^AD��c�U��S�ҕj�����^)�f�# ����k*��?-IO�[�'M[6�jw�6ֹ(ͽ����3#:���m���|T�KV�V�?z=�d�:�]m�l�[z���!W�k^1��)��"+�%tnJ&�fl�$�V�|*����`����P��0��"j� ]��0�GJ�μ�����;<�ކ�<M��׆���G\$����i(le}���)c�[�y�������[|ZR������C��p�w
�=���<q�%NO_ӯ��x�29e�gWcI��ړ��Y_[�,݀S3�&`�@��<�<�:f�2�Z������@�?򔛰�5ɧ��6��,�`�@��hL��l_��.-�H�����#�0�}��i�z��}<�����GU� 7���{�~Z�V7�?�ޕ�A,��EYJh�5dY�����r��,V|w�#��.ʇ�~R�6T���Veǭ�Sˑ)(�dÑ�\i��L'MbZ��:�Ii��5j�~��Á֚��br5	K3�33�D��nٲ"���e�[*s�+��=�����hZۈ⾡�Աi�E��2F�j8!.-O-wù��,��V��5w)��(-枱���ǠQS�����W+m��b�N������v��Q)��d�ٴ޼�"��T��o-=M�:L�k��hH�Ay�ҝ�D)ݶ$Wk�9|O�h�h�)"�G(�U�K
Q���%r�̪�A�Y�2�����i����xdeRa��|�jN�Q�ʃ�sU%�U��j_8����S%��}�z棺�5��ҍ�0�����B ���~*�t��K3�� ����e?+��Xⴶ��9M,[�֌ƚ#Ua�]U�����P����{�38wK�hz�U;z����)���M+�Rv�2w�,�f�!�sʆ6l��淴�)R�O��7H_�PO�S�I��K���)��RnYn�U*UY�=!#]Cŏ��>�1���x8���k׮���J�j)ݒ/�ǖl�j7>J3�v�Q�Fi$���0ƚ�F��[�	�vw%��v�*���;��,���a�'����hl囸�x8�vؖ��]i.�aL��,r���}��=� Vɨח�t('�O`h!XĚ�����zE�w��P�`��\ٓ,�p�tቼ���dԟ(:���M�wY�D���b ��V�(�ǲ��g�������%\��B{M��t����s����ey��m�0���+7�N*���:wN-���ұzـ��Z�l�ٓ A���)�j�g��;��!��}�����o�&[g�,qM��di��kșs$��e�7S���t5s��Y^,��`a��cu������׼�d�2u�D�b��e�6&z�5�X/*g
a^�uƷo�ֲZt,�����l�W���(\貥Q�Y�jW���]S�a�͔�L�~T���TImL�	j����MbY^Y���2�uӵ��$R
(
�.A`�7e	=�$��U��qQZL.���n\�6�f7lɚl6��İ�q��������@׬�,�����`!k+kX�H^{�5]�6�جP�њ&�m�F(L�bF�li�BܲU-�J7��a)�����֜��TW�X9%��cK�b�{�Xw:f�|5;MX(+��HbX�ݠm�	im�\2���W*�z4h7���=k翂�R��rEӭ�������&�>#�O��6�3����w�7��M��N���O��ER&�3sn��������5���L�̭	�l���?�4������]ߓ��&��5Yi/I�cx�V��@B=IjuZ��>;��g�ؐ�����Lϣ!�r�BKL�{���2|��d2���#C@ts���O�ܰ�\��f_*Mδ,�Zؚ??s[\�*3�9J�uS�̓�ʖ�x<+��Z�����F����ll�P�`G�b���C|�c<:<���*̫��l^H��:���Z�1��z�TZ/*NQz٬E4��|e]8icmm׮�\�<2��'H/|>?����x�(��ma�.;Z_�i`�Ho�:Ő'-r4J��ƳyrK�_)�R�Ga�]|�%	���^xI�V
c;#5�G:�hl��p�Y��M�g:�;���r��L���`ʃ-%�ngE����e�Ξ<z�Qy�⫲s��QZ��{$����R�#��SR#�����+ɚq��ha�+2�t2��+��߹)_��o�SO<"O>���ܑF��J�yj�.h�5X�_���e�M������(�}���y�]���ؑ��ѝ�xAç�]�I��Aw�/=����m�:���Row��˗�k-��"mvee��NX�A�ϓ�*'U�ncd�ۅ�pK�f�ş�zXk�)2X�Z/�R3q�X����js'�c�����}�=�t�bln>/ӡ¦v<��U�♛}hQQ�S-��Yݲ�]���5�-I�ޑZg�h�T�M�sPy4����l�j }�����6���k�T��i�s쎶��?>��	���ߤ�ft.�`��eB�ݒF�����ђ)h4y.��V��%���Za��pf����X%���ּG�{.d�LO�Kǲ�&�\=2\S*��2�Q�E+k�^�¼���m�Rz$�� �����{[�rݭ.��w����n�Vv�{������:�y�e�V��V�����D�5�\�fK[�~�#���wQ�m���,��Ge����@:������7�1~7�I��T���r�2�3P�4P:f�1��ύ�XSM�V��+@cI+����r�Z�j��^/����uSM���֠Eݿ��gu5�p�=��,E���v�l���t��W+�U��yК������ʡ�,d.Q���Z���<(A��kW%*M��{Z 73 �v?���E�%d�}(c��Vm��]��V�i�9��p%#*O Hs��h�գW�,��g-��c�p�לzj��
;
6.���&���E{T�ټ1ɿ�q�)�ܛ� @w�]�
��Ot]�?6���\�rM�����EpcxS�QOV���A��w���r�ʊD����Ť�^2��#_�r��,����O���d�^�(����H�4tQM���0z��IM���K�Pw$?��
����Kca�ڒ�C�NW?s�eL�2�XYY�ҝ���p�{M4�oymUn�9����AQ�~p�9�\�I�n/��M $@ۿ�[���dEYb���n��2���|LQ���9�3o��ܛ1Z�j	�W��q�v�ݗ��G{r�ԦZ�����bW��Y}��T���z����%%�Zs��EY^\V�FR�׭���)��H	T��ie���g�k=���ns��b!�b�]�NY�����Zh�Eg����H�[i���Mq��u�r�܀�㹽� �Д��e<7�̾�f�X<��T3������Vs�^�P�����U�T�`�yRMZ������
���$Vn��L5����;���t�6�TʗzGX���f�n�2�9_Y�^X���Lhr��7�b�N�3��L����]}�$�N(m�#�a�ܼD��;��#L>ci'���W�a�$�$Ɯ�6X�6��R�ֵ��(��w���P�s���1���?�MA;�r��k�f5N�U0���Mg��sL<��ʙ�N �m%J��:,�zݬ�ڈ��L=KLT��g
���,��uUc{��>���]�O[��p2/)����ng��b�m�0P�2c~K���F>��1''3חV1�ɵ�\u;��PT��L&@�d
|�a��Z����*PF�Yպ�?(O�^1-�4+C=�|��^
��u����<�����n��'��
�/��ȘÈ
V0f��e,�Qo�4���^ם��8��h���[�b'O��3Ot���<�FG;��~�8A�|Oʜ�}�Ё_�z���d9��4��<C�#]�ލ�HVA(;�r��	U�7��"gN��ߴ���dxl�p�Q���tπ!�:!�|�醮��}P��}�s���lo�tq�L&Ѯu���괴􂻛|�+_�O~�������ԃ�ً&���n�H�!JM3�������eʚl2�@��,� )�,�%i-�^ݒBQ�/K��,�� .3X)H�*���a�B�Ai�@�=�� ^"�Э���q*�%�u6����ۙ��>TlR��H='l� �Mi��+�XwK�;����vL�w�~�cK�q|Ua��Zkh}�Y�g��sg���ӰX͊c[O� �H���6��22��) �\s��猦c0�H#�5<�?+y(��b���,��sS`1����(?�����}��'?-�ݹEZ��iӽ�Rl9��h��lƢ�P�2g�k
\U��e�<�I����p�oפk;MLI��Wf�[F���Uz�1*�,����WetU����W=�uS��u^\��R&S���뢖ub^���3����WVK���������1�(�sVY��s2�s�+`}�yh_���_Hl�J����_����������W~�W�h9&�x��LS=hy7�i�!wU���������;*7�	d0�A�G������iI_��N]�P�.���bG����]}��E����X��Ҳ6
���s���� rv�0@�������Iys�:p�k�G��n꾵3�B'�ғE��h�c�z�c�\+_���<oB�~��p�9.۽����z�w[�/���-������A���^/�%ȚGJ������~��G��~�|��ض��zҒ櫍r�����?���c%x�-��{lEnt���&&�4Q�g:�;���s��\t�$�c�w\�o~��)��z%��Z��,�n��;��ܔh<��o}\.<x^n^�,�/��}����0K�$)��Bz�w������{
�a(�7�Aʎ���2�?�'O���m�0���^���'�����O������������s��$$�B��*���I$��� |�d<�x��2A��^^�>�0pVrC��qny�;���<U̴*-�(SK���[��A�'�l��eN��ey�Z����:/�cY�U�quO*CZ�k����ٗ̾�yBN�-c˚�\�b��%�t)�sn��+�\V�a%=�<޵ybk�lUsYXY֬ov$3���
*ԓ��A��A�2yP����-�e�dxZRt�_�yC�P�T"Þ�:���T��w�
�[@�����z����L!<xAK�h�j�y
l���pgހ�V;��h�3t0���P�:�+s�j-ԙ/�%D��������n� ��y�ñ΃��	�J˸�p��&��s�Me��+����sH���Myi�!���YIi�7� ۱��A���}����"Ҍwz0B(��7���i��c1P)w<����,ف�@',w�cb]���C	so��M���t�[/��BP_���ٟ���W�^���[����rp��K;�z��$ ���E.�y6��Nx�8����׮^�fD�q�9!EYwHK�JAK��7K ������T�cX��fG.�ti�,[^;�������ۅթ�
f���iХ��������W�Rg�AZ��S9Em�0ِ�'c�]�\6,:�ۗ#(4W[�Fꦣl^��Ӟ�Q4�UR#��>=] ��'"=T?�Y�
銍t�{�&D����M�E��ח��O�^MA�h�C0!T�A�K�~s���J^��K{�8��C���L~��g������]b���]���rcZ��m��~?q��I��w
��ǣ"-�����C^�I#�RkCڰj����Ң�`���r%Hcb4��֩9>�me#���j�1�L�a��ʋߑ�<�fiw�rp�i�0� rh�{��a��#�F0��U2��՛7�ч�+�<"��ߕ_��o��Eƺ}�
�u����S͒�49O�<��h֬��%�J����.�#�=._|Y�,�u�W�n��T�E�X����IK���S�N��Զ4���|��%9��&	��J�oYl[�rc.�ײ�]Gw��J��������%9E�Ԛq!]�ui#P��_�5o9iI_���.�����ɆT����v) ��<XZR�S10����Y��/K'�|�r��-9�L+��4 �VWt(�g�^E�w�n鞞a���!M���v�fw���o�X��#�ϳwx ���g����5+|yyE�5�.@�Tض��Z��>�|���0mS$�z%�TǍDZ8o0�^�d݅����"�^�s  I �mؒ�;���QX,�k�RS�Z�2C��Z�fIy��% 98>�Y���G�O`J�H ��{����~�
�)���h�"�ttl;���5k����3�/�Z���t��>L����5�&I�z]�Lx$�i@�W.��м����/�+�-P��9G��ǚ�׀2�u���=���[Oo� ��ᑼ��d����Ž�e�����-���y�[�K�&n��PQ���Y.{ֲW]�[@�� ]Riq}O�>����dZ͑�ʜ%qE�e0U����pO,�����s��]�j�sⲛ�H�����]�� ]�qV�8j��@��oܸ���{�����P���ޫ1h�&h>+�j��q�^��SC�וi���7�``=pO�MϥV�Py{�^�ߙNw�u ���Ӓ�����V�Ah-��)U�k��p��́Xz{{G�d&���z����`�{U�RyD<1>[X\�u#��e8�J
����̹a��4s������;��Y���&~+56DHE��� nҗ���)���="��J��D:0л��ץ�_ ��Yjk�KB��LD�i�S*�\;�=x���oߒd2����P��2)�� ��صr;K�5GӉD`�-�vo^�'��/���޺.)���['6��934�g���ca&�P��R( u�Afé|���/�?�9��/=#��˿,�n�&K�'���78�qק�� f٬B�W�xH���C~�ԕ!�s_|V�Mrv�)x2�X�!��d7s4��2���u��*�2S�CE�A��My�ŋ2����S���e��1�Ė�� a}4Ks�2��kV:�/?-�K���zpÉ�ݤ�C�՟T3���*;5A(����j��P0�����m)��tY�9�V�n%)[a]��_�i���}\�����*�K�^�g�yF�
�D�  �M��nm�Qe�y�Z�#����ߴέ1Y��d�w��������b����{��&�� ��f�rUr�I�M&�EA[l:��g�[�%:T�,I�6��B�C��{}{��� ��cD"p]��XϬ�K��@5	��,����h	X���u�,ҿ*�e�祥JE@����y�l9�TF�������r�x�5����@�7���1�25E�P��N ������6��>yt��,�v�3�NE8�?���j�x�e:�T{7�����#�؟7��i٣�5����8�]`���p�8֐*ɬ��X�I�E�ߍ��rgo_A���S��@�j[]=��hd
�t��'�k�ӴNIﺦf���/j�Zh��C��|�Y���Z�gz�>��K�@=h� h�L(3f�[���Ώ�S�)��u�=Nn���F�}�Ħ�wyЬ�e�Hǆ5�W� �@����L���X;!6�N������;�44�^X�L�X㳅u V��Qo ܒ���,��R*h��),i�)��cn
֬���'��kus��������|��o��S��ec�w&��d��APw�@�@�1�����5k�������]�q�Z��mY^j�}X����v�҅LD�f�6� �cW�)~g�8Nf~C`QЕE+�^5�(���?����7Hl�ehs�0���5��<���}X�~��D��Ɗ�Z41�n&1_���RYY�����ީ˻��<݄R����g>�ek�6-`OK�X��������)��k�V�ƺ�������7�uQn��ds�������\�n��*��qRa}�lD�aq�֥k���� 06e��Tn�_�x*#��г�U_r6�����-������Z,S��͎[ז�����־�����|wOkŷ��UJ@t��W�1n
 �-�,T�h
�nmZ�Z��u$H�B^ZY�hz;(������'��O��ё�������\P�������(@��TQ�뵘	�Z����~��SW��t��9�B��ţ1��������h���y�$��x-f������uo"�F��Q��=���	^�2�hU	�Y���Z+Y�6�$hBg���e�XT՚��<�cb+ز*�}i����>�Z>x����`[�#���j���J
�����bKN[�%��:��%��cW�ݹҒ�,Ϊ1q���c�t�����+ �܊sme���t��sg�%�M�Ro�V{<��ey��5NG��i�b����sA����&lW����v[,�r"ܻ�tD���qc��8�;�]}զJ��E5��Wfֳl�e{Z̆&Rm<��\���f&{;hwZ&�L�bM� _�1�(����״�[Go��3�k��vaa	���v4�) Ҍ��r�r#�2���9}��U�B?�H����A�Nٓ��̩ ����4�8�i���j���>=
P�{���?t3&���l�1,r���gu~��Zu������74tH�$�dX���\�S�=�u���t&?���^\��m������q�)to_j�;��i�ueT�m=�ɧc9<�!��Wey�F}���3�j�-/w�o>YT�O���Eg��1r�Ȟ:�%_��/�ç6�Y�K�em�S���-�Ig��ȴֆ�z�i���Wd����\�|E���ք�7�@tɔ���K����_Ӥ^���յ�-R��/�������Ɯ;y������2�%l-�v�*(;K*䋲	KQ6��c�i��<ֈ߸~Y[Rۻ���O���ݿ�_�,j����Xo*։k+β���e��ي����H��͗����tRN>(��{����lk�Q��n�Il<���M)�:t�[+V��K�@H���`4�ض<�ج�o�@{�S@Gq��!|��@]WFS*(wސ���4fIK�.睽]�\�P�¤
�/�K^���_~��PY�e����
�������>
w��Q�--PZ.���y�Z���ĎzCuՏ�}M�Z]^Ҥ=����x�Ca>��Ӳ�-�z���|&�Ъgrύ7Ԃ�~г�=�m�R&�Вfܒn�%С�C0f�y�=������{
h��UX�d�{Qf�[��<����O�MQ��&O���~?I-w���*t�Jё�5n��~����}w)\��R�����Jw��Pȏe�PZr��t���mN��0�N��C����x����:jS(LƧ�:s�*��3�5�����Q�Zt�l��jw�N{����h7�}��e��*;�""�դK�� �sP+�C1�I��iR�� (���,KԸrh��Z݀���͢o�[�ˀ�eb���������Tx��S�Q�{̰��΢�F��\�(�ֽ�NT�p\�u�:sc*�(@�p��A��Og�{*=�9=�4��dr2�
���`8P�{��ZU_�֫.�������yLfLR�T��&�x�:�{#�����{<��f)4"N��|����zq_��'��q�)�2�p
�l`csMF��J0uX�$P��?T���T�.5m4���\�9.۶�B�u Q�V��V���YI�c�:��x��1m�tg���s���v��":���t��-e��Z�NU�b��l���7^u�BK�;1ﳟ��&�,��}���jl�j�!@)29��S������t��%����학�k�!�M����r}W~���������Ӌ���s+=�Px���Xv,�?�F2���`�׶w�ӟ{F.�<�0�-i&jo/�����=��SM(��8�Y�a.Rv<3W��s^&�ini��b(}[��M٫���9�g}���j�l��[���.X�k�<W8A���r��Ui�,;��ge^��Vf��x>��Ϩfv����_�lp*����S�p�:uN�oc�TY�\Ӥ*�S��ɧ?�)-�j-,kw�P�k��;�!�g�}mXA�����QI�/�
~��w�����X�6�䘥[f��剷ʃ.�����gl?++&��y.3��1Oa��hVR�m�%�����+?��z�(���F��.�naZT�Nն�?��e���;ıXs�{�G�=ex�6�����T��p�Q�	y;�=�v��{�m���3�{�o��W�����'�$ӲDN���K%x����:#O���a���f��^��3���{�fWY��?���5����@ �HW@�)`=(b=z*�sQ�
��D��	��T�I���}��ٳ�^���w��w}��/.�W���{�w��S��װ�[��{Қ� 3C8���J]C-+Au� {¾D�%t�������c�`�:���u����VK�qf��LO���k �黗��*5�:�L��G?3VUc�>CxSt�*���gE�%�I^6ny]�s޹"����A�bz|B�ܠʙBU�\�Ϣr�uA�{��^_���^�U;����j^%�4��B�l��"aI���X� �?�g�/�.���ܕs�|��,'?,�S�d'�\�V�p|�l�ca�\���ww핃����T�7�Cw4P�E�y��`.\8_�r�I�wkf�"1>y���9IW �R�S��2���yjuш �z�ٷ�W鱹��0�9ZS2��>3o��X�-���5Z�c���em�-��FCZF���k�<��-�M��h/��-dz������<��Z�C�,{V���M�	ʊ��佀T�#Iy)y��F�[d!NX<5�2>6�����Vt�;w��~u�|�}�#�X( �ʔ�P&�tcej�1���z�����M�e����揳g&(�f�Ѫzb0��쒙��S��!f�f���e/	jh̥\!�08��}b9z�p������8tF00pd�+ �j`xD��fAP��РY�$���L������{�Ѕ��3�8Cּ�V�����tǌzh�Ϛƫ�΀� ߫ϔ�4~�E����{YVh����.u�5f�@���z�լ�mŌ�3��_/��!��l�I8��K�C=�N	�� ��/�H�����W�������n��c�Y��P��W�\�����| pA��G��������qN?�� _;찊J�������
����p��0���%ϙ9.�3���� x�Yz�AԸ��Kw/T��0�L.x3����u�M�Q&�ݣ�1��bH�|���,W<D��A��g�� �%[A��{�s����Ȱt�@��bMC���S���&�>�|Y�d��A&���+ \Q��rF�־ >��(Pu`�X<!g�}��^���HJd]�u��x��m�vY�n�t���"���t�"�f7���/�--�k��9��G�`�1HGF妛o�}{�K�@���N��#����+�$6g ������H�����J�5F�5�Qb�{g���f1e��nVΪ�>s3h��<7X���x��`&�K���W���?�p�K��L#�m��c�|��5\����C`1��c��EĲ���������Ћ���6�3�[	�*%3�A}�@��2T��j�'$��,�p����43P�,���0�11�V�LjҔ+ߟ����X��Y��Z����푚�N�[ �̙m�Q �bƎ)�!�6b
[����J�ne�_F*�N'�܄����'���"1p h��kz�r	543��$����%�7�,oY�BN�I�dA��e��J,I�}J�hrJ^ݸY���5 ހ/� ��c"�$�e�f��䄭 ��'(���rPU͌��OC�[p�ְ���M�UQk ��7�MIss+�+ԣ��Q�a?/��^Ѭw�!�HOo7�i�H8j�{R�NN�,}iD���K�N�������$�Y�j 8y� x��m+~ϧ����	��۸I�.�&�9pz�4�>ރ���sUu�fd*dX�L~s������;��wY�rv�F��u���uc �e���o�N}���?��@el	�᳙��M��st|0ⵂ>����({5�c��������錤�#�A�L*�Ȃ�m��Dd~�/ ��w�\y�}D�N� 9��V���dT^#
�-3����z��
���*_��~`M��|L<w�ӣ�PV�~v����m����53e�.|Ş��Y	k:�:���r۝w�Y#q@0�V����6��'u���J��`�+B[��˯����;.�l���?8��>�H=�a���ѤlذE��;�����el�d �Q�w��t9�]�u�_e���'���n�a��!pv��x�I�a�qY�0>�i��D3���N���f��НG���ƼeC���C���\|��"0Գe�A�����W�14��Y��T�%I]�X�
?�)�0"�!��P��}�l�I^����С$[�Ԍq�[52l���8D���i�ޡ��ե���B��Q�h�B�j|ri��Q�]�u�(EST�\d�9>>*��ɪ�E9WIuU��~-��c��2K3�Be�J=>�w�@�����Á"U"c�Hv��L�,�E�e�idw��F�^R���P�u+{L�7q�]�Eʐ�P64 9� �[%��>�W���>h�HQ�X�+Ã=���O��tтi��Iscy�GF������z�HR�S�X�Cp�qJ�BF���F��&�T��0��z`�E[�8�E0 ��?�p�ާ� �y �N%{'SU@3��8�l�F��{X>��N��D�Vg3�:�X4N'��\��9��x�k!�����^$MM�>�R���}N�Pf�φ�KN�i�L9Y�rS>7  ��1o
��L�D�(�����%f�Q֣��d,u̌9��Ѫj����3Ih���QIOg�� �W;�O ?�m�ݱIcL�f)͢��T��x��?�}�Q~sӗf����x��
~��d����g�=�|�Q��'ؼ<�����R�8�k��%�q��8�n�˥YuA�xUO|Y�f�Ƕ�Ď!��t� Y⿩��6�;H�#F9���Ǡ�Q�F��s��e�l��c����T���<�����C�F�|��-
��r��@4j�r�6�ЕC�CΪI(L���wJy�f���0���ҙpJ!��7Y�ҭ�[ Q͆׼��� �b��gp*��"��\�s�w�S�'�`�Bڲg�_+]{�b1>�,�EJF�hw���@[2�Nx� P1>��c �w,s�eMI�<{�k�T*0�B�B)\� X��S�#b�D���X)y���l�EZ��Tq�����b¥P6�To+�-�xJ��;��|��z)h'z�13��Q�S;�a�xC<�H��h�8��s��͚m6A�<�ʈP%м��� 1me�L/�O��eE+R���wZp�y;�a�DXnˁP��[F�Fe�qo��s܂
��G�ec�%���5�_D�8�%�Y""Md�9�b����8����ׂ�#&j�S�#��	J�ۃᡰGWl�� ��$��!� c�gX,\ �z��t-�$@f_��cB3��:�foz�C�j�b���N�Y�M%�L�	" �Q�r��A�m[��e3��:�
�`��a_�k�m����X�hgf�]�<J���y<��O?��č��ȭ�����v�,��y�GF0� � dJ�3�(N�}pC�Z.HOw�lڸE�>z��_(�*�M�T�����쿖@�1 �,�)�Q�	�d�g��:K����{+O����S$h�Ufz���3��,��MNJ]u8K��y�ZC�C�{��)�Ƥk5*�p�XC\'� E�I=|���f�'���Jp����»^���0*�nא�4�`�=�1��T,(�C�hU�Bc��E�a?F���|��άZ��yF��%�1ѝᢧ�Q��W�b�:�������}m��0�,C�Sjq��(R�d��
�)��!^���W)���1[�3����`���9��,��xMP���牟���������5e�A�v�..M�ul	 Xt,oy(��C/)�q�s)x}����
���H-��� ��@ ��pq&Ѣ�N��~>���u��/��hXyN���
�c�����Y`*� �_9lFyQAd����^k��= =4' �T���Ӣ�?�3�ϻ����02%>�8����mU7H��ܖ*��!�@��o����2!�ɑ���¦|����B9�������4�	0&�����L'5���j�s���%�-��,�7�B���X��%`�% @���W�6K��Qcر�f�v�~1�/�N���:�I��ե_�t̝�2��M����p��Y�y([�0�
�f��J%	^�Y�-� d������+zi(e�(���y@��MQ�gT�����<�á%:lS��[2��0G�*QG�U0���	��C�M�����:��tun7���IT7	�A�UD
��f�U-@/ ���(u�����,���,
�k�q;ʒHD���Rd� Ζ�YJ��� >!h1E��:�A��K�cO��_�$<x�:�՚Q7�c�>!ms��#ZG�\��m���~���+���Ǿ�a�WG�K_���v�i,o?���|fcc�,�NL$Yy�F)F�鵧��<pRÐ7h ��(�UFx����Q�'�g��0��[(�W�H,ZE�����|�]$.;Ԥ��Mg���eӬ����r���UŐ���f�Ӓ7q*W!"��A���U�s4�=K�B-ҋZ9���>�1������� Ɛ�����H�� ��̃eֿw��{��i`��k->��Tz��.���K��q��l8�����]��t��)R��Y ��}�k"���1��� EA���:R�
�"�B�NϠ�TSWO����yϒ�� ���y>7��O��%�����2��H�a�ےb޲��-��?෾�4��-�\5pzP	�g���:��k��E�P�����C;��+�VZw�^�1-3�@��f�f&�cp�#�-�#�T�!�8��>;/��r]���6Ԍ�I �����GȘ��}�9R��W�r�w�&� )i�e�\Y�kj�	�	@T�����Ρ�O�x�L��~*��Z�wx��}�fG�%��1����f���)˪��D#T^��k�.4�T��t�5�蓪�_|�2��٩���%��j�B�R����,��^�Hk3N�Yx�f�}ã�=2,'�q4{�������3��EnD�m\��;#������z�c:"
O�rP4D#t��0<�=0��@L3��4���FfQ�v��#[��SF��=�B�gb?pH#951*}��t�����ԩ�y�CÒ��VG��d�z�U���+h�s�)�I�dl
�Of77����s�Oٮ ��I��2�y.����,�,��}�b�e;����\Fv��8�tzB~�˟K����'���{噧�S8!�t=�=k�n��Z�p!9�����RW�`8��S�� �v)T=����qn�h]�u��V�&R�L# =�xTzP�G�՝��f�"�Z�f�n�B`�͚�L�-�ӌ��pHG|q������s\'Z-���g��0ͨ@���{H�Q���@gT�K�-�oC
�,T��w1vt¶l}U^��m��!�5�Q\f��xF0	������qAI����wN/�L� H����X�/��yj��n������ɋ<T6�9����جߨ�y���!N�X6EruC��1��<���z~������S�ř`��JӢ2���c���X�����Af��X��"�Rٱ�a�!�֢��:H
j�5D����0�~ qKA��㧾G��"��H��t5��Z�Q�=F���(��5H��E6��������>�7���Ǥ�� x�y,b1�FnզhG��=e��=Vx�P�ϔ���p�4��<8aDih+�(s3�v�,}���k�./G�b����
W��*Sά�:�FQ~��NYت�װ\�a0�:4� ��z�9t��q�|�&P큱�C����}��,!��4�fR�+�j=�׮\�HYt�F�)�%@iK��� ��X%����m,q��w��`��ԁF�k�0K�"#of�9#6����E�:�d(���^zQ�>����P��ڦz	'�1LO�9��J��k��'����VsV����}=����~D� 3MY�D�a�h$ �����'^�������Y���$G\�qc]��kTgB�+u�S����"*v��nii��s���ޝҹq���C2=1)y��,a�FHf|L<�)�� �NM��wɺ�at����&��NI��:=��=z��^�)u�9�%�$jN��ɴ͠�y!C-2�Ʀf�Τ��Pň�e�.�yy�/�����.�����~�۵K@�
��������Mh���XOR������_�x��޲��6��5SG�Q[�h21�yp����ߖ9m���s��H��t��w����wj�Uk��2��3E��_�yʦo�ָA,��*�00E� ��b��w�F��/l�p]� �2� 3��C!��m� `���D�q��=q�g\��b�o2Sf{�������Ir�J�)�G�tԑH�:�Es�P3L�xٟ�ؑC�R��G�����+j�lvg�c������3��O��)���L� `�A�d��W�Ǽ�Y��I��� ���b-�̯Y}ysnq�1�Y�#x �b���ʄ��L�%�5��/ ��B�$s�9�1�� [��	� ��xM�k�L�^���ې߀�ж��L�JE�{���p���}v|�� ���A�M8�Ǆ�an:/U�& @	{Y��b���QM<�f�6����d2�}��cJ���F�À��m���������$��І�� |���(ׇ�n@)�č*��qJ�N�㏎i�-.N�8e;�`��P����{��n.=�<��{{��6f��C������p����y��>���(�� M�Sb9�
���4+,���`7Q>T��ƣ��M:w�z\�Y}U�b<�f�c᩷m�?�$?�?(Y*]{vɣ�=/'��YMw�ni��mz�荡p���n�щ!�;�+k7m��'ǽ�T�T#fF��L3������֨p`�M6�ɕԱvʜ��ŋ1 O��H�*dj:U��n"���`���s��O�����z��\+�5(�M�F�\�H�F�(��ԩ��r�4��Ѐ�]6n|�Ս�X����-��_G�����������-s��`�?Wc]3�Ny������:�@LIks�&�Q:��XP<	�b�-x��sE*5)�hL��fYe��[Y���:md��xD��}�oPJ-���j��k�^f���3o��f9�mo'�"���l� 9�HY��# ��eG��&��f�8��f�`��$���f�?��/䥗^�k���A����"m�s�?.�,�����=�>w.���D�U
�c��Xr4���<�L[3��.�
45��#Fґ�j��Sj<��OO� Rp�~��_�	����#�o3ʎxq��&h!� ��NT�����7`< { �x�i\]j�CP���,�1�g0����U�S�� �]v0��_�դ c��R|V56k�s��� ӥ��&%#/�OR�}r��F9N�A����+|�y?���٬۰�Y5=L'�mFg�x<��햐�s��,&	��j�������\DK&�7��'ا~#���E��  ��?���(x�����{�H2�"��4+B.I�2U�Afu)����bn��̦,�A{Q���� ���Wѯ/�qP��4�:	��Z8�j��Xu���c����O�N螨�ϱd@�T�<K��pY��L�,pұ�IE�,U�b�J���ת����n��r�;&0 7��2XiX��n���ep,z<g�"����dJ^�w6�=�C(E��V��μ8m]�V�������"R��"�}�z 0{^�<��y�����tR�us.<�0ܿW�}�U�hj�%sȤ�`��\�0P@;�����@�WF&'��o�w�y����ь?�Yh�)%Z���[:tn����n9
�,��L5�����U̖h��mg5�Oy��e�VШ���I�5������SD��F륩�Z7j�m��xӎ�-D�á�y��k%��y}��ֵ]Zԙϟ�!��~�V,S'1A���5�IBؖ�V���8@����1�4�0�Z�t�ɨjO��UF�s����yS����[dv	ֲ֦��(G��=�Sԁ��,u;wn7����+4�Æq �_1G���s�
�;J�.�㫯�*g�u#�m�����?]�	���?��>�/ o��C}�B�;�p~�c�=&��2o�|*T8�s��.Y�x��Èt��/�`8#`�|��׃�
��UEtx�l2@d3��2d�ܣł-#۬�&V�N�\�[+t0V��R��8I�A|��l�\�ك�c�!�`e���i#y���.�|���q���3�c�K�h��@�Se��eey���Ԥ	����خ�,��޺����B�l2[(����XA�D��
����D�ϼO��lC�rN�G�S�j�I������h�Z�ͬ�׊�`���X}��5�n��,C�#�IN��Ѳ1(o �B�PAO�,`vC1=5�f�e�l&��ud �a��o�(QÁ��.��=�7X�|�+h0�@��ɑc�#q���S|_�7�GSDy)8湃�-��{�������@2`�G��Ũ2�OTq�#��.�L��e��O�����X'��=Ҡ��!�*.��8Ro�I��	�M� �X`" ��@��Z �yMۇ|��py<�y�Y����L1 x�(��l`+4T7���m���: �b�� �����T���A�n=H�`������^|zz��1��*&�#Ժv|e�=n�p�e� �A�xR3�̀��Z-#M��G��7�����R�khlT��iiTc�r��d�
��6��"�&Ub0�c)5���'#&?���ǈ�q~�\�`6�q��#j�TI�O���de|����M��!�	��"(�=+A����!���%O?�4�·5A�)����sȏ�gg'y�Wq�tn~Mҹi蓋>�!9�S��5�˼�v��k^��aF3˖�V����/Rz,���3��,���ԂΙ2z("�3�(���^p�5ǓAxr��'��Ed߾=�_�\v��A������4����S�C~ء��fX�k�d�2�cٜ`P���
 N}��E�/��vtt��с;Ne����'��6�ܐ郌Ƌ�4���h�G�661n�KE��(^ĳ�S&�#9PԖɊ��ٷ�h@G�˔0��&�'���B~����I C@��`��O�(Y��y<3�qz��(T��bplȀόh�'tok�<�8V�� �'�I,�=�hƀŴ�<�,��	U�@�ᐔ�QN8����/#�b���ދQ�$P�M	U�Q9	���rO��`Fa�������\���w<;W\	����C;*e�N��@2 *��R��Q��k���sL��ˌ��-���pHP�C�'b�S�W���l����^`E�bM
P"����rh�� �C���f=�Ӛ8��}�-�ƀ���KT���(z��2 t�s�]�w�m=�w ���ho`���dtlXb��\��ɑai��&��<�m�hg�Z�˴�F����VC�k�:��#,�ψ;�,���R�f�\@`���}Ҧ�n�M��`��R캤c�o)�m�2�ʻ���R��z�9t�Yͺ=j�g��Y' ~ݤsϑ�-���D��Fh,G���! �V_##��^EN��@�VS���C'�J0��KJm�F�y�-�ɔ���+S�Sf�7�G����FPo�+���V7��\�L�z�q���Q����x7J�K"�	u�,���Kb�D�Tck�̝?_|��Y�qk� ��ꁍ�o��᤼�n��M��2�/J=����m�e��.��N9���D,���X2-?��lX��fm����x�w�N]�:7P���x��e[��z؆�qhww�Q[[���Z��CY$g��t9�����x�I���S�/���ɽ.V�Dײ*ed��QG�E�aJ�4;�ƒ�����bQ�NO���a���~�Zv, �:�n��yi Ɠ���z�*Y�a�<���lܴ����ٳȳNv9��F���.^�b�1�n�ҥ���F���p#C�%���eւ���|F�,zQ�?!����ό� �G�c.aʛ��ZZ[��r|R��������o�۱�j����a�{5\e��h�e`�L�7�.�����#��3�m	|�lc<G�P���iР���X`�B
���L3��Q�>�,�ů(K|T��%�� Z�� �i��뮫��J�eF�ݠܥR&G�5F�h��"�>sؿ#CCl� ����7���Ag>s���'��xn߾��Q���V��%�)�d��"�z��SB��q�S�3H�S� ����:��ǀ� 9��)����iK���L9lYX�m l��՚�&��[�����4@�?uc]=m�	&�
��[�PK;e0/F���M�(^P���L��$`�B�Vp�/���e������1�U�m��lm���^9�mo����i��^�����N��3�~ �:��C�yfo���aY�&�<�G�'�1 eQ-�ހ-jh��~'�qٴ�����x����#1e��>�v���R���z]t�����s�d�!P������2���!��<W�_�"���t�&yHZj�қ���2��r�*����s�c7�1=t�")Q���B9q�Ӡ ���m��n�������/�NbRwT3�,4����w�Z5��P�hʏ>����Ñ1��� ��!��=�Iҙ���j�C&�Z<����.�75x��W��i�h\d�^W�%��=x�I�y�ʱ�M��G,�@'*C#��xg��1��9��Qk��W��`�>u �D��t�L����C�p�:y�͑���b��Q��Y9P��jթ�4���H�/�/"!�emK �w3Ռò#S*����"t������hF� YS[E����H۝����}��[Zi'���c����A�72�����y���A� ���D�I���Ӑ7j�:M%B|��_\)ɕM��7�N�瞗�:v����dx(;z,'9j�� ,ت��?z"mj��I��0�e.r�I���?ʓ(���Iq�z��hmk�{g�O��ֲ�y+�f�"�1n��7`���㰼(�dG���0�����S R��������ՈիW�\a]!���E��=Ҫ�i�R��-z��<�Y�ԛ	L`��ܰɩ��uuI��y�9�
��[�2�?�^�ͤ��7�[��9���������	o'X��c1�ۙ�5��?�������wɢE�䥗^�'5@�({�_*�x��7�
�>����һ�(/�����-^,��[�mN���6��_լ6,5&_�N�k�����G��{�4γu}c��$5#޶��#��e_9��� ؅@�1}��&h�77��~x�|�S����T��ȁ���zvA�}���]~}<'|M����h4L����-�/��+�9蓏�����O:Y�bq��뮻�����z?Y,w�qG�m�>�d@���d�ø��%�"{����ADz٥�6(zzY�JN��u�1��|FZ[�e��3�]G����/>��C�}�{B ��v_��� �応���z�~ܰJ��Fxޒn�Y2�U�eD�j�jB2�;(�RT�j4}P��,����ҵ�-�,�Q������dVbԋ���f�@�2��l���@��)�qe���<�J�&)r�$ U7=L�-������g{H �v"ƅ<�و�����,;@ ٮ�d�΢t�m�֦�,�h�ͯo��;%^� �c�dhxJ�-Z&s�-�J���HMm�n:i�h��Pǜ��'�@�^h:ݭٮF��d׃Ý���_U#1$s�g˳�>#{����WJ8�QI29���9J�~н���t8d�e&����s�%l(ȍs.}J�ғ�<]�62r�K�8���׎>�����ǲ|�r�����-���g���Y����!X�g*mʖ��Ȋ#����!���V����
\Dg�i75�p�P��3a���,?�;�����0Cx�;W^)��匌�w1w�g��&h;1���K�I[�a�נa:3%�g3ڰ~%�ϱ�'��^[/O<�� �R�2d��Yuv���Zr�"����/� ^pp�w�lQg��˯�\�R-N�� ���L���J��{�gQ
��$'{��*��Mk0QW[ǵZ���_�琱����t�[5S	�?��:�nI�����S,���T/'�|�|�}�`eĢ��5C��o�M����B0d�M��W_v��!S�i���_s-n��&:�o|�r�9gɶm���ՠ(D��(n�Z\g��1��㘵O�D���{ｗ������_��đP�'��
����"�A�=��9�#�V,�˾�9�˥�^J�X��2�_�Sʼ�5�\c4�>�3�o�E��g�{Zf�w��d����d�Kk�-GEb�+u�s� �vD�-qc�ߩ��X�CR�imu����3��w�a^~y�lԵOi�̬��,�QCp�e�IjPp�i��ӟ%t]���~�ߧ��*�A`���?S��G��=��c��_�"�?��_����pO���Pپs���!G�ͳ� ���wH���&�w�L�?�����Y�|j��s�&T�B�NK���`�|�;ߑ��[6n\/{՞a���j�J�ʗ/�K�>�=}��˰���m���*���t�8'�5��}j���]&\:_�P�]dVV-[*�-m����h���9MR2Ƽ��h���475ʋ/� ���w4��t��e��BP0�e}rd�X������������ذ��FT�_���@@�4�=�����:R8�;�h5AQ�e\[�Ze��%���N9Y�unֈԑ��{�~�f�u��Ï�$1�r�wD��̙�$��UR7=/��B�m�8<�Ǉe�������P�B[Z�t��40�(k_y�3�E�xC�}�Q#�m}i�ٵs���T��v�~����~�cP�-���n��`�Z)*�13�jqQ�~���塇b|޼yҥ���@�JT#k���P2�U� zTj�aܰa�l�����30���H�,��"W�eVF��c�Lf�F�MT�rU�ܙX\;��u�ֵ���: `^C��H�1���h�[7P� ����挔��M�=g�B���Oo�A.X,��C�P@��у{��'���<��_�>���[o�_��K��?>����ߧ�*id5�LO����;w����?�m�71{���~�������IN��<�5׾��4�nrex� ׏�
��oK����>�ӦJ��=�ϹxL\T��yAR�'?�V־�F~��1(C�+_2�k7����_���g�Rz낾���K��}��v�mr��,��|�袋�����,U���}O.�����t����A���M�|I������gk0�����+RԵzL���?�Ij�,�cϺ�]5�������pV]}=��{���_.��B}�4��?��s�d��-ë���z7Է��.��|�s�'��]�M����}�5@�կ~%����ѩ�$*��ό�cv��m�|�����_�y�;�� /��G�ьp"�{?��|�#���`[�
]��Q�L����>Dн,`X�R$'zFP���C���X��e˖�W��Uͪ�����_��׽�L����ˬ��k��]�ws�As<�)�v2z��� B���a&�����O|�����@��Na�#ீ�<Ka0~�� v��}�Z�(��V�O�d�Ο�}@�S��O���3��#�w���Ϻ��[$Qe��`��ݡg
"H��Ge��C4�X �>���Ҹ��a#�bH�K�cpYof����\��Ԕ��޻g�̭���-���Tʅi�QJF�Q��A�9G	����������i��4�R���P�Pf�U�|��Fs�0� �@V51��*����ѫB6���5�(/8��B�4V1����f����r�����1[������E����lwL?b�F�5*��Y�!�g$���>p�:Č�I�-���+/����ʦW�1;��ye��O<Y�;+�Z��������h�Pm�*5U��`L���dLdfm>s��.Ģafژu5�X%f�6�&�5��/�҈�V�wM`�����@f53��0���N�r��2�2�%~͘�y=41��X�w�~׀�
9�� �Mi�����0:�F�UW]������[����Js��f}8h8_M�$���9���e����=��E��ׅ9V����*P�d��#�=ʯW_}�<�����7�,�xT�uŷ��w�Et�-�_/us�13��f"�q�n��/_|��5s<���5c���j�%����DD�}��`�mָc�X�Bn��w�g��܎v^+�lQ�mj���;��>9�ثh4����1g?5���]�A�ClD��#C��}�N��_x@�$)��7#�(IDP�����ɬ��c�=!�~�y�/����&Y}�ѲJ�;Z8�ࠈ}?N4 �mhd�]W�H�u6l50�:�v�j`���4g�0��=�k���3c��o���@�'���`��=�K��o��o�}�=_�u�Y���7�ɶ�dr_�~� �M�6����k������?�C`���:����_�n�Y��x\m���/Ӟ�-��SO��7Ƞ>������9�m��)�V�p��Ls��[z(�������o]!'�x�|�S���.2��~��u�=l����u��cK�"��'~��Z�
��S�.���Xi��k��G�'��_�t�f��0KG<졋a��E6�� W\�=����o���7(����=��s|nhI����`��	�r�t�a��>� �؛����d��ax\���N�GǓ���h��6 6I}��r�s����4���HW�@�i*/�	
Nj��������|�?}�a����<6�N@�WPN� 4xv$I�5HT2�Ǎ��`��p�J�Q��jQ�4a� �\:A��<d��,Za�$��P�C�'�~L�D�&r4�3�4rvV�\N��p�R�ΏūF�����S@��M$%�0�ƶ�6^ٻ��5�YP���',����=ʡ����>��%�Ռ�J!ʴS�$b�}ON���|�C����ww����VЊU+�\q��;2��)�ca�q_]#��P#�����(g;��7��-=��{����A�˃ %a�T����@���Հ��� �cf���� �*�2���=����k�q��\8@H�B��}��L�RB����ҬN|���LA2�?�q�4/>�����,�\+J�p�pX�}�r�f7�`�ա�٭����	�� �k��Ș�wp�1^y���Q_}��.�uBv�'a2�Vc�%����	8��=�F��Z��E��Z@CvQб��s�� ���T.cK��r�;ϒ�n��̛�Č-M�`�3���M �@���L������o��죲D������a��k�54:"�K���f����z**wP�ۼe�|���t}��ϓ�%�SN=Mv�ک~!dHH�E�L+�q
tT��II����b㨾5��vG1#�`�|�^��ڗ_�3O&'�T�P����3��}B�Մ�}�"��on�h��SO=�^0�Vd���P��GǆyޑXxt���	VD�L�@S�ԟ���%�v�I�X/d�U���gm�F���z��^.������̡$��נf�HB���8%�xl%�ـ6AF��^����[�n��r�O��g������O��M�=����߶}�<��c��A��=1�Y�e������Cs�d^g0e�B5R9*R ���k1k
.b	��� U?:��C6�R�z栄XY���W\q�چ�Sv�*w��z�>���g?��M>�p�o�AZq�[����7����+O��&}M����޷H���en��N	g���Ş48"�F�$ЇڢY�@i@7X��l ������ ��#%���-�~����0��n���p��N�I5"詸R�@?���X��l��+�4��"A^/gs=�e���imk�Q����i�T������&�-H,�W� :�Ň�����-t���AW#�}w��hPP$o6������@�F�+�Եx����d��ץuv+�y��
a42�N�����-�돲^p�9���^�#6t��J
���T�5(H^l�1y ��8uj�i���J�=!J�0*��+�;��=�t\����0��>�N�ȹ�F:1��A�j��򶷽� ���r�f{��ի���^�١��/�Q�cP� a�q/ ݐ�W3�}��T�q<��5�������Ge�dH�*�7�IF4 
{_�f�p����;���xk5�>���%ґ������'�|ZV|�R��G>"k׮Uc_'��9��������4��W&g�l0�	�Q��@={X�=�=�%�0jh5�� ���~ �J�f=�"��0s��{�a��'?)G�Z��#�"��D�Z�>�X�6_����"�(�X(kyI���˚�{�[嚟�����3�b���O��Fj��<�W��c(h��`	Z��\��կ�ͷ�� �C���|�I򽫮���sz���; 2!��P��� ��\���6ȱgX,� ��O��E���� Y?� �@�޵�Kz�C�2&G��# �*e꾁~����V'x���p]v�ed!�B��6>�����9K�_��d��]s�5�Z׽Z����6y�'�]�{��u�9r�]w�g������í�>��Q!����׽&��r�\���j��ΊF@��0��㣲��`B�����ZD�S^�����X�:�:���;��}���}�@ �l^���Q���~��r���~��h!����w���]�M��6�-������:.	�<��]�S��9��Hm8*g��-#P�[�y`4p]v=\��>�q��,|�C���e2=�g�O���oI���~�#�㟗h��-C#cR��,)��=9;go�t���3_�:8���4z���lcZ4	�?��nl�pՐ�߳���l<Q-�7��2)j�8�r� ��������<�SC8cY�`�#�"�Ñp����r���P�A�q\�U"��ل^C�Ω�p��@�l����R�l��)�ã�+D���7"��Tth�1��['*�_�)���½#jO����%��:�!���Y�h1f�e���/��{vHc{�E=t�G}�<��qS2��*嘱��`��+�{�ctK�.��l���,��U_���ո|줜�<�n�Θ��k*M��〚ga�`��(Rv�d�p�x_hR#0�ԧ?��3Ͻ O>��f�r�g�u��(.��G��s�gy��3ϖ���;����3p��{�0����c%��UG��O�4ȗ~��w��{-���ԟ�c�:�`�۫5�6�0p�.;�;�-5 [�����%���	�kh����c�������'��w�w�+���ƴQ3��d�^�O~�9��K"��]�(�y.Wd��4����q�8�Tt�UuR�$4�A���ñ`��	Y��wܡ�|��}��}��[[SO��m[��&�L;5��a.��N�@`���� g�~��VU�-��=���R�L���#�YF)�JfG3O�[D���R���ģ?��|���uM���[@�/=�S�`��^C������͙83�J�x����>� �K���^fn轖��0�YE�>�hXKh����47�ľg�>����ʑˏ��_~ٌ�����c�>)�Ījm�E�ԅ& *Bp�2������:[�lbK
�Gu�Ƹw����o1@���n@u��(sj��)�����`֨��]���?�*����$�nū�h��<���_4!�nج�{J��̓*����M�~	ɕW}G����^߯�i�<��"� �«c�B�S{�q���h'�N\�cO<ì;Q�� �d� ��$P甮�C�}@2z�12H�X��%���aD0 �g:�L6��AΖ�g��W��X�g#px��qM~f�n���)yE�h^�[г?���B�R�X�n��|��u��$��9t@Q$7�FiްPg�?V��H�LdEz�S�}�~���j��)��vgFѣ۷���c�[I&;)Sz�XJ�?(�#����lbU��+�G��BQ�/у�HQ8�Z�񢿅�w`�Y:�:Ȃѻ��C�	�8� H
z4H@�/�}C���.�<�X9��p,L͞L�F�Wc�e��CUR�8[��=j�։'Ҭ���K�|��S�]�C�%�����ݿ���j�5�a�5��&���q�0c���rk�,��� $-8�j0w���N�b�������I Y��Q�_� ��9\"�Mf�
w�ed9���S/�����L�g�{p���$c�ɐ(�������K����O~���I�s�.
+��w@��,�cs�x���):`�aTq[;_���z�|����ڳ��풯��н:�L�14����/����z�PP���A�R�J���NP�)���h�e��n׮.�x��Y�3d2�*���]3��o�Ev-����=]�я�T���- P��
|*h��h||�k��?>�1�_�Z�A��c�&]n�U-(��a 8"��(��~�5O|]s��tO��s�3�y~�GѪ�uI��W��֛oe�<�A�-��4s���,1o�B�Ώ���r�C��������oZ�Tz�e����D��#\?�T�����d�s�2��9�+����A� ��+��Ї1{/b&�&���Z��18�	=�~�R�982.���[Z�e`p���EK%Z@&됴X�2Tނ!b��۲�s;�X���=o��-��3�ɟ���Ĩn��>Ӥ50T�^S��8-�̴0����i�:-]H�b=jKӚ	g��Y��.p���ڽGvl�����XM�K�C�<�����ZE��I*�J�;��h����߀Y{z��k�����:V�h��NW�̫����9p��h ��7�hz�LV��N�LL�R�r> ��XF� ��Й��r(H �����2���%�Q�"c�æ0��g��I�d*��lD�*h�K�/��]�����g�
 �A��1����VIM�"���=�2:��YMU���M��C�ʂ�6�n�-�?��BM���,�^_߹����{�8.�#��K �a��(�>歲s�nyi�$+q�Q�ʓ�F��^�)�a�,$f���!+Cu =��FrCãv��?{���1.�r�̝�PB�2�l���$��-�-_)K��W�8&�}Z�����W��%Gɍ7�!!��;ϑ'�l�Lx��H�F�ý�6,1	�5<>���=@C'}�C2��M����� �CF�.�]3��p*.���c.�n� ?��sv����]�Q��V��������a0����̟���\zTD�$h��R@v���-��>��/��l��Y88r�Y/��Rin�c�}f*��=w^̂�`�(Q?������*"z m�N�#j��d�~���D�ׇ �\��^Ȥ���a��Lv;5ܤV���a��GaZ�4�m�;G�43�>+��9�ʊ��a.���Ѡw�}�5G3�Y��㏗�� ��G�ȣOH�� 3�\� ���h`�F�����$�AI��7��)�,�u�ev����z����@����Mj���/}Q�z�ye��A�Kb3v����f8af�S���~���1_�Niv�LD=F��I=�-1�B�Q*DOy=��(����\��E�PQpw��[d�� 1}(���^{�EG��ɶ�3�jвo�.9����+W�ş�D�����Բ�1�j�NBʔ��U�p�H.Z�̕��i�7P�x��G�e�l�i�7W6o}�<
�i�>)��Ñ]��� j�"�m�t�@zi`(��9u`~��#��2'?A�IN��y��t�鳬����7�3�c�C5`�H�9ZA�d�p�8�H��[��O�'9��� G�~�	�M@���ր��F���)iҲ� ��_t�<���b�<���}v�b��Ǽ:^>�?�L�GG�W8���{߻B��I��5ײ�9�R �BU�aX��O���C�-���K��}��cX�zk0��	't#��24�'����l_4WZk�r�.�: FFF����Q����8^���q��v�<�ee]��s4@#�`M[/k���H^�!��Y����I�A̶��"F@@u�h?���'L����-��<0](��u6�Ȝ���D��c>Q�૿�NHy�Ȋ凓m��y웭}�u��/���VJj� S������S��:S,�ȼ��:61l����w��ꈾϸt��=�-�����;��ӟŜ%���Y���>�}Z�\��XH���X#g*j�|	�u" �@��1����x�4��Cw,��_	H�7�m*Y�{��9{��`�`� �2���GЅg����+V�)�/{���q�O�{��0���'�̱P9����k��7��������B0�����o����N9����sϥN�]����+���X���u��$�	�D����T��� �ͼ9�[j<�؇Ϩs��]6�f�� '���캭���c�R=�-����J2t�Qi&<o�r�������6��� �'OF���P̴Ur����Z�`�4��C~�yr�;ޡ��"���sɻ����~Vv��Kp_����& D٧Z� �N�{�6J˾Gܫ��q��8�J`@A�Y]r�2�ajz��\7 �^�~o
(fu�'�Kg�X�'��Gf*t��f:X��A��ey�.�e��̳BP���4*�w�H�@���Ի�j(�g����Mr�}�˿}�By�;ϖg�����G~*M]
йs��\�R�Qdj"�2(��ԧd��L(���:�J�а����W�.Ct~K �s�5@�ǥ��躡�)��d��Ӡ>��=bE��TL�*C04v�����~I:;�˃���$4��)ź�4hEU2͉�V.���=D�C)[�Q�mD���&���̦hZv�Rh�w��Ǥ�[f�~�W�*g�u����Z=��|A���������<&��؟\� ����cwM?��Ҩ�qQVyP�O#�t��#�S4m4�����8�@9��C��/���0p�����a�L%'�^���#���@Ü�*�P1:����yQ7C����q�~B�5���2Ң�xZz4Kh���'(��B���9;��L3SG���o@����O���3��`�B��hs�T���@��yFd0�6��_vl�#�씑�YP2K�Au��%�⾇#{��Q�վ@z�%l�$�-���ʒe�k�Q�DuT�j���P4D�ôF���xO�d2���`#�7��G�����a���0��D�%J���ۀ�Ȍ��/8\�N���9��0077l2m��%."޼w�)VF���p3ms���4Jn����X{�;�:��h-<��\�9��a��ߣk<��[,��:��	p �g��b[ˎ]��G?��s� +br`F�a<�~�s?����7��?l�r�ʻ����[����w��Z6n�J.��!��������[��V��������İ�]��o��fٶu��5��̼��Qڬ�6�����[��)���C�"�u�������Ih�IP�:F���{z͋k��w�/�.Y,�_�	%"�s�3�:�4K�uG���k��P$�);���@�l�I���F�� ޜ��eÖm2�z'�z����jCcKԵ�@&5�(���u�����ydbD�K�`}���5��e���:F��<���z��(*j���'Sz���c�PA����5h8�dO.{��{���g���G ���f�	�z�p���(�9�{�b��� ����Y�CFخKj����.���!�K�In*#����5����ߞ���1_.p��W]C�MX���Fpz�����ЬVI�Gߩ` eꌋ(wQ��qh����dP(� �+�{_4Q��A�N=ni�o�Sj���x�y���k^0��{���#�Ŵ��sy3��&�c2�IpPH��յ5���Ya]�b3��%���?���
?K/�m�]r�ѫ��o~M���ˬ�P�<��H��8�裒&H�H���ԵN'u��'����K�K8�5�+{X+���7K���U��=A��� R�=ZH�y#26�&�b�C,����L0k�����-��f��Y�Y���-}���I��Dm���v9|�rY|�!r͏~,�P�|��_���[��#�S���T���h�bgLk���#��;N};�U�H��_��׺	3r���Q�p �/!"����d8R#�Cc��*�}Z3̎y(��F��8��9~�hE�xFR�]"�7D$�N��e���PE�ǦL&vđ�Ɂ��eˆ��ŋ?-+��53��f&F��PNkTif�á��p�2���:�pл⼭��YO4� 5��sT`48�v�qMYyN
1P2��uLZ���>6Թ�h�G#���'֔s��sp�)�F����l_�B�p��pO��Cj�{0��YD�f�; q��)��<��Zin��׭��ǭ��F3�(��I�\:�	����2�� ���K�K}K�L4;m��������-ݽ}��o��:$Ḓ�YO>���rڳ�s�#��o���� x�#A������ݺ�S"���~p�~v��X� x��LN��x�����S)����b�a���׾�"��܀e �P�����430#8ҥ��2"z���_���A������=P���C(���w�iPUӵ��_)?��'���X�g8���P�Ek
�5�M�ՙ<I���ߑ�a|TV�Z�j�G>�Y
"5�5p��@��PӁS�S���j@^�o@��Ɓ0������cU���ƒcIc �m�J]v\vX���@АH�[/韍��)_�UU��1D `����u ��
Ջ4��u-ܟ��ɪ6���zQ,��E� D�	/�\+8b�i�tgk0~�y�ʷ��#J�&���kT+�����Zl% h	�\���z�z��L���� ��^uYw�ߤ`5�x�%'ALfk`�s��EPC ��ł�7r���愃*[3iac'V��@�69��Q�4A ��Y����X< ��v�~�\Y�n�465�Рy���GW���Oq|�1^���$�U�Y}��_��-��?�Nbz�M	M,���?(�{�|�S����Kٱw�}QL�Ʊ�9a�{+r�@ ������p/�k8<@d	j(Z�{�� �B�%5�L٨�ԱD5�-������O��6�BS⨱n[p�'����%K�-=x>�4U�j��:�40<!O?���O�P���'��~�LFFǙ���p����&Fsш:B�����"h���R4Z%ɉIl�c�Sup8ʕ-xDm)a�R_Ck�A{�0�a�BL��zI�\ٱ{�Lp�D!��uj�2a.Ԓ/��Y��Zb���^�����+%z�����vI���ׂ>�}qP��k��oE���i�G@�l�0��ZєK֔�L�+F	�1��3@�\�Ku� ��ei8]�w���i�.�����ia�,�T0�����nnn�1��%����M��g���er�1G˪�G�+��'�$+��U@D�NX��	�գe��` �^]�Ǚ��t�igA���G�
��G���	![����]%~�C$������i��a)��	�x��CG%;2��K���~��'q.v@�]�C2enu���k�1G*\�(OC�j߁n�J"����!EE�S�REI�m� p(���~��mۤ����v��9��������J%���s�;zݸ��[�r��ҡ�n�����l�/KΜ�Q!�(�+�Z)
y+��`�e}3h[%��1Y?�˰�n*�֩3#9�h�N~��e��x���^��h��ƂSC�j���v�|�c���}\�m�4���$@�T��5��y �"p@EN����;�zP�8�ly��5<C� �����Q�Bok�8^^�܂1���Uv���k����l�|��op����<�y&+�Y���x�͙u*�P��rL�ZU��5x����ݺ�Z��k���g�u��Ĥ��߾L��_ɆM���Ε�&_���4����{`�V�\�}�jS�>6:� �������o}Ku��5�X�A<�#Uu�c��Ǘa��s����z�9�b�s�^�!��,�N�FӼTr�����NF��f�e�0&�x���F���q =,�K0��LZ�#�ҠQq���_~��]�=�}$5;? �h�t���$
��r��}�">0��`���^~����%1u20��bV�d�:�Z��碟��V,�Umz�$n�H����^f4҈VM~��` �x�ٻ�K3�i��m��n�dP|e�u�@�SB4Ѝ���Ɨ��UEÂ�H�:�|��7><8d2p,&�'i(\`]��0��2Ǵ�OG�_˨:�10�Y 
����3z�p��=W����΀A�Z�=S<�'<ZT;�rpW����k����@���ij��4�~�2w�|Y�d�<������~F���>��p�ҩ���u��u��5�w�yr�m�Șf�>x&S#���_���<p�_e"9����=66��?�u��n���q��q��e����r蜻'���$qDP	�
"�+⺺�U(�����k`]VTDP�40L�9uա��½��<�U�=�������ҡS�����9�G��[���c R"z W9��\��cG1y�de�z�$moO���,�3C4�<��g�o��˿>�P�͊J����ȑ�� �j�WV鬾�X۬m�H�|�wư���%�L�Y^�'^6�������L�=p�B�(�=���X��$1�1���/��ΰ�7��$/3�������|��2ޓ]���?��w�9�qF��|�-��Gmۓ{e�7���jEP9�\�R��	�%j�H��=_��7�0��"ӿg�rT��w�߯�	$��ݣk)jIی���8�"qN���Q��9�2Կ7Vm�1O?�r��{�׎�;�y�n\������oGBl-� �������H������׸ۧ6�wқ��VL�(20�$�o�/���܃��>��X/A��W�c��y:��TT>[��C0EW����r+�~����?�C���{K����_ ɉ��~���%{$!�E\[(��c��g��n�X���?�?>��:�A�F]Ɇ�X�R�n.S��9y��,����1� @�;0É��r%K
�l���IfL��:#9I��}��m��;��MDk0wQF��	JFZS��y�b��i��
�5��������۷�sdO�E��؇"*����̵MnEu]���uvti�gWU�(�
=�)s�f�#:t�b�I/84�F�de��m5ڰ͢��eY��5ω��]mu�>��M��#�G]z����?Ѕ`ĕ�pP��)fe�=�Wa���J��Rd��_��_7�`����Wͬ�AK�,q���[3.q��;5Q�<N:_��ɊE'�@ǭ�Q^��/��$Adk��g����󘉫��<��Q	ܘ���,�zx����5_z�i��]�x�ʼ�v���_^�7n��Y������@#���&�޿�o��?|�X�d���deM-\�P�uw��x��?c����S����gFLo�JqTjc�K�1I�Ԡr��@8�r��j�<~���"��c�&*d�t�����ã�&�
LjF�;�1A��Qr4���� `BNT\���u������p��E��G��OMr� �ؚ��N(�Y�dM}�o����5h�Ԇ	fڻ:��	>T
�������h���d��V?�Κm�������Mo�[zO�R�}�Wx�r�d�{���r�vW�)�����8���&[Հ�����{�v��T-L��=���mU$Uu��߄'���f�~!`�z�ʝ�*�1�����|�[�z�L����iξ+@1U�Aτz���Q��0>Gן	��^��Ai�ft��O�)R�npTM=a��T��Y���F��	��3zh�����H�m%�o��װq�+�ɞ�S#���T�5(u1שS}1�h��pp��q�W��/}��6}�j�O�๪*�;��w������ZUU�19aR��!�x7dZ�5羹���СK�`�+`� 3�ͮU��,��r���.�,sr������#�YFu�9��D��(��t�Nޕ̹B��^qln.�jV��v�D6>���CSC�b��y���𮫯d�U+�T3���q$�puu|���ó�OS�n������O���x��
|1D89da���<|!ok�͂A��a���8��SZQ��"3܉�������eTk��u%Ӭ�|+T0(Ɯ�e�hijՑ���Nc}�)˔Ɋ�N���G?R֧d�)�ssL�}8c����ʘپ�=�Q�)F���k}R::q:i��?��O'��3X�������]g�=�X��]9�)�#N��~(p���8?�����:�?R�e�mr<Tt��G?���
<��$�\�S�4�km�����%!eO?�t9�e�<�ȣX��jmC�>������9�Ք}pTR�������8.N�pm�%��݀�*l��2��̨GF��HR>��1�	DC1�<�
ò�G������&	L?��KfR\S=�G�u׏�����[�09:6��i����s8֖�9u�Gfo�!g�?����U�/58�%E2�ɐ��W9�~�H�"_��#癕�0 f`�z��R���J�c�E�|;�&����j���]��[Fn�߹�V��_G��S,g��۸`����pDs��HS2ƾ��q
��B_^�w�HB$�8��|���
c�7
j��`E��Bes�����y���eD��)���N]�W�,��ZŌݯ�Ԓ�b�V�*���txpHlVѴ���,��-^xV��&(2�"&		?�(���X�\��[���{��ս����\�/5��-*�����y��	��6�N��5k�/���K7s�4��I�{?��?��$]��$����rՠ�`*���t� ���Ρ�ŷ%�K��n��Ѝ譊 �/(�e���hE� �ő��'�]�{,J>�9ڏ��G����t�;��O�`��dˍ�����@�B��itN>i>�\y��>�>�tC�T��d�A�	���|c����X0g�fC3$<��g�'���DrE�s�r���64�4�)��}:qn������� �M94�Tcw�>���s�75:���l~��A\á�r�d�Uⴚ�Y3�fvM&5���#�se��9M�7�90{f�94��`�̆�Y�y0{fߜ΃�3�y�i�h٘��>����}��9�Q,[�L:�d���gP��le���@14��3��&/��D���e��~u���/��R	:�1�y��<���r��J�qC*l�B�����r��z����g圞Ew�1CS+�5)AgV��k����DL��K磉�m��k���
��9d��dQ�'B*y7o��5#p������Nl�*�{�ZɲJ	�/<��J��ݥY|8l�ˊ,��o��n?�%n"�����T�1�m�st��f�T���GK�$;��>Q���K�;{�J�C��Ɉs��t4T+��Y���~,�}u�Ô�/���4�E�P���J�� �:���#���JoY���g���-u���^�\�K�U� �c�ԃc�M�=�C��ʺ��b��*�u2�!:ݵC��
f�]��4��� �������N����c��;P^}(�X��^K"�T�Q�k�|�̵�ql��O����K�z̖_;q�}n��?�a��T�$!׆�oR�-�W\P�68bB�dߑDR7�F�Ł�iHTW��ѹ ���^�B����?���oÇo�;<��#x��ǵ�Ñłe@����^�0Y�J6���ϡ�~ϛ�}5���y
Vi!@��h���&��\���DYؑ��� ��04Ѝ���4��ni��ކ��c���a�n�p�؇G18"%Q�1	eq0�c�8�Q�f0kr"V��w��������,h�hX��b9�F��Y8�������ڶ�f��s	�A�Ēj�G�Қ��+��(��~x�b^'���8���;K�����E�$	�LI��[4�*GNAMD�s����я:q�\�$Ka�_���S��С#�9�$�dV��ݥ+tn�P��N[�N�y�c�&Ӳ��K�>ȍ����ϥ���{��0K��'���6f�4�wK�,(g2tc8HB� �����+�&��h\�ro˵d�r�����g֠e�$,����dťx��?`�������a�D輇�j����s�M%�<$�8e_M*�i���G0a� &y�,$�mV�H�9YOpY�^�d�fG��#0�D*Ӊ�U(��Ȍ�x@/*��za�y=�����x�k]t�CA�1�Jո��?��v,.���X����\hϒ���W��u7|��%]��Sp��?��dg�8C^�4��h�ҽv���;T�;�kwn"j����,� �����r���6.�����<�s�^Vh����}���ݽ��PF�,�g�z`<�����J��Xq�=�wd�SB%jλ��3� �K���>f?��j��19N�:9��j�z�uתwPv%nz�*��UY�dt��y�SP,F�x=J�������#�:`d0���^߻t\�'��Œ�[va�_���0���t��c3p�=��$����Ν�����۶nW>;�(���O=����z%�� �E�_4ɉ�-�Ѝ��@C}�~� [Z����6�:z�G)��j���ǡ��Ϗ�:�t���[�W�P"k�id���+:U�N�B�С��f��7W$m�w��}̡���]��ꚧ��T����L?jB�O�ԨF{����O���?=�2c4��&���Tg�Rd{<FB���@F� ��d�A�a�������ںJ�E�U���%���
�m���cd�M"��9R	�$h	�Q�OTz��h�q�)Ji�(��ß�&碹�QБ�%s�r|%SO�@X2�Q	"bu	�3)�89n���}�g͞������#
?p#�ӝ�1���\Qe kt�$eQ�ב�f�t���i����zH�qR�r��sb�B�s��ז����?��� ����q��Y2��W�O �F��R,����f��I;Z][�dRΘ�x�c������ŋq�Ec��X�n�����v���ͪ���!����vu����	�:P��q.yNALL���b���V�e-V��{�a�tu��k�EU]-�؃�p�y�d($�q�Q	W>� 
�3���9KGAgN�\���� 5ȶ�|��N�o��rFq,*{������~��?}�<�V-�1}��7Q��p`�+��.ߓ:S1+�k�e�>��������T�uP}��d3T���0NO���f���alt	|��'{��bO�Բ�6��P����(}��bO(ϪK_����1>5�qT����b���l��Y{�1��^�o�iy񀇘g&ȪaXEA�eWNw��ۀ�U��P$�!�F�?� ��0і� � G1&`l�T����h�9����L%���Q͚�L�m\s�mV��8㪟��{���u�J���r�s44�b?) 3({�ƛR�K���S*��� eXwx�Lx*?~H�1��Xΐ� \YR�[3?�퇨knE/9$�HT�y\o$��0dB�3�If%��d@�u��I�nٗ����uO��ΟիQ�$�XL1д�涿��_�Cwǲn�v9f)�!��i-s,1�aeҌ\6E�s������J�l�l���v�5�C���ݘ3E��8ށ>�
��G�(�b���:�![W�XF
$�ye�cb��V�ŭ�¨L�?�B��d�s*�1�I �~h.��Q�J��I�R������8��v�r&�(�qL\�����bɇ�B�B�He��\�0�f�.A`�,ޖ)m�=1[�瑽�%}F���#�ā��>:�љx�Ί�Ha�d��|gTF���̛7}�=E�]1�X��j���1Gsu�t�t�>�����!3O΅��3�j���i��Y��k�P���[T3cTM$:K��Y�{0;߰a���������٫V	׼�:��$<	G+��~J�v��j;��2A��+c*>C�[U׀Ç��?�C�#.�:�VYΧtkB~>�ޮ����C֗X�x��~��H���Ŵ��8u�\����D�7�4wt��ނhU-�m܂�� V>�,�r��q��|V>���`�H<�
ff�ε���\�t܈��g �c[E����df���ٞa��DO>���>��VE��;����h)ݧ:_"�a�V}���BYԟ��\��w�"i�8E,��s�'?a.��M2��#,������W1#���N��&Vt��)]�K���;�
�~��$y*�b?�����%#�NT�0��a[��$��s A�nA�̨�O��z	n;�;����HD�1,��@_���h�6��~���5GiQ=O��d'��m6 S�8�
�d7��-�����-ss���R��}�xԽà�QASY�������4x~�s�8��@$P*�h,�v��G`1�G=���$�L��q��%��Ƃ��O��]��R��{��P欳ߢ��6%)�"6(XS[���K��9��cb��+a`Z�Ԥ��B�%�uZ�ID�_W1H�����+-A���'"Ȋ��
��C�67j;��W�H@���aMt���H���k-�<���(q�&u=h�朱��B���!��cda��J��x1(�7%U��\cdr���Qp�=�P[ia��V�ȁ��N��|�iqr�񶷾].Z=�z�5��O^��@����\����P{�d�Yv�Ǥ�:\y�
�cx���q�iKu�?�ܳx�����ם%�����& ��%v٬Z���XW]����2Jq����ut�����|�|�;�(�d�<�p$����3e�b@"};hX�:�%��Eˆ[��mmM�5;��3��p������������vl߹[��јD�CcxM����~��3}-s��K�4t�9%�0���;0�[����ѡ�����_n��m<v����h �M��N�.�O���R�:*%׀�`<w��=\���u�K�kX���ى��f�1� %��͡ѣ�w.��D��u��{����j�sT����$+Yue�w6��-����`�0�q�=�{�V�k`Wqڂ�8�w`��/��܇3�.�M��lܲ~�QYi�:�Gԉ;vH��~��j�ڎQ�c�j�|gU6}���x"I]g�~ci~0Տ�۶+��Z2%3���jDG�g��������ŗ�i�dr�(-��2j���=�ԕR�~�Jd��y������y�b m�:<3��?\�Kf��2�Nopާ��a0z&�.�������t_'�Μ�)�Z�� ,�>���,���� tfLY�U:�V�vnݤ��F	 gΞ�U+Wb��I�ıw�6̞5�gM�Loöm���6s�N2pOpM�|M (s��+t�Dʽ��8��Ӧ�z48����ʔ�,�V���l��xU��!WǱ����]���:|�Sߐd�Q�C]M�^[�צG�t�qޜ�ZM�$&��rT�#g7y)fϚ��nU<�(gH]C�$�P�o,��t���޳S�a����p�M_�+/�*	Q��l�S�{B�
.�͘���؋�ʉ�w�^�Y���e֬}E���e��O�$
T5��� �[�����ͯ��w7N?�T���/c�����\�-,���=4��v(��?�~�M�7t���ߏ{Xe��7�-��o�z�1�W�,�a������9�K��l$C����@0D^�	ri��K�T�(EO��D6�E2��E�;{&��I֚��Lmm�U�B��V�y�9⤧c���:�44ډ�7#��Ⱥ3Z���Fe�H�fI�܅��[��I�S8�G�����k^0�Y���p,�x������-���y�de-ֿ���$gbGp��-�ڰ��Z�ˆmliñ�bmf��Q�ftcq��ƑN�%���S�wɜ�′Zj��l�iؿs;�D��!U	�s�F_������Q}�c��ݿE�&�y��8�޽�չ�3�Ӎ����Ο���@f�/�E�u~t����u�8v�C�i���QSPCT1GY���3,g�b��*�$���@�ѧR��Pm�<#-ƖZŉd���W�}�|b$��lVcF'W����7N���-Y �|��AA%�+ &�#E��\&k8�����(-�X6�lo�����R1@r�����̩���h׵�I���n���p%{�={2���+YVZ��/rޢeX��v�@��\�^���6��Fo<G(�&K�&�la����mO�s����o9bg��L���|R���<�$3�:��J#�=�,F��3���V�6��+���)N�D�zٶ�������\����M�gx���E	�Y����]x-��� ��J���$�v�[qݵ�5�V�P�˩-���}	���Wo�"f̨šC�����?<�V\|>���7��*��}����J }��$�o���������gp�W�"�+7XА@�W������R��O|�S��7�͟�,.��g��e����ō򊊗5k�d*<u�j{�r���G~#V�|������{	ګ�\���1ي���(~���]�"Nw��sTWE�_?�6���r�w���	���W����Ќo~�&��850�9���/	��oaӖ�:��x��?�[7o��T�?=�0.:9n��K����5i`;��M���*5\�l�0���w��;������G>��x���j9�gu,լ7�i��23��m�S}����O~��iŊsP_[�mr����=E�*�*7�@!P2q w��Q\F'�f��e����z;:Z3�1�<�N6y�����8����B������F�����"�<`;�WG�{i���������?-&:��"�X�\��qS��GX۲mB�#�u��-�@ �}��u��Uȯݼ�Ɍ㍉` �8[>"�5dFj�%*Q��E�d�$W!�*��ȍ���#yLn\�ƺJ-��bl'IV���*�f]ԊH �~���Zښ�6�+W=&�F��aqLM��P���U�Yv6��`/z�P��a�"eI7"�v{O����9Cv����%p�SK A^��c���b�IKq�)�a��/"QS7����6�5OE�,��гG%`S�1��$D�ǣa��9D~q:3_�l���C0��ղ��u��Ĥ��a�hѩ:7��ߡ�l��X#"�º������OSG�e�p�͈H搖�3f���6G�XronlR"f���:���#w_��N�����m�A��%�Nz����o������:�uCTb*&��5�#��|��fɏ�p&_�O��PM��4������!�b�Z3���� �^�sD�	[�)�ylRA�R��t��v���8Xm���<Ik&��J��(:%�YY�:R�hgY�"�� ,�x�Ȳ:���z�x��XByOY�t�n�B�X�-b�MU
�M���n�٥mƍ�d�y�K%r�}�dD�r�3Q�'� �ݨ��c�>�|���a���g��*=�1�Ʒ�rg^�ᛆ�9F��!��9��Gn,�o)8��������}k�(I�Y�c���� �-ύC�
S�z��ߋ�	�}�\�;~�s���Z\��k�[��o~�_�Eq�����t����ŕ��|�x��]��'��s�;7�o���8��N���M��A�oQQۀ
�b����'����.|�K_��s%��*��E�li��6i{���Οގ/�V�}�Ϗ�PD�0�?'�8]\˴�6���].���+/C4f��{�����*�t�=`�m��$���z:�c�J�|�٧�g?�j�F.]܆m�ڐ�@�e'�s�ᇻp����e�;��e2�i�-��Qy��ڐn�0�;�TY;�{�~�r�R<�����~&�m���+�����{�zNY7C�A����?�������ߣ�_��8~q�=Z�ɩ7s�*EP���U�$�a��Ů�$Ps���EhoOc�+kq�����g�Y1�L��൸8^gy�go�!�0�R(d.ۼyù�H��o`�2`�Q�h%�K���B������F.�<��#hTn��y�[�6���N��X�RVVK��e�e�=��T�p��(I=��#�6` �񅀇L���h>+aĘ�f2+�1,�#�39-��ŉ�`��ݏ����.XZ�"SH!��DMU=�E�v�V���s$�ւ��d!���٧�0��}�\�����)�')����h���-�ɒ�@�+,w�pq03P�Q:rThÔ�#z�r��;��?��.�b�:Ĺ��m��1.�@{�����K�Ɩm;1i�t����C�G^.��Y>�<?+���!²�%����m�p�)s�~��9��Ӧc�8,ABWo7;��kVK����y��A��#h����s0s�<q�9�)B��j�υ_[[�N�뀙.Ǹ�JF'��^�b���Ѩ��\g���g@BgF��S/���\G���9��+����SiT18V�"�(n>�;ȑ�ȹ�SN]�ǟZ�=^*�%UF�])H����g����I�H�'�CE)��v�)z��!��^r~fvĨ_��ؗ��b^�]��|�r��9�.�+��z�w�1JpfE�,�0#&ǔ��r(�9�al�3��rxZ��'kT��ͥ`���}'c
���6et��쳬�%W?qկ%��虼�zk���X:�f��+|G/�vQʈ9���Ht�f�$�F�ˋ拙8�^��fZEiTi"�N��¥��6��Ȑ���a���ݶMn��P�[���m���:~F.Ɏ�q�B��8��v����y�
\|����[�-���ظ�w��/�O~��Z��O���Sc���7l\�D��CG4��O=�8���J���/`h�_��ʭ�ޫ�BAL��׼���gdoO���֩�ِ��gW���@msl����Z�P�JǴ4L��V~ub.c����r��v-�9�dIjپu^x�}]����=�����;�9����
�{����o9�%�X�`���X��#������_�UO>*�-���Z�������]~٥�`������v�c}/�ooG�D_{�b�n|�#��#��yܽ-��yu���Λ7G3�-[���*���$�~�o���[��8��d�b��_��~�~���� ���7�����̓���a�j�qb����K��*���GNT��_?��V$��N�ֺp��&����m�di{���lIb����|��;���e���>������Ff�an"����,��2�c�"g�n(�+��	qs;�E��ƈ!�EŘ�u6UBq�����w$h,�W��|�QB�Y*U��L�.Y�輄�c,q��4�N��M�K�s�����0:(��ӧN��m
z���B`^0FG��1ʪR�0=<��Μ�-�Ytaۖ����W��W�O=���G�{��(�*Y�9�-G�D�Ӳ83�#G��Li���{t���hk)�X��ѭ�n�-r>3g�m��3�Ş�[�i���}H˟;voAg_N;�l,Zr�ܻ�s�e��m#f̚��\���x��t��*����a�\GX,EUG#a-��AZT�.ҩ�r�)شiSQ��w�:g3�)ׇj{�<FF��}t�O��Q��b"Q�H��� p� �����mo�[��Ԓ+=u�WG�:{�5@`5��?�:���lC��4�Ռ�t����bFP�s@��Qيs��X�A9��V?��}��j3}�Li��56��A�P�'�Cݍ׶����<�em�5hh����=�P]߆��sL.��@o
����[L[��5�����v���A�� �|�8i�����9i3#�ε�4�����R&)�%�/�� �]�e�\&A��ң�:T�$d����S���-��^��|�(�K�R<��#qJ�-~��\L��|��Y/Qߚq,c�,���d/��A�=��H��-سᐂ)Y~^ AX������������.;1���qxq�i�����D2�3g)�����]Ԋ#d-!��l���秞�6�rSs��89s���,Օ���d����� �<�T�4�bT���)STfJ[ڦLRg�j�Xߠ"#�	QǦ�3��\�l#^��l%�by�0B�u�0��Vy�I��a�Ν
�[8
NZ���-ȥ���W�I��ӗ�ȑC��!��J �p�,��%N���$�d�����S�?�=����ǟ�=�L�k��֢ן����.�Ġ[�1�a��J۬u�Ƌ.��������݁�?�.��b���Oc΢���/ߊP�����Nׂ���>(A�/�x�n����Ϸ~Y���m3���L�0����y���w��߬�ڮ;�����i ��1U�؋�Rc��94\aO�N���7�P}�~?ѡ����o�����:9����ず�2\�	����`�-��Ė���/��ı��K�X\��MPtXz�|�u�J�R$�Ք�Gu�2���������1�ĀW��yۣ:�̲8{f,GsCQ��Q����zV�r2ω#➈�H�"�&bz.F#��NխH�!F�}g�s_���⒨Kn��)31*��k�n�7܈��s<������b85����@P�"�YƯGʌ���qy�~�s�A�سC#c�5m�l����R,����p>��Υ�y����Fu�W�z	�����#9�}�o��.���[�{����٪��f�ڊ$MĒ�3g�l��/��eϞ=ꤹ	Y�9�'��as��T��=����`@�Ϣs�����U�T�k����=�T�I�^TL�F�PU���d�+�J�!����:1d��<+0��8"�;�%S��VެYκ�iQ��!f`�(�qʂ4����^����-�`�H�o��v�:������K�Z����E����,X|2��g�̛1FGIbX�+W֑#0���)P�2�h԰l2�y.��D�z3� ��P�G�_�b���&��D�� �5�q���r�[+�f�Ѥ�i[f��Z�+�u�f ���}a?�w�~��y�a<���Ky	��z(��Ql1loZ��z�D���mڋ������H4c$�}
Z�h��2��w��GCSU��c ��5�9N���>k��Y���Ｄb֔�C+�z�m�ڞ!�#���0eR�n�=x�><����۾.�<��Spl�M���얽q&�n �m�Ѵ���h~/A+��}��T�\K���+�����K.���ԩM��M�{@w
{vta�$�u�x��O�>�����X��W=.P��GW� g��߸qN=u��'�ūtJ�����YsuT���WAx�	^�"������A/�s�!h ����H2�U��Οa�������G��Y����=�8����^�a�,������&�/�}r�/8�\\��k����F�\;L\CЀD� �A�c�����3F���p��e��0Z��E�:묀/]�)���.�8���g礮�.143�5���Dg�b�m��r��K���}�h>��#���wJ���0��6v86hs��2�rm�Bq	�Uw<�֋���:���
��a����f� 7�ԭ�I�lI�scɄ��qF<��1�b�}8B�)��I�A6
9��:��'�HC�PP�S(�R�Ƴ�Ӎ���q��UIQF��76����=:s�kU%0gѭ`99a�kSk��g�u�f��C��2�\)Q}]@�Ku]����twJ�٪z����$���O��߲�7����S%��SƤ��J"$���aR���z��by
�:�����'~r�m��kߋ�}���,Y쫛��L+4�^�a���l�y�-Ǧ�[$zߎ�� ��Xq�%*h@'���Z�G�A���K����ϓ(~�4�uM�:�2GN`��~���J�C)F@G�H�;g�<�8vKT��C��+�+���_���D��0i�����ƴ�������%!�����2q�-YC��F��)KVG6lڎ���U��%�rm��\Cc�v���D����w���?b�B)	F�0�&MGP�h��[�h�*:q�(��1M�j�L�<�6�f�1`�K�`��53^b���eHl���l{}/��ۮ��l������&F�2�i��5H�U1�-/1��P'�9/H@���J�C+s�ni��u���������Ş:�Ɓ䊶Λp�^� `�\���z+�<'���$�Ϡ��^�[?.��"��wX����e�$�Aj��[$+ݲm�d����O��e�������a�k��CJT�_ڞx<��6�Nl�9ZZ�d���I��;�,��Y,[C}�d��cr&�1���k�!q�$J�53���S6��ɍd�l-U�T�!����c��݈1�{Ǫ��˔L>��(����Z9��W��w��
|���S��u/��bG�vr�����Ź眉UO����/U����69���^�Ҩ���$-b���qe�R�Q�\l3[�b{�� k\r�=�c�z�olAjxO<�,z6n5��@�Ev��~�U>��/[�������q��?�2�����x�����t�F���Rɞ؀�We�e}�����wH$8���T�" �3�tt$�/��P���KkɅ+:�)�'�&)��uc�9`��9�1N���x�����q��s�{�!�}���1��c�_'Nl(?�
0�<�#��[��R�5L��1.���kefF#22jX�R#�0x��!k�j�m�v,Y�X�59K$#ΰ$�Kz��WQnpX#r'�rl\L����M�:��c m&G�h�j��D�m�g�/N"��	�}=��D�|s;6��%m�T�R=|D5+��I/���r&�6"38U�r�	�SϿ�f�c�>#����ؐ|Π88VKB8"AmM����� �5M��ϼ�����w]��n�n��g��~X����d$#'p���l�_~�v���R��UǷ��~�%B����a@��j	���]��<̾���%��J6ެ�;�͸�Wj H���"�)@�y_�qϸ�|G�'�S__��O��/���	��F�z��Yc�����̍�ɊJv���^:�FF��Xe\+!���a��("���{12{�m�d$e�$�s�t�D͏da��5p4�Q��Y���Q9V'Y���&tS~W�{w� 
����"&ǔ��ǐdH�����;:���`�{30n�˔��RtrF���,��e��/<�����,����Bg,�����R����|0�HO4T��������:l��l�7�ۇ	�ׇ/+�����������;�D�Kϖ��^0,jht��{}��Uē�R@��ņ�/a��˱�9x�g���/��5����{ju��/�c��Y�N��7����6t~z�O$`=Y�Qj��uf���۫����n�iÒ-?GN�&��ʯ�������(��	b�ށ,m����u矇��݇��}J�)��9�ǐ���$�BLd>s��Ū�h�>�YshB�r�Z� v��EXZ!�k�۱e�.�u��8�{ ;�nÆS�v�X��#?�e�����~�3�>_���%Y8�U�W��w�]����dV�J6�7+I]�� $mQ�:r愣Y	���Ir1���TR��q�3�$�#9��7i`�QY�,�l��s�Ӂ���K3��`�J'���9sГÿ��w�{�Q	(ek���I�lC�<�|����v�͹��Q	���6�z���x�`���X5�"�\��-�#�p�_��6��=����sN�sG���ާ(�g~_�x<�rQb�B�M��O�1~��I�X�l%װX��Z�^�9���\���%ji7�z�޹�&X�]��_'�������^��_��#f��(9����j�A܇*�RI2r�g����B�o��i3�XW���c
4��6��+$�g������S=9KOa0Rm�h8��ӛR����1r����G�5��=�)�Iq:bt�}�Q�~�%�͐���@����4F�^�Q	*8_��b��U�2��T#b�=�Z��H1�q���c��jgG\	{9?��F<Y��z^{-�Q{xHٛ|q�!	*H��<'�y�7J�݋�/��k�G^���dT�>�
����i6�O8�g��AP^㌙�>�GZn&��2�=0�#zQ����D�<�$�VH c>���3�dT@��0���#Jq��a�Z�}X���:��p����pRǋ����Vvr�d�s����M��J�O�l��Y��Y~&R�g���/2R̰�U��aƁ�ch���R�Z�]����3����l�U�+���'X�5��� ���0� �_c�g�,?�>$��̓mb��/�@��޳;
��k" f\���V��̛�.��ba]w͵�\�'��{�y?��ļKt-�����o�>�O7�{���g����:l޼Gmѹ眯h�����/)���I͞MѦ%8�o������K�){�����ֺ����Y�~j����9W���x�d�G0�,U������N���
x(wW�P@�,�w%�bi[�\R�XEM�8* .N2(�neU�$6i�1y��!�߼��_�5�*e񦭻��+���*�������/\�G�xR�0$�F���Mhg�/_G冧���4���b�oh���E��O�G�t:���c�	�sx��C�������g	\mlnCzpD)��bK���0�w�w��Ż�}�.:Yl���|�&	D�x��m���O�@�4k����6�k���e;�7;��8V��h��s�31$��Ks�~[Z�'�b�������E/�e��X_��Sj�w��
	�?O|����K��s(���R�I'�����|�������ϰ�9hd��̫��QT�,�P�3��Fᰕ@�B��4q�R��d�7k���cQ}�X܈
d3��0R锞Gem��ʫ(|�e|9��3��y�$dd�X��Dl�J32"t):2��Nٌd�ڷgFdwՐ�=h�j�%�
�V�NQg��ȡ�w���'?�[��lz�5�֫�?Ѝ$���1-O��F�d�r�)��m�22Q%��)��H�UJ��ඍ�=7I�02����ND#	�6;���}��?�!���:�b&A��U�#(��et�/�x_p��$��a�s������;��В�>/��*ƉQL�k�C�'���B9ԁT����Y��lW��ɮ4�  ��IDAT�����#�3'�f�1	N�G�$`�F�f�����m2e:n��pԘ(��v��X����&����E��5\��ҋ�*��}zֲ� �:̮7��ؑ�{���#~���{$ @��lg�Rј�^�^�hǀ��w^�P�s0Zc��昿�+���7~���?����+����|-_��k�XkcǶ|�#7�O��-_��8r�<U�S�����5�*|��O�m��;$�'/l;.<M��갮|�
<��&<���/ނ���j��ѿ�G|�������Z��t�޻~�oq�]w�e�'��|�����4O�(o��>�Yͮdl�ڃ��N9�Ző��4��� �<�9�%[G�6���/�
�}��8&v���0Ϟ"Q���	J
%qow�;���_!��p���Ɲ�ĦD0������J���'�S>������:9�#�S�!ɼ��0���;!{�:}�G�l�\��e�ӟ^GǱN���M�[K��%���_龫;Ƒ�x �h}R�M
Ց��F`�C���uÍ���b߱Y�����cu/.Ͷ�eMRS>��f#�f}X�R2�\*�{��uT���@}
x�g�'�=1�����O��O��=ʝK�`�)�3����,�������rQ��S��:������G�P^u(?~ʈj�m���A	6B�l�."'�=� K��n�Ƣ�X�af���HVS�dq�9���)��i�&�6������T,�Ǡ2�^��d���}ԁѡ��(�9 Q��c�zx|�J�m��`��_��Lɤۑ��cS4 GD�@���,��F֝�4[����_���͵67H���/;_2�9
�#r���(�I�OG��@� ���Y�
BZ��y�t��z���W^,��\-�N�5/�]��{B��^[���;�����X��%����V�`H4\S�)��Qy]��#cz�H���\9�]m��kk+�X7)V���i`06�E���Ft�/��ܔ
1��(|���cޜ��� ���* �XHg�)�;�<�B���������np
,�Miݵ��W{�F�2nU�*[�va���\{��P�-� ���wy�-0�G�Rց�?��f��3��uZ^[+*��٧r�g��Y�}~�ϔ�~�I:��W�i��lJF&=�ঠ��U'� ������?b�kk��A�gd��/h�|�G?�w:|� fϙ��s/^�u�߳��V�O��/|�������ŬYs����y�?8�QY]�'_��W=�D'�Ǵ���O}V�/���R@�2���R�&�zCd�c�\���H�ɚ+x�ì�&)����p�n������~��۰c�.Y{I����J4{����C}����]+h�P���7���
��Ū������ӏ���_�2��5Gw $��G?�]���E��Y��%��ޱe�[N'-���v��Ok���F���+��8fBJ��o�N������:�q�dW�ut�����F� C�N4Z����z�y��C����ǐ�4�`B冹�r?�-��_��|-�sy�W�iTG���y(�����4ug}��'8�"Pn����Й�2М_E��lb��3��?AI�*U���u<�a���`?��T�21�PI�\��ͺϣl���?_�`� l����A"3C��A6�w�R���@%֔�VY�RJ�eO��WA�����6UC�%1�z�,�;n�`y� ���tVAx�`He:��r)�F�F�("M���&)�Kv��pg
�ըm����~�e�S �͌�?�+�X�o�Vlٴ�@�ϒl��$�3���FTI�~������c���fa�Z�ĐA���Tn�&d���k���/E�@J�p��|��+p�Y��֯|�v�z�qDĠ�z�-��f��w��3�\��Ί�nƐG�j�%�����`�=7�R����Ց��&��z{�Z�VW�h#+�Ci���������H?"����8:Zqt���:f��%��fDb	����N�����ɰ2�AY�Q�I*����5UP�Wٞ@Q�������������@פ�S(�6Ԡ��"8�_��7�]>�j>ʳ���������\�>����ް��Z%t�ε{<p�?�6���َ���ܵ���s�ZD�� t���hl���~�hH�Zj8%��<���(�ɿ�� �r�;�����Q�c�{4�S�@�I%+3����r�C��^x�դ�ɘ,��N8X��صw?�8��p���}oE/�ۖ�2@�rt��)�9�K�|�elC*{�ŕk$`Y��~��~�l^���'��0*�k�ۡ�d��a%1�)���� ,{).�xH2�g��V�.�2�;qX�_]}�ڢ���(j��t����?H02Il�V�:}342���Ftu���NƧ>~~��G��S+U(��>�8%l[��-�$B�Q+��D������.�U
��q ׮�p(�B�ع��j8v,�F|��!;����
��u�T�����dE�[�;���#(���'ܼ��N�#�/��2k˲��%ި���č�?=�s���h�r�ݛ}�Q�o\t���}C�#7K�4���������Z�x��X�����."�(XM-eOIl�H��t
��D�g�y��A��,�ΐ�05�sit�-�[%�_BU3C���ϻZ>��֦Y7��x�R��A�A��J���gFh���԰E�ӝ´i���Z)�� :��Q��Sf���S���v�_�?���{~֩������[7�������<ّ�D�c����ӟ�$:����X�-S���O��H�J��-���o���X��;6c���h�4�58&��V�����[��������������]�GΏ�htA0
vT;�e��Vi��2�*�J�c8�BD����R�A��P
s�O��E*K��A������_fń#�uu��}ȣ[���dV�j#��s$��xZؽ{�d��He�X�p	��#��թ �u��^R�UNq��9�_�>�_�^���׫}���s��9`���ʾ����k��a��&�j��rY(�>�[�W��J���˞�����_ǝ�?�;��u�����]�(��Y���Lv$=���p���!�X'�=�{OuE�ұH�5�V��1`������\GZ��Ti0T�+�N�B��p/����k]]=�={&�4�d?�:Ӗ���������H4��F*��+����s:�l�Q�Z>8�F �b_�T�{�v\t�i��3���/��UN�(-�m�/��yܕ��&�
�lke�rL8�e�5P��������b�����}�"0pg����񰂷G$P:m�bH,�d,��}�&�$��AN�'W�(Yڂd�Jj�����$��	��	@8��M�8Vy�j�+w	ߋ`8�K��Q�-A	a*vt`������U6C5�m�o���fQ�\s\H����Xܛ���7*xO�����8�j��O�(w�������N���q9�^yV�;����j�?���w��cw�����8��cV�R�r�K������6G�B��1B�#J`ڬٳ�q�f1�B"�<9�V�3�򣨠p��e���V*����c$x���%ƊTX6N%��D�r�#CE�=��:��ټ%>�m��X�	j*B���G2�̩��Σ��G2��ض���T���J�A�@��<�+nx7��ݎ�v�;��W9���=N��xm�?*��w�w� Wb@"�j�0�H ����������g�y�V|��?�s�+�?'Á�U\沷����aē�j48O��Ysfc���@Ea����*S��n�U�~�k��(��ͫS��`��]�S��Z�Pal�������ث�/�Rf�\�0�L�� �/�M��I�6n�c�Va�g�pQw Rݭ	3g6`��VTTM���l�����c�V�����ÖU�ެ�	{c�Ͼ�-�������^A���U��OL��o����:�l�%T��������g�9V�?�c�g��9t:ÐUz#�-� ˻�,��!���أmZ˩���1>(db x�*D��]^#	���+�+�&�#xO�=3N������ʡ�.���8��� �?��ق9���]����Ǉo�+���y��#�K����җW�u���T���s��RU�R�WR�9�3�ɑ���W�8��j�Y�QYk��]�|q쏀9�B�����OX^�}�9�����*����d�?Yh�k�'�W�}o>(��+����He�bػ���V����|�&�c'��\���SϮ!N�(~�^��7S��dK��+��7�����E}6':���zFr:7�����K�'zL��OT>�������/v_P���>��;p����A��W�:9�h�����s�,?�1���s�{��@pG8�d��
�K�Y_׆�X���*uH'�=��
�<∘8���I	+yU̐E� 9�
,G�|�˚B:�@���T�D�հ$0�\W��a����h��Oy�c�*W>yș����e���&�TԠ��1ټ1Y�C�:c�����3�����ڌ'�� �{���F=O4Z�4	�kk�ݛƒ�����Q7�N��)_�4w�-3)��/}��g+Y�2H44G���{���k0���%�a6��{�3f�CGu4��5qM����x7-��89Ό(�Ѭ�����]�tc�V�4N»��@2�lް�*�hi����=�I4K�Q1�I�q2��I У
p�q��a�r��RS	{�<L�@`�xi���-_D��i:�`y��}�ʐ�<���< �p| m�x*n%�ߓWyR�dm����Re�u�����ms3aJ߾|i�w��]����gF�A�}��pa��%
Y�m��F��u����� �w�qw����N$B!w�@�u��ȞȲ� �B��'d�RE,�yA��)��q�'�1ol�OmEC-�\��%���N�u�:f��Y>߃��QJ#Kb�@DeZm˫�X:v�G>��g��Lt��kN޴�֧�J!�r�rNf�Y%��	
q%���[�.4�A7�G��%QS׀���,��y��ɧR�z}�����	�Drz�o@���B�CFƔ�8���>�ik�m4�R�/�M��o��;�ⵦ��Ҽ��(H6"���2��A�Ni�{k�r̾"�c�$����	���Q����M��-�����)O hUl'�fQ�r��x�e��1���[1-EE�*Q�N�vխ�9ۉN�����}����lNԃ>Q���3�멗�g��M,���n�B�$��r:\����w��Ο� �������C�ئ��Q���tc�,<��P�ǘd�v0��Ū��H���&�,������iɔ�0��E6������F���_U6}V�ɞ�~�� K�O��77U��SOU�I6G��~%cٷc��	
8{Oz[��y�d��9E�6����F#*|RK�j;S�G�D�,:{�%c�����̈��̙7W~n4iI3�5̒:3��@�ʜ�;*�#��*Io�1��o��`a�jL��1�t�~%���`?&O�����
J����r9���R�)^�#4��=�{� ��q�a�l:�w`�_7(Ih���y7k_�,2J�BŬގdR�����jrs�����g.�ϯ��M���:)N�]�Q��7��"8*��-�5)���`̟9���U5ĥ�/D��Ͽ�*b�J�}e�d)������5I, �����L޴]ry��&�U��p��-����k��u=*U��y"�ĸ�F�D=���W�.���D�>��5As���R�=ѡ�\r���H�f���x��-��}�Kx�4�/ū*d��\��A�w�7�y�����BmK.���ؑ�Z��X�А	��ޫ���`ާ>�y�|MYU��V)Xۻ:Q�<
�ʀ�$I�e�5�'��J9��7�1K�|�V$�\�}D (�ĸnjk�p��1U#p3�5�K�83��,_O��1:�������V Oyu�Դ���/�%��Z�WzC��ن�S�U4Fq�86��������by�$hy��:��>܅���E�jPj��6j�_���U^5����K��OF1�1�@�.��&ߜC�f���s^�O�_�9���&�S\�;A�Ҋ��2g6�]��KY�_r�����r���o�Mq����� �<����z%��|�r���?������_N�Q:w%��ps2���H�k����ܘ4Q��X��Ñ{0g�t-�_��t�ؐM�V�3麪&�y���8*5c�,q�3��!lݲG�v��k���z�Z��e�!eA�Nx<^��>�KEFc�\��r��J�e��%�P���D�QGK�TiわUV��gg�_��q���.�T7���J63<0�!���5�#(�kqb /����h�1q���m?��b�ң��K�l��8|�|˓�@�{��d2����I��N!!���V2^�Ⲇ��=��̋�	Eb���#d�|i���p(=����dV�̘J�v�S?t�'/i��'/]���!YL9d�+���E(�h�r`��\ό��&��;zw��iKN�ʕ�aH,���S�6��UuX�a�8�$*%�!aP0��P�5���`ɓ_��!�8�� ũ�l&�H��f�����:�w�v����s�P�_��Ė��9��� �7ãc��e(�L5��'�K_���.�ϛOb)���4kU納�L��o��f�|^��A4V4��'�"�U��L����J�U��UG[�ܨ��RY���Hx��M�Ӣ=aچIU���i�6GmBU�F�ݺx��
���H��]�b$=���*�p�S��Ъ���ɌیT���dmQ�t���S!�Q)�+�ICL��y��2P�q�ެx��>��ce��13mb+%�~s���/B�_��X����}��W�8w�݌xZ�N��U��$�Ŷ���X�J.��(X�2b��ت~�׋e���g��o�1QV!0>����͌�z�^��[�ޅ(�Ə����&�NO�i�ϭ�h-W��G	E�F�a|�^���.Z�������8�ŕ_�(��U�]��e����X��Sa����1���K��f��B#r�3��yf��,tL�Wa�\I��z;u����~��݈M��(�Ecc+Z�bزm+2�v��NuBݒ���"�|�8��.�SG(�K�Ú�^C}�d�}�Ɛ8�dEFFe��fn�ԌÇ�*XΊ�� ���75�����h�<IEC#��5����Hg/Έ�;R�'�yW�㝨kiQC�Va�8ef�Q��e�z	��mb��}���m�#�������cÅ�dr��CYL�7O����G�{�IVV���{+���ꜧgz"0���%�PP֕]w�uݟ(�*��[QAA1��� C����tO�\Օ�}�9Ͻ��z�}�x��S�SU��}��s��|� �8����!?�89��D�� �N��8W����2lh0k�()������$y:9�߁�W���x�N����0`#Gz��A�+,M*|�V��cسgT���ɋs�
�oo��$)t���ȠԱO���qև�.�������xⱧг|y����z��^9�h�KG�����p�s�Շ�H#��ۢT^1(H7g��4YQy��re*^��Δe�E�d�������G�)PZe�"��%6f�s%.�#��P���*�W&0��r���y��M���ِ�7�����W#|l�e���s�D�^u$���w�D����'���� Y0:��dv���2�9�u�}��T��)x�>8h�e�a��<܎�[�7�5b0Km �����k%'q��"C4F��v�~�ȝ#�cs?�O�M�'h�KYeBZ�k�%���م��0"�'��e�t�1�ʑ���l�Q0�	����TwѼ��S�L���M����N3����G�(�Q�%.�}奣О���tKo��\�!H~k2�zAWp�R�n�9���Xq�fx��N����/8�nC�6;��&�R� u�Y�[�mu��0�����]�b���R�J�x�>z��K������h������i�竞�폁��Y[e��C+���r�p<[��9�B�������sV���O���\;�d3���=�b ��%ǲZ�:I!I�*�hb
�\���"��Vr��Ys)�Тw��<�{P��qɍtm{�J�c��M�9T��N�g��O>����qKG�"�D�` ��=���q��CR&�ڡz�g�i��y��!��#4����tx0��G��L�^^��>�A�۵w�ǲ�K��w�~76����~i�X�ڂ�47�:<�ѱko^{s���?xp'�}�y�����o��]-mشy;�9���v�����ދW�\O��&ƐӮ�y����^7IIe�{�����XQj�ȥ���إK���[lټ/���x;ң�gG�<�7@����NTi������sX����3��OYq��D,.��`�Nqv/Ɔ�����ǹ���� ��'�j\�݃ɱ0�^�ĳ		gfM�׳d>�4�ظ��U�M�}6�r}f�Q�~V�X}l��
�[�=��R/`��qT��#(��[��
�%�KĥY�����M���^�N��)�"�ɚ���-(e0������	�Q.-��v��%��C���ũg��կ��PCKu���>�'�x�W�(���g$?~�}�I���_���:n��f2
���+$�����ӓ3�����ݍ��#dD��OK���q?��Gp֙����.��/����z���.|�[�`ݺ5���N���5�\#��'?����o�Q��}�����>�яc��Ÿ������!��8v��,Q,^�K��Ħ�g0h�#����E���
���Y61��ڬ��&z��ʳ�a :�^j�Rܶb4�s�n/Hi���i�{��+�_`�ctX��P�Z擙�ac-ovM3���/��o��7L��P�۠�<,���W�s �j����P�a�c!�9d+SL`-Z]��S��:� b���.C��y��}����7+�a� ?�7ֵ��7�a��b���\�6k��@�R��Z�ڦ�9suվ��p�ݰ�� @E��O�LC8p�aW�>��%�g���Ԅ4C��^=[�5�0���k����ۨ66�ctp�����$��ý}��b�{��o�Η��� k�l�	؊��#h�������/��^��{�IN��llĢyZ�#�A8�	�ԑ�JJ8BJ�opg�z2��Ū�oa��bd*��[E�������z=������p�8<�f2A?y���Z����g��l޶�.��6R�3�~|��;�a��E�3RcK)B �}��`�T�x.~�L�*�qYd8HJ����T���$���%C���t��O�:r���|'�8��w;�ʍ&�o�.�F>-i�$	���G"36�%�io���$y�3�$<�Z��Y�������� MK�sφhmiA:��=��z�f�03c��M��gw3��[R:L�+���H5�%H�'�V��V�_�X�o-��p�V���P��.]�F��S[^>g*�|��}�_�<�Q-�1��4�U/*w�9s3H�@3��w�$b��'0�O'�c����׾��y�n���?��)��Nt�]��_x�[y.�`������Ia�<kE#hJ�����x���I=�k9��g>v� ������.:g������~�#\w�eX��ÉK?����>{�58v��;��u/V�x,���$����� 2���	�{��e��'>z�TPl޴۶�å����ػg?#Oњs��wksƧg�7�K��1wwQ����2�Dm�*�2�-oe��/z����4�4[ɳ�
I��P��Pd���\����p��fX��!��z�bĚ瘬�iP-Fr�L�B��������E�r�w��\`�ռ��U+W>.��R���Ԫ��*�o1�>{�Y����+?�K��K����ػ��|Q�Zƍ�e�Rey�䭔4���(�镞��.�����߻HH�M���4aҙ$y�	Qچ�N�&������W�m]=��H��K
y��v�L�D8�`m,Z�C��$�^S��6nڎEK����(jC��$0:�����i�f�5�ԅ�HH��Q�Ј��w��X�~� �؃e�=�]�`�om����a����TxW\uv�܂d,�Y����`��c�Q����1lܾ/�~Y��6o�0��$�r�|͌�^�^W+&F{��S��gFw'ӯ���Ķk���ϒ��'.?E�q{G'�>�����?'�7�N2Pfq&�R�pLړT$1.��!��X��'�w\���8M�D���l&!��u�>���H�w�t0<6NL��6Bʺ=ݝ�/?�w��8?�Bv�x���E�0%��[Z1�?�$
��{\�ز}��.�9GB2�@�0���-"�8Z�cr������)o (!_A��i.&���B�0�����DK�MА�A�}�(p�ZUK��9�|����(�0�)����o4�C2��3���\4�-�e��<��}���_�芁OEW�H�>�~�L�����ظ�E��^�lٰVZ�|�<����;��x��U��⋱}�2RX��M\@�4ײ�Ȩ{�'q��T�f9�v�KH|����T/��#����@x2�ukcٲNl�̝�j��oк>/��Ȫ�{'�x#6�? 
'���_����^���V+��p�H�w�b^OɈq447�㟸��j�گ��=��O?S�q��{09r�ɖ$�$RSf�f����XS�s�f�F���i�x��Sx���
r�/t#-��U^[���|��[Q�|��R.�����ӌ�2P�U��w��L	���"
CA_Zi,�]++�r*��n"%Z��3��Eiy��`M+�-j���J�������ZG�x���V��@�^G��u�jщj��o�3�l3�	e��Un����=5��M���ȃ���S���$f�Q�%1D6�y+�(O���1#�K�L�|��ڎ={�!��-}ӷ�9,�-����a������)���,!\.-����u�!lڹ�<���]��������
W�`jM�x/\,a�C
�Wmݼ���	>=9��y�x��p�E��w�?��N���p�"Oы��{���$śc%�>�2"�25f�pxm�X'��8����w�9��}�xm�vi�^>��[;�p��G�.���}O>�^x�A��ݻ�����.�x�^�>!��4��^�|��%ʹE6��[��hN1o~�.��!��hxϽ��{I9�����0>�9����Yq״�N;��y6n�N
=�H_�}�����sϦq9PS׌��q:N���!)��Y�ddq� #��~*͈������h�5K�En4��H3=��%������?.*Y������c����F�W9b�;F��-z]�������G%�&����G�˽�6(�2I�t�qؕ��?~���LD��u�M����W^y5����j�}<��W�Is��U �c��[w�\ػwT* ����ʳ۷�(����陏={ ��w��	������q�ݿ�>�۷o'���ãxu��޹��������	����/�A���A�m��87���!�Bw��[��� �\������u'�0_(k?�ѫq�W�7p��o����ں�>����
�\b$��n��i�3��Z3L��Ѡ�I�S0���0#0�L�yC�W�Z�!Q0@���sIv7� �"=�I�2���/�
9�^6�xL����{^��X�%'-�J�z��-�ɰ��#J��?�YLns�׫!֏�R��̏��+�,sQ���Aٖ� ��̀���1w�*���Z��V���Λ�D��O�d+��n!��8Ag��[����$�	�Dƃ�'^U���tJ�����<��N��fr�D��W%��u�_���I�5ױ�NJw0����1�u?�꛰x�8D�g�뱷wP��#�Ѣ�"�0DJ����y���u�낋��y{U3j48wFc(h$:C
��P/n��6<p�/�կ܌�n��,�����w8|X���k8B^C,��E�#�0)ZV�Q2\׫(sI�f5�RYV����F0OX�d9G'�s�A,?qn��7����۾�m�t��B�82:���i2��җ�C�5&>S��&�+�w�̈́����cЄ#�7F�3:���}4�X�h9�dh� H��C�=# ?�j�'��H�(p�2� �|�~/Fɐ _x�����0vKT���.W<��+`Rq_���[�';��'�PЇ������p-	�ֶF���Zlش�l ì0���퀗�.�4M2c��G��,V���K��U
f��
�nɚ�"���~;wȻ���r|����w�{�2e�r�t�
��A�W
^$3A���< L1������lǞ]Ø��g�	x�;�f�^���{�u�=.[�12����Q$H>�JTw�)�03%�9�֮y�/��N�����S���C�?��UG�L��(�O�뮕�z>��@��k�u��y#�\�� ����hRD��]�F�'Ҙ��a9�a�f2�EǼ����o�Nh� p���_���r���K�.î��O�ܢ9�"�=�f��I%IƼ�&�� ����r����|����J��^�P�t�I������J.wPass��?�H)o3�B�"Ĺ��j?��0r*�4mF�c/�]�����l�� Ea�
�7�ڲ��	c�e�<$������C-�ϵ��Sh����GY�%���>o�e\�im�}UB���d+Ĕ{����l�a6�u,I��6�y��q��*׳���#R@8���K�$T	�ؖ�o���ܴ�Ə��	��I,?�DR6��MA<�d���A���֭n��yS����n�Cp�����ǁ��e���@�s��
u��.����f�νؾ��r�B���"FV����1Q����8,��e�9w(�D:���q�6���HK�&\��È��w�]�����}������[���:�&�z�r䒼0���� �HB�V�t��K�1+�X2C���<�$�u΍NQ,[Ҏl<��@&'HB�w���ӟ�y��o�ߎO}�:|�×K���� ��Ο`+�`�Z
)	�J]�Y�j���((5n�z7�>��c	z=n�"Ԑ0��N��a���Q�.Wm3�>q�q���מ�S�n3��H��8�ۏ1����1��d0�{��(2d� y}A�rn����&/�+5��q�e���Ϭ��Y+O�ƿ�pol:,�*�-\C�(�4y�\�� Df�2�u"�ذ$��*2�5���ެ���T[�PƁ�}9!�E(c�V�ס�aܗ��`!��Oʉ��^|.qe)%�K�8Nk�{��h��6C��U	����8�Na(��/'�����x��''-��P?�F�0�Ͱ�\HL��F���%ዤ@h���� v9��I7 Α+Z�hnW��{�3�!ɈDV�gv2vmn�H!���ƕ3Yr�� �)I�C�HG#b�st�fin�]5H�г:)�Ze����`ҺF?&�&$�ewHV�zI:���+���#C�����������N:$Bk��й�C rLj�A2�&�T�
mr��-kL����݌Y@J#�P�Z�1g!��Y+�|��E`�:�^�:����"*��%%k�茮J�r8S��	{��,Ԭ��*��-X��|︪&gS�z[u���]m�R0��u����f�y�R�*�[%ʻ4�^m��͛W��u�U��Ŗ����>�� 9���[)Mu�`Q�hf��;{�R�J��E���^��b�n����{$o���SV����؇C�F"'^��2eYΈ�^R���#����l�0��FT�+�j�&�X�9�ӊ�$ν�]n�C��`���,I�0d��U]=Mh6���f��è%�T��btp�=�4n��p��IN�����c]��w�"!�VT�vaQG���ڙ��db��2W4��c$0�QRS3 E�i���?D���^z)�]�F�(���8���lڶ�ƚ5�x�9(������۾������Y�y2�Dw���&���q ���w��� �F��� X��;���mh�>j�����\@ {�yc���jz*B�Uy�!�D�V�[�L#$C&�R!?=�<�*3)!aJJ��;�ϟ��;�hn�����M��׭���8O̳T+�p���Ͱzi�lUXѲʵ�_i��O
�T�������z��{�ئ�m�^�}u^��f�0�&�T^��9�:@�1 *��a��n��'-ü&�Q~���Cx���i.kH�\�-:>=�L֐��B;��81�M�4U�mY#.�#&u�N2��ϐ�DU��lZ�8pS4��S�O|� 99R06�g,�4��n'�!J�@�)Hk(&%h�>�I�GF���I�,�y��ւ��T*��Z;c#d��E47v��>�_��7����;�����k%��3�A��&쟘����\5G"��&�l,>iS![KqN#��q��5͒��>��_p���G3m뼳�:��~+�7����
�kd攏���'�):w�+`�|֦;�=fӎpUo��+�j�mHr�f�n�b��)�P�H�<�^�X�Ҁ�ʱZaj��4p������j�+7��ˢh���T����F%h��>Uɷ��ǵ�e���
=!7/�l� OԫJ�87��&��p��%�ֶ�&S,��+d��L$.S���]X҆Gȓ����0��JM�a�'�+gz�זzdvP���)ʠ���\�S��|��FHq�t��u==1)�˕A27��]�_��Ex��M��G�#/������h�#%����#���^�ޙ�i�:}�%o%G����y��l�E&9-t�\��\���듅uۿݎ�}�����@�7�8�%�7<�â��d^n�P��!�P�;~%1���^pU@6��t&���x��]t��$@�)d�����M�����a�� ���W]~�D8���I�A���7y�:2��x��g`������b*6��%�POF�t*/-t��
H�b�� t�ϼ���[p̲Exu��xr�+�E/7���lJ�5��	�Ba��BP��+[/s,�b�#4��ޝ,+����j)?�׬#qfWsI�̒����2�<���5y`�>|�����]���v��m�A�;�@���F6!t�y���tӨ渼M�3j��/d*� &�;�E��t��̨*����cC#��_'�tn�ʲ �v)z^���ʘ�8յb��cI!O"ӎ�)���a!7j�n���%+�������'S�m�6����>v�196!T�:�]w��{~����cㆵ8�����څ�^ێ��Q�}�\����dZV?�S�f&�E�K�-J�e�Vb���?�
���PH�m]�=RI!
f����1�{ >{�Qf����jG:C] x����^G�]V�q� �+G�J3o�L��r�\W�V�ڧ�⮆>�[Wͩϱ�+eպ���\[����[<Nu.�JT)���;�<�S�9DYd����+�C��z^�Ê�LJ�K�?+����x8���4V���f��D".�2]OI���Al۶]]]�Ahcs��]�St)ᜪa+��>7�G�d�`�^&&S�2�-�T2*�m���g���I�Vf���['0��'>v%���"���ո�{��Ʀ�tF�ym���xuLN	Z<�����Rx�n���yk�1��� <1����F��8�Ɔ�����#u�L�����o܂[��m|�#��=L��0��(���Vӽ�ѵ;D�I䧠��s��799.B�K����p���_�	u������y'�{�3H�t8]5����r~&�Z�q�Ò��p�|���Ni/��,v��!,_.z~Sa\��ϐ�7��	���D�t�#����r�9��%��I���t��M$<���q�}��{I
hj\j٥�=X���gX�jX�l%Q�<�B�� ��@�ε.���a�S��|����9��22\s4�l@�:c�����yg��w᷿�=��o?D���M-��ꄻ�%HY�y���%O�$�P�(î"��j8#��E��}f�ǜ��n��02� (��"��=N�0�$�<ff8d;a*2��P�Dnz�nG#�zSjB_ߠ�ʹi�յ�a2<*�k�a�o�S����\a�Q=��p�>��G�k���TL�6v��%#�n��m�Ž�I�xs��~����>�=e,c�2RaQ�W�
}�����K�����&�
��?o��8gν��0�:�t�����ǎ�HD��UOF9��Q`�L^��2v[�]z�z��� @��	��-���9�j 7�|�Q��n�r`Y�2�P�ϧL���Q�V���;~�Ҷ#o%��*���	�Y߳�:�ty5�VV�4�g�Gq[�>��
ԼfN^��9n��x���q�Oq���
G6����B�3��㡅���d�������kR%Y�[�||�g�\���2��A���k�mLfCf"K�7 hs�`��e'�L��sIX�]H&"�I���:T[C�t��Gq�U��/�����hi�C(���g���=���Nh�-�k�n�G�$���	ᔎ`s������ؓBzt�QO��5W\���_�|�|���H��c������n�]w���>�@s[y$�����Y*޿p13A�X�&���+�˳c@a��GjŹ�[K;c�s/8<؅��H�p6�I��L$&���<�����z2\8��7���$d$a�D@)Ŗt�`�K/����Ź�\����	v�+F>'	g;]k4+5���i48�
��K���0	����)ŋ�� s�>GN��p~��9]�k��U�9�Rj�X��
`��2�S?*�{���*�ڦ��5�v
��μ���0�M�l*(ˈ'o3M��C�=��p�9�9��_Y���$h�8�O_�O�`������ʳWH�I��YCB⒟�*����yac��l
!?�|�Ǧ��K/r�Vʶ��<��hǺu[��?�@�xh�E���Mc�����qr�&W����\�m;�a�>��b�Fh=�R$�Y�%��c`�)'��`/�;�DƤilݼc�1�%�G�7�5#��6�A�}���y䩳1"Cr!G��!����OO)��n|����_h���[�_�p�������<u��"T
�=dE���%��W�����E&)�����W_�B�0�X4)��ˣst�o�-���U�.����`��/\LI�0���x�r�n;�b�U��/!�я ������c����m�9�?��2�N����Q������uH)tVƥ���ɏʨ{�ि�t1�%�f �=,˝�ta2 ���a7��e�����%⤱�sY$�	�����[zk��lh�_~��#���ܵ�$C����1��C���tZ����0E+?���F�=9:���~�.͸��ts;l�$�q^g�8�4<��u����&e~���Ck�w�
w9ϗPm=y<砫��<�"ҙ� ���gP���4�F�$�77����� ��C-yޓc3r}_������������-_����o��O<�	�Q,\|9Fn�x������!(p��i�s��!20��܇�{�A(<��7�&�8-]=H�s�k���ȓ��^�v-�8����-�25�=+Z�K\�ǆۦ7ף���w�	��kɋc0[��S*?�"��ꐊrȕ���%d6\C<==I�T#o)$�s٬���|eC���|�P��DZy���f�.�kE��Q���f-��0���V"�ف�rC��&Lb�`���hX��}�lzk��y
^\�
��<������ H@d�'�����O]q�q��ڇ�[v��!4�9]��DpX���w	��������lݴ�����?�ŋx���������׷���#K��g��J�/���#�ĭ7��X��2l��	;"�Boi'͛�Fd�ǐ"��O���K;X�$�#q4�2�����x��W�{�̺`ؼк�&����xk�N��o&�`������X�� �Z$��NY��J'=�lR�"����#9dՀ΅�ϸ|^�D_��z�����6G���X�m]A��%DaAZ�ٜ[�-�9�Jj��`"q�]l�C�[����ޜf����E)�u~T�v��̡W���>+�	�[��<o�I/A��
�]��r+k%�Nmf-d�6f?��7���*SˉG\z�2heA�y�`C��uV��H ���O���e�Uf�b#�,ߔ�p���떅�{&��/BT�tH���;)ؑ�A	�דbf��tB��ڸ��0�7?lf����D�_V�\���M�{�(tn�!/}j2���{�,���k�Ķ�o�#�~-�_��|�[��#I�އ{_SS38�g>�8q1y�6���I'��K��t���aYTg��xZI���gQӲ��7M�2�dj���4]G �<�Ç��3�㦿�;�wwc2#e6�q2\���
��s/�����k��CG�LM?���E�M��A:A��&�̹��%B�����8�4���7mí��w�|B��sA#�ˍb2�1�W.�g���	Ͼ���݀���}�y�/!AƇ'���`��`����bߞCر}j������ݵ�@H��9ܴF��H�lI��87���,୉�i��q{�@a�qbbL8
��e���Ն��yG�)�K�B��Q�V{��"d�c����*��9�+�KsӬ\yQ>\Fj�.�܄��󊕧��k?�k^����U�?4�Qwm҆$��S����$��>�rJCQ�s���*�θa6�O��"�B��\J�6gƹ��ڗ�`~{ ��q\r�b�<?���d$Ng|^���#Gs�Kkw~{�[���9gt�g�<��m�T��i^�8��/9�����)-52�i�E!���\�	i��7�������R��Y��}�&3� ��Hf$�b���hl��{?�^xy-|�2ٜt2L&RU��J�MI��o���0?-���j�RM����S2�W�a���)'���>��sPlF�3�Y�d��g�z]/���Z�O��N��(*��J�����J��Y� V
��4K�0�jh~�\\)��О*�?²���J��f��H[���mE��rS��b *��[i.^�AB�����T^.�K���ʛ�g�Y:���
��D�J�4y_|����B�Z��G��������T�.������q���+�SyeE���|�����������iX�s�p/���/b%	6���J�z�Iنp�����(C|f��,$D�uݝ�?��<�}8��E8q9)�P;���]yꩤ$c���{��xb�DH�3K�˩�}�ߍ��]XB�����7o���R������Ix�bxl
g������i:IngK�xd
vo��.��D(4�q-'Z*R!}�ɠ�{d�g�?0"=��X�x�]� &'gd�x�.�azܫ�<s���x�ȣO�G���2����݋$����,�Ã#hnlŪ�_��AǼ,b��$<J�r=F�3��Se�~�6���IШ��p�Z��d�Df��F�������EȰ�����x��T1��էla-��m��˜�B�Ô�9z�6]��+O_��O��e�a����D`8C䕳��$�5!��X��RZ 9Ғn�ǐbt;5�n�`�|Km�U�iv���IQ���t��GI����[�kΉO_��ݸ�{G�%
5Қ�eN���)�T|	���w�����^�����7u��I��@�������-���n�σ\x>��e+uтF�۷����;t[t�Dɀ���K��2onk��`����,�#�:���Vq����o�����Q�G��s;x(F���0d<� �1��k��[�]�&�v��W+�\n�NL����zsq�o<�]�j�[g?�cl�c��'���hb51m"KǮ�?��_6�I.S���]��:ʛ�T����
/��$��U��<G���}���x�G�*#�B�<-:W+�����Y*�:>�ޔ���);̺��Y�n��:���e0y��1�H}}�p�'H�����	�^��q�*/�d<O�΅�~���X�$W�ecY�w�2�on>�i�z������{z\��b-�~lh.�j���ؽ{�p�����k��1�;��<�ȟ�_=��uV���>�
�p_]�5l�l"̦&��Rw�Q�ǲ�=�P8�s'�676�A���}R��3o^�p�V�r'���Lʩ��Sc�$X�?���$B�=�ęc!�F�BC�NR��R�O���fx�<x�ggP�ə3��E�����0�%�����2��[P�F������Z��l4/�C��7fsؑ"����i�e8���u*�j�x��'���.=��p�5��܄;��/����g���MȺ|
�Q�CVs"�m9�3b�_�w��v�^3��a��h>��g��� 
;�#E?M�>�׃�i� �w2X��'#�{���`�+YAU�w�~z��+������\�{U_�a�A;��Q�ٴ
�z�����D>)�Ű�"x_��lX31�')b�~�1���ش~i�8<>$�4>�K"$ܺ�ɛ\,;hN�2e�� D�� #��Yyu�qmHĎ���t<CFp����!07x�		'��L��{́&|����[�+����R�d��N㤀=b���t.u@*K���t����ڛ�L�y�뎻�y�nLF��kj��� )�U���KpӍ�#K��'��ӟ����]h� eD�p����x6o߈���FgW6n�"-��i�]�t-�s��Jkeln�[i:��1@K�y�3�J�8��fJ�SZ��&/M�tx}���13=F�:D�\�l]O#T���,��ZD���������z�s���;�$�n�[���n�/�TxW]|�E�.�~3�L0S���mG��;��U*�w2��1U�G�>�޿�.l�pVj8��d*{.;�kEt?.!4@�84φ ��rP���N�8w��<���\|y�mhom�[o�C�<�F��t���053% ���mr�w������ۆ��>W@`=W\��׭����mR��X�4y~���|�4Y�����صe#>��O��{��G�Y�M[&��F
��Gf����������z=$ ��ؐa�K�k�R���)��xw{�3{0F��Sr/�ɋm
x��t��"�'*�~~��WOG%�����֏��j��#^�֨uTSƗHCC��B(�:�1{W��朧U����r��R�a�h� 	e'�+q��P.=�,�ՂE�;L����Ò��$U�n�[x��.��8x�	���sp�Y��g_@�����2[�.x&��{f����W���dT0�]�;��q2�Ô�}Lˀ/�-fp �Xxʫ��bڬZt�(��;�J� ����J�RC.,�\��ő2E_� R�/C {x�_�җ�*@b�=s*n�wl4�o*S�ق�b�p�.]�`�v��TA�	4�Pt��gh���z���cp�߇�?�G4��`��3 �1�e�l��)���D����5��i+N@s�C�����ޟݏ=��9���u!��#�8�T=��S��惒O?�=�����o2NF�[��=� ��޽�ګ���|��O���e<������t�P�-簐�92��;}��$���wE�]��S%�g�Yî(W���r�������ה�d�*���E�������ږn���Wכ��_۷�Sg.}'�Df�^Z�R�ڊ�,Nd���$W�̷�j/ݎt+Q�3��p�׌�E}��S������`�CW�̏f�^�	��̰�e[�k3J���F3�8t���ʷ�Y�si�ϸ�_o�T�BB�
��u��X$Ң��s�6Ց2w�1���,�YcS��	�۵�)eڿw}��
yD<>��;�L�ן��x���$:Z�pՕ��?�)�ǆ��gb5�z��`��U�=�k��0N;��D����}�g���-��BrB14��K�x�C�pl�$�\��"�=>'��q�o��t
��Z�g.��hb|DH ��kA�ᝂ����TS�E��c���֏�Ȍ(�LF'o#
���y%�|
�u���Sk��9V�"AU�H�����L6oVah�yrC�� m�Uƨ�~�;���C��wp�Ƈ�HE146��zf��04:��?�K1�8���4o�<����4�1t�%��OK��C�iS�C�?W:+yj!#�)%"t��nS.7��/���odf�HXA6�8�#$&������.F#WQhU�K1�Vd�R3���U��<;©�Aq=�-�w��u��S�E�l�q�nܜGP�lܱWI7��&�gn��=�<��#��o~CϪ���օ`1�~y��������y�,����$-Ygh̗֝_sIy>.��Ҷ���wlǞ}C��7bjj�t�c,?{��,_rY!���>��Y��BxG�ߍ�^]G�����C�Z'^z�o�=�����,[<=ݍ8��e����d�(�)��{EĤ�pKk'n�{����yX��rR4��0C�+���Nf N7�wg��������U�Vp��rfyQB��) k��܏'s&6J)���:��l�ţ1�I�򼈐!5�H��=�Sv��|�������|��S���H� d1Tp�W�̜p.N�Rֳ�<�RE]-�>����[h£��J�_<����ت���އR��w����(K��/׍1��W�85�,o]�rº�
��%m�U��Iǥ]��/�/\^W��V�����AB9�֖.��p������:�Tg�y�ݪ�Oʇ�GFuׅ|��ᖯ�k'BuAa�rz���s<OX�sh-N
��kS���&q�=?������')�C}�^I�~Ý�b�,>^[�g��2:����Ix�Iie��b͆������`���)pSi[w�񞆜́�׭�q'� �k,��$��5A:�V���i�±(�5�������)�Z�(BW]�7�
����!lw܋\����W�@�rfo�3w%c�ϊ5K�yV')�R��'���C�F��Sĥ�28�v��гp�<�V����~Rklڴ��8�"Ylߴy�qr�9K���:ģ�r's��/&�t+uS��f�.C�Zi ���J�Q������$�1�y_�K3��p��-#�hRks}^�[�WY�e�3�{ke��(�t��=t1�$,�q��(f.Elk��ȇ��W��\��^�x���D�����mKY��*	��>0���id�뢈hT�����$z�9�,�>�/���S���~iR�6�61æ�r��3X�ь���2-O<��'�@��ܭ#/[���������ֳ���Y�G
�|�o%�v�łu�Һb/�nc�vžx�w���!\v��x�͵�~p�,�%g�UⰘ������p�г�R��DD�ϊh|ȳм�>ǆ�]��M2��+ωK�m��X��d&zܡ��~���}�oz��3N8���IA��.{7��(���ҕB�4�BN���EC)�"^-�Њ���ʕ�u�������zN���5��1��1���sF��s���U@e�j(Q�W�����^��M��P 7+�]��к������s�r��l4E+ɔ���8v�ᩰoN	s]|3�y��3y�AR�\��%Q9n���6�N	��˲L��4���!����@KK�dd���!�u��Qm"��;���8T~�E��TQ�/��?�ry䍈��a���&,Z܃X�����zt㗿���o>�y�k��Bchu��7m'Ex4�G�y125�8&F��h!/~��B��������ڸ	!RV���K
j�,�Ǟ~�n�����^)�Ӥ�~���BԪ�qy�V�����Pmf��&!O1�4����&��Y!j�/:S���q����Q�ѼIrɓ�3O?	]����~����Ec�K/�Ɓ�}8v�
<��?�p�u��zh��NF�S��9��sƦ���eb(#o
=#ew�5�R.QЬ��ˏ��HI���fB#�Ԋ3�
���r�VG�J�\td�hqŵ\��T��L	��ܣ4�Y�aYq��VH�|�^�n��ʌ�a�a��	�(%�c��F<��Ә����L9��pМ���9��?c.�4�Z�3��D�QCy��rŠ̋�(Ҭ�����y�M*C��'��7�K���z��/ï���=4���k�s@�E����$.8�L���$ٺ�s��98���4Nk�W����j��0�`����yص� �d�z�x�rt�'����p56�����Y2�kh|�#����A��y���9ͤ+����^x~V�����b�%�ǜc?婗�EmEC*VC8�虛���/�.�P� �S���K�PW߀Hx������7��R�����{e�Cןul��]{�yk��[�����|V�W~V��r	�^��l芁�|d�sUF�{��k�e�U�yW�١@�Q���������7�}Ӆ���RC�j�*�q2�xR��G���PxҢ�scRRܭkɢ4Yl8,��<��5m��x�����4���s����Վ��~���зm�*�m����*y�5�&�}�[jm�}����J��8���w��6�aR��c�Oؠt�z����e���L���C��&/�?y��]*��n:�������{��m��H�p�����=8�wƧ��Kk��(S�v�7ʸ�ƢHE�ƺ�����Uʛ_��E���/zfj�/Uԛ��뛔&�$��)o�pߡ��R�(n=��!9P�Y����%�"$���p����j)�x�LL D^�W��U4���g?�6���O_�K�?��j46-������ٝ>�ӷkn�YUq���b�f<ep�7C]�w�0('�L<��K����I�I�&מT$G�����pu��+��ն��&��K>ڭ�G_�<���ƹQ�e��ߑ7�HD�x��ǟx�����t�^1���\��M��W��$c�қ<B�}S�'Gz�QP���Q���Ŭ��(�}����J�n�I^�o��/~S�����پk�lB]K�9�/vB���*��� n��E�:��Թw:ÑS\n������p�bNҚ��}b���1�=Ћ�]�ho����;��I����ؓ,9��p�g���.A�'������7h[���\��LS�Zۻ���d�;0�Y�\y�ּ����yI��s44[cH�e�f�Eo%���+6��d|t�d�3�ѓ����t.��;t���G�����'�<��Hc��,ӳT��w]@yV\��-У[m��V���B�V7Ա�)ZU�[�:K��j�1{��+,;�Q
"�|�e
�Dї	{_��sɘHxK 2s�f�d����:�۸*Nw�)M0C���_~��%�m#
8�����Z�~ �O8����p�g�'��?�N�1��a1ln)����h�+���1��a�񡍼|�ML�$MP�ǳ�?�yB���?�dʆ'�xNX����y7ڛj��{����d,IA'N>����"K�dj&�y�Mm蘿���M�1>��w�^���?N��1��&�U'ew	��}�2��j�O��F��M���1�5Go��1���w�6�iB�˭WU*B��ܸ!���L��@[sn���8��^=k�����O��#Ct�<�Agp�eW���{IJ���߃��ڂ-��h�'�K��c��`]�;evg$
�SݪUJ�� U�Q��)���JN�d��B��,QD��J(��{cէ[(q�U:
�>X�����������d=����I��H���8�X�d��H��v�{�+Η������sO?�?�s�H���f�f�p�
�)�+�j7TN�2,m��Y��]7=s���9�/�'�x+�<+V��N����k�}�V�5I�3)�,dճ.�U��i���{����=~��)����4yr�8�$&Oݩ9If��\�W�"��� ʑ�l.#������ͦT���p*�/w����S��i�l~��@�ֱ��_S���CӘ��s�2F�Li3�� Yp�#-��T1���^#�-�}4.�]s-����?�ًk���N�kL�r7�
D���|q��ٴ�L���˙u�*s�s��K-p���yyH��%�u�Ŷ��a�|�j��+���mn���A�y�Ս��y����w�;+��)�D��_�yAF[���@e�i�Y��)�,���9,�՜��Ԕ��6��[��Ң��Z���M�Y�}�ž}�0:>&���8r��8@�s	��� :ڻ0o�"�O�P؅��f�����d�J��3be826��>u=�߃�h������uo��?�C(M���#�J	�-�|��W��/���� �ں0>1�^{S��
�lF<e ��������G����ٹKP��W����p�y0=:������5���2��t�W��CW]��|�C�����@�!��}����0��)���@�P���X�h�%[ɺ�(5~U��ql��R��0ϐ���؂:�SC}��
c)��NZ,eGl��t�Mx�Uذi>���15Ex:���Q��v�%�a˞>z�Ch"#(��Ѽ�d���8%��$R��`+.����A�����
�H$��T����69+$��d�B�N�_�h����*�s�@��xG�ck&1�)W�2G���b@�N����Z�92:i�␚rfdR�N�A  ��|9�|s������1>έ�k$���.v�����t��؉�C�+��D􋑤ƕ3+
)����Z4�W�������܇��o����Y>����?=Ec�(���C�,��3�eRBZUC�3�Ksc=y����>RMI+^Ƥp��T��kh�oD�\�\�I�K��T�qf�~�q4��!��	R�i<�裨o�!Y4!�9�.͊�" В��"�Y=òwU6C��ǜ�T��K#��9%�jy�f�]S��bJ����cu��7���|)o�CRO�bfZ ;9c)z�Y�ǡ��é�|���}Ͻ�����~��)]3ޣr�6�e�rf8릔��5��f1I����}��ly��Bwj�w���0�B�Z� ���T*�։����ceK��K_�8���~[��S��m�֬s��?��bg典�A�P�Z3��T��Oܪo��&���<��S�\���̫-���d��^z�O��`C,�U
�=>�ۮray�yK��PL2��=�w�<��s�8����ɻ� �)��]N?8DJ����x�ŗ����ѾL#I��'���3r����j9Ԕ�q����uX�r%�w��$���i�v�s�#�s������74��{~������_���>��|ɞ�X4���,�y'��U�Qο����{��w�(�,#��0�<L�����1�����h�L'�hv1:!<��}��p��g㟿y�oۍ֎$�(��d�8��!��y���o�T��8$�bz���ڑ&�&)��	���`�	�Gd�H�R�Oyjl��O�A��Ŷg���V�BK�[x������ ��_�2^x��ܱO��u��A��p�O�Ǫg^F������s��O�#E�$"����C@�����H�^0zs+	�0��ǥI]�����5`z���2��n2F���FQo�)�
�|���5�Y�}�V�0�4�xw���s��(��e����U���=�b=�58]�,�q6ĸi���;h����SO=_x<ֿ������D��'P#t�R]���i�0_���_��F�[�rcDR�z��'��_SK���f�pR�L�"�E����4�,�aAw2i���DS�l?0@
�y\{���{)�˱���{�4ߓH�G�y�1bH�#�� �%�Pe��=�n$�������R=��q�y�r#���A@�<u���3�uqs�����.��4r28�q��Jk�G�[���q�5/��dT�W���V���#�� t*��\�����
ƃҝ��ƘF��g�o�������`�4,=X����ÜVf��P�C�B)fz��2�T�R��g��+Ƞ�qc]������L"��N�۶t�����gk~kX�h�\-�:��$4�:}��
�gy�s���f����X��e�0Een�ͭ1���2
P����*���/9f�w�c��BY�[�Z6�.��ٌe-�0Jĕ��翪}a���"��p �211!���x�+��g��T�,U���-C��f����i��m��"#��7)d7j<LC1�L�:��={U�?�!+���r��-g����y�i�Ne��Q�i�ߨ"5���zq5F���������_�w|AF���t��ޜ�����8���;��\xB�����#��6��&@
�%�,�����~��9aE:�~�����08�}�c^O;�/ ���_�կa�{N�֦�dƤ�%el��Q۠'믅e���vy1<4���x=��-�@ѩe�i�(���
�y6^��%�nf,���{8��Ex��Gqұp�g��G�HFa<����f����'���ؓ��hd3=7��ٵI�Aw��� �����^վ�U��4)�D8�hC����|�S���G��|E'A�ڕ�-�T�Z��\�ٯZa�67i�=!�y��T���hbQ�eTe�0_��>��v���6�I�PM��L��"p��y�'p��B^m7M?)i?�4�$�g;l��f�&�3���ӊ"XWz�ˡ�C�}��Eɋ��1��3�v�Lp��&�"�X�����Lq���#	�� ��>��=fN=���{7^��/@oJ[f��ǓQ�R�4?�PL� �t��s�Q�vGFR�6�kb���33�q9�G��AG%�@*�j��>?� )����q��q��^�Q�,mC�8u�X�z=F����>������T4,kU��M�g�-yn>g��&iE�f9��{
Խ淅�[��|c~a�ߘQWNi��uӸ�%$e�+�c�e2o�C��kYi�*�����'����h��X�z��t�~�������GO[��t�!�U7�T�("�5k��[��@i�C�շj@6k+�^����R��fy���{���JB�G*���J���B�[� �/	�i�җܚ�&+'VH\GΔ��}�D߱Pa�׳B�Q���\�Y:���؜�R8�aZ0c��X�l1z�`��C
m��b&2��O>�ƥZ�Fci���(�5�2�P�WDf��СC8�o���k`��������p�Gh��q��R�L3������ ��vn�����4l�ER�2��`���y��Hhz�d!�\)un>р����i��T[x4�4��㇏��'W�R�q�!�%#6�&ለAH܆
e������3���}t]q�\��_�%��;
��P���4H�L� �wb~G�9R��.��E8}�2d�N��E�N���D+O;�_��^]�u�w��uZ;�Kۄ���ܢ��x66s�$&/�� T��pASK���DB<��V���om*]4;�&�_h����fC�W��Ў����Y8Z,N���S�1��o�c��S���&��3Q�8�n���e�V\}�54���m���s���2���-�n%uF_�HY:�N��dϐw���ܯ��4�;�&������-/���p��<�q�ٔ #�p�����w߇E�9��V,�|�6�E������2)^��l?�ܯ��������xs�^�OY9�������5q��I�䡹�����9ˇ ]�v>�h�4�����>�V��h��zE�-Z�;v샧�/J��H@iTcbLl��k��T�k�ai)dKgY�쪾�\��T���5yFJ�@Z��&	�Z*o�拥�Q�yk>I�߫�"1�56qqI�1����u(|C>K���t%��%[�~"����_���k�8v�5��B/�CW�B��(�k��EW��K߿S�j���!�K�;�B�ɗ�_P���+*�⹊�1G�	����ǋʴ�˝_*���(BŻ6��4���E�)tk���Kj�9T�J	����&�Y��E0�t&+a��P��Cdy.eF6Z�-dM/=�X��`��t�9�0�MOプ^(
���o�_Gg��&R ʡc�ӊ�I<b3��/~k��n��×����Y�o��u�8U���������hMM-X��-��w`O~Uޣ�� eε�^?ӬF��
j��e�|p`X������=t;�8|��������8p��&������5��r/FgHs��)�]�3�KȌ;D�P�w��;��0�0w��f�k8%����5a�mM�&�1���݊��xȀ�ۃ�z �#�hiiO��q��%���W����������������g�y�Z�{}�wj~�;ڤD�;�u��}#d��y�����ܜG���E9_�Rk}@��Z�G�y�u�v
ZyAYX��ӎ�s�b�qUF����N��:��>�{Q�%wc70�$��CB1�� |L'$@p @�	z7�܍��ؖ�dui�Zm�����s�{gggw%�������ܹ��{�s�sL��[K0�Ր�K�mo}7����������(J���dZ�&D���܏|����^yb�� �|�c�Č(��z�<! ;�B:_Q�J0ƪ���&�q��}Z���/�09����Mrm1<��>�y�Cx�/@f.�׾�5��F^ε( �tؤ�%a̱�i��p���Ϲ��x�܃c�sr-!58
���r�6q�Wi�g���"���СC&�%�7�=����p�8����#���?���HX�ٌ��y��_���)��G�+dB4�&W���A2O���02�r�vI���,G�õ�C]�u��}�֋	U\���FO���/R���D:��
6�n�'��g���e-[���K��~58<^��tny��ț���&������k�}�Z�N��U7��րhm��''Y���?��jVw��V.����v]�����b4\C��ʵ�H�z��h�7�⮖������\��K�$�-7։�;*w��9�^=�;��=�5O���I�i7k�R*b��|�(�8
���&��xva^�q'{p`�>�/� ��~�(ģ�ۿ�[Q��aC�z��ΰX��l}nT���3��,n��V�亟㑇�>��>�߸��<�D���.�S��f��T5�k��G<y�Y�Ae=5;�ۧ!6����U�~:�HT������j`!����g=�"�ҋi��kF:�WW�&¹"��n���l�
˧ޒ@(��G���-=rH��i���������x�A�i!���v�h6�>4��Xg�]ZS	�ȫIn������G�H
����_��=��o�s�#p��gZ���/������G9'�<��G�mm<(	�4�t5���Q��P7���i�bޮ%�h5�:��\q,�����і�.��Uk�-	���i�~�պ�V�j�W]+?��ϱ�g��ʰ,&vkK�v�0�+�4;��d�T�\Ǣ��f���㦅�ʏdF~+sg]���Sh�� ���jB?y�ӓ	����F�'S��:`L]t���9���<o�=/��s���/�y�z�yj�3Y����W��-���O���CcSx䩧��y� �ߌg�s���� �п(k6'k'��.�$�>1�� ���~1Bv#��>�����Ұ���r.�ĺM]x��A;��_��-QL�����^��*E�9U�x���Ӫ��^��n!��&�m�<��nY�9!��}C$�Z檷+������Jݵ��#��bA9�INU1�$Øz(�Գ�����E ܲit1���]��߽��w]����\��x�x�]K�m�G�RNd�O��/�� �j�}�o�c�7*��^��n\�ދ9��՗�9������]�-�z�>��i���ն�i��K����^�f�����D��������'ƮQ_�[��_,M2Ɇv�k�� h������ZiTT��X5�>E�G�#֤9�^�ёy�y��4c���5���e��W�n�L���n^�|c-��T*���rڟ[sĲ��wb\\��l,eab�ˮ�(� eO���6���GG1*V�8-u��L�Bsԓ`�$���/e�S"I2��ׇ�ьh��/@&''�~���^��k�RȦR:���X�r<rk�þOh�1��ʾy��P����|ǰ��b]O�˹#PBڈ�%����(�&f��(R�G"�Tf���"�.?ikS��u�T�i�ET�bn.�MX�zrz���"��8�b-�a5���g�k�Q�l�kU��L�J]��*k�O⟉�p�;�\Y�/����?ρ㝨�Vnj�1l&�)��7�%Zb��	�G��Lr
c�Â�"��| V�h�Æ���˼<�(j^���4~�����@!9'V� POHt�W3�SI���p��'c�I[T�NMqt�zUS2�y�W�z�`�cXL`���ɜ%���o@�F�s1��.�e���%��`B��C�����s78^��/��w= ˟���JG���٫@�kqa
��w:�w�s4�a۵w�R(k�F���
X��u�iC�L��� @�s(�<��d̽.45w�e��yl����洐`ƲcרӶE��U�!�Ly�
�FS�r�ɬ��I2v>3�Bs�ZGA[u�qX-�3��C���m=�^��}U,��0^�(&����B��'Be����
�=�O,�jᦻ
?�~ɳ�Jf�V��s�o��w-Ok��Ďw���N$�Z���#��j5kU����*��͇�l�J�V{\�mnN�]閮�TSz��ʇʐ����S�Fĺ5Y�~��T!�*�P�O�2p�G�hh�S���Z��Q׳i
@����}3�=���$�zj���(�2����JG�J$Uy5�#�7��>8p ��8o��V>8����M��qv�ʵ��b�DJ\�4�����&~��ݚ[[DaGLL��mALj:�Ҙ$y���{0=9��cg9�����c���==5��"!�Ef�'5�������u\��q���ג�|Ny񙱛N&DH�Bn�����(��I����ԩh� c�n�5&�|r옜ǅX��G��.����,�y C����k[�S��2���8�S����ħ?���9W��b����}:���%Q���g��%�%�mwދ@�^Ļz��ъɅY����ȦX��Y眎7�����7݆��Xy>L�O���!�YTR����BǃU]i=��fy��۪ᴺ���G�ǰ���6�s��,�%�VU�N���U���-��8�H4���P�Y�O
?��u���oG�`n��.�t�@E4cY�眀��?d��p�����"6xq��꥗�_�*ʲ �\�,s#J�/�Do{ ~�ho�j���ݥe��8����6e���5٤�
kH���z�{p� �-�ƿ���\��'�]����V��&�����|H�Ȧ���׼
�o} �Ez~�|��("?���o|ݫ���f.��S�!@�,�Z-9v�5��D�z�q|��O���<��7c1[��閯���U5F�&q�n�[��pP}�쪇ZVy���,;�N}��'�\?%��)��y��ː�ya�����hQ\
>�OU6�ͪ.�ճ��S��ږ	sn�@.j���&V�4	df����	�����^����Nϒ>�[Xu�K���V�Xi�e5?�{�}�R��q����5�c-�ڽ�\m+=��H���'�v����r��3���5�]���d���j�ѱ�{��Ӻ���ķkI�jͪ�8�mM����B�^ͥ��<.�B��9���~��E�ݻG?c�yfjͱ��y�+�w�}J@���k���b��z�*��>����^�H�d�UiK�(��i%O�5r�͊�H��g�*JG C4�u�U�b�b�3K��f>_@�Ń�YnD�e&~bqZ,���([/�ɿA~/�����j�]島�,�l��� �����▅Up$����������</��t��b�T�BgW:s
�G��_��9<�l�{ߊ{�ُn���Ø[(�=�\n-#�:�$M�G�����E�^���&��Lj���k߯���;H&�"h�*���:۔Տ1�Hss�<���U�k_{�<=���S���k����<e�uR�nmW{��2o��,�Z��\{[˓���q-?����D�X��'��?���3���A0nX�ȁ�&@|ltx�{q�s�C/�Į]ص�Ʀ=�f�n�"V)jYi��r"���d�k.���7_�
t�	��nO��-ʿ���p�˟�g��A�{	������%�ɔ���� {,���=_j��!�dY�C@��p?��v��m+�sFʹ
E����mV�_D����ø瞝x�姡����X��6�j����絤���GGG�z����se�� �[n���4z����S�:�X*�q��׎���x��x��G�7+��$R�5ϐZA��TÔg�!S�;�j�Z6������n�j-f��$�]K����$~ڥk�#����q�3��R��.�|��b���v���#Ͷ�cN�%�I� ���|��������|jmS�h�&9zP�-ܟ$����?4�U�]�{ܜɉ-�7X)�9�+���Z:v���z��3gOi7���7��N���`V���Ƀ�{�9�Q\���sb�e��D�0�
�Q�ڝL��8��sl>�e�"L�S�Y�,�ZVkŸ���
7+1Qv�`�B0�ևIӨ�j,q�|�}baA�z$@SS\�ҝҰl.���XO�Lo9�>�-'��Y������F��s�R]2���o�qX�H��`jr�hD;��<>��s��Sb��eF�	�l��A��Y]X,�#xJ-�k^X��l6-�x� �#bi��/�3v�|_���7�J������pp��׼���7ԍ�ɏ���/p�o��K��^x9~��_�\XԞ�`!Q��-����WJ&v�g2�XW1�Y�Efn�����b~. h���X�Q�u�>w~���05Ɩ�mh�{O�N"�+-���(x� eQ�������.B�q�lI�\�|�2AU�����ҩ1��#��c��O�<Ib�ͮ�@���H����#������a��i���y����JdD�W�
�)f�+)Kue�q�.�̪���<��w�oW���������˭�����7�T��4^�֙0_��2�&7����*�F�o�-.�ybq���J�!�,��vQ��ڠ2]^��t�?��M���e�oBJ,�W��p�e`.��B:����V��g3����x�ɽ���	�K�h��TUɱ����Qy��f�,źq+��L
?��-8m뛕�(qaN@���8b��13��߅/���%���F]�����x�%�$2��n,����F(�A!�'��;�㧿�	�~$��U��OeM���oǳOq��6㳟�WM���u��ڥ�N�)�<��\����1��F˦�($�!�{IC>6̱�m�Dgd�G-q� p`���5R���Τ��Dd��4���P(�Ch(�TQ ��(cc�PR#���:`�
��pXv7MNyZ$�I�%9.�9s��7��$�b�/�;[�##�rK��e�P����e.��%ɖ�a�/�
�z䔥,w�x����+]�u��۞)�^��,o'�k�����}�K���mU�e�2�?��ֹ�zKݴB���S�NABdƤ0�}�?�;V�|���N}z�2��cВgi�r�G��x�{��!�`ᢋ.�駟���S�x��_��ﻚt���+^����+�)͎��ߴ��ߔF��=Kvbh!�I��e��c�t��d�r)�%��5��_�"��ݏu��-oϾ}����Ռc��E͋�� ����&���駼PI:\�:�"��i��(�����p	T3X��"�O��_+c!o�{�� �L�d|�8�� ���K�Y�%Ͻ �\��O<��]t�>�C�Ī��kt�%W?��uho�aӺQ�%m���We�.׿�0��
̔���RK�� ����s���L{[�X����[T�0�Xw�&f���kEk���J"lDХ���׾�O}�}����7���8��}:��1n�����z��s��ջ� ib�0_;�خy���3Y_�Y��[�+���ϗ��N|�Z�a/�#C�E����KTrE|�������r��m����V�����<�l���1o��>�_ė?�I\r~�ơcM��9��j@�^ԥ�qE��¾���$�%t`KOS!O�̩91GC�82)������N�\��Fs� n��l����U� �(�d���l:y��׾�}�o�i�j�hӦfxJ��g&6�ɫat�׾�_��w�ڷ��Z��F���2�� c6ikf��]�ve�<:|@���ہ�61ed�K2��F%W9�v!&�"�0���_�	���Ȩ54*I��
̨B�X��#��3�E���>�A�)�Dsc:N}=�X̥4�����)�*��(����t*�9�Z�U��=B";�[~N {hY= k��)*�?[v�]�|9WdV��S�X�LU����F>��>6�,����In{&Q��]�0KN��R�WOe�(�I��Ӭ"�����D�?E���X��Ev<��L��f�����C*�<��۪������%��\�UW�VY��[}�>*z�Kw{�uO�<6�(V���J���]M�����2Iv�tڮ*����f:�8����t��D��G��_����g�����5#}��Q<8�K�bv*+\�#�
�ё1����vUN�60vO�H�TLJ09Ӄi�RiN�'>�q�����+��o|�r��}�1��������T��n�@bqQ&{	���x�Gd��0�Ձw���X�7���5�Ͽ������#,�7�����(k/�b�"d���Q�E��s7
 "
�t'o^'��G�s9Ə���O�s^�P؇����U���K���~䭸�������r��]&��(
�~Q�MX?ЋB2���fxeP��� ��D�KU2	���Y���H�ĺY("����"���j��=����}I�YSr��`T��ҳ�h��ӥI]<6C9��8���~쿕C���V`7|Y=�Ĭ��kϸ�q�m�e���X���8�嫎\i��w�Y[��.u�1΄_��״��Z6�.��<
ZbZ�O�/!^��g�8=���qX�&�X�#3�_�#c�2�!L'���hiħ��*6�w���|6l@kWno�S�ny�C�w)��~����D[�r�h�����w�ig�h�ER�]Q0����[��VEM/f�����w�&�uZv�;�)Q���z�lƞ�G�,V���)|����������W^�BS M�&g,o���w��=�?��n����af���Ee'l�
H�BO�X�� >���ų�u:F���<�X0���<Z�C��B��ط�il��I�7�"�tva_�ݧ(c$�u�HP-W&�ƚ*X߳�n=CʫQš�cJU�86#��[�[)�Bv/����w���I���c���/��Y��W�C�;�Ā��#���܁�o����cc�t,/[��ݐ�gSA��h@�^�<1����%#a�p�Z�1=����j�B�[��䋕�b��S(Y��^�����e�U@���?����<�
�M��ˈe�&����Ol�Z�[+]f��WS��$~�8|=Z?^LoY2�*�Y���Ǯ���\u��h�;r�CQ�A��YM򞂘qؼ�y�1�(kG(xd�3����L	��� E��,&�M�O �>����HX]���WW���GT�45�h?�p��b�7.P��鶢�H.&�^�V)�4�M����Үc��,R�x�ؿ����c�֓pˍ�k,�eX��¿��oڐ����=�h�]\����|B�>u�?�����L0���G�1c�ϻ�%�|*-�z\�K�*y�Č��+('|4�G�P�kf������<���W���}w�?��p�M��8����+^~��v���W�?�~=:$�i���q���M/G���SO=�&���>�CC��jGG{Dk��JT��ɽ,ؕ.�ٳG�1'�~ljɬ\wƍ�'1+�  �&PYVD���<�f�����=����,VF
s�3H�spf�S��g��tu-�J�dWL��|�JM&��-��6ֶ����r�v�֘Ժ�\���q�5��������(�vY5�bJ��6?���[��Zp�-�`릭�"
�֛oFP���ܔv�#����1?'뤩I2۳����������Ǻ�}h�9��3�^���E�N��oj��+y�������3��羀��v��z��3(s��2E_��^&�W	a"Mm82~���_ŖM�{�~��{�� k��/�sJ2����~s;�o.<�\R�u<�������plbB�j;
3.���yK��u�*��ʜ��>�Yܰ�6�w���"s��n�����+0�ӌ�c��=�L\r�EJ �\�����ty�-x<Q� �0GDdD"���ܱc�:���7�������E;BF徾��o�<"�dg�v2>~�[��������W��|�����ԍq���o��z#.|��q�٭��!Q��T@ɕ�6�u�`�f~��e2�*4VR"�Z��l����Z���O�����]x�tggg�{c$,�*��g~~:�㉝�=G��Ʀ��rj&}n.]\��|a�R�h(�I�e֫ەT%��]�v��~)ɠ^�/-9g�/_��Dn���*Y��kcl�ѕ����Q�����b-?F#ǻu�{r��9�rE_=��T�TV�X
���n�gL��c�}YK84�Όv[ٓ,$#S,�r󵴨�L���!Qˎ������}}��O:	�G��#�'�O�g?��bE2��"�Q�!�C��\'����NO��z��V���h}�e�>-(:'����*��U �(δ�G։ωe��Z�l2���,.$���G�d\��s�ry�Du6�bflB�Uiv�Z��!c�k����+��%&8[�>�� y*�trˇ΁A%����T�Vf������a�ob��w`H�W�������E�:?��^��E:��{��R�k>Eo�_� ��Æ�v��?6�Ύ65Lf,d��>�_{�gGA�����pthN>�B�}��/��mL����� �����y���VK]}�8����������6�A�3]����8��Z� ��!`2����5�e�.{=8��d����X�"��!p| ��_.�}�<�ʲ��c�ZZu�!ˊa��Cye��JY����[,�tw��o��q�r�=ܸM�� \f������D��IOՇ�ޓ���	-C���������,�Ɉb�-%���bS���t�\�Lb[?T�r��Le��{E��㱧��={���3�)[ry��ᖵU�����܃Zi�r*�M�����.Ě��D������bo�iEX��k����Ɋ�/�� �.j�K9��I[�����	br|�pge}$�舯��䤶l���|��� ���<��&��
��9�W��:��y��w�ET ��c����cW�?z ����)�^�8�O|�ø�SI�m���/�1d�i&��x���^�����2O��q7���f�����L��lr�Xfa���/>�{o{��^t�����q��]��������'O=04������a�W=U+�k��ء�u��j �����J�"p���ku��3���s#����ZR�N���}��s�s�5-���״����������b�^�Ejc� _� y|&E9M�?w�}9 �L�m����Ě���#�1Mx�gYS��Vi�뽀��YY�������zח��%X7؏�>���
�M���[�&˸J"p*K��X�R�3(0q��ڣ���?.�h��'�%룵.��q/9�"�msT��*���ο�(sZ~OQ����:�4̄�8Y{_̢��U��('�ב��{�G��g������Ca( ��"����7,י�����i�D��7�i�%ފ]{����뤐-ȵ��qp3�=44������WLC�@�X{p�駫�Qe�u���֖�(�$�'�g�@
�Cs
�ȫ����I�x�Z�H�Oat��֥ҳ��ԃs����"��iAV�L��a�=!�In6o���`��'5��V��0:�sΏ�lw˪_����*Wk��㭛����|�mE��a�����q�9ޫ����jI�˓�̾KM����ɞ�����N�k*L�]r﷈�DjF�<���|=N?S �͢����㲆�hn�cxK��=��1��� ���X0�X܃p�M<���AΚk1�RF��eߨ U�v�H��ydcvgGz�)�{YS�ZX�O�Uݪ���.fgd�th�"s��qNX��O�]�����
��L���[A���&�=6���VY����-o�
7ߴ?����Ӄ������YE!ΧE+	�L$�d=��;��q�Tř'o�o��Q���-&qp�8v�:Z�PI�>?g�\�j�b}�ǽ�>��6��
pZ���:p�mw�z�)�-��T*���}@g�#��'oڈ{��G�'>�a|�c�����"K�f�0(r�*��)T�yص!�۴�-�L��ۖON�,,L�l��o{�;������c���gp��2�͇~�w���9���=�wd�*��[ᨕ�9@^V30��^"�-��z��Qg�׻�K]�H}g�ot��E[�~9�]}kt�7*��	��߯v����k�����*Vy�X����?��fj���)V]��P��s���:Z�V^���{k���v�Wpa����UK���$0C>���Yg���n�>� �Zڵ����Q�=�4>�EY���cOa�c{���Ȓ�l����"JiH����1��`���7b�w�,�y��WD��L' �f�WL^���`_�
��]ޗ�0�1�%I��,�a�	A��G�o%Z�A��.��]�����E����M�P�O`o��!�,�ydD1�se%��l�O#'��'&C��)!��c-r�M^
��Z#�˖񜋟/���5��翾�s��Uf.�q�:�L�jY����4qqL����X�C�861!�nVX�d<��S(2K��YQ�\����-T������GQ�s%�����.�(���Q�Jf<����f2�+�hLݣL8r����^[Ku������WW�רPW[��V�����ꪲgi}�����w@�j
]?/W�v�.s,��vV��(R�	V���X�)�~˭8�`z2��C�ϻ@��.�x���jk��:�Păb)��a�~����{qF,Q׏Gk�	��D�_$38���AV�?P�s�Mu<�����C^�\����v3tU�ZOd�����u��b$��s��\�E)W��hR)j�r}�`��Tr9���\ǎA���}��hoc�奸���S��;�)� �Y$� c	�`Yݬ�ih�5�&,�:��gk�@��DUqO� "��Ք��(O�</��n�Te͍ܫ�`� ffS��ʰ��看n�V@�z�]!�X�a���!9%�4+���V;q��7����߼�=XL����BH�i�MrB�+���P�*��v$,�%�R�L�W->����_���>����h�v��'LǞ����l��?�g3o�x��2�P|!�W5ϳ���3�c�3,p'��R�v�q����`���쏍��o��z5���k��9�s�j���/�$ˬ.4���M�P�&X�DW嶺w]:@�����ٔ��t�Zs�V���]��%�%w}��-�7�G��ˉ�bi	k�Mͼ�KB�.�����u�)���;�u�6�eB��ك�Ͽ�=���� sO��iB=���yRu�2g��a�SZ��[Io
� ��V���I��g�P$�������}*���"������ƚ��+�+eeƣ�B��E�Lc���f�s,��b���Y�,wa���z��8���пn��s �~��(��^�m��b.����af��Ӥτ�&�n��#�+�x��g��o��������x��6���`��!L��s�Yk��"��ji�.�	�8���S!�ԐX'o٬���:��ٜen���7�9��-�\k�J�#(��bA�!]�s�$@�r+f�j���M[k��d�S��d.&�q��嫻j����]G��U��	ֽ�[�WΫ��՚��"�]�*�*6�]=޽����p�V����+]�|�C��iŴ�+�Lw>z���� ���:$�y�����cذi>���#!��?��7��-Q�m+�̪��vq�LKfry��e�g/�3X\HirR���L�a�Q�X��GP!�0[����J����]%s�r�ͱ ���$�89�#��v諈u���ĒmuiDN���a�2���nS6;~���w�̫O|�j�߳7m���Ț�G"+V����(�hk/2�C`GɹY�Q�_�<� ���pΖW 1�T¬l6�6����O1)N�~[�RU��J%���a�d6��(���^�����_`Ӷs�����Q��!t��z"�:�\�����`�MW�b-͸���W�r���o�s_����g3���]�� �������%=cBR�G�9����Rf��˯|��H��o}��G>��~}�}OlZ�'�v��2E%䄗Q��𔝖�t���2-�ʖ���:���KV}+����Y���X��Y�Z��ěk�Yj;����v��Pg *�:ۥ�,5��]�cm�����2��\����F(ee�Z"to�ܮ�  Gz�xx�&.��D	);P���EA��H�I�b�i9qc-)Y�����(�g$_��#=��Q}���X���L�mE�y������vc~a��"���E-�?!h<��H�gw�EH��&� �T�&�ٵ��b(�c�� �����K��TRr��(���X�mM.�h����H�����l��ʟ�o�� �|��*o
TЧV�Gv<ޤ��G���E!�S�qGR��5*-pv�
�<G�>�&R��Rs6���^r8��6���ߢ�������aL�MMϡ��b���2��/f�bc ��7q����s��՟����C����И�5��6؎#�X�~G��f-�N?K,t�g���6	E~���e��9*e�X<=H��2����hj�W@˔h�{~F�n����1e�b�s�D�l&Re3�*d?A� z3z����� �y&��~�%>���V��x�4$d�_V����v��K�Y��Y�PqR��kUk�⯭Dː)��ot��vs�"�F���=�X.�V���N^신�(�	�m����d��3f��1K�e���xt�U�J�J<5<2�+_�\�*�u?�)ڻ��N��#ò�"c\����r->2��m�Z�i���y�c����Q�iK�\s�Ó��r��0��#��*�QSO7��rF�'��2�.���G�xss�hi�c}�z��w3��Y?��a�b��"G
2�{�ؔ�OO�U��*���M���M���?}������|2��'��Kd'd3)wP#{),LM�#�Ʊ�Q�c]D��R�駝��Zd��L���]Oଳ�+z�Z�n�HH�KM2A��fe����C׺������O����<�a,�������܇q������w��/8?��;�"��2��v�=2�o�h;�z���x04�$^�bZ�V�Nd�ύ��S�[E$�OL?y�9�n������̝��/:2����G������4F��+8A�LV�f��hV�-͊�d���6����F�����^-��D�;T���_8�R��J���7^K�Pb9��zr�v�Q�5k��P�kXV�ᄎ�}>vP�2c3W-��R�Z�a[ne/�~��i*�#����p�}�Ţ4��ڛ<�Lo�n���n�>�
�Q$sb!��y�28��w�ua�9t~Q�Lؚ�M
Zu�u��o,{#7<;�5��)P��P�����9��ggTA�ejKK���&�}��JGI�_���?��%�oF�p*����`�7���V��t��y�H-&jnc�b����s�5�t���$�L*���@��<���w����ǰnp<$]�G�-��ڟ}vnN3���	\������at�blj��_����=�@����v��F ڂ�v<����M-�6�8��c��G�[�ǎE��E�y�������$ ����F�V~�v"�ԃXs7����'�ގ��������D)gd��mL�̊\sY��Ӱ5��9����N�Qτ8�_�T"P����/
 �1�h|�g�b7O�S˩i\7N{�M�2͚q<�䫮����%�J�?���a���7\���m7ծ��be���=Nb1-����ce�K{tr����e073���Z�����/�������u���S��##���,>����e/8	?�l�����+�ϻq���W�G?�)�r�)���^��q�>}��<\}�;�r���n��������l�͓���|��·[nًk��g�{>��w`Z�ϧ?��شi#���+�Q����ۅ���w����ħ��ӻ��n�6�����]�v�mX����"0>!�@�m��1NN��b���݆�]�G*�EB,�HЭ���X����`Hk�]�6o��0��|F��i���u���gIǾ�� k��q! k�gp��&,,�p�^(묨Ի=�R9�׭^9��|��kq�g+���~y��GhkmG�D.I�"����H���0��(��n�ie�37!P����.g["�߽������b{����gnx��}c3���ʛD��Uc��?�N�:��L6ザ�^m��ǘ�Z_�>��T��K�y&n�g�lW��|-�]�^�X�����V��~ո�D+�J�3ԁ��k�#�����q;t��Lu��ܧ�����Z�[�|¦��S	�r�H�f/��1��\"!f#�CJ��/B���/�B0ք��y�u��<Z��4�ҙ�)4�"�"_L�k��B��@n�����HD�T�T���4EE�K.�Ё=xz�c8u�VQ���^X0n�b��c��=�b��C�[�c�NM�����9�:7�3Y� �xT=]u�>��-o{� �&��}�C���o7~)V���'U�55����`�c���F���wxB��!-���p�M����C"��y��ZƮ]q���޻^���f0+J��2>̔e���}��2�{����׵/�Æ-��nw�FǓغ�\���[E@?O�;*���5��P�[�]�mH{��@�Rgw�nP���+C�os�zTѰ�KBS|��3��_�Gk$�Zj˸�>_���n[�ڝ��WmM�.Qm�i��5�����R�\u��%�PszS!��� G�RZ�+���"+�n�7�o]�]����ᡇ��������a��h\%�ZzTF����iFK�3���q��D� ��@X&����X��m��F{+�|P�J1���$Gٲ�_���
�Z�w��mho#4�\kK�q�����4�J.��2��w�CQ��;�PXAF� ��*.�f�kF8%[�j�D�bN����1�D���C�ə4�Tl�z:
�"ba�(�Q�P8�y���2?��)Y��S#�U/s�E�������7��`�b�?��Shi�@쒵�B2#k=��c���#�SW9���fh��ۻE���qlb3wܫD3.��4���;����Ɔɞ�<�B�T�m�����7�`��M}s�=�{j��b�]�����`��E�W,WZ�Xo=W��֘��e{�d��7+?_�'��/K�i�l����s�>ֺ��K���|�5R5�^�J��Z��2�Y�v̸���e��2�tV��0���` ~��5]�"�M)�!����E6��g�������&6��5���ړ���׾㓳xr�^���b���ǘ^IiJ�?��t���$
�K��^�i��\�����wzDY����0;9�͛7j�����I����ڕE���q汝�}�Mk����9<A��}�)H��2�=�����%;������+��^������c#b���q��AX�p	R�z�����CQD!:��w�g����n<���H&	����������R�������d��|����%�f� $&2�ծw�HL��C���0#����7�k�����Mv�}Zo˸+W���rT�B,��V�z��{����jB���[��,0*J�� %ψnE�?��`�T�|w|��V�Y��������?�j2B��.��n��$���W��;i?l�Q����@ݡ�5J��q� ���܈G����.��!��wR��&�3_��o㞭���1w�_��q�Y8tpH�[��ݟ����hE���~���
G144��bIr��+�ф�_��&LL��_���[����{����o_�����8� ��x;�6)�}�{X��G�j&�£�������x�'������/|�{�?��dw�o��Dc�F"b�W��A]Ӝ��5�j4��'k�Y16Ƨ���Ş�192���SNވ���&�-����lA���?�t�L$�:thH�Eo}�{D��ٳE��aAQ�|�"@X��BR�SM�n�J�SA 1t��\eK����ѱ�)9�U&�M�6�*��uϗʥ�'m݁?����t��G�>�B�UФG���q[.��N��x��c�J�jӸ���Lz�]������u�x���5X�g!׶��k`���:��#�G����\:���u��q{���j�>Ӆ�^�W���t,���U��2*^���-���8�R�V�Ӑ�Y��EόP21�J��Y�u��떅qҖM���s��#;d�̨U\�urj��oĕW^���ާ:]�<�b:��x|^]�s����f�R��;�/-f2�Q�2���
&�T~�� �o}�[hk��=yE!��w<�K@	�MC���6=�&��rvj��A3o�&� u�O�i���\�����P�2
Av�{��^��M�N�1"�`c�<�}��]�Y�%
x@���`����<R2>%Dcq��+������X�I���f3k�蜜7+|���\eva
��=<�
��� �W�����$G�y$҄\z�X�w�]�TjJ�+/�zPv ��ڽ�����.�����3�[��Ͳ�U�1�ԌfQ �HXKz�;�A&ye{M�k�k�����u!r3ŝI��0�c���^�y�w+ַC;[���іg�/5Yrb{u�z�K�[�5^	z���OiLs�u��bZ��S�Eid酋��?�Óxz�Q�aRFgx���˳�!�Ԅ����J0/ @^��s_��
�֖A$e=���{M"���h� n�������jY�ѩ��Û����\��翡!���A�r���n�5���u�~�G���ڭ�y?��oP(��{i�* d��� �l� �>�<Nm��1w��
n�*+�ե�%��cT����+dS8�]�����Oba~M�禴��d�A���[A8C"��ɱ�Nd��*O!�܁�7�@S�6&ʈ��4����S"�z�ɼ���Tz~�Eʓ2W�Vo��m����E�R�x�]��yf���rj�My������Uȵzҹ"ף[��������mD]�8�+��p��^:V����k��]��Y�����]�jn���|�����Z�Z���
�J}�P��)�1h�D�g՗�9��yP���/��[�R�¡u�AK�\����~��+S��47��a�WLv&�@o�����8�Y�D��BRӝw�U���Obl|Z�$v>�.��>Y,�
�I��
SS���e�"�r�2���T�N+~r|T�aA�ϋUHƳ���=�쒋�w�crEq�h,�ʚ�

��mI�=n��)��=�_둯�F^�s�r1��1��z�/��MmNK���X^,ײ��f�zE1��]b����}��3LЅd����A�~뼷Q�$qY��Tk�� !B�0�A�r�==}Z+��8'֑�hyA�b�FEƵ�mP�0�"�i�"��<����J���5������1�Lk�AKs�6��D�E@���y,�d�*��y+r�i#�Z�V����a��dBK�ܰ��&�)i�i��l'������_m����ZV� .�_�z-#?V��h@C�"s��o�cAR�kd ���3�p�f���{�L�D�d����s9-���o��h�~����S�pm����w���|OD��~H,�P��3�&E��C���M�68��b�<E�A�d��!�+�{�-pxBE���z8<�6��c�JJE�D�.�-Pix�9��f��s)K ��+I�I��V ��j㯪�w��G��Ɓn�wSh���9�[.�bgJ�\���w�q��m ��,��8�	 EV�����h�5lij�q �Eh��em�1&����P&ۦi�E3��}ʞ貓�-C�̤d��̈��C���4�57��'o�+�s[Y+o�������Q������t�����ޜ��ǧ�1N��v^W_x��4Ii��.�����8���l�5�U�j�W�,v'��R���u9@p�ײ�B�)�J"���D�t�fe��P7-P�/������z�L�tV/���br�L�LZ��(F
 
�d"�����8�����Oj���c���$:d,���(�����-��w�s?��v6���uN��=-�hԸ�[D��4�0/J����-*���9�'�	L�kk����8�ۅ���e�.��~N�$��<���f�[B�V*j&�9�é��˜ni'I��S�(���c�D>�<�yQ��t	�|��/��G���>�Y�y�z�q,$ @��M�6��m۶afa�� �)}�=}�r�uH��ܿ�idi3�O�O��U9Ⴢ���1-�	���x��GC2�]��6%VK4ޡ��XA�'�d�R �<����)�Jښ��Kƾ�qR�ӓ��V�J�T"�WRK�_H;Iql;�;5#��ȹS���/�r��|؄Gj��a����"�����w�g�}���$��^?��/�\����ќ�Ɩ��x�%�"Vr�'T�.��̑W� 1Y��-Q��ńڄ(4�<;����Ų$CcR^cv���"i�<���AL�˹U�kY��\��Ɋ�EQ�\�Yn��b=� ����<���ч��)�Ԛ[�赒ʖMNL�4�Ld�r^vA4���jQ k�	��ENÂ;o@�·���[�iB�<?�=�9�3e���/��\zM��26�X��_{'T�q�����)���ȉ��ϋ"�f����ًc�3Y�\p���#)k6/����)Y�~�vp��L�A��M)+BJ���Q���.�᫯L:`N��3F����j�],,���\ݲ��e���u�f��wUҝa�)��ZJ�2[�+mg�ը[��V���k���,�Վ�����c9h{���m����-j�VRQ֎c-�%���/8ѧ�gխ��ҡ�)���k/�q&|�@���nO-ɩ���Z�n�^\���m8�c�v>�[K��^=tp�7m�ig��J�V�`�F����[�kÏc#�����O�* �S��$#��e��K��٭��J�����V;]��3z�d�ڽ�	����nA��},Ԅ8���1���&�~�U�̨�+�Ix�|���ͯMG`⹌A��!;�E2�P�wE�S���ZG�>���齇eqq�g��6�G��cw?&�z&�������kӘx�T�m�1y���d5���g��� ����j]Q��=���kLΉ�%@(��1�N(y���ϣa*�K(���u���M��Sf�H8���1��0{?��j���W�%/?��̤�:��6.X��ʚ.S�Ϭ��Z-.�2�X�b�y�ֺ!��i�G������+矂�5�Ӓ,:�Bw�k��D=���&YS�_3�ð�>w|m,�*�"**;y��2_����W��Yy�Mj���̙��~�����1)�?mV�5�0!Y'�bN�R�C#�bQ���N	��#r�քH0i5&��������&D|�J�Z*��1Ѝ�q�x�[ f.���f������+=�V9��D2cDTY3M���{L�HQ����٥�
�.VД�P֦v8����y�&���Caq.���턃�6O޺��7���7�3��F�zTdO�ֿ��/w#�&�;EQ sP9�xV ��a>eJd�I>.�>�Cf��KE��5\��Y.����
�wP��
ْ�M���įo��5�ك��3��)Y��帏5�_��P���w�Rn�b]ý�v�\eiqۘ�4,���,��$��l�s�Ɂ�r�.k��}���$e���j2��X�3��1W#3H���������I����4[4V>	TX���;���1!���0I�0rtT㜹BA{TsRi�5�������Ԇ(l����uutt��c��z/,maÆ.��y_S���Z�ꛝ_ӣ������xf��4���w��L�T*���>�mw(E�8J��L��bw7*�M�6i��2W��Q�dw����U����6Hp����vzȓ�ɉ�s-ۅ�!�C݋2v-�ļTl�1/����
2��~�*�{0r�M�z<
5"��G��˔=��jkk�BG[���w�ڭ A�j	���Z���U�h�����Τ��W$,kZݴfrȈ5���C@�
r�]�X��EoW�zk"2>��cS�J*�09#s��s�<U�
��F1!������>�4��)����<26L��v�\� ��������z� �K��H�2
N=�n��l֣�n�Կ2ٰ��2,sv,+m�Y������}<�����܆%]�*k���ɾ�����;�.%��o�E0 �bxߵv�j;D���֞�U#���Ɠ��ﳩ,BL�,�pg(�����=̬f��e<FS-kei'=E9����������\$�[I��_�DQ���3I��`�^v#=�ښ��k���9]"󥜲&2���e����R�y>��+��1s����e�m�V(��h�Gs�yP���94�����_�}�Z���]���O��[S�b��[;�}L��%�:m�)����K#��,��(שּׁݼ��R))��eb�Eۃgٜ���UJ�k{?Y�@� ֤s)0'�^5�Gh�b�_�T;��?�,7:�?�}߾p:���8�)Oى��X�e�J�d��<��[f1;9"d%�
��ߟ�F��x������~b[a5%�|f\U�\����6JɗV��ε��"��`�Ήl=v�4R/j�ȸ�(}�$E)��dY$�V<ˌ�ɢF�YT�xƲ�<�`�n/.�h4��cl�0���^Y��Vu��؈4��j&f����܄�&n���� �������Qk���v*<*t'�M�Ck<���7���X%�o_���3���TV��&6��cMX��R���|i�;��|V|�cE�+�������sȈ�@W����>D�mxx�.��?\�����Zb��u�L�a�V�軺��a]�X�q�ElO{3��,���?Ѓ��	�;�����P�M,pK�A.�Me
�,ܧ�H[�S�<���|�O��{��n�:U���M.*%oW� ںz-Ⱨv���y��hkmB��u
�&&��yE�-�.ڨ&8:y,���R�HA+���Lm�Y��Qo�Y�_=��R��y5	r&��rrLL��FS��(�F����z��jy��v�׹�-���HH�(}�����t<��W��ֿ�1�i����c�t����P1��N9��nu�}�ZˍAm,���Қ8�
K�y_X%SNe�Ϥ@�:��F(ъyn:���L1\�b7!qiwĪ���#������UCŎ���{��x����*���;�q�4�ܢ�I����n�2N:i+6�
 .,(,Argk� dQh>�^�xn�uHE���'�|���|����}�1�*i#"o0�A�~aF�
�[�b\�T��_�	�$�j�H՞���E�����ܹ�\����'�ff2у���[�Wz\n3�n;��A���t���L0n�^���XEy.���_?ÛXK��{�R��\&���8�s�5����x������ޅjM��Z�[����X,���ue[��$(���Z�
��J+>���k�=juRq�Z���#�t�ue�mP��k�C^ÉNŜ� !VxWG'H�$�� 
����%c+�X8�	Zt�{�m��y�A�,�a��\�+*\�'�\v(rQ������R&�
�`�����w.�Z��)T�+��{S��ј�&��4�G]�^�F��Ȅ7�A݃��Zڴm��^�-�O������X�>U���s�����7��\�\92�n���҄Q�ݭb	�/ �8��]t��abbϽ�9x��/�`���Ǵ�CR�3�����D��)Rҋ��S�S؍��N84����DGO/��ǰn`����7�Z^��ߣ�G����թu셼 �`D-�rm^7��Z��x��4?r��9f����������w����;4d�)H[>�+N��5|�:9b֚��V:������^J�=�#�Tז�t<��+�����+l��ֶ��m�l-�I��R\�V��T�G�7�P۠�Z&9��BGA_C����hoU����w�
����-�	��bNV��<�j�;<n}���V1T���Y�&�Z�@�N��*�rD,�*h�&��A�ZA�*�j0�|;:p�T�R��E�\L�a��bb��0%k��Q��z\dc�<�i&$�L��kU�/�p�W�%C���P����M��A1��-������.;�~܎���mEYeMY��#����ה��ϼ���>�Ɨşh����J�K���v=f�V��J��4��?�o�2�5ia�b:Ѷ�����3��xװ�Rv�珹�����S*�䝚ifSq�� K��PKc쌯�ꬥDe:�.eķ�v��&E,��딺W�Ū�&˘R76�iɉ7�|�.cȊr��R��D�4M���E�Ǣ���;�/�Q㯭b�ӍK����_�b������ܶ炛���Z�87��~���sؼ~@�3��U=��*�,xA=�L����[�g
��d�&��-����On��>�w?�o�C��f��d�Ett���c=�����9&�1=1�������ލk>����t�G񊗿��?���x�[��g>�U9��3�"�|h�@K��p�닊��m��/�y_/��vd�	��#h�mb&o���05�_�q�e���۱���x\�y;�؁�/�L��ޏ��8±0�,��M���Y)�S�l�KtΖ�P�������W�Td`�]�9,r���sS0�2@�j�Q����N̪Ը������C#0wTJթ>Y���R����\��{w2^�W�>��pe����Zy��Z�l�Y�� �m�W�31����i�;ƕ�����0Qi�j|�ڐ�ᗧ�0����J��7J�sչ"�YŖ=�H_F^e�!���>C��8: -F�	�Jv���ĥV~�I��B�p��8JC���z+���z��ů��W�#�į~z 睵���c����5����yM�+��Ȕ-�ϣg`#���h�E�G��,���S�m�+��W69Ta�n��q�T،G��U�/�3B�߫a
FR�>_S*�;��[�v��ձK/��s����ܻ����_��WOM�����Tŀd6g)ի����2%�7`\O.���mP썖��n�e'\�d��}��~��ھ'�������f'�ZV;���,nY vԥD����J��o�X�Z���0��1A�j/Ms����8.'+ǂ���86s�L:Z)�OY��&&kN]LdW�x-d�ͩD���%�X{WW�(����ڬ	Rl��L,�T�
�	�w�f�Y�	�97���sOw�LO֌$F�<��E����&[�	lN�ew�x��^�`X�`��YB�QI#M���9���9篷��;�ܞ������ÅQ�N������z�.�t��H���R�&''�{UG_�G�Hk�S�45�%˛z�kְì$B���~�=�T�׵���Z�=(�c��dM\G�i�M`����!�<�"t "��O��3YO��?�'�|�9��<��MG�8A/�����C��T�����`�#�?��_��~�]���)G	��'���t�7����}��@ǎ�@�P�����J�4q�8sM�^�QvTI�Ϝ!�G�����NЩ�Z�q/���<Ha#����h���hr6����d�����R"��_w�r�u4:V�;��:��J�eZ����Z��R� T~��.����K�P��k���:��CVZ���n�3���*jZ7-�g���0��SZ��|X��|�+Eߤ��]�;���ݦ�	�7^"Du*�a���23��i����M� (r�hW���"sc�"�t��U@��Gji�.��ID.J�]qā��-��=���`��S5h9_���5eu�P`(���Z":m���vF�HX,s�]��L���2����-�eb���n�������)�a:�YI������j#/��ϊI�>��������5Hi��<��Mf�@2�]�Z[��i�k��WBh�%w�_�b���gE�Ό��~����4?�(�o<�p������ᱹw���:i�AI�8tk5�`�������OsrA㺚��l�cx�j����67�j��Y���AV���bY����__�Um�[���l�!|���Ȝ	"=�BSB`A{�dZ,��fiĞg�6�zݓ�5OP�R����u���{U$@Z1��ƌ��Tu!�U�tL� oK�����ܺK�JER��d�]^$R���t�����Z�:t�?�.���� IS���J�R��{������8W�ڑ��� R�`�K�.�����2�|� �C���r^M��zɺ�1�ON�R�&�Ȅ���=��c�̎�[��7��+/�D��z���;�>�aZ��C#�*t�7���o�"N*�g0�|H�A��-ѹJgN���Q�%�W=Ai��ǩ#�>�\�H	Q���~��w����F7��T+/I{���(����r��-S���~���Qg7Q{w���u1�s���r�fGzh�1�j��Bv!�g�{H���k�@U5�D� ��-{�}�t���ʡֿ�ܻ?���S�k�����JZ�Ś����t6���
o�>���z��[~�]��q��{x*�m�\��di�Gj(�>^K1"TF �K�5�	�3-#9M��0�7^�T����@������u%lUs�MB֍���Y	5G��m�/6��}��S�R!|J:�����sbZ��,(>�\~���d']���Қ��fܞ�o��vl?�{��²>=J7n���0}��}��O��m���8u�YOs����œm"c���#�NuE]�d���F�;�V�\t���әT�[�^\��������꨿�ٮ|n�|�}���o��_~���R��?x���=r�Sc��\���E�@$� !�FvX��*W�M��ڐ��:�V�&�8Wt|��j�֠Rܪ,W;D+�v����|5̡�]�J���y?�Z7'���"��Q���U$6D����h��T.z�	��:G�J�e����H���a&ua��AAD���w�������R�E��
�a\�+"F;��!�S�^u�"8r��1v}t��(��N�sh�ɩ���OOS ��\-�m}uެ�&���C��O}��"�Ǒ������Y-_A�Cď��a1�Y���ߍ���7̅�(�a����!K���¼ҕg�w��z���3B�S��VZ;�tŒ�p�<��J�E)���g����˴n}���C|�~:q�(�+�@�_t9��/^L��g� y��I�$!#�DN�ؐ��&�)?|r������m�'�p�ex� �H���e����m�ɑST/.S*���>:|��ߤZ�p�N������{�tg��r�O�i���Z�#t��{�_�#����V��x������'Dg��ϱ�V�9l�-s}����Y�j�I�s��?�n�x_ӵ�Z����l!&�m�����{������Cl�k�7�2�"p�1�DU�v�&e�!1��&@Xq1�k#e.tʠm���~C]�W]4`��%_�T�K%�����U�Z���fxz�$H~��3�7�r���R�CW��Q�E�8�`���������'�������5}�?�$��Ko�w��m��C���o��;v�E��nx�[hdf���_�,�k�m�ǎY��{��������J?8G���Y�>���Xʀ�{�m�]�҉�k� �7����������a+�~��~�_���4����u=��c������,�+��d���0� �����p���"ZhGe�q�f��q:V3d^�_�U��Q�����H>�Ui3���T�Y�z�L)�%M��$s��k���wݺ��úw���j�ڠ뉓�����IS�g8�;,+��Z%j��B�PMK��� RM��*J�pĝh�G~7�����������]r�N�5���s���̜D��XZ�H�u�_-m29���0]w�����E������#��K�^,Wk�rG:��2�مpL��qLx�1�7��uk�mT�}�Ǵg��������J��[r��?[յУ�,���0��pÁR �h�ۆQ�Պ�ݢ66�`��c%��0mڰ�~���Q8����ez�ٽ���J��x�k���8��� �H���O�����/?�{t����������n�M[�
1��+vу��!m��@g��|F����|�V��ؠeSQr�yo�~����&6H�����&�{j�hM�[l�.����:� b�k��ٙ��=��ߋ��/�}��<Lł*e��|!������J��!c�Z�ի�q�,�-��g=[�J��#N�T�7��se���g�L+R�����z���8�@�	m��[��6�/�����yy��������m:t�"��u�;WGضV u#�s��� K��_E�bƸ��sF^@F5�K�&k;9�;u=�P�P@m�v�S�2�� ٫��#�(� �F�ag������M����z�$�x(����g���t�W3����<}�Ѻ�������޿�|��ش0X�##SbSE6`�E��Cm��#��l(ʏV�� ��MB]��#�"�6n�t����8p�[�]��阥�(��x$���ۿv�C����w���_y�MW��Жݣ�����|��{v?5���b��z��.��49�c�*1-K�^	[^�1��IBw=�����f
��֔!�47��ҚZ>;J]!�ڠ����,��h4kd�+���$��N��v�
�����<=J�5���PZ�Q����p(@R4��R�JҌh�d��ia6�T���s[��y�E��aJ6P�KOj��V�dj[��I݆�� ��/ _�5\����f�cV���:����N��0Em�������t��@K3	v��4�H@��ht_m�0D9�|9�f�wQ��%Ǳe� ue����O��ߤhB��A�7m"B�9j���U�R��T����j|!�N�E���7��#�i��<o����d8(�U���A�!�Q-�gY�,鍟�[���������lٴ�������9�ce���������_}uv����O>+�i8�*%Z��b��>CGG�f����������F���:ƪ���%+�������g�������׿qs߷8�Η8��a���A�b~��{��JFitn�2}�:t��g(��p��k$
�����`�v���MGN��Ov��s��9)�����ݝ�8
*�w|J��X.�a #���I�[�Q6�=̪��t�P@t�tdH��2[�]�I��:X�
�N���%><���o���:V�mvA�JYAO;Z��o7���ƭE5�d2"~pc �⺴@��H~~N�a���@�Μk��pv��i������������{�����$*�mD���v� �����D"�_�����1�HTڽں۩��g�[�D����Z�*poW)E�_>W�6蠇�{��f&������/�E<~�,=��n�����{������k�����6����8=?O/�?@_�����S�]��'/�!'�b�r��!U��
���/`���X*)U��g�=�ke/�O)p Oh�vUx��˶�$k�]�R�j�#B�%6%���*N}c���|������߽����ï�|�L_Oi���τ��Zhf�L���L��/{hxt�ƅ|����s^݋%0� u��W� �`�kX��d��Ȼ�JV�����%��"���z��ٵc����<V�SW�V[63�jE���h7���ǹR�&�%�����5���{���Zh�:��i������z�J�Eu{��Bт�}T���fې%�'x���� ��+Eq�XLP�*����%���ab���1����"��D�4���gBf�9b��(�AZ�8����uȍB/=Qd?�$]��������)�����l-р�"@?���@�('4��7I%��1�ch�KЉ��Ї>Ď'��C�����i��C[brn����3:���+��a�P�OI�i�\S��D�|�n�Dc��M����O�����}���/���مy�0{f���R"������m�E��~��e�]M��;�Ž/ЎW�G��������Ct�-o����6z쩽�^�ə�s�Π'�A��c������Щq����s0M�܂� �"��xܧH#_+�ݿ�&�
�!�F�^:x�ΞAܚ���yTK�Gׄ�`�|�{$�!K$����=�6)6*c ޸�P7{Lp��j��[�u+��e��ce���[���fHiBv
���������L�b�(�d����ym;|�f+�a�K<m�ߜ�PW ��g1Q �J�e��#�@��D����ڞRps���9.|��������^qh1�(�2�~�ȲU ^SW5i�s2Y�@��[k���8i�Rz4�j�����>FV#O���k�ګ��O��	�����>����#gh��}��;y���U{-)��㐦!2�B�1)�#> c�Q��M��Pwo�h���9 ЂX�=��+�{ȵDR�H3(�K�ֲ�M��[	���G��ٙ�K��{�M�O�N�Bn>��c��Rȶ��J��Rs�k������U���+�o]���*`͑��� ��:��	�']�Z]�f����.��Fk��Z�xo����m�­��-�zZ��mM�k�k�T�8IS��L�g@�]��G���� 5i�D�H��Uz����ԓ�� �BY4ܔ���������O��*@I3�ͦ�l�#��D(qd2�D	`��ف�f��i��{�$9%���	�D0�svn�&gi�ŗ���+!��:A��,����8�b#G仴()�%:yj�6o��-.2�(͠II���;:�Ƞ���bD�:21F�[�ny�M����pt~BƇ�[��je%኶��E�!�����.n�D��W�$jG�g\l�r�$R�p��s ����%m�����o߾]�4�<F��4�8�竴������5Kг��R-L�st��!���~����
�`���ջ���e���B���W�＝b�n�M�X�?>�%��Rq��o�L����A��=v�l4��gi��Aϐ`�(��X+(=v��8Jǎ��(G��pbKwQ�	���,��	Q�����.C��6���A����G�D����"1� # #��:�������u������] ֹA|�C����Y�ڣ�~Ʊ����f6�Q�������,]G0��G��h�
D�jrn�t�I�O;j�ylr�~*_��m�N�����_�H�*��v%Ŏ�
W�=t��@��|6�c�TZwITVd\T�t�F�����юQF�J:۔To���t��o�D]Iz��W�k�o$������O����W������˿�t�ko����#�������\��
�gՊI��V�;OX��DT��/ؠH;���Z���-D_��m�߁L,"LS��SR��݇� �l5H+lE���̶����Sw9 Ȧ�=�T�Q��X�8n��<'��OG\�� �j5�fJ���w,���$6[��{�P�\���4�c&��a23u5�~��t�+RA�ս����D�+7�o�������*�*_�X�YL�Q�)p���<X;�10=�p�oF�+ltMD�k&��O�����0�R�Z)2i���{�LOdI�V���A�w�H��jRQ�i֙q�	�Q�s��O]}�ƫU��q������𰤒�9�Ä�r�Q=&����ť�;���UW]%����1�񵯧CGG �$"��tA:a��@��1��z�M�B���F���������~�ﾝ���Sai��OU���rĸ��ln<�7T�ܲ�to8d%��~�JEE�(S��(_�A�:�
K����	;������>ڸ�~b7���,;F[��:�����Ԕ�$����E敟��k������cg�%Y<�9ʇ��h�3���E�q����񓔯X2Z�Fqz��):p�8s����w��PO��uX#AF �>�L6�ն���T�H1�@��^Z��)�%0���Yz�To,@�=�D'��I�.I7 ���	ْ�7�� ���ΙL�ٳ+�������-:){�����膬��w�	�W~��������|?{njҺ��� ��D4��W�5��fV/�>���L���������M�n����+7?��������A����VnI;�Ț��J�Fɥ^.K��>d�|Q�|]Z���]٫~9F_?M�HE��vv��-/Ӎ7�H���M���,-��|���G{��(����Iޗ���ki���hi�J71x^(4���'��Z���Jl۠'�H`�ĸm���P��-�&���A�Ŷi��]]�mK�FMׄ���фd� �#!ղ�z;��dTq��b�T��e�<�e�_ר5"�h2��Zkk�ڍ2�W&BY�hE�s��Cf�3\#[g?�oî��
7��x(2U]����[nZ�o�\����M}%��оM�9�))-�h���֋��Wi�&�_PV��4��S}���-���}0��D����6V*���r�E��o>ڦ��kZ�]�Ul�/[�����ҟ�{��B*�D�x�Z�؈��r��ύ5[�t�9H�&9J�bǠ�=lܰYf}�����:y�ES�m�F�ze�x]E�gF������-�.��?����h�c��}�>�nk�Լ)�@ Ƭ��3�t�>��O���IJ1���?M���$� ��m>fOG�c��(�|!�>�	��{�Ej�z��N�p�g�[�I9u|�>��O�����P�y�
#��C�K�#I���a�U���LMQ��ˀ+��.����^ą��Bmu\Ѿ�8!�_��l�v�:��b���uq$�,)=��q�H�����r��_F{��N
��Y��ə<���l��d3���C0���G���2�K<�?����5x���JbA腴�aO`7��U�������9S��M���W���o�i�k~��aƄ��j"�����8z�� �ke��8x?�]��ט ��Na� ����
۴�Ճݒ����`"�w?Ut�n�W�y�̔�����:��Ku�h7�>��ߤ�Nw795O��G	 � �JK"d��c�f0�p.��q���X�����vWf>T���="��2{���_~3�]/ܯ���~�0mذ��Q)�˳�Nɺ��Gts#d�ɤy�C�*Ց���ѿG-��}<�?'3a�W+EY��;�}y�(}�zVx�Z!�P���&�܏����0G�giYIQ��Y��!����# ���jɍ�k8~� ���-s��U3�-���ڳ��!ʒ�\X����?���h������^� �_Y?�n���7�c����7���ͥ�θ�j�h�5�D��sZwy󳛈�8Y؎I��*�����W\�ZĴA��f2��T�u�J(Q��O��͎K�s��!q�!q
�Ă��!�ʄ�ʳk"p��iLD�t��ӝ
�^�x𚅅����<�c��{�%��Dn�X�+���_u��p��,�����<~r�:*�49=G�B]�^1�	=u�� ��S�xLq�N���$[Zҋ�0?-�"���?��N�mj�y7t�sj�
ԧ�}0�S)���q~f�ju�=�p���=z\+3�L�D,N#ã�������������u����	Gh.��N"��[+�`�Hc�Yq��	�(��R\y�|���8@&G&���p�0��TB`}�|�0괭�_&��P~M�f��F,cD�T��.�������}��s���(P�(�LI���!�Q��ɒ���ATkE��*��	�?H��:'����E���f7Ip_� �0����Σ�xE���"�s�}e����Fr�+#�����y��^ﮰ+���)w�h9�Xlլd�y+�]K��?�Vgn����U�DGpA�m��Yk��$b;mKϐ��_��v��j`�Q�bx���������IM��=d��M/MV��o�x+�
9Î;��9uf�*�i�q=G��`3G�5����� w�����׾���Z��O>Gw��r�ͰM�},M/�͌�9��#Z��A��g��^K�^z)��k�����+K�9J�w
O ���>����*�j!ҁ՟`ۆ�2���&p �T�M�����Q	X҉�؉��^��"�P4?B������3��|�b2�O��SM���,�� [�/`��E��e1�����E��bDP<�0��V�s[�e�P괻/|������c
�N�%�|�ѫ$��O�3�Zʱ�'�y��$�<6^fY�j �bA�XMY��I|���,��K�S��!"��9�vf������s�0 Ą��`"v�b9zs���cT�E��^G��!�.�Kr��q�<�*�51��!O3�Q	��H;��+|�1��X��F�Ȧ�y��eA�p|���&�dGT��8�B��s�#}��'��lG�h�c�a�!��Xv����	�p���%Pt�Qn���v^���ۼ�����)�4/mf�iA�L���kF�^TJjZ&T8 �h�e#�ѐ^�L�c0����Bmis\��2���]��K����S[W=��#�/��i;m۶��H��!����!�M�5"i����q�, �ax������H6F�AX�1P������W�|@���@�}aa�K�N��ܮ ���ubSq)���r�9��ɱ�v�:ٵ�"O�?|�r�1��uJ���dLF�b�*��F�̑H���=�oS�ݒn���oA��GZ��Ag*�P��F�gy����8�Z�iV�׬w�N.o�|�?ͨ�d�����P:Y��W+U���[��8t�9b�����$�O�eYOHi��B�A�X��BQ5�ur�a�F����
R�oaiY@�SsTǎ�
6��1J��U�
�{nI�[3��hԁ�f�_[{����S�����ӧ��.��>�~���/�d�&Ɔi��f��{���/R�*Ty�Gy'Rl�R��CԸ����C�|Ow'�띷ѫ^��so�o��m*3��֕Z=�gq�$ӊV\�!�q!�S���H�$S�^EĲb��*U���uc�>3�,da\�ץK]D�tJ���b�0�AN�BYN�!u�hnJg2�N�'6(ō��|��٩t�ʵj��U$�<ӉS��0���z���!Jۆ���R=Ix��%��ns�"��j4�C�������c=��޷":�4��s��Dgh�H�.tֆW��F�\4��4�P)�MOO�5�\#(lj�Ƽc��
�,�%�;����	��D�$iiG�6lG�Qc�j�S��@z�D�u��������Ը�&����6����0!j�b̤3ғ	��U�a��4�KyIS���b�)�0w����;�nZ�q�� �����a �f\��6��E��LZKkzӕ!I��m�r���}�kD���RP�ý�C�s�JMXG���8�x@�	��x�2���$��w;�ꆩTD��ЋƱ�V����t�����.�?�����ٯ-?F��,G�)�f��i�htj�Q|V���I�38��aF�PZ������đ�'�J��e�=y�K%�zψ�O�B��;t�^�M�CQuX,���LN�Z�^����5dP��P#�k\�ҲV�0�8&ÁO�1�96��s�SG�ZG�X]�*N���=܃f��V��;�opR5ݥB+��Z²V��[���y����Wg1~��Q������ͮp����ɲ�(�Y��,�R���G��:]�_+����r|��
���<j�\g��HOúA�0̀{E&��S�w�Ly��R8t�����<rP��.�C �D:mxOb�+:'P�Q��?�U�)m���i=j<�M��N���|�X��`���L"-Ƿk�մ�#&���|!���	%���1��-�`���y/S�2�IDp�8��6d�"�ј؜<�5��4�����7\L{_���|�����b�5;J�\���2u�tK�k�R�@��<�"��s�i� ��M��n��_x�Yz�ч�7��D�}� C��nPJ�|m�l��a�����G�G?J�r�}BU�{Xe�1��7D��0�ѣ|�v�޽;�c����ӧ휑i7���� @^@p�q�R��_��9r�0����U��R���L���k�Qc�Wы�K	�YH�ScA��W�<�|�~���`�[�=��0��!�=6Rè���jj��8�������0��P����PO��p��1�����޲�F�:��2m�_���I!=�� �g͉�1 ��c�˘6����l�,\�T�  ��IDATET�Z�ː��'h``�6m�&����G��]�!��D�=��b���q\��0���y�B���P���(�͢�$��XC�Q�S���j�#OhKm����n\�� ��.�>/�<$������5�����g�t��jV6���R[���d����7i|�� @��6=�]$f�@u$8?��P_0�{��+���s����!�����5�,�����^A;;d��FK���$=��3TsCMey=g�w^�V��Bw���-��0'�Mx|�I6h�h�<��V#�l3�Cdb��g"eǏM�9�0���q���8ow�V�-���K���T�D�l`����*y�4��i�ګy�ڤ�HuJ��`���/ ��^Y@�V�5a�AER��u�<<�
pZR��չ&!���׀��W�j�ЁѲ2f���NT��>��T=6V���q��җ<O��{��J��H�DTP�O�wU���s��W����qr����n!����@-�'����r�ڡ� ;���a{q��d��*&8ԝ��[)�ض�K�&�� nq��d��k�����+�R&�����#S�����Q��c~n�~������Q��F����F�s��a�S�s"��v�Ư���O�]w� =��~*�h��:Z,W)˶k~~Q4�!��ݞ��ǎ��[n����KlGJ��*�l���mt0a&:�,�U�-�ˀ;U(�=����mX�z�Χg��.�������}+=�؋����.�p����������7�%�n��/�іmk��g���az�m�H��i�_����0�lI�; ^��;�TJ>��	����
%���8�H�����#K�ƈ�.	&g����@[l�<IӄBVȰ!���6���Y)$�7�Ϩ&Xi ��I��&�dg�Rm|,�퉃oH��B���U4�:GG����B*<OJt2�n����ˋl�i���I͈�?j3�8�)�D��mٴJ^zy]��Իf@괩dF"K8C�\C����&��7>�͔q���&B�H������.�����Iv0o{����v�Lr��A�����_@�T��v�-�қ�P��@�lp�!��Mؑ��k6Z00�;��8?6�xH�h�r�Yy���%-#�a����樈�	�1�J�37�R���� Q�x�f�f�z��o��9s��~�	�9uk��Y
,�cnqd���Ñl��g&yU�t��A�֯Ӻ 3b{�zفϊ����G���1��m^��9�K}�Qu(ÿ�������ŗ�lE��R\��#B4C ����T]��箎n��]%�Mc�Ċ����rm1�%�D,"��ohP2*5�_�[�l��uk�\��Y���XX�&Dq��;(ǯ�HW��q�nD@�쟆R�*�ʪAJ�`�_��7Z
!�Vh�K�SF����T�ԕ:���Pӑ�jmO2%��6���޼2��-)k���|��]�$�[R�ιj�/�Eq��h=����U�>[ ��������z��X�'7t��w�do�y�F�ne��_o�~i���S�=z(��g�ޢt�0��"S���X�jx��~X�%��os�ppձ580CK����j�ff�i`͠NQ
2�)d���;aN)(0�?I�t���Ob��s*�m�V�a��kʔ]
{Q��S�ҋ�����Dr���ˇ������)�8� � ��-�P�锱x��y�=�t�Q���o����h�Xl$��	Jģ�c`��k9?~��n\O�7pT�:3|�������_{+�>9F���率n��>��ߢ�[7����O_����Ӄ��O����G_���g���_��+#�'��űLT!C�\ D����f�}|pp�α�3�db��۶������)���C
�P��[��*�oؘY�F]�cX&`�����C�˗�r��=��e-�⣅�!��,O�}�w�J��:�1���*����	� e<�ֆ�	G��J���@G�d�0NdDx1vV�,�~q��x��Q+Z	��8��&1Z	ʌAV@�Cg���4,�>�'B;.�HR%G������$�Lq,�/<$jo��r�(g�cT��ԞD�0bY^��]���L�e����,�}ｼX�e�O�:MW��z��]��_�S�� e�h���݈��X�$`����f!���ŀL�[��щR��葩y�*e6Ԉ0�5�ꭕ�*#�+5q�x&D'�T p�	 5%��6�ƺJ�B�ؒQ��p��s/�Ls���/C�,%�ma"\���� 4   �T:+�Q��;qL��
����a�F��|1'`�b
�|,�DRR�6 �Au���'���y=G9J�Mm�����uok�d��Ϗ�C�0hC���&�Ej�t וʅ����`qa^k1��s�����mRR�A���c���O��DL^M��#��T�J��SL[�����i����`!�(mJq2aѧf�nc���2�zġ��q�_�Pfhh�:9>�I�u��9�A	���#�S2#��t�S�V�Z�U;6�q�j�?������g�kW�ן�i-ϳ�nyo������F&-%��u
'"���(7J�MaE3� ����������\�)�e��Ƈ����������s!S� '~}5\��Y�r�$�0/�l���o�m�Y%�}����+�E2��,0�e?�{�T��_X���q8�����ZH,dH��ϛH��������C�<� &�ȅ����H�U��u����<���P�����:_�H�ҙzi�a��_+�*�@K�f�;��ZQ��De-�O�QOo�(ϲ���sϋ#E�.,U��s]��؏�� B.��T��w�4�e;�:�r�70o�v@yqi�}�a���Ɯ:��_����[o�������k���dV;;����sZ.�٦8|��h�x��0*q(���x}��U���?p���%^��H"\��'efY�@CT-�jĪ�J�g�_�`�7�[e���؟�Bbn��x8�vHX����c=V�U���pm�f�.=#	Y�!����Cܰ��j�0/�\)ϸ ���H؊G.�[(�Ѫ�v@��PlОCOC�u�/6$�4�xц��Qs�J��"Gp�$uc
��<;��]��rI���|���ГO�o����Ӊ��2z�3�DW�qh ������.�z;�:��a�2��&��zU�8Bk�{E\�W]D�Ss��g^�K��Z�k7�;���t�5׋�R�]��fq����Ȓ�*>�Z�Ħ��5��FU�H�˰>A�֒�5)��Y
���9j�°!SյP\\��n��g9�:~g��==�y-����>P_;|���[�L��Y:}�8�{�e1�u�6�|:9�]����;ʠ*O�]~8����c�9��^z�.�����k��<$���.����>>���0�mxl�v��RZ��N��=u���������xcq���Y]i��(�jƁ#��z,)NU��m(�=�yv�T��Z�$��ľ�R\���q�΅z����#����iZ9&�rf��%�d�=��m����=�����s��8�F�������n��Y��8v������-�.��%���d°N��>�4��	��g9U�@��\Lu�ܬ���kZs�n ֕ C��6/5+��s �>���9�7G��,��AGW��D�
�S1�6��=����JGTE�ڠ���܀�\���E*{��YtK���H8C��d��3��]����H�(�'�Us�K�G"�N���AEA���ͩ�i*�V����$dV���ao���:a�
���?�a���U�d0���7r}�o1^�epa8�)�
����aݕ}�t<4�_ڻ�2|��]��8��x5}���JY����cl{�5�5��d�&��n%�.�8���%N����b���S2�����LJ�g"���7@���Cꞣ��K|���,_�d�0�-��IT��Sdw?�b�t�;����_�')���;w�{���ŗ�r �@���|�����Tv��]!�O��5NaY�=�If7+��n�:F����nݟ������^��¯������O������r�zw"�!�Gтo��";Rd��~pl�5����(�E!�K^M����@|�l�����N�:%�y8F�rȁ^s���فœ���W��b��u���p��eJ&24�0���B�lM�.��̬��غY��xD1/�I����G�h|�)��[������ȶwS����=D/�}����; �0moI��ޅG�Qowg�����*D1v0P�tu�!Äd�`~#1(Lk�Հ�%��m<��ؘQa�V$���W-qBX�HӴ�NAWw���QXB�V{6�N�@�O���S'Dyn��e��w�Mk7Е��H����B�v��Jʗz��'�ï}-�/ѳ{2Jβ���%�$h�n�u;�~:r�(�������ٟ������������e;:��{���ɰSG֢��W��[u����eץ�1*ߛ�<!��B}=��NA��VH?FݰN�|��T�ny���ӑ��W�ߏ�?x/��G?��l��޹�f�������N7���숣��ӧ'e�m���U�.���32�2�@4�	kB":��ex �`���  B��|��2-è�1JV�e1^`榑ꬔ�t��������ɗ��f���ރ�Y��H��~�15�7�jG2Y�v\)���w����Ei�^�{��?s�ZZdp����T����g5������x��z3~vem��,Q���7I��Z�f�0�M�>��A�7�0��(p�-�Nl|�#:4`�u�P"-����5k4;� u[��%$M#qŅR�E�x��֎ۍh����ы��L�s&��J�:�r���!s����������i���T^^��LB����{�V�e�g����b%; @���!G�r���G�v��s������-Oge�Gy�V�yQ�� �IpnM"u(�֪%�fQ)�!=ި�hvz����S_oT���Ķ��� ����k�����(&;ۀo~�2��Cw|�N�0��g��C~�G�ۨ����7O��H+�ۨ�r��j?	S��g����e�d�?|L�������7�-�bG]���cbU����? C��ŝ��I��(U�����..������{dS�egU��i���/����`��;���GR8h�A���ӻe�J'�00䁝�%F�!*Uyq���)���C���`2�"d��r2.�C]|��������ԓ2�$6d��5�=S��1;/�aHC#]��+ݖ��$�l���s�����^�/�ڛ��&�<�� ��B��S�Q��сI����LJs>$�G����v�ʈV��Ϝ�6v��'�m�Vzamf�޷�:{i��ћ�|?5ɿ�-罚�E�~��stzd�Q�J��R������I!��]��{�y9�L�&:xl��0�j!is�g e�&��͓�"@k &I&6���RKm謅j�te��(G�eBi�P�I�rD���0��E�2}��>H�_���w�#����P�K��w�Q2� B[շ��G�����^˭N�Z`P�����GX��2�>��W��y��:{ya��XP}�!��(T�"�� Rb��rM��c�6�V�͚F)�%�hq��{��������~��s��`�2�s�~�gO�qm���j̎JIKǦ֔�M~[�|�,�O����V��'T�����J3� �l�4D#cS�z6�pP.�*�Rk�}���v�;��e��9.�jq莖��;�q]1_R�ZԄ|��j�� !��.�*�
�жZ�I�d���@������)�ml3*ұRV��]W��F����k���Ll��±�4CZ95}�*Ȇ���	�95y1�J*���g�gxb��ȍ x���Ҽj&5�S$���_�U�9&��fe{W�,� R�_��_�x:#��<|�-L���萁3G0+$�����ό�i������ҹ����o���_������׿�/~��w�}�2��o��.��r��_�����+��6>��/������x�y oxQ���'�=�MF{%o�o�H��T�͡���ա�����_��e^��$����7"�Re6og^T6zѸ�s�����c'O������Q�ZXZ�h��z�{�����:ڴ�6o�]�������B�o8&)�6F|�_��=65#�N���\�ʱ	1�R�xx6�O���%���<�Nq����5k%�A���!5����m�^شh�HO����i�B'���za�><2"��'}�!(�قpM��U�Z�� �Gz�Ǽ>�N�M��%ՎI`x�0j���a�ф&2�ⲴqtSw�F��EްQ�ɳ/�s��c�4"�����:t선�;>�q�����u;��_��Dl�3�6<��َ��A�4>Y`@����Nã�5�Y����١�bp�(6�MA��tp:�f��� �O�uk�-�F'��}A�����d���J�ZʙE��7]{ݸkU*�N��[h����=wQƫS;ߠ��a^Gj���z!G(7q���b�}k/]|�N��w�g�E���O��_�����tŵ�d`�O��%3�`<��:�.aG�L���������;QS�sG�W��E���B��\zE-u�.d�Ԏ}������ZkV����-��O{��܋��>,�	¡+9fd$ %:ђ��t��Q7��]��\y1�p�մ��h�q�Rz��,Ȁ(YH�qV+R���Q��4�OW;����&ƩR��~I���6#��SO�1`���=�ֵZ����F�* )���i�'��P#��`��`�i�j�4�x����I�V���@>�*�3"V���̇��%��
pd�R���{"{A�N�U��1�>솒�n��R,����y�����q�G���6*a�;��r_,�D�-,�ʔik���J� ���;X/*��8pw����ꠋw�/1�0���K%l����O��������ߢ+��B��Ga[���1yoY��f;�G��z��w��Էv#ۻq�^�����&a޳�U.�~"JS�G�ҟ+�0۰l(�{Z��Hf�D�&$�E4F��@5�V��5� I��rI��kR�̞��F\J��x߬E����(��5��n�F��J4��0����ECI��ˮ��.�U��3����W�G7��,=��E��4�'��X*C�JQ�K��G�1��`;⽖�K�P�G�d,l���ֈ��r��Q�9 Kuf��;� ���sd{�����N��|&����Ex��7.R�!"t����Ąu�S�!���s�q�,���*��Ԏ��9�&zX+;�(2�qM��i46w�*�� �Ju��'��Y�Nav(m43w���#ߺ|V2�-%n��8��h��I�dXر���Wu�Ԡ�������~J$3� ����i�"Dd(��J~���؉G��BҎ�eafMc��"	)��lN�Og#Q���1�ܾ���9�&]��/��e�T��� ���)�t�i���^��%}Ks3t)Gw|��W�����y-G���!��8����߃B� ����NIB��t����	�C�Z5\���3�ټ�1]
�&�ۯw{~���V������LH\�2��?�ں�&m45�u���Q/[-K �2�M���^}��6��հ����y��nZK���f�Jt�5�O��^�\�������4�K��%��H8lQ�ke��6 ���[[���Ԝ�-�b�0�!����R�|�%�/S���Gٱ�bHW]!X��3���d�-Z����)a8TQ崵�(�>W+g��s�K!A���H�F��9��C
[�S6�Wm�l�ع�B���495͑(lCT��2g��F��'c]!�B����A��6���X��\ԝѢ�=K5K�u�8t��	��@X�M����	����[�ԺKmI��n��]��m��7�DC�T��dк����S��LC��=�m�#�����[��vi�NW�5t�k�.	v�z;�؉Q����8@k��?����03M#S�!Pe�8U�
ۺ�e[T���r�P�U*���������4(��x�Xc�N�ŬV@K	�X��RX���p�F���U�JiO<����%��P���6m?O�L�=����0�D�^:x�Fx1A��k`=�.�I�ꨑ{W)��p�h�a`j�B��h]�9�V�Le���j����υ�%ڨȋibD	���S2�R��A@�@��jie�~7o�A��H7\u1��u����C�^���n�?����vHo3���Tz����d�Vr�|j|M������U.���a�`�;�z嵒�t���Y�FH�I����\�zSg���:��6r�kT,y����4���!Z`Gecc����$�/�<%>�:f-�s��J�"1Q�6560��*���s;��"S�q�=�^9�~8j�w c���鋖�ֿd`�Ne���Py�כtn];uҩ^�E̳1�["I�nݾ����z�)F�|�.��E�p�q\�tj|�7�2�O����Y��Y���U&`#2�v��'^�h�����E��h�wHZ_(fG�ZD��	^���n�F%O��G�}x]�Nz��c��t'�g:�ԡ���k/�`�(�)] �
���%�=�N�e����	����g3�a��\ �o�����g۪ �,J]�����z��q��|p�5�8�E�����L�����&���0�a,(m�hu�|X��)��eLD��}i\3��S�jR겖,�؛Y������D!V�rM�r�겁V�
�`�� �"-���=Gi���r���ȴc:_�Sp��.G*P�~��/|��tA��ӃZ�Lis�&y�!V���w��i������]��Uz�[o�Sg��o}�9I�S3��`ъ����! s-��K_8�4ʪ��.�${o�8;�9�|���0t���Kjܲ]��ʰ����M2�YP�Z��3�cP��!�if9��w����v
���r$.ba��>(�w`M��ܻ˞��$3�jZ���BH!1�k.�	V
r�L���ꥎ�5c{X,��[OU�A��%��f�y1Ȏ$�0=?_��Gn$)�c�QS�x!�J�x����t҈�nv11r{�6S�v���Kt�o�֮�ǟxX�<�����u���fN���a�����=��b����F�L�'������ZH����Wg�d��e(��5q���o�U�i>8M�G�&A-R���/-,�`�Ԡ�ك_��Te����/e h�o۱�x�ӳ{� �o#u6$q�:3�[�-�IB�U!l%Fb���D�h����(�9�Rs��+lBa����� ���%��B�7�5+Hh6�N��#�Y���9��c�vu����5g��g@$=�":��Z����Df���#%���Hq�29ɕ⥪4$ K��.6TW ��LG�b��;�Z��~��mF�k���L{w�0����������BZ���N=�|XZ�� �+V)�ktml�6\]T[�J�N{?/�J��ü6{��{��7l�W_������������ ������A�%��,�r���X'�}���кA�u�NZ\(�5�m�Ç��G~�]p�N��ϋ!�g��s��� э)��mN�/�(Ε+�"��Z��ǹ�.k�wZ�ns�z}k\S��l�v$�M VҝKJ��;-/,�Z�}h�#�Ji�Ώ��o�E�w�$�?xH�8B"�b�Zp���Ǭ@^�V#���u<<��	>��|)m�����
�1�=Φ�_��W�Q��!����>��k^Y�Q<�Gj���@*�Q6�Jp�ٳ������O�ys��V�YXd�>)bW���-�u%.&ѵ��ݪ�?�5 ANMJf1��G�l_ ����f����ʟ������-[���G�A*1(���i����D����]ߠ�G�'�b�[��	Kv6���L����L�\� 6S/O�8A�DZ��Қ�Q:f_D�)���Z���(��vqr�#���iK�s��)��,wt�ۖ#6��?WT�p8T�Fc.�0���G�>AI%BqS�F�a���J|q;��P��ٿ�;����?�;��S�r����;hbb�.��
v]t��Iz���h~xq4DL&�>M�DZ��=ө��\=��E�r������6�.���߆���yGw��!2��O�fyC����$hM����w~QZ���7Ɓ�'铟�]r٥t������u�Rq���9��1+�)�zX��������@*cX�~��f���������/jЌ>�~��b�;U�z�uÏ�dX���@�B~��n����N�@�����G)͑$�"�w4�I��R�r����cokF�����}���9ⱡ�#�ĈG��-B*��IWj�h�Ni�/@�R��0���)z����uW_N;_sJza�M."B�i�\�{��� 9�(85��n�F��h|bZ�sˋ0q�8J�Jգ�}�����+1/I��V��?h>���H3:!^����i*10����(�S8��ݓ��� -��c������Zyp��zj"%q�Fj��x�OS�7A��p����<
�ŵ8}�~+[���+����u��_D�2� C&�LK4��l���g�%��9���N�������׀�b8#� 	�u���c�}Q�r����������n���[��/l�R��+���z ��F������Jֺ�w?X�X�A����/��(��{Tuc��S����9�����em��W_B����t��5�z?��T@R` d��FJ �m����DR�rq��QF$�])�֔�]2� ז�E�a(.��M�"[��)��_������:��>j�$ �T)+���T-��b��zץ5E�%��H�%�oM����1��:t�C��T<FI�h/��x�֪���<?'}��S�d1��"����s�rA�a�E�h�*R�7]����L`0�e�RfgX-D7L�X�'����1z~�Kt�e��Si��w�#�=M��O��܂��d3���Q$���t�-�d�5���aTo`���QM�l�v�+�����Y��S�aA�q�,i �Ņe���aCU/�"m�A ����D�l�7�A ��"zuM.r��d��h���p�T��&�I��V�m��6/;�pL3�s�%��� !���CY-���U����J:�	U���*[��!�������1l�+�� ��ܢD���x-827^;q�Q!�s_Z�l1�8^�@h��Aa�
�_PG����B�p��^De^]���j�/`A�@��+`Hj�ܞZ�������mt��zy���<C3��;��H�457+�Ď?)�!�w�7O=��;t���{6m��N�-�ڍ�i���Jœ^�j]�b���u�J=�$�&�)�NO�C����i�e6N N�-���?�U�������c��aY�O��Z��L*%�#�Ǖr��&@[������W���<u��q�5׵�k��I*����=o�gVp�s-�5�^��񴲙y]���T�r4��V� 8�K�g���S���6X���zC6c��E�,����Ĵ쯬ŢD�9�D�~B�jNrT�kE�S��2��7�$0����u����0�$���1�d���dXsm�?��#�*�*���*#	�S�Ewc����$�� ���3�:D���_�e��D�I��Vq�e�rC��Ҫ�*ΐ�A/J^:A*��Ș�%��N��2�p����z�}��g�$�ݜ�W���^�+����3t�5������i��S�M���-�]>19gD�J~\)E#`\X���А�xX�P:�_潆�Q��Ed�0��_;��VͥS�STlXtޫ^E��2�1ض<�¢'�l�ϕC�CI*�	�㔄��v(3�-�Ar�j��|UE!���KӚ�n�$ک�����6�43�S/H��b�ff�Hd��Q;j�I6z%����t��ܦ�������k=~�r�)9y؁�F͔�������77�4�RN1��h�:��u�e�R�!rK
U���-�|I��+5��<;��[�Jz^�CCz�����Q���!�?1�dj������s}#���bz���Y2��	+�g@�@�b(�*��BO���i�F��إ�0t��6��H�"��#��C*2�Tw 28H}�N��j�n�d"ԝ`ď�s ��(���f}]M��uF��;��ya��P`�I�()����LGMO-���@E�Jf��&I�"�����r�(��<�z���#�Xri�Kh��!��%v���|@�C�,��Gj<.Z��0B�&�!~�|�on��\X���7_�i�>C��;�-��'�m|]�Y�24�g%�|�!;�G�k��}tM���J�䒯������OL�t�7�oh6�hi#�rM+�dA̦RY���ԥ;�Cw��k�e��4�`�Q��F#'O�^��h�L;�޵B�*V��U�1���\��gi����x�{kn��j�L���O�3�J����W�ݿ� /&�����`]_}h�[�����oE E}?�m��*�����֢"�N������]��[b �����T�K�3�v����a.ZK��h��4ۑ���j���&e�/���6�s0�r�sK�.HI�l����f�=4vb�m�ƆOQ���_w#��կ�)�k��>�s��`�P��& ��
PY�:W���5�tp�˺��$6���A&Zd~v����z����"2�q���˼A���ϕC��۩�m�IG�DuVH�Lj�5l�r�����g��Fn##(�R���1Zfg�q�v*�x���na�{%�}7m!��#*��k*�fi�	q�*%�jMa�8G���2��.�<��������J���OPqy�#xF�N�����q4���c�)�HK�g�����߸�2q�&��pԿm�>�<�[�T�ela�Ru�s�6�����J`����uwd2��#vK��#fF6����) h5<~SU|����qڴy���ɱ#;�������4������&�	��T�
��J��Y�2�[�p��=�#��'�/�������WG#�6Q~/�^I^@�	���4�[P�����l�mb�ZUB�Jo�x��u��4���1���d;^_n�&C&��3iQ�C�e�}�@V��n����.if�����(��oW&%�d���y����<���(6��ّwf�yM��}�������b���_�^��� J�o�����H�R��V�J�煉i�W:�����{�YrVע�NNݧ�t���(�F�eIc�s��ml8�m|��{1���� e$�,Q�&����t���^�:�3|������:�TU����kY�S@s"��77����x=�n �p�uL���"H�,,jV��'��ʘ��}=?��R�GD�Z`��_Ν��� 4*nP�4����n�h���3���
hfz��|'��/�����;š�*G{���V���'���`_��ҵ8��l;�����<�y2966�2�i�	a�=��5 ��u����v�"��Ҥ�,'�Lޠک���_7a���5l�kG�M*U]1���N?r��;��k�#wJS�� 5,�x��ٶUn���q��-[d|r�{PS;�����!Y�z���/�`������ZD�l��Y��[�0��PD6n\O��NVB#(���C�O���إ~']���E����
�U�˼���r��HL�m�LfL�`��4�]���k.w:�d�����q��������]}�JZZ�2>1�LT:�e��: D8P�Cf`I�/�S����g2�e��7�w��߉;$k��;������a�Gr
wF�1:�Z!.Ҵ���\6-ͺ ��_%����������:\& ��Ă�����O�!?��̼tw��d_�"N�΀���fj �@X�B�ؠ�WG#��� ��y��D��F�����ZQ�������⃬:Fd0����Ju�+�d\P�W<���!�|2���)�F�p�fJ�Q�
�#�1(����c���`�V4!�<�(��G�d�Kp�!3�c�Wc ���"%:LRYJ%Y��#�ǏI,�A����;��&q9tp�X�֚"is����,4�q�.4�,��f[ejA��ꂤ�!&T3�6dP�@i�݁���M'��X<(�6����Y YGqQ��fI67ĸ2Z�5
�̦qMB���0��:����1\���6I�?P`zb=�K��L*.�ݛ�:<��Ľ���Yr�����b�[�8��nl����{�|�ׇ�P'��7*;5 KY᮲�8h6z^�֭��b2�MI}��?#����ePt<\�(RzE�FU��qk��YV�;}�'/w��5��x1�P�9�;��;/U̽�kｖe�v�dO����(��벨�m=���E�5��&��җB�� ���:ԡ /:���%WY�k��)d?�)st6�}\PۄJ!dN�j4zm�H,t�Q�s�0N�ʙˑI{��`a>����^I��]r���B�L�T[5#/�gعs�\w�u�۟���ڵ�-��~X��_�K���V)�4;7M���n�B�԰ �"I���t}-Ȋ�~�K��MF:(�|F
�EJOװǂ�	�Z�$g\��`˭�6F>l0�2d�Xl��&�I�J�DĤ:,
(L6,DM(�uw�dAo, �Sh�j�b>ˌ$*�`b��������Kj���^��ŷ�ˤ��ʇ&01Q�e�P�Հ=s0���9�jdp��T)�PDy�(�\�y�[�(?��o��};)Q���5@0k �����ŏOLU9w���IU_czn^3�E!�r�Wǔ��&q��Y����B��u����ӄ����JQ�L�F9�G@���-��!����nP�GB6�N*7?Cֻ�:ʱ�òn�F��0������9?1.��v�A���l�����̗��#�u�H,��/��BFT�����\��TzV�F�j+��&(ъ�	�-����N�1
���,u�A}��[*��R�rN�����]o������I��Ռ�&�+&t���6sa��/�v]�j��ě5��dz6/����9y��������hs23�uTI����ٙ���Y�k�����OOʵ���<xX�>.�3j������"�c<�����,5��0�� ��W��L��:q�G<��YƆk}	���>�l{���2t�U|�2�����O�u=I�]�@D�ԡd1�D4�u������l���%��˳�R��:�x��; ����bhMq�O��/�1����G�\������!Y֞8�x%��K=�t���>w�k��3�%دz�Edk�D*a���M�62`d��K�	̒ͤ�.Wmb[��� RG뽟�}��Vg=?!v�ƔB>'�D��I�҄=��L�(���)ٻ��A0FgN6;gir� 9���fҵ?��f�5�����it)#�Cu`\O.Y8��Pz?���,�x~�Ԕ�{����������亏�&�/������ȁ#C�}���^��t�uHV�$��صϰ�f�@����ԙ���@t�1��i�g=�"V��L`�����Nج�(y3��W�ɂM��#i
��u�:�#\&����gx!K���U�İ�����kp�M��}OR�d:~W��%�8�r��b�ɖ~Џcan����Jy�5�\zFz:����mr��^i���3bi���)i�7Ig{��w���	��9!�n�@Vjf�G��c'ث	�B$E��NQ
731vB�oE�l� _��?��G��=��#���2�k�E$]ҍ67I���d��\�H�S�ߑ�1��Ms� �Z���u�-�}�w�}262�l�E�J\&����薣G����J�R#�]�P2Ց�%�oA�����HD��\�~�<��3�_Y~&(�V���ޓ�imo���V������L����t����Op� sF�Qsg�-�)�z�7���A8���۽�9��h���S?������g?�	Y��M*r�X@�n�z9#�ɪ��!&�����u�2�ay��������>}�%c� Չ�&���$��uC`���������z��s��'?u�l�`�����W�r�<���׀kq�B#���쯫A�(RQs�����1`Kg	.���u[U#R���^(�_���\�Ñ����R��k�{#m'=h�{��N�Z�>,# @�R��$g�ɶ�`VX5��ǐ���q�9�U�r*�4�/���X� 6��Hy�����y��n|>��m����A2]�s��	ͺ��QzF5eZڷ����%�'?�T��P�k������ǃ{�c�3_�.^��:.��1�
F��V�X���#�G���H��Ax'-B��@5�8 1`�k3��'��Oˮg��G4���bN��� A��������(���>0,�?��TC�(�D�#�1hFO�(�{�H&�6�J�1F5�������Ǐ�V��{��[8��E쓟?�8+�ss3l&�5�9����&4[�ģ�n�zr�@�ྃ�L����Sr�<-��~��`T�9+jT}�q���;^��q�F���x���S?[~�U��d������1jDI�%e��E����G���/n2�-,ZSN��T���`�N�XT%HL�0�(���5%[\��<��}q���c4֡0K#�� dq��n�3�
A�Ğ����#G�]���ޕ�۞�g}�eޕ])���Lg��4K����1��_��#��8�e�s,�l���IM�~S� �cllDJ�E��ҋ�����d��0J�1K.�`+7@{G'�>��=�Չ����ʞ>��:�!���\���	��G~�,JǏ�]�o�"��g�������^����l޼Q���Ԉ�9oݸB�������dl�ע����]�A�H_�n������3n�%g���m�J@d�:�={�J[P�?��޻G��<�ѯͫ����K:�R��gv3s-���,s,�e�圭[eb�?rH����˯���|���+�H��s�&�n�Hz�����d'��ϕ�|@�uNOHA���]I���Uo������<��ۨLH&4k�赘N:��p�$�^@�`���.ft ߐ�{�#J�U3ϋ.��r ��Ygm��?��b���t�-��C�������i�M˧�NГF��?ؽ��B0�q���Dc�,��:r���K��S2���TP�)q�\$Eu���V��a�����`��� �-��
"�t�SI��= 
{瘯�Q��Υ����tr�x�˩���%0���������m�~�F�$��3]q�:\�*6����A�/��n@�`�[~�@�4ʕ��� ��E���☤�c�_V=�ߵ�^lфanvT}�nI5e����}T?CP�����>&e��=�ӿF�_x�� �T;�Sg�A��חD9�C���m��j�,��+d��;�F �6~�Tv0�%G���#�����0
X7�/@C�-}�3�<c�;��kP���Az�_������ީA2z��~bMf�r��g�C�����#}_�2�3�mC8Km����������h���Da��v�f����p舒�uBM��X���e.
e��M����}[8�X"DG����|�ɚ��� ��>_D�(��L��#.Ч.e�H1�,S�����	�����b0�sB��p���j���a)�j���`��5�$wL�iu��iu��j����n��2�<�Tͺ�"�A6��'>�j`2��%sS�R��H�f���Ⱥ�X^�uY���%�u��=���D�5\(I�~~���T�KD}��>��w���eY��������.J�[�n��g�
N1����<�󷝥�n�<��'���!��r�9k�7oA#~;#o���T�ʅ[W�ֳ�Ռ����_�h3�Z!����]��;��>y��.�/�;n��x@r��ɽMw4�+)X������7������������D�A��nΑ��4'c�/�5�>,م)	Չ���9&�zY�K@�y�#�BF��Ӊ����߳SZ�ZeQOg�]*�g�&ؿ��l���Y���;K¥BV��p���moe����OHT�:z}�)%M�����s�~�X80����>a-r�O�H�:L-Iu�xmSi�7F��t{ɩ�ʷ�.e���;|���y�S_��Zܦ%z゙c=G �"���j <77k�5U�F�K�Jc��49	�:�Z��`�R�v%��`�~�WV75/X1��CE{�M��Q��e��J w��\���q��6 �WՖ������	�L�/���y�{�����
W���'�b�b�k�8�`ِ�}	#
ɛ�r�lXӫײ&�-r���v3�^H��8+/�< M��y�v��џKLg�Z��"r��F�cq��,N��-gKnꨴ%Ze~b^"VDº��{zehhH�:B�T��ş�"^h��s�9�yU'o
_M�V4�.28;�Y?��<��泶s�AL�䪖��n�7���;��&pg��p��L�� S��#���h GI��2ꊄD�L�H�V�Y����8�)����{8���xذP"酏G�Z2<�a5��fp�g��TdA�DD�M:Cu��K��v �=dh��T�jY��EAq�6Z����(��1��O<��ņ�F{G*!��G���W�7$ͨ�(y���
FH{
��m&'�H �S� =��e>����26~���͛��k/�D#�q��u˃ܯ�|��>F��bn�%M�����Z:��%&�Z��w˦�j���	6u(t�fv�YcQ3���>�D�����{�N�~�4�\��"����u�dllH�o��r:"�m�n��ܤn�fܛ�N ���k����jt�l��������,*	ُO�Ⱦ����қ�˪UmX�J�{���3R�]\Zy�%G��sQ~\Hg�	�5u��{�V���H�9>||L05V��M���)H�@�,,f�8zO���kB��c2B�2�{���U��R�s��Uҿr��M�I1�N@��IP�`��ߋ@=uL$<�ȓ��cO�TeaQ�rԓ`�Jґם�Q̲L� ��]_��X�r��u@��dYWJ�+�"��g13������8ܥ��4Y۫']9�?���<2md��(�_���4�d��ՠ�*���,��W�����Z�&�Z�*\�����4�Q��tKHq8� ��!Nq5��KԹ�,#t$�k�"�<~�M��QQ{�����^���I����Y�W�3��kL;ؖ�P��q���4=n���՞mܼV^�K��..Ȏg����R�������[��m��������7��R�����S��7R��o`�G����G��5"{w�=L$5�kք('y�e�;�f\��!���@������D��o��1e�S�cx`��~?�o/�����$�>!S(J�؉�;��2lFm�Aa|�9t��7�.3')�y�|�~�s�A"��
�s��k�ӑT㦎+�@v��>�5f��p���%>?�[�B[��M�� �]>�e;O�]��*����֩78�yU+P���7�3�ˬbL&�9q�`#lTT��Yں��fa����PB���;��@oS���eN83Z;z��{肋��� ���j����( 0W���\N3s�et|V�֌�J@a,�D9�s J�$�5�c�Б����̒+*�4��q���~���4� ��:Hff�Xb���	#��ᇂ\�Pz���s�;�=7l���s,
��a���f�r�hs4'Srx�f���D?yn~���J� S����A��%]��5�m����Gc!u�>�br��e���eV�š�{�X+��ԴDۺ��eFf��� ��2ْs1���$o���ܪ��[4������x\^{�2�[U�O�K �&Ǝ��kO���H��H-������<��~���i����}��48�%�y�/��w�J��|�}D$䖛o��e�����iY�i�9.=�aT*�1��4"� ��u�qm2��r�7狤�� 8@F�U����C�'^D(IbmP�,]������!4J��;�����`#
}Cf�K�ݩ�oYM���7��D��@k�:�(��V����@S����'���E"]�TsR�u�ԫ[�ʡ#!�h�p�/�ЎAٛ�L�l�}�:f�5x���IdS-,�|iΌ�6�ԉt赫���g*{dK���ǩ�׻�r�xﻜ����9��'[���]b�Ɏ�83�4� ���ڀ�󇐉Ǥ�3D����&S!i���ѽRq��=w�/+V�Ƴ.�����ԁ>/�O��>L���u�l�hA@�O��W��5�Ɨ������a�G���,�M�(����a}�IC� <�Ƚ`��1�6��&��s���I�;3w\M8Ȅo��M2���a��\A�C�%��U�3͡�+d6re4����ǹ�Ѐbf�_(�4�w^��cq8Keq��Kt�03�3,+���p͸A#��+yp	D�sb$z��Yٹ��?<�Ө�A�#1�U[g��?�s#Q��C��%w(@��;�L��V�juIE��_&���iT)�y�����{�������u�압k���w�.�lX'l|���:��h
�ohLj����o��6�cO=��FD���hi�Y�n8�x�Y�(����ww�S���������QJ8� Q%9X��F�)��$��9�)R������f�R�;�4��3F����zP��ԍ*T�u�I�����5�*i r��!F����Q����yݔ1�q�'��5��B��{�����������f�$Ë�t�5G�ߧrҙj�P�/O=�[��Z�z��iKyࡧ䬭��K��n�^�?��%��y9o��O��?{X�����/Ȣ:�|�O��秞ީר_|�>ɩ�� ��������i{{���5����޻��E#d�K�Zdl|X�5�
�5C���ӳB2� ���4�Wj�ۦ��(n���=F�������a8
��e*TH�#��,��Ş"�l`i&�����Ҧ��3�/5���5ʝ/�������4��%���E���x₮��fb-��o���q�b������7s���L��E_�jےחojn^F��{[f��vs,j����ͥe�eo��;�s����_/�v��ܼ��:�7F�8�.~���a�l����~��ܘ7S%�����@�D&��jv^:R�,�́a�� ��������?ˆ-Rs�a����õ�\�g
9Y�5&�A}������׾&��?Km�����tu���������E�~���#@�@��s�`_P�ٵ�t�AC(�����Q	x�����'[S2:1m�Ӻ��CrL,���:2�eˀ�jzӪ�N����=a�c�Yn8 M����r�y�Rʲ)�2�s`P�1_\�JS4�FN4�k~Q��]
Y���u3�~GW�t��ˌf�O<��L�O��F2�M���,�Z?fب��Y������ڎ�9�lӡ�a�7��o��|���ݙh��ՠ<%��������'d���J>�({��`������_�8{���4N�֯��y�xTv��ED�HT{��~�H\�۠��,M��=�eﾣ���[���<-;v����d3%����y!���B�<;���0ea���:�9�f�ɀ��{Ftg�F�S���.r.u׾C �aor[[����ǨP7tl�:�}^���)��У?�7��J�����|&/#3�f�:u���|f5+���2���3/쑞�ղB��GNH��*I��V�H��W��%0�+1[��P,��/�ebdBڒ-���,uGA||H�A�<�� n��y���Hzv\F����t���Wv��I��c�˕�x����WI�}@�xz�<�ϟ��||LVm��#�z�Kz���ե��/=�mT~:.����Ӭ����+�����z}F�hG�q�Ϋ�7�)�H��6��:p 4��F<5p���6��fJ3��7Ǿ�'��A��,F{�x~�@pP����mw���6����ӑҐ�N3F,��6���ў� ~��g*�����tŒ-�f �?X���f����y����h���q��?�x�W�YwI�|NPb�D���={������Y3�Q�җ����0e�q��͡w�U���Guv��>����V��S`o/���֋_�1�K���O��x88�8q˛Pp�ު����|v�"G�����q-�U��>�.�e㺍j�j�ؓOip^���6�֍�Hd�D��5`�-P0�e'���~T>>9&����I�ڐ�}���@#�c�JL�dK�`��k�R�^�y��e��X,��!�g�&0s��21:&�o� �C�i ��ƄJݧ��q�B��qF9t���}��j��"��9�_wٛX��M�d	%�i-�r����I4h�X������ CB���H����L^��EhނM�'�p�ݷ����Fԓc�$I���V`B�Y����_~-3���� P�3�^�͞��N��2r�/��
5"v�E��g�a��1�;�yH���.��M�%�>(�%}m��F5ب�d>W����f.(��4�B��k�H:����K��p"%���nI�S~�Uo���~5�m��<6<.�^p����;�p��m�iW�yp��5��(,	5�7���Ї> �N��=�q�Ξ�����am9�B�����;�y���O�S���C�J1D4Z�{���<��3�_}�Fփr�7�[��^8�L���a��ټ~����]p���F�7�������h��.50R��f��XNŦ�3�P	�XA@�Н�0�����V����w�+��~�:�&���������ȸ,�Q�6 B��x����G9����n���-�R?��:�o�M>�;��BF�����1����5uօ{� ���d=�TPn��n���4б����G�T7�d��a�13�Ci��ll���o�3��`���lـTI�ff�>>Y�IKn�E�Yf����Nפ})����s�Z�~u/ f��q�?���EB&@���Ġ�4 Iu����@�*�2)Ɠ`�;;;i�!��'�]�ܺD.#n�@��[a׺�p䭪	�3�fѠʓi�� I?WA1'h04���/8󓮝{E=�J4�/"��{ �k�򚗛�-=nnB���8pP6����ZY�����ell�I2�K.:����4I������l;�{&1�<b��Ё
V1Bd�=7;M�����哟�]��w�Q�n�(�?��t��&M�3��� ��1�B���/��  C���E���t�M^�4XH��.��d�Ή�I��v��y	�t��½��3��^��ԍ�[D������I�L��3��7���rԡ`$-��@\>�7 cWŬf,vQ�k�6�^	 5�.�+l�do�+9V��/���.�l͒�xJ����±&�����̧?!�n��펍s��I���qЖ������8�[�`��>: �"��"�lWg�Vjj�Y�	G%�/s�3����� �
����hc5|Qu�P��R�Q	��,.�z:c��0���ՔL�{������}��eܱ�L��j��AjYT:�o�� f������n����!P���X��ſ2���������t��MQٵw�:>��:��<��iK�&|�}�`�bN�%��ڷ����wq5�y�����b�\�(�+��Oȅ۷K�E��������80$�k7�=�q����u��b?�?M�L%˖G�Ϸ�YbP��Q��$���E�9]C�Y�8g�9Q��*�T/����u�H�����h��q�����:9��CH��~A�~*5(�?D>��?#��ǆ'�9naJ��<�a���/�ߺ�� �㻺zaZ>u�2��~�a�b�y�� ����|�8��3����#���� ��/�\ AF+1Z\���$[, u¬2Ȓ�Q�[Q�	8<��e>�7�<#_����Ig#��q"����hQ�Α܈3�aC����A�@kR ��@;���:y3�TAYUx���u��
f3|��fx�e@��@8�Y�g������K��.ؚg�yAn�Q�\s�f������CSp9z���\?K,����[��	z��/<Y3�>���^��h���m��/^��(.���c������>��ʺ��`��8Y�0H��](�ҔԿ��;���<��C���G��iw<,Ⱦ8�����S;�%6dafD�mU�!r+v� 1$�QQu��G{����Ȁڕr{��^P��~ͨ繾�` I�FCLT�i"8�L#fᰱ�Pr�1㛨�f��`&'��SP�!����������v�0�����&�:U�)U�[�q�}*����*5��ቘ:��R��l��1� �@��ĉa���M��QC0���Y�Ӹ��S��*tBp�E;�+^Ϩ.쏪қ��'�J��ٸ)@S�ǃ�+I���fȃQY�����#�H:�y�z��u��A������ �!�5 a�:� ��>r��}Q�˨�)Nu֬�����]E.�1������YoO.�`��HC�@nR3ː�p���d�i��!�Yg鴹5�����,�P._�?p^�܏Y�@,(��I�c��}�v@� hy����n�n\�B�dtl�փk�9M�O�	ͤ�tS�Ob�3/3��rh�>Y�jP�:��\ͨ3pT#��-���x�����p�U�։_��iiь%9{�7���
�����.X{UrP	\?3�NhP����E�������fa�f	�����麁Z�9�M�$�cj����-�6f�(3�Z��ƣf\
k(���#��d����2�p�������HF%�'��z� �x�[���e��(�ڥk��=�ʞ!���VA�CIB'W�$���iA�*�)�Ѣm��(Pi��DE�bWݬ�gJ��ՠn�����6=r�|�Fv�9��j�+ȤB��
y�<�䩚�N��W�q<�"�hx8QT���cz�1?�u�s����¸�J���{����!������Ao"�>?12!_��w�?������`�����X�^�=��,۳���rG���Ϋp�/w��ܩ�s�9pاP6>�?�����Gy��w��o�K��)��s��7�^h�`-!�oפ#�IׁCJLW����Qx��h'�����3�����[���5����_.?��d���ٲ�AR�H4����c]@,
\�_l F���(9֔�Do~	����C}*T��F�$O�u頮�T�[�qX��>�3�l�&f���m��sl��EG�\+��p��'�g�����������o��U�f J���_�Űj�j����Igwi�j0�T�13�9 ���@�r���s���*U��7��w��9t�����4k������Q�W42���1������$�eVD�8?�����q#�G@YD�?�3r䬨I��� )[��t|��Q ��v\���D��k� �A9�mAs�����4SG��(^�}#မ�%�s�lp]�@��P����P޵ɬc�+��#����s'H���p\�Z;���lk2?1+�)�/�i�!D�T'jyF�4�~���fD�Y���h���pl>�|iҟ���M/���O��qނ��)���`�F e�B~Q�[��a#�6��^�i5꘰P��w���9@V���PDX2s���=o�6^�y HY,H�P�#'*\ϽX�rv#Eҳ��_�A����	I&[Yr������v<�f����i�����v���`�H��_�j�Z�ā���E�>v�����[Zu� �����C>@ ʹIDc���=I�% �ՙ;��B<��k�
�j�Q�R;�FVg֡x���Ŷ�2}j��?_����1�!W�v�`�bYZ�)�y+h����#�7�<~�o���Ai�u$��'4��l�ZNA	��bt�Q.��'��E��~P9��ҮAg|���-R�k���S_��s�"���h��-���d~:��Ws������t����O}?�g����?��N�o�#�������xB2?��]{�K5W hHbqӳ�tO(lT'�d��` ��������Aw��Ts�ۛ؈7EerbFң���OZ����P�Ab!;�-��G�� ����Q^�:h�k��R��D��p�9X'��3<�5��F����`�Ŕ�յ��8*���X���9���|�7 �M�3�b00�_]�:9����l�mut9�� 3�[���9��0��,`Սƻ��e�ڵ��:D����h0"�B�=��V�@��C�����l��tn()�|˝r����(�=.��X0�LЄ���P9��|C�R�����J?0�a��+W��G��n�dg� b�g5F�tu/���a�# �eV͘A�P��R�Tɩ�T�!�^9#goY���Ha�0��k^�Cd!�>-��k���ޛf��%���icA���Ϭ�H���&8�(�!u�(�#�By-��D9ev���}�~uZ�n?��M�3}L�n�-�V�H[I?o�i&(�<�y�����K�B��������	ȩj�������L5GcU�s�4���/mb�d�4}])��~]�oKv�� O��l?o�$��y0� �IHNP�A��f'�Q�.P֠sZ��<�p�1�L63��|��[7�s.��i������k.��*W �5%;����Te|��m�p�=q�k:��9\�;ٲ�%��MF�iDb�STK����aٸq�|��]+�z-o��mf�ft�;�%��9��5〮��:h���R�2����,m9�{�Е�{̃��'�6+@��TÍ�����tT%PI�߲u�x%Ud�x.��z_�&�P$�qXz�"�:�D� �1��|�Ba3 H}H#x�4��P�b�+��z����c�/��c��;l�	ۜ`��	]!$j5��7K\��w��r��Wh0?��rqO�����=��[�����ڂ|���L�L��=`��@��7�����w�M�Of屬��M��\�d�x�{�(Oc��H���~v�B�P�w�3�����q>n���A#�P?�W!���իeB�5�/j9�Z�q=�����з&��@8���F*���~yh��Y�:fd�p&�<���cBb0q��
�w�9g�|351�Nb��}����I�4�>(;w�f�d��<d�j�mK�#>0�3SR��	�
�&؇��a�3֠79��A)�Hv$d�,ۨAA|�p�0D��Z��d��0���C��,�TMv�r6�AI���<�'�h�� �qz��"?[�Rc�X��5�r�7zԩ��^+��>K��8�sjI�\p�A����1~�E������{D	�C�e�nz�5Ww�6c�lTUe��57�zM���? ӓS.�JX�"U�F�p�/`b�C]M_#ՉѻN+$�X�������M��)��֞>�G|�
���)��
��Tg����9ÞIg�k�f^������6�����.��������T|���"��z�*�h+�reH��UHE�Nra�2��y���5j�h��yn�\��D�Ct��_�'iJ�ؒ�Q�$+�}���k�sV���pQV�j������ww��t�-�ɇ��	���v��Z�����P!6s��8c����%[��$'�q_��S0z�����y�l;�d�,w�{��?0���LmP�z�af�]U3��ڲ\���0GҔ�O����B��"Q��z��SE�<[3���d�IYn2���G��S?>�󅁶����c�ە��1" �2��GK��V���FP��Q^��k���c��
F\���;�9���wv���u�qǟ���h�����З�c��%^��	;~����fPL&4ǈQ�f�2�0'�&��M쥟{�E�n�
�d�6�W��z���Y�LQn��^Y,�5XL��ni|6L'h�`�>S���A���?��;E9.۶�+�=O�1�xB7��jܗt����ҳ�px�̳sF���HĠM�}ԤAl�6��|Á�d*0��J@��Z53b-�&�y=�CA���V�6��\�A9'�Ͳ<�y43����	��U��<z�׼�=r饗JO7��06q�րx~������H���q�hD[R25��x�f�&�/2w��%�R�8*����FK`�Tk3˦�D�udy��%rxco�Ը�߉}�E���w��� xr$��Uh�k���x.4v���ɽlݐ�`a{��E��eu����j|RɈ|���L���;"�òM�:0����%���<3�L@��:%�
IKKI��7�i�[�},��%a�9{��u��M�&�ɵ\iD��������]��s�����ƍ��j��NH�f��:���R�srh�Q�Kщ G��z�Ϳ|�\}�er�}����c����Qck5Kb�V٨�36v!���z!'�cѳn�@gN�O#�����\������k2��A���^"�A��v�Z���4�����1^����A_\��z�p�w=%��}r�k��5���wP�:������'��4�z��}296$���L &�n�
�����^�&��o����SY�j@%�(��N���2�ٖ!�1Cq�5p�C�)��@��y0�vC��)Q�����M����@��'L֣�>_̸��V�,kH�f>��Ջ��ӕ�OBQ��I�V��o2$5��کS��*\p�Yu�蹑��9#y����~�
\�Sɯ�D#�L����=��a��i�d�1��Q��m(a�D�����H���,��_�����/⤝WY�x5�5�F���*�;�2�R�%�qh#�cFr���ֈxka������8(T?@�Ҭ{՚c��~�d�h�������'%���f^v���}� �\�1�F� ��]� �BPK�l1�O��?�2��H0��_��d�p����bR�V�:��@ f8O��<�{z�9t'���O3tu>(�Z~�Y�P0��`��eN�0�MM�I�� �z�Z������R����ب���S&g'��%!.�����?�O{�1}�Y�ܶq��,�ˤ�=�N�ʍ[f�\�:]H���"K�~��Q�Q�F������dv���a�M[�L=rq�DB�k�����%8' )Q�(�3�C���(��e{�HV�������KW��52f�詪�.�P< &,�e��C6oZ+��ݏˣ�'�'��vu"붬�cG�������,���a��XIs�ȲVg��\����`�a@�6JN�7���6ѼG�� ��S���3�qL��6�$����lDWH�_����#��,u�����ɇ5:�ށ���_�F���s�o���c�?%�LI�S�z�J	�<��i}����7��Č��h5�s�Q��h�*Ő%kV�ȝ?�Q��'�{����RM������fU�:��4�ҡۣ������\7�����t*(�0cޖ��o�EοD���=������dz*ǹs��ܿG��_�IJ�y]���ӿ�I��Y���>&��,%�p\�{{$���g�Ҹ`s��@����5��g{S��5{�:*b�B�LWՈ5�o~���+��cǆ䉧�&�m�%Š��l����AZ��r�I�[n�ɞ��J�K%j��6��U�`���n� m2�	F�#��nda����^���D5 K�a��,�����bt�$A��5�XA+{Ĉ�~�X�i���o궽����σ��_B/������� x�����{9���W
�՗~�Ҳ4[N�WWZ�}i��F|�v�и^��T+�(�׮g`4|b\z:�LƀmJ�D��)Lw���*���6)�6ey;�v����h2	�D/<�*��Ԙf�a�I�݇v��p�G��50FK�8�A�t�F�ճ]X��p{�hEA�jQ��a��}��j9x������m��:�$��I7ġ�ı5��;	�=zG?K��+�j������l#٬N�'���4Ni��?�&ɖ�LN�����Ɛ�����P�v��#F(����v�se��u��Aw̪P��ؤnh"}��r��A2�V���YU0��$�L6p�.�̜~�4��@y�s�Y}�	j���b�hZ� ��d�N�iS�����9�0�0�.�K�i7������x��/sJ�V-�{]�W\�Zy�{�&���@o�\��wjƲ(����d׎���S�S?�sp����F��"���L���\6��� U����_��l�To���Z��ݬ���!��`p�O�2�l�y�1��9g�-�gI���>�rW�9�z[��He���=�>��Q�9�[��!�_�F�__���r���?��ulY��-;v���f�K̀V�������?��M�s��������jND�:�M���;��vI���������ほ�5��C����܂lذA.�~�ft	������N���<'����^��K��M�����}\N�XQ�8+@������ryٟ{z�|��׊/�$7�~����S�9���5��>�_;��<7F9m��9J�a4��WM�C.�h����U+���	��?~�ճP4�׻Dq�pS����YE3�d�tE#����`��Q�ٗ�"1NЌ�V]42Zq��!������t�.>�h����F 	c]s�
^�nK<3���5st�UE]�����9��v���6=Y���Q�5�JS�w^9�~~ �z�)v�i�Ա�Z׻���X^1�-�Oj����@o8.$0��Y��#��`S�;J	�n�Un��;v�2%�*"�'@<��"+"�SjWú�sY�G��l�a�x��A�59��W���<D��#��ے]2=�ր������UW]%��k�&��z+�?��Z\��}�H�t�}��
A�k^����y�x���|�����y�Lk��Q�n�s^v��XP"!�p`8�Z���\����k�B䭏�Qd�]�G�Z�Foּn����������4�����(7X�|��p���[��M�����ɕ�*J#���$�%I�����ԒF����\�֖���s'��=)u�\�e��$4�h��-�c�m�H�̃��/��r�j����oX���"��4Ш[u�r (��CZ�%�����Ɛ��7,�+�u$ }���hNh��g�������kF����gٸfP>p�{����Ѭ�c������,�q����R�bx�X8�e5HCp=a,����@O�?�����@�g8}S�5�:��h�Ɍ�����2YfYS���u��1F՞q�kO����H(���{��ٿ_F����G$L�W��m)��F����ܧd�� G�>��+5+�=�����db�&ݱ2u�0��`L��Dz4x��������D�+z���L�jf���Y�)�,3�)9�H~r��2;7/�6����HQ�bY�]w�%7��5����Eo�Jr��[�W\&���;,�]ݺ�7IkGH�J��S;\�r`7C�)狆xG��?�w�#ܟP��,<�aI����:EK�
x��1ޣ�-������@�D1��
%9��J�Sw��g��/)�⢨�z ;��ɬi^Ay2�*�>����L�v��0Y�@YQ�uP��!ڄ�:(��eA��k��>}M�Ђh�^ThK���p�Ñ�"��V���U����ߝ��]F��4s.'�����T5.Ų��Rǩ�t��9�W|�[E�|�H��$��
� 2�~~&���i �0�U�dr|B�b��i08�/'N�mT�A��.�>8�.q������<z/`��]F�k��]n�ס��χLߣb{��~��|>�=�>f]��U%���ׁ�:�kݺur�e��B�y�fy�o����p��� 3�?�5��q���v,��4)AIU��Z�3��P֪;�|���?�|A������X>K0H9��4��ŝ7�j��hnmf)�n����iPeB$j�y��5����mWO�#>  �H�r���SzD����'o�����-C�G�%�����9���
,�:�.���sb����6��@�;�v��^��zd�D��cT���%S;?._���Ƶ+����jy�\u��埿�O���(�ȇ�׾�}U�v`�P��;K#N����nubeWw�E<|�B6C&�֦f^G���`31���@LZ@��*����.�
��Lg�t� #��
�2I�335�����f��;����cc�~���Y�ܟ|V�AX���?�����a0� @俁bsI#��~��{!��)�@{������ ZP����D,�,�Q}��D�}�,�f�{��n�ZY���#2�ۧ�z@�zu�n���&��?���r���e�/��y0�8���3;�s���0����$d8�15��hF���ci�DQJ�QH	#Y�)Ⱦ4�>?���.�ۂUF�h���vPs �Z�aR"*&Uݸ�Ь�9[�����Gá9f��cG�W��i@Í�}�e�u���YH3o\8Âh�.oɰ������J�t�Χg	�*��{�pl| ���?�ܶ�v�:�K�ʱ��7���9u�|i����r}�W
��X^�`p௛�WJ5���u�L[���EE�1�^O�U8��b|���W�g�7I�GHd/@�}j�xA�8���#Ң�i����G;�5���>���X@v����'�oS�&(0�.Q]?\p�>F�L���o����g�}�`�t_8׫63��)��Q�:c{��_:� Y�k)UȐ����$��Av��w� �S������a�afzR�(Y�߲eJ�;�锣G��`�H�ـc�x�j$��U���
�/eR�V�+t�������M�2̈$��w��`tc���U�{~������S�`�f���c4�~C�A�2E}x��G�4ԍL�����Hⱐ�g��o{����?�亮;Eg~�M?�ǎʿ��7e���rx�n@8)3Si����ȅ� 8~&d�IS�G�seނ;Fd���8'<>������b�Ҝ��^�%��0�H@�U0�a��BoNi��Ne%8���e(x��v�ʕ��keӦ4��׭�ݻ��?�ӿ����/�SO=#�<�����ۥ���5��Nn��.��b�J���WM�"Yր���E����zݤ�L�b2>>�k%/��m�n�j����e`�Kz��(��X�������q{������y�2��XȮ� �>�)y�����T[L::�ȼ ��?�!���r�2�e,Ue+'��*`4P�H3�Q � n��R�]��K"��� �	����� p�wؓ`�3��Ս3���`$��&:Ǫc�n���hv!���W)����O�{�Lo����X�PP,���ĺ��Z	�+����̚yϸ�2����T��ӾTkM���T{�;�h&X�E���s�=Cޛ�7�5VO*���d�u���q���0�myN���+d��.�i��+�l�>����8�@��J���	*������I�I��_�������ft��f���G]R�
�k?BF:�3�����+�U3����
T.��@�W��i'f����BZ|���(@ q����fE��5�����ͨ���<��ݻw3�K�� Ne||\֫=M��˚5k��X��=ỳ+j\s��8��󅬀?��$��s�h�2�A��s��wP^6��j����W�&�1�S��H>  �	R�6���5v{��e�g�,����BJܐ\���4q�/�Q]��!�+�X�"2�"�Q��2�k,����l��oQ�J���+�ҋ/Q�|��tU����py�9s�"�����1�l���(�v˚�J�PoE��귽U�x�)���/~V�{�I���_�w=G�}�q9z�t���I�J��[v���#ǀP!`�����y~. �q�s.��(�.ʸ�Gv�7�x-�(k.������0|s/�FU���B^��)+��
Y1�QZ\�+΃�5(��Ip����רs픕�rӭw�]w^.���"O=�4G�n����w��O70�~~��g�N�P���KJ3�yijN�~��&�0#?�3�/���|�Iٰ9�`-��bF��:��ML�I�`�<��}j�*r�5W���̨ƿ*lߢ�.-�=�������;����*Y�z���ʫ�p�̤�E3���M����2��^o ����e2�C��q5,Vc��>�r�,g�!a-�s��+�+���9[̡s����J+�������0�s�O^��{��#�X���k8n)��2D0�\w0��C�2�Z�d�����6Œ2�5��Pf�t�������֐M8�^����߱ 8]`	�M��m9�3��3F��%�:��疱���[����t���W>l1�#v�����]u=��S[��I[KB�R�b[�|�%w�!XM-��
8�r͌�Z�S�'&�9�0�UB�1����Sws���o�4�Ô	.2��ep�������Z���� ���:���qNS�w��d���:*�o|�ٞ�������Af� Wg1"
;۸6Ι��5ۤ�U��pYR�W����`k� ���"(3������d?C&��l�k��!��܄ �?���׽浤�<����?�d.@ s$�4�7ٿO��dfnT_kNb��0��R;�tq�ca:r 2�ۺ�@̓l�` (A��:΃C_��x���1~n(�A�j݆M���ˈ}w' f���%7��T����x�{5�y�%[��?��Ҭ��]?�C����)j�u��eQ?ߑix;5�#���fI����@������c\�6n��s�ݫ�d0A>�F�8�2d�N8�ӈQ?�Zk�\�<������8`0�ϐ��uӛ�(n  ��X�[�y�U���ϱ�s�5W�����9'6����V9�V����S���;���/�[�|TVm�&3Y)U5��e�����;�J`Їӯ��$!YXX���ɡ��$�)��W81����d���NKk�I��<�����f3Y��G#��:�O�������FVɟ����n���[�f����I��w>���b`�ſ��@�����^]�s4RXo�f���Tث�ʑ �Y.�΍�H��ڢ͂,�����G��`���� V\���w����>�ӈZ������Q_n.9����S,�I?5������R�W�&LJ?��P�@�WB�\5cz�;�k�����+��k`�3�=E�"oʼ��lN��,?��h+�Lϟ��F_��W������d�\�n���{ٹX��5��4��r,ʟz�_�/�ɢ6��ܜ��Ao<�1�E��7��4���]����.�lV�Ҥ�$K~
�p��rj�`�)�re�+(��7���Ԕ��e �}����f�C�Զ��Y'�=��ڸn9rdVJu�q$v���(��ٳ��{��^
���kǣ���ǚ��@`�qU`{�X�����w�E"&�n���n� >����8��c�}N�+�Y���l�YG� �����&�9�y��J/@FoٴV.�p��w�|�ɧIq�ȣ�?���r�Yg����+r��ˮ�;��]�p`�
��`̡��ӓ��n;w���&d^���c��t8���G���h�QP>bfӔ��E�R��S#�x2)�}������%�����F���������eeq־����5W��;n�U:Z[�W])���n�Z��YI1�Ӭ���e�իWs��.H��`��-��8������ģ,'��������#�@�Lj	Id�!�ْc6�-�<���詡��;:v}��^m�ԙ@2�`���e�^"?���+��.]~9|�tu�4��7��
���g���+�"w��$u��eݸup4I%��k�@-�e�P��$h�e"hCu��8F�ǥ��]֮�Dހ�C�253O��.�V:z���qY�f�|��}Pn��F�֬�{������1����}^�q�5���!��q���G7��}����_ҙ�^��d5XF��F&%���
d�3F|��in�m/�k�p�J�3@�h��Ao�d�>Y%T��%�q��^�j�d�/���a���r*�_t&��Yrx�q4���U3 \�D��BC�- (C�Ɖ<�0�g� �|�,25Ԙ�7�2;*X���x�qԤ�`��pT����`��䆨�b��f��7��+�����S��~�,�SG}��d�n�ᘵ�s5�D&�zݭ&r?8фdҳ2�����	�/�J��6yh�æ�Pz.W1��n8tϑ��o�5�m�o|㛲�K_��|�7���jDN?*ɶV�B=;��&d�o��w%�U*�%�4�$Y���Yr���La����wwtI����Y�}��>+�tҵ?��m7�Q��o�$a��`�lp��A'�_[kJfƏ�	C����/Ȇ��`"�,����t�,��n��u�[��ѣ�����r��Q���F䎑+�����M�z�v�����:�����Srp�~�z���{� �\�ƾe{G���3�iV�-qJ���Og���ҡ�AX~����D�XG�q.3�Ζ�<�k��z��Sq���\���s�٧���/ٮY{�N;ٜ�4+�g���vuq��y�r��1�p2K�]�(tyQ��'�V]JÔl]�h�p�c| � ʹ~J�Ny����ܝT?ù��Ȁ&Q�m$ɑF)��hi�r�ߌ�����4��`nzJ.��r�n��}�cRÌ�>n��urbdN�:{妛n�7]������ݎJs�C�̓���ҡ����U�����F���}2������8'��?H���?`��16����8g�'�O��z�X�R~��7h�_�/��ۏ��os6���p�����ƛ�#C����^�|�5&�A����@�$y��T��)t�f���/˥�tܶI�������S]n�k�P4�lz+7n��/��z��4�5q����~x(t�2=0e���QN��O9N|��3ju���&:wTʝ�@�����#� r�B����S(��@���"�ȂK��K!�6%�/�d����������,φ�s��F�޷���ۺ�	�@ 	B �@xzH �M/!!	����ӌcp_��z�����J+�V]���s����sF�-v�_;����4�����u_ł�p
�A�ɨ�ݑ��,Aa�#�T�cZV���;�]�A�;[����=��z,ͬ�ރũ��9�GO�Vn<�hU���D��prB�Z.5�/ۄ_}�͘�>��\3�c�j�����܋���L�d��oZ'`�^v�� ������qCG��G>�Q|�3��������$f#�9��c���>�e£�������F��.�
�r�/+�/��� ���L���v��a��x�#�jY�t�ؚ��	�@��0$W9�yL�WN�jZd���)�%C*(Ukؓ���J^�oġ���o��������7����i�i�1����:��"&��,��H�q��mjIJ�ԉ�.�(ٹ��lZ�/��f�쁟`׮��9��g�H�N�N4�dP�����Ȗ-�$�š�`l|�̸;�R.hVkz���fv��Ln	H�P..���TS�5`ٰn�j��MO��+.S�����l޸I�Rܤt����hL&M���]#��Xznz	Db1
ajW%ױ�Hg>�
H4�}	r2��Ȉ���(�gC�D���C�FF�Qa�^��K�u�-�,)o�k��xFuݚ�8qr���#Gɪ���|NW����c�sr�G��ӁGF�ʓ	v<PRR�Z�0b$"I4I/�\���N����7��J5@T�:t��4�!:++d��Ljc�7ްJ�{��ŁC�f�z\~��X'�ƞ=�0r����=���_�Sxr�#�ƒ��i�5�^��w��ɞɠ!�|5� -�c�&�8��U3V
4d�P���N)��T��1�q&8��Q1VCǎQ*����ktO���Ƅ�e�̨�k `�������c��Ѻ}��Z�0�X�z��@-��]ԍV��;:�P�X��W�����T�� =�ܸ�BzLmY�Nh��6�L�.���3&#�½�3���͈&��KIxF�����[Y���k@�pC�-Oֳ����;T}��}
Ԑ��A�i�D����`ܩ����t_t$ͻ�������_J�c85�U�U�*���1��6�?�u˾"�����ɰH�+�|th�=��C��?~��Ӷ�k�)^D7�ً�
!�'E�b�����S����'>����?ф��gwbՊ�j���W�n�?�>���M�~�Lq��+�1�߶wtbp���\'�HI�lҳBҙ�؛`c�j~pr˭_��+h�Ev���G��,=�AE�k�Ϊj�HI�@�Qnb�P��)ƱW��%pH���׾���]x�G�u�8r䐖���ڍ��v�ɦii"�!��ɴf���$��4
��D^)-���t!!p�~[�R2*�_�G����]��.Y��MQ�!�܂4�,ӒBu~!�XS�8m�>8U:�R����44Ĥ�%Ȉ��̜��f� �G�ӵ�a�M�q�<&��(-�M�������%0$ƺϿ�W]q%�gR�����CX�n!%e�74֨Xi����uk�;���1 ����S�g�ٳ%5����e�L�ߐ��m������gYwAK��?�gVʋ�wǮ��y�~o�A�ɬ,up|x�v(��K��v�z<����Œ�NN���F{W�IPG�2<2�_y�d�� ���Q��Q��b�dvQ�hg�����::z;q���Ka�%�#=;�-��Xz%���7߂��a�JFΙ~f�y��������GP�o��w�s�&	�d,��+�O.��b�<���薠��f��J�)�Аl� 3/�/{�m�@�*�����
\cV' '����u6�Z�ZDK{�<�\�ܗjP�	����U�F���%�p��^����
vU�.�� t�4��+:������Mׯ"ycWZtf6�C��`4��/����T�m@s�r��1����a+�����~fj�O�L��$�	��c�uu�<)g��s�sU��?>��3�`�̹}Nep��lrt���O 3A���ieN�9'kFP)9�ٯ'�;�qTo��]A�l��
9�Se�|���}N^�����AXq	E�'�+P6A1�>c��/�aא����Ή�á�9B�����_��{����%�[��(��!����&���h���Y^'NsttL�f3S�H��[;�䳻d�5�a�_U�� ��A�cV9b_�VT�/��ܐ�������?����η�?|�+_��}�u<��Ƿ]�A,|�!r$�E;�s5tw�H���)���3������Ԭ�}��)̤g��߅�M��5�����l�B�������{h��"2�5�m�*��cg0p,۠HY�g��S�~VPa)S��ߔ&2��p�-�5�Y�V���>��7�ǣ�=�e���u��_B�l�g�z���r����\���T���h��^��ة���ᆛ��X�E��2��i�1s�q�ˍf����$��,�?#�C��*���3oH(:R˂r���f`�'�@���rӳ*aՕ�4�c	�h�*�hP�\.�����{���'��4��z���4���k*q�����*e�V��G�|v(=�r�h���ѿ�\�|Y�# h�Y秽��]���Pؾ��'*l��0%8ҽ�S��>(߃�"�[�@���F|X2��5�e�eӔ_lU��W����:5�����ͯ�����'��Y�(��@&K(�c^Y���״L��ա���),<){�)�\�;��.ttu�;w}O�3>��������g��w��d�̦敂��1����,�' �����8�=���"��X�v���K9tt6Jv9��%�ɩ�!H�R0��~OQ��|~��r��S)/2��~4��3J��ݳ���G+,4Ǝ�V��/Ж�KP[�`��G�cB��w�ga����166� ���U�f���'�������}���6�)h&sc�� K�j�p�X-;#�g�aQ=��;3u��y֝�����G�8i�j�i�NDGs���C�{��vYm���$�����Ri,`(��=�y�[�M��� qgM�g9��q�3����+
�7g���H/���
��w<�\�ͺx��q��g��%U5�=�"�I����|�Z��
7uR)V��퍊!�b�)�����w!5=�U�������8֏��� ���Z"�� ��?��o�L��Li��mW?�kg���۪��Q�ɤ��[)��=)���iE�fq^;��1z�KvY���np.<icr89���0�*��T���B��DP����Ġˡ�nC6����.�\��\O<���^�Ʀ6mلG~�R�����-C�ʕ���2�N���Y"��/�V��D�=�8=*ƸՒ��{UV"Y���L)��;)gdg)�)�`��9yҙ�h����2O�$fϊ���us�:}��Xvd�Tuk�t���7�4S$�l��SCi
)q9ߋ��=I�z&F��f�k���$\ѸK�m��U�����w��;�� ��vW�D=�f|���J ᚹz�u<]v��'�X���3j�QuN��\CV*8���14�w�,�ќ �߳�q�L!%�E�l['Bl��ɏg����q��W�?��Ϙ��h���Ù��,��(���3�Mb�x`Iz(�B�:(s!���mbR�F�*`���O!Mbt|w��uflb�?�.��Fu$�5���Y�;�&����K��t~tb�\u����a|�# �7v����]���*5��LnQF�x���f���8Z����z5�}�z��(�p�3Ǯjc·se[��N�Ì�����6������Cc̈�L�:���I�c˃���hml��؈�:{�5��=�1=U������5�:^L�r���S׿!Ø�U::`:���	ؤ0��%5)�������]2�L��g�gj:�mm-��T%,��C�
�do��>��y���Z�k����¿�}�^�'^�8��^��s���{>��EV9����|��QI2�X��O�uN+G^)�{���1G����G�ֶcA�"I| hr ���y�p��\6���w�Ǹ�ʋ�������q��>��d��z6�:CDm�qa���_O�e�ޫ��� ����)lf�u��$i��cyb2j�B%����Wm����[R���W����m�d�@Y���2��K�ނ|-����W��*������sӦ��p׷�FKg+~��O�D�HV��ڨ������>O���Өɖvd%f���I��~(�A\�up�lBf؍��ᘙ��9O�O G߂���HLKB�����]�DcB���\��-�|~!+�"�97�A~��h4i��j�Q��e���*��=N�]!����dF�*x�Z�&	��Qs�-/;�{�QC{��O����Q�����p�\i\���dDk��Ѩ�����`�RO�,�'\����h�_)kb&��}�LV#�,ˮ�-�I1�a���4��p*�}�\� �Y��>��U��`d���o�h��[I�m���ıW���R"3Y�����+V�П3h�k��)�>T��~z�}x���+Aay�Q���W�:&���-�2`DvW�`�Zݍ)	��E��my�R�����>g󯸲�s.��f-v<���!��@TQ�s�*�>��5[����A�}I�R�J�&�Y��4�l]�`~|D�|�8y�����س��Ԝ�߲v3.4)Y)U��F�!5qA	��'Q\��[��#�ա��q����0�ňRg{O~���� 9������/���މޕ�qztԔ���@�p�D�fW�f�r��~_�GMT+ � �b�g�*꓆	(g�N����$��N�#�y�r���8���y�����S��s��{��c�Wa0x
�}����Ne���^�C�������̌��V�^��Q\}�5��m��ǝ�d@m��kyS2�U%�m�Z��+�I����Ɔ���c�� ���g�!�̽������&��=cW�3�z{�W%is�ۖ�ۉzgPX���d��G,S�T���>��|a�ܭE���8�Cg���Eq�pt�A`,$Y��F�O�}��Чv<�DK#��с���MT���9�V����N��mm��?���Y��Y1�MH�]̧�O�	`��P�L����ظq��/�ڻ1xrH���Of&QT�����I�b��AQ�i�_�U�ԏ?�S�����o���̋���y��k)�T�ͮ��u<��������(T��8l��M�����'šR��IQ1���D���I�,$`���<�T+��A^�0}YT���W�T���%%w4f��=)���L�a){৥|㖁�NfgQ�H��c���N�>���}��,S�^����fU#j�g���!Nڲ͈Qv���J��i
Vbd��q�؈"�e�� 5�Zۖ����q��j��]�����s�Q�D�E161���CI���g�ٽ[���Ï�K_�*r�]2��v�r0���2NQ�te��5��. ��d �l��c;�8h�1c(X�����ꂣ{H){���Apv�>�l���GMD�x��bu][����8�@���n�r\{���>�:���i]���b�s���~����>=.��m�����_���2ZQqa;!YRc��B!=�Vq��E�x*�KG�[VΓ�:���qU�{�,��A��Y<ւ��	�����"�<�ln�W/�ɓ�r(B����FU��Sc�P\PIЛo�[�^��|��N�~��(.�a;�Y�#㩝;�b�s���t^��\Y���K��M�?��p ��!�;�F6u7]%ںZq��m�����~�����S����BF�A@���m�*�E�A��HP��k����b��������^s=�zd?"L ��f�;�h,fڡK�/����'g&��2�4��2L���õ�������
�c"�ܳB�K�ⱜ�d�O�dk���s�c0�����>�0ԣeW�Z���CbLG���h/���yq���FZ#%"������H���ݑ.���ɑ!e+��Ќ��o��(�����ถ�9[\	%ѳ|��&OON#/N!��+�S��C��������O�F��q��+N�]������#z�5�I�ߩ|�=��F�e�6��1��
� ؂�gn�\��*kY�*�@��Z�3c]�?�2@"v"ʬ�L�%v���,�8#*E	+ȥj�R�v�zQ�_1�A8�3������ޡ�cQ^$�G�Z���߯���x|�N?����33�%_=>xS�4})�E�`PG����n��ؾ��iΨ Eت`6h�x��ϑ
����&"�Y�m$�I6�)�<�2�J!��&~=k�o�h�[	هyU"��ʁ^��-"�ZU�kn��mR�a�Z��[�x=�z�����z+���º�1����r�/�QKJ�z���kȠ�s��8�x���X�v���<��#����1��H4��C�10������>X�,3\�Bp|ө����܏�/����K�rn�!,�H������]xRr�)��������>��]��y�/a���:���mسg���/����c���׾���lۥx�+n�׿y���:矗L��/�� ^���T�R81�{.�B���[s`JK)�bUz ȹ������o|�m����%�<�h�)�ĩ�2�~�*|��"Y=��w>wǗ16>���n,\C��#kz�����8�ۙ��|%�}XK�?�#ۯ/��;Ŷ[,�\��?{w�}7^�˯�Em2X)�uY�}�b���T��g�j��W�4���>N�������A_o7��G���ӧ�%�s�v�
������:bJ��/�ʠ����~nۋL���q���碚1�~��_�U.��!��*�Y�i�Mᾢs�$�k����*�Ҧ�������D�F����]s�Z1\%���uvnG�Uu.Fی�Z��MO��9� �|1���.-1�h��R��\!��g���=�Y��ۑ����4�$@sSV�]'A���ʟ2󞜝�F,l�E��d�V
�;N$�Q�ʆ�sR>���3צQ��(9��u�$��{�|�r�?oIeW-�9��#���Ū(�R�͚��C�X�a3�۩T�:W��)`�筗K5�a%2����e��q��?����ǔ*f��ٖ1�U�����h�t�Ji1cw�Z�^C�s��
j	�lUu���T���"�@���+��}��!�+Ƒ�}���l��+��L
�L�hZRW$c�^vl���+:�e2ZVy��$'���(Ū��0;� |�K3wb��-����bsQ+,��D�Ɉ�����c~_��CgO+����%c;�",�O�رc���i*� 8�A\Mn��8tz�MA�"N3,[����(���kh�U�+T�����'��{������X�Kd��TU�X���(JeL�l^�.�=��\Z"PB���.�P����Sش�df0|� F�B[�����W#�pl�.��D05|Tň�NQq��y�c+Ҡ�O�B`/-3C�F�b<�����8g�F!��$�nL�05=��]H�M��%�w����.q��u�xn�Uؾ�IY�9u������$@L�fѺu-��������|*��r�4� O�GŹ��������sf��=�� ���/2�����yn���$(�l�6]�[o/b�8ڇݍǶ�B�8c�q�h톋��ы�S��|�fL8"{'f|�>Hf��d ��h+��Ը�����:ɾJ�<�n݂ɩӈx":�"�:�?["Uo^�/��;�z��q5~>*�m޼Y�%G�����$�u��\eB�� M��sl�v�u/8�N�ܪ������3A�s)�l^�b%^s����#�s#oG ��Y�c��D2&���cʡ������ҭzC��zt>�N��e�Z���� ���Iq���V�Y^���GT��P�d��Ƒ,{V6�m�z���g��".�����gǓ���5>�1Q�d)���ŉO��~g�r��%+K�,�r��DU�qH6N�6G����g)J�Hj�'v<���M��|3bHڛ����+��Z$�d�=�`k���P�Wu>�S� wA�t[���z�<J%Z�S��ԕ�-h��:?f�v�(���c��@}�� �+o���ZZ��xrzF�⠒$�0o�)E�d�l{��)9\ش�"�����GR.Td�8>e�~�rI�@Z��f5F�S�H�3�kWGo\l�pZ�	5�>-h>��
�ECJ��'������q��ʹ9��H0A�9�?�^}��T߽��G�id򮖋5�r�C4� ��c��iz~^�C����$��s�[ӣ`��P�LTT����g�bZ�xD����}���Ls�!*��'��ǰ����y�܃+/�(ge'��o�ᵲΫ1tL1	��]�Y.���7���[�H����mـ��4N�S����>�O�:�f��(�8�0�@4����F��)���q��FYT�'�ȇ?��
l�YՃϪ.AE���$~�������t7�����,[wq�>��~t �/ڊ�{Zɐ��d��M�I���ښٖ��·{�T6]$�Ϲ�O���p,�s���x�����R��'O���'�l��a�5X��Rq�Jk��ONVq��g���bqLU���f��X�b&=sO��E��&gdu9���ѣ�����V'�(�Ū.���������W)j��(����ӃmW\�?'���oքqϞ]�p� N� ����u���}w�Ρ����Q�����7��RE��#P�+���].^<JJ����Lp|Ԇ��NU�8s3�b+5 �!bј�`� ��C�<�	*�L���B�Z��X'��"w~��H�	�4�P��Ł��fAN��d�y*=�絔S������GW�2�����A<���J��̜ ��l�MF,&֠�_2���f4�$a���5%12r�ƨD��Rn�$k��s���Y�N�BYt.����$�Z�`v!���G?���O) �<�dFb�Z�B(~#_��MZrg)��7h��<4~�=�֌���,��F����G�J��eD3��HF�bl���#g��s��AR͞��{Z,S�� 6��q�a����1�#�?�<�=������ν8%�a�M��0(�|D�(j����&ѽj�����dKh�c~V���wf�9%�	��&��}@w�V�q�'�'�$�]��������)l޸��lشQ�3���+vY�TZ������x�/��I������?�����)3���C��d�㚖�&�	ئ��}�q�T�y<��Q��Z!��-r]s�ֱ��"�*�H4��1{�|\�:7�`��!�$������s4ֳ�,-"�)#珥�h,�ɉ!���^��]���q�|��� #^6_T��=��O��V�%���gM�!�`Ҋ�K�������7\��z�{7̾xPI]�N�>ԡX%��������PN��N�k 6jga�TL���	��Y��翆7��
Ժ���ȹ�*��v	�5B9��-�}�K_��Μ�`�5/Ξ�1�Qmo\�Bu<{Q��|�|��O\��V��9����w�6V� u��N
�qm�_*O�N�8��gKz~|�vD�\g�g�{a˥I>������#�J�K���M��}(r\�=q7޿��k ��"&K�L�.Z�eX�LIEt<nr�����,�3��>���+Q��8��$�g�k1��If�'���	}m�[��J�+�}v�|���P��H�h�k��1����[Ӈ���F]�F|F[k3r��")����j2l�5�(�J���譹�I�&%P9���k"VEB"uru�C�J�k����@� ���u�%�Y�QO��^A��"b\�H����)�=[$r�S��.8�j%$Q���3�I)�0LF1��,[�V	6J�E�f� ����h\�<�74󱜥e�3r�lt�4BM
�I�4k�aNP�d~��>��<�s?>���S�1�DW "Y�Ï?�-��K��#�d5s
���
�S�����T�3�f�(n�oF�G~��g��~˷�ޏv�Q~��6���W]/8���5�����x�{�60S�rC` �]�w$�xv�.�/��ַ*��W�;{�z��9.� ��O�Z�}L��Q4��k�l+;`J�����~�jV�+V�|FZ�,�d2�c�������t�]89t����u/�qm�oc�S��	�]�����m8<0��}�����`4��a����O<����}�c��>���5h�X���Q�������ګ���=b O�#�q�)	`v�����1C��S�Gv��ezA��S����z>��Z/���߷3_˧,% 1��su+Y�H���r����	�S�ػ�y,Ƚ���׊���z�]����XL���' ��1�Q*\�$p��B���BzƐ.��JE�ü.�߹�Y%�L:������cSe�Ԉ�DS+*e
!qd���p���������/*1���B�Y1�_"���N�Q���*ׅ�^�V�+�g�׾�ͤ�i���fw�e2d�:��K�*��Z�#�y�rr��^���<�̀�N��xU��G��%��X�$re�ł�U��0.A'�2��-[�G�d�;5�r�����Wtc\�'%�9��L�Uk��:��ؠgQ�C���VB��Ƨc�2;�y�餙�����I�Zں��3�VV1�S��(J`� �r�Tv$���ľ}�̿%�6���3"�4���C��>.<���֮��G���3K��"�C,Ԉ��V�7���#�S!�>q�?,k�}��x��/ײ
ˡ��,��bp��,��D�.��ܼ���{�X�+7nAYR]�(�\Q	$�r8��eIv��֋�d=}�؜�ϕ� #�c240<ň�e�Ӓ�V(�"N��-�SL9�0�m��/H��h2�yB a%[ �(O��h�)���y'n���صg/���(�xkG3F�F�z�2,[�����x���W�p=y�I�r�uX�q=y�I\s�U��L���xH6� �1�}�v	��C����iwhHyp��X7�/�Z_�r=dn�đ�X98R�E�,;���U��t�~�HT��e�E��,�-�#�ٗ#�z�q%y�g��������寢��[>GH�
NO��W�z�b��w���t�ZvY�W�V���\�@�E3�0g��/��a�#��B%��/,�Χ��ìd��:[P�̠)���}HO���`��(JE	@�y%��s&`;�?�����x�m�Q�k�������q)���q1��n���BaM�q�΍a��!��{ށ7��u�����ێ���Ajr�#���+�� ��_n�Z)�.�~Q�1�Tk���^�h{N��g�~�u @��c��(.��1���\A2�Y��]�~|�ڱ==�i�hW�G���i8ipmk����%6a���X����܁��N�797�7q
�3�� t_UK�e(z^ł�����2RV��"��)��M	C�0_��J�g`�V��8!�$��
�$�y�z�YXG)����T=�Ib<e1�3��AZ�>�үġX�8��u����+[��J�Z\�F�Y��!�Gfi��b��B1��kW`bhT�톗�$gyG���J	x'&Nk�kŚ��8Ǳ�ҋ163����VXL�sE�ZF��m��mp%|��O��@g�lIjB��ڮ������N�\�b[��$m��:k
�	�p����U+q|Pr����/�\�2=�����f���,BM�%��s�S5/�Y���z�VZ�6�Jc����)�⡠S���7Zί��*��K��b��`F��.�vA2��5ƞ+�h8�5��8�K��v�N�!��8�,���s\.��J�)1�,��������b\�Ĉ�*�$��`TȨ3,��4��Lx!S��\V�MT�}Ŋ"$9�\����dٍ�,?2�|�k_�^�t�6�}~?v<�mm}���"��\�lj�=����7����C����p�ո⚪\׬FJ˖�D�;
���.8�c\�⨘-�����>I٘ܰ��{F�A���/)i��9y_�I3�{PK_ڗ�����S�UzR%Vk�j�Of�p���C��+&{" �d��G5cb��[��.�۷���K�Oc��M葌���O��x߇>��.��8�������J$-����U���_}��74a���㲶8�l$�+6�1-���Ĥ�P��B��9q�l�Ь%�{�'5p�3�^�
�H�tZ�8������b�:E��K�ޅ�/Ə~��NW,_�����ڙԌ�/����Ú��۰V��+W-WB!rP�©�T�z�gI���{IEĂ�h��I,f/��}�����&�\F̨PX�b0�b���{��%�m��W]�\�I����r�>}Z_��<*�w����0���/��g��)�@v|V�KV�ȧ���(PHh��W�h>P���'�:�{��99��փ��1=�qq�3Si����)��AoM�Ĭ�Pɷ�h���)�#����z>��тz�g�4'��a����v�+�����y���J�E}���k��Zc}��o��Ί����`�,Uš�����m��CC3��}\am�86tE��m�nO�ƠD��F�B�SIk*�<��B��������_Z�"ۯaoԗ=sVyv�ء{���M�]a�ܗJ�S͍�i���!u�3��$3��|���.�Jhs��#ӵ"`E�Z-��)��5���D��Su,׮CZ"p�F���`4��Z��.��f�Cj�4��k"$M�����#�Z�Mjۻ:�1G���mزa��F)Ū�r8�5��~��$��N�-�T+�$�8-��	�	�1ٌ91�Qɶ9��D`Ȁb�dN+y�E�T��5U�&''���t*��r4�e�MSh�őBKs� ��T��=(����v�|-Z�s�(
� :��@Y�;����>���������O����&N���IFۯh�m�.ǯ��7���"ז���nTn�8� Q5%'f Ց�ݗJ�!e_�\bśɴ�T�M�{�.�����dωY��}�������e����c�'�r_����bÆ���6�o�����O)�륛6anv�]���,�� �p�0#Q�~�#8�J��̱e�ru�=����U�����q�������ơ�G1>9���N1���O=�S��ǻ�������mƢ�p����#ã��JI�`O����hB�ü8�F��_|Ri8�K�Z�0� �|�@F�d\�D9�� .9.�X����S�oP�����q�8���U^p��jA�ɘ�Ke�@�3�i4��1�y糮<�s���.��ֶNmk�-�m����fQ+���~��n����N����٣k�{���e�89^�\�a����Ɔ��'.�����٣N�s��8�GZ.�eX�T�qB��B���H^�xL�
�"z�$����x<����r�5����	ЪC�g_�ocR:g�i�Mu�J�dȝfU��l���o��֙�(��ޕ_pΩ�yO�%�o{�21Qd7U$�p��!�1D͒M��vq�MW��Ν�m�����O~����4���M�Z���+��Y�t	�J�C,��SVŮ���a���z����+�r�y�h���A{�>�+������2��{<��	!��c�=�A�ͣ?� W�ge�W�׎�~;тB�:fk��t�
��ٙ�"Ԓ�OkK��)Yzru5����Ŋ�f�³��^tIr�Q.q<i��ѻ�˺���Y�$�B�d��EW�2dK�-Ҁhk��-��o�%u1���d{ݘ�^.��eS�A{��$ja�^�z,D,�y�YW��%N,���SS�m�(��\eՠ�	�3�!!E]�zBᄒT����aպ8)�)���݋Ӓ�D䳑�<�Yq���ܿ��}���o�_>�i�R����+�r�z�!=tPu��,���%Y�hnI��e�N�� 9 ���Mnff\���"���}��OZ��y�`����{�Bfs�=K�;�w&~v����ԛ܀A�ө�w����}�#!��[^!νM�]ny�ex����>���7m�'?���DK�
�9����$�e�ő1$�\{�^,��^���Y�T�#-)'�n�(�e �:�Q�|�Z��Nu$��n��r���+�r��(�M8yzQK2��[����7�ds�d/i$�&H�bv@Y�R��4�h��ɉY��C	94���ߴ��Q٪	�M��TQB��8��;_8+#ǒ� �YA�|��`F��<����}����ӄ;����.��G��c>�QřԌN�p/-��Q�JNt�R�l� J���`�$�s&�E��}N�5�S��}W�N94=gM�M9��+�go߰��
U�%+���R��D,�A����;b�~yXec�j�:��)6 4O�&�3��X�@���I8E�Q	�L2��b O��]�q�񲗚D�E'�Q��=�kR��S(^ϞV�-��	�hk[�I�_�a��p�k���,���`;��o܆���r�h)�2̐�S1@EǐmK��}�v��{~=�=�7�u�c널��	hu�g���"�]ϔ�6f�>���������"���%���6+�Z5�}�� 7D�R.�UEX������Ipi�hy}�V�3���E�5Gt�cnf��	�7�t��˦��[��3,�`&_В���(²!5��;xrG�p(�����d�Pf_K5|]	L�ϫ��o~~���b���w �D�-�>)���f��|Ϥ~�!�(S�`D��x����-�T�~��g^���x����]{���T�=����Y�jT֩����:��d#<�������������?��Y:rkV�P��e�_�+�ܦ4���!0�m�ͮT�b�X"��[���&'��m^Ai<�	#�����g�n�ژ9���6_��QA�3��������Dj{�S
JI��kРs������PĤ�w���7�O=���o>�-_�|��:5��u�ݑ�4x����	M�~��!9��`h��d'���hE� !%go����K�y�2<��O�w�S�蒍�45���ݻ�W��$>��߸�[��Y-�<�����^oVZCK��hG53���� �`K�ւ���j�|�V�Nʽ�#75���e�F$`�%�;���Y���f+��)*#ג/��
W�E��m�z�|�����-E���ciP�7,g�%hr�Yz9mԠ�i���n��?����9�9ߓr��K(�C����	�
���x`���0Z�`nvZ��K�PG��8�\��/*���4ek��]����<�,�lNE��S-`��)U�Sp(i��Pπ����O�a��f;�?�h�ʂ�mŀq�JTU�W����K�8xA�o��o��9��������%�_�����������v�����R�H����^I��*}�7���!���C��޾}7��MML�yE�܇]#�[08˨;�N�"q<��vl���x��i<������Ϥt:�����*����m�?nK{�������ʎ�K$��w�����i�|{�B�S��A�P����
���,��Į�x�O^���G}��#j����l�S��qh�N������+�drbZ���d@ɖ���5��Zn�67��|֌!�W�l��-W���'��&Kh��y˖K���ߪaխ�n���xb�s����ܪ�i�>��☙Q�3�F��"�[�����;&�7Z�vm�Tǣ̔�sӳ�G��M��I�0�<�4���(vc>S��u��э��)%?��Q�����S_Ɵ}����?�=���/c�C��ݲqV�\�&Y�\v^Q����5�02�	�ֵ?&�1ʪ0�xi{(T�8#鰖�cJӘljQ�!DK[���<���2���������},��O�%k���תJw_�fl�&+k<�?}���>\rٕ:JD^�~�pJ�&&Q��lZ2^��>oQ��4�8ц�[��{���/`Ӻ͒�)�U�gf6���lzR��r+td�u����=J�/GK����F���8���>5�iɾ{��#��>%���c�$%x+ʽ���)��L�O�\c17���nL�oi6U
�]=�pcْ�h�@�ɱB��F�3J�k>�n�bx�­�p�3Bk�W|�|�3�����=vTR������4^u�e���k���*�c�,c�u@�_��ک�]W�]f�DqTMy
�`�u�P.�5rO�`�N�{9��}u�D�kz�D���\�٨��z�dU$V��@(H��JFu�&1p�5���3�􅈬�R�uU6�8l]��U�l��g*��w������=W�Q�]99�z����X���Z���{-��<ry{���@��,���ȉ���>��U��~��u��P���%?�����U�$������VL˰�u��J�� �&8mY{��S��?��/��oǤ$}�b;�T��.r�8̄��'rF��%m�U��Ϩ�
�Ln��=<�"턯,ɳ!.j6����N>-H�7-�"���ݥ�\�C�Ⱦ��!'K��`��҃��l���M���G�@���^/T2��i�\�Q��g&S�I��w���)�G�dXdڲf�yo�U���z��?~�� :�-G1��\5��sF��`����+VB2�2f��h�(-U�Ե��!�k#y^��=�X�1���O�*��<���8[��JZ֨�;I6�}7[u�]�!��d��"+y�K��ʥr�s��Dl��I1����O���V������������'pZ���ƸD�1�B�m�<>>���G��x_�Ȑ*)��3f�vtj��4#8���Y*�h\阫n`�QpP���4[�C�#�[3pT��a��숁&�����Ø�Ia|j	r:��ek�ů|�}+����P9��&&��ա���xDRְ/�r�B���wn�wa>���]�aT�����,��(�%(W����r<rHǫ�$Hb�{z:��c:�Bmv��~�[ߒ~-ړ��y�nlCScFF�%;mA��ױ�!�0�:�D�	S��39	�l	V�L"��Q�,��$�`�QP֒��<CMm- �.�w\��U�",f����9`�%���`	x$���y��>�<��0[��;��K-e��Q��w���?��u��䊛������%8���H@5�K.�L��S�.��3=��S@ܕW_������n�c�]���{2���ƶE8�Ր��HTB��؊���gO����%��1�/𱴜� �܂����
U3��`����D�ƂX���Nb8��U�����q��{��!ׯa��NqU������Ue�N=����O�Q!]�{�a���k���_�fN���J���S����]���bש�Q�[ډXSBG�X�PP[��9}�S�4T�Gr����eO���~Mt�a���g��/x��5���!�l�z�lڀ��59�˱��=���/�V���2�9Z� ���<;��.h�&{����)�����-���IdS���H��,g��>�
��Y����F��>,rs���/��'�=	2b�&UA{v�Qq�sXёD�d��۵��i��D�Tdx�(ɶ�oRæ���HM��";b`p;w����)�M�eP�����{����<���	|�����҈��9�<�c/.�չ�ƙ����o���*�i�j�Y�qj_;�j�N���\^���8��J��g�M���~o��j���?�elY�7��e����ߺ'R8�w��F�Z_���hlU��$�8R� �e��yT#�ꗕ|v1��Y��p�(��s��+�Z���Z(j�X��=5$����LZe���"��PS��B�̽�vɖn�x�x�;�${��ɑӸ�K_�l�A�i��F�����{��|T:r6�B;���>%Q�\�a�NO!/�fl�������j������1��;w��������>���yݿ'� ��ׄ�8Nf�v���t���*��[�+��1���/;>�Y>c�����`q�v%���?B�B7�C�떽�	_|���<���3Q��<�W�]��?y�QT�I��8�4������r����nĕ���dؗ*������q�_��~m��M�g�aEZ��C����7��7o�]�>�t1��m�;�}s9	f��cF����Y�����}i�|��{I�Z+��[�ǳl9?a2���'m��pIak@V���j� �#{h�ICJ9^�]̵]s/��]�sе�Q�����)�s9��8<�.ʞ:���z#�UA{��z��%�ɹA�/�T�@�Â�'~�\�썡����]��j'D�H4����� T|Y^9��$f9m� y�ڵ�J����'��V����89<�=��Ӫ�U�[�J#�}+���cVMG�s����aR����ܜV���7o�H	f~d���̦�+�$ �� V��*��Cwk���i�������6�!lD5W�s/���Ǫ�035+7�]"�>����o�&�y^@2�@<�7���2�?~���\�zn�6�89��ɍ���-�
rcΛ������)�iE[�:zF�
ƶ]���bj��rk�W�4`�=�bցZ,��x�-�fR���Z���9�i@4����%F����@��J�b�xa`��6����-�p�ś�j��ش�%ޢ����){�8��kDX��h��:I��!���,��s7��ٛ�x3��m�
�lAi]倒���n��a�u������ Wj�u^��^%�)98u�4���v9XOb�Ġ���|�F�Oҝ�ڑ^�?�����E,�z��E ��Yg�s%�Q~\qv�����d�m�l�lU��'�|J�Q�c���M�E���h�C�&%�
#Jv�\F23%a������%ٰ�3�w�W�{������R�T�j/�E���߳Z�O�q~��iy��LF���t5(�L6��_�Pc�r#�ø��'% �GN����)N�%Ӳ1�?������hr���VV�M����~��+��g�fb]ص�c�r��W*Bz�2������6-����|g���R�9��.>���r8���s>�W��T=�2�v��g�Y���nKq
����:Gn�Q���Fp�ԑ�$/���מ��;�ť{��$���Y	�EM�j��u�r�I��>��D�N�ș�.+mV�U�D< �S9�����0�p[׭U��n~%Mqe��ţ5.�?��YeW���1���}6��5���af�����%@�Z�����6�'rx�Z�����Cׇ�����8��%��e�/���Q��s(eRJ��bٔ��Dy�q��(6��Q,�敾�(l�>̈�C4��3���x�0f�3�6uh��JPq
�lAgI���F
�5e%K�K�
P4��	�xc�?=ji^O��/U6��ԟ/�olJ���V)�7����^�)}1Y
&��G]��5����(L������ރ��%Eos���>;�A������F$C/��$������x2���,�RǢLR���7?�:���&rq���?�Df���+���o�J 6>9��h̺׋cPA�̂΢F�	WҳZݩ8�=���$��R�kF����f}�ge�U˫컉3��Kq�-�a��U8rp/���;1;=����+תl�G?��ZU���՘d��|��{06�Qn�2�xX�L���b/ t����z�56�3z�"y���>H������z���3Aru�d��	,E�Ƽ~���;.�W(��̲�7�O6!"�2/�f����<?�՝���k���q�B���
�(Y!�AαCw�Q�=95��t��sGC�SZ����R��ھn3PRt�a��k A۬��H;1�hy�y��y���Tu�^�U����)�__6��z�5�x��Z�裶���� ����/vK8v��p7��F���ҸE���2�k��ү���9v́W��wAo�ίi��h�ӫ8��a�޽N���A�n*GF�\FC'FP�{>w�$rs3X'�U���7�۴ڂAGq0�	�tOLMI�T���`U�+��JWY�Q���HQt�:ђ/���e���AO�Ф+�C]�Ⴅ~U���! �t�S�Kv�l����� ��U�$���A����U%)n�R)ɞ$��X�\���Ĕ���B��/	�9�lAѶ�Wo��̜�SڑBl�It�w
Z�uܐ⊎����Tj��f.��x�c2e�ZZN�<�������A5Ʃ0�z�D�,����x�ƸWMo��r^@`�}R֐l�V�Aӿ��z ����|�YX��
5�d(�%�g�P��JP�5	!�Ү����+���
�ь��9�Z�Ca� /sd��YLP?���ݭ�:6eb����6���/�Ґh�-�U���ΥL��2,�˺E�lE˯<dV���({��3�p&�qj��:Fy���qt�6�1j���kW����s�Cxٵ��~(��[.��3���v�rX�`㦋��Շ'��G��`4��Fdd��q-�Qx��tݳ���g�'4ш���2�g��U�;�\�ʐ��tŽ�b��5؄��h0�꩞���A�9�Ԏ�*�'_UF�*�k�E��S��n��u+q���dP�6�e�:C�����ɺR3+�i	�Jy���n�2:t�GĨ���ՉT��M�Z�C�w�{�+!���OW+f[~���kdֺ�!��mѷ��1��<g����<� (b��Σ��:S����y���T^;KK�g�J�E�R�;�������[n�+�꿯�j,��������{�g>�:�2rU��H>f����:�[��*u�䐙=�t�\�4A�e0͒�1�*�m����q��Mb���8>8��7byS'FFFPv�b#He�b��*��삜2򁉜F
�"[�(E7��%Ay,n1K�Y[�zՎ$� >˥-�����e/��� �U3[�&t�Z�kF��M���(ʱ$S��;J%#���0cJ-�h"�{@�H��ؕ$KZ�e�w	�9w.OF��pU���O{���"Rs|&���	Ee��5�%�Y�%���W�!q��2豢yڔ��z��uY^vnim��l��[��WT�gy���F��F:���� F	M�U&c��=8��Xڷv*&*�a������P�Q�p~ޙ�q��@ROsgښ����$&f3���Zs��R�U�E־C' ����lF��cz���o�<zG�ZR�㜰ikؚ����d�S���Q#��P@�Fec�94� Gއ�
_�{�����V����"��2�f͢:��$�(j�&'�c�r�Hޱ�p�UW��˷!��K�>�e���nLNL�O��Oзq��B[�J8��*��đ�AC��\+;uz�o����_^S�{��U��/�� 8�}χZ�T�޼���{eҗ2���\�,��k/��s���9��
�4�#�hkƛ�WQy�+�A�=��k���oޅ�����?�y{≉1�t�����k�+�߂������1<>+{�x�bB��%;:��ߕ����5X�8)Hb�{��t����N�7l�2���R?k��rPշA�U^�O�cR��z�o��������,ZK_tI��R��������4�W��u{R�S5�;���֬���)4{J�����imiT��\9��(�Q"!�B�B����JnQ�/E�[�bW[/&��50��C�A���ک ��� ����W)�+74�+���r���f�e�`\O��Tc�܅��]���`�Q_
4��ԣ�( ���,<,�dt�'�y1�,��թ��cl�|�B�"�Y������:&�����ʆ��;�ԢFU�f��77�f�u,eE�zi��u�Q��( ��Ic]]r����%��=7������^��Y�2�ׯ�GD�d�U�!#�9�r�lF�'1�Z.�-p�wjV����嫔����[�����R(*hP'D[k\�t�0z���d���|�ߵk�]�Q����e,>G�Xֽ�k�O�]���$����σ��Ba	��(���r��}|��i �k^�D��������9t����EqD���xz�N�E�\s[SD��C>��?�T�+����~
�h�?��(��($H
�J��
�q�ed��X\/f}CX��X����Ƣj稶[��a�i�u9��S�OH��'i�:��S������ש+o�TyV>�6����z.�+��L�W_�j�p�:=L�:�sp3��]��D^�Qc�W��]K������d�	��������0�T	ڂG��9���ީ��҇]W�6�zֵ��zW�n2g�[��Dp�`Xh���cl�=;>�T*kub�]��t��q �[�r�����U[wSɱ���}	�n$��jX懋V�u��gV��9t����j*����W���}￴��Ul-�2�
z��=b �H��ULF ���k& ���hk�./ϗ�T�|{8�x"���Q��Z�K�e�G�4с<�$LV����ל'/>F^�\0d5�4���	Ș8�v�=�� �^���*J���F�s�9t�rjg�<^|s�����uBHH�H�dډ8��g���!5F� ��R�G�������8E�U�¬���#�VL����5�3@�@$�cY
��8��������5�s�^"|Qwen-�^<�>�m}V�$Bׇ�Z5d2����XV�a�{���K>�Mo�f�a`b$P]E�<�J%�PQ��ʎ���ӉD���yA2�)�d���IN�	p���J.j��Tͬ��Og�^(��9t�α9�)��:t�-Y�Ks��WzTy�H�Ho��̩�/*BY��9W�Y��W�(��+�����hu�e]X[��\������#�>6��{�����$���F�'�N��]{��b͝b����r�J���H�$�>�8�o�u�B�9�3��m�w���`�|Yi���<�U�X���@�����;u;�����<����浅�@�tAQ�{y߄Y�|�+�ȑ�kanR�8�����zD��㓣��jS����A�ٟ��>�S�M������7����;1:;���d�e445IvUP��zn_p�vFk���ώ��	 }��0G�g-�#~Z�f�_����xTm=y�� ����q���؋6ª�R��E�k׮���n*B�N���<%w˟�p�-����J/���|u�y���j�~�/5+\�V�����m�H�����W��1s&s�1�LMh%�ϥ�N8��i�'�l둿g�^P{U֪��F�WV��k�����B��f�\$�y�H뭇�Y^�B%����cZ�l���	�����C��>���rᖏ�v��z��6循npMΞji�
*5d�����XB6ǘ�Y��E��=�[�h�F�E�mnk�tFg��!72�D���"�M���U��^�I�D=x����~�do�D��dy^�R>Q�pk�z5֢.<��Ҷa������j�!�Tu���m%�imm㕩r��>����iH���qcsTDY�yw�H�(Hd����D���}�4���܌dU���*ɉ���PR���e/��q��UNSE9��g�5Պ�b �fݴ�Rg���6ص,�ր�\&��X,��*yq���ZG�1�&?m�g���)h�2ƛ}�`��}j��ݬD�i'������S���P�Q������!q^�^~%6l܈c�=�\�n������M�S CçĨti��2�U4�Q�Ǹ�cR���ln�B6����4�±��`�����z}^5^^ۃ<�ӓS5f,�[X̜h�BIs��������x�����Y,�[uc�D����UG�>4�Yx��g3��J��r�2'�e�Zlٺ�+z153�����O��K�������i=���61�4�6��n#�Te�;���u���.Җ֚��:|gX��ug*� ���+V����gI�D�d����V��hJ����N�p)�k`q���L�;�z*%'��ꉳq���i����a��G՜��՝�����-/3��Z�k�x��{^���Yz�EjD���ڴ��o����d-�Y\�k;9�R-q�|)����kpH�`،J�=;�����@ѫyj{�=hlhCS�	�ӳ��V �4�%̉�k5��{�|?�|!�1VF4y��j�����A����P������U�pT:�k@L�
��Iȴ�jk pA9t�]3��t�X����e��v��rr��w�1�������s��Q��W��7�9"��7Oz�%k���ٖ'�`pc�.V/S���V5�������*�Pn�n��La�e(�@ld<�,k�f�'���r""co��g��7��r��/�t�̌��w�w�}�!j�FQߙ:󣴟1��9U�`���
���|"r�M�������6��X̫�$lW3ߧ�z�������f��L�$�ᰮ�a,���=N��2�Y�����zYp�T*E�@��	1!��Up��lmI-bzAS��^����|}� ©�n&d*���4�n)��U��qSKGj?�!3�L1/�ǐo	�h�{v�["�f�i����t�xt�a` o�met}\U� �ɨ�����C�#�����`��d���E4�j����'&r��1�dO�m'�������ſ�)��3U�����LϤ���ͯk�ّ���oˏ��� �[]�����ŗ�ht��6	2��y�����d�9~���Z{���o ���:q���È ���P�D��{�w�4V��!��9 ��+Y����7�uB��8�Y$��WƜ���^�i[�HQ���)Re���x��[�F��zΪH���k������*s�Y�6Z�o���Q�JuEZ�5��t4�ڵU�kv��d��i_�g3�(��1��5�?��5U���:��Ϡ���'2��A�v�������!9��E�&L����:t_z�>��D�t�&`'�w#`�sP�����D�`�ʜ3�a	�g[?v���~D�(�Ͽ��&t
X��"�0�`����O� =��:��!�>4:��@j����ڀ���?e$d!�o�����!����)�1�ġ��j��|$Jv�pg�D@`�8fŊ�<��3d���EVˉ�wl>A���͠Kp 7�����p��5��k6v,��%�ME��H#Y���3D}�;ӏ��RZ��w��Rc�5athS��#��b�QH�]��([�mh�	�1��"4O�N!F��jj�2i�fggd��r ���v2cZo�s���:z�'I�M�H�׎z�C')�(D�z��Sג΄�+рDE�O'.����sl��5���@���{���i,AԀ6#�7z�s�{���d��Ӹ�}Aل5�;P�6��2�LT��Пy�F%=���ڥ�%�l̀:{\zs���ؙ��z"U�(\5X���F=	G�F�)3�r��^l���K�}��R���_���w��xᢼzmY�<Kv6��Uq����dw�*����k���f�q �x@�2
,��I1j����}���7,c`@����'��m{0�ɸ��|��kS�7`QB�岎��!8�����٠6E�>��>�OFұ���q�K �X���c��>���Vj�k�f�f����ٴ�_�x��g���(�:��81�\��?��?�������m=����ɩ3w������I,;&w����c��_;?b�hi����Y1}h��%Dv��$L$�W�Nf��{zM�� ����{���uG��  ��No}�]K�\j�m���r�ͦ�;�^ϔ�댷�ᢹ�+a�lL�)�2�9����;.*��У�|?��q��A�Q�	'^suFo�,+��(0��X:��S�
,)��#��	d	�ECs���~
�)C��T�tiI)�z	پ rf�uz�!�]�`�B�A�1>#��!0��7�Aw���4飃��������U9�K%�j�6S���Y_r&��y�jc��ǡ E��I/��|�!�bl�B�z���Lz��N� ��Gz�X:`t�L2�)�&RuM�8]���!. � �.�I1�g�kw�2�p��/Ms�IR��객�]���s��>�$��#T��Q��I��lm(M,,.IJ�ӄ �;w�%A��K��M*ҭ�u.6�f�AH�̀DcKhBR��1 �BQ����F��j�0����6.�?��X���̍:F���s�Bw2�|�LD�n��u�bT)�#��r�Шivz#3�Zυ�Mµ��0��A"|:Y��^mSȳ����t�;rL��7���T����%���NԸ�����'�}��M�K�(J��d��]q�b�rɚ��U�fD���A �\���f����H�03#���v��dD����Q?��bRTX�	���q��ǧQRc�A3p2�ڄKdA�#D³�(n�˵�]����I`�R ���_���ujʑV͕��)3r��5y��r��+���$�%���+��/M���L�ȓO=-՚��|��T��ړR{�y3P��'��w�?��d7^����۶DY������c̀�̣=�4�#�5bgJ����m_�k�� 2�~ ��	d��2�0�؞	fDn���_ ���ޏ�C�>��1֔ܴD�8�#�&(�������؟���C�>�����a����Āe�s<�+��l@��$i �a��D ��ed
���l`%�e�Ũ�@ȅi1���]PB�T��lk�K����}.,�X��:܋AB�i�}t9�}̀~c7!�]b�w��<�PQA,�Υ�/3S���v�Y��g��&��'z��m��::(]�[����G 0`AA�O�k� ���GȾe�b
B���PeUp�1f�b@�~$�<jLӿ���6gZ=pԴ�*'�ҁ���Y�ͧ{<+k�W�б�6j�� ylK5i��>��x�=�iD������������α��eggG��\c;=]&��é)��M�lfkmM�Kc��gȤ�0���#�<1-*3�yr!W���@p����؈�o�ރt�nF7!���|[��G�dO} i��бz2�8������u\��ƒ�$�	�L���#)a���fL�ԢUh���T����e��a�r�|���I#ǌd4�}�dژ���b�,k��\^ߑ˫ۦ�&W��=&�>�����}��D�ԜL�ΰ޿��FY�"BZ�\�i�ʩ���H'��\�r 3#!B���-��D� &Te�l�ꑂ'���ܨ?�W����i���o/W`�X�����yX	̚�:Mb���|�ԃYCօ���`��Ey�[��  ��IDAT_�{�]ff�U���ȩ;�ĉS�lt$�r��>�9��/eckO^�xE^|uE�_.]���O*�	kH:��U{�����5*��uB}��f� �f֌�u�쁨��>}�O��B-�]_D�)��QhH>#�� ��N]�5CKh�ۑ�:��9]�3 >�]1���2��������l^��f����l�3N�D{���Ε��ۯ��n�y���x)� 7�/9'��+꫘�O��~@��Z��a�'p@UV�ы�~�0��ɤ�	�#�  @�c������{*/�J"�FV��R�o3�E���]�\P2�?�0ُ}�񈀦�Y�Ө��rS���/V
+�a������KK�W��H}Cz`��ƻ�T4��t�Rܔ���?U�o�J��T��kSKߥ�&af�F�� i
�:�zkÎ:~�d0zO#�x�`HPHV��Μ�֫�w�����ԩ\:ͩ>�$�rMY�/K����U9s�y�WT�/q��U���)w�f#�Q7M2L��R�[�.`l�^��¼�+%���  	�^,A�$�F��/�ߛk˜5WGc�2�ٕ\�?���f_.�鉙S��+��e?���@R�!��Z�v�[�0��6����H�iv��4F�0h]	�����h�؉c��F=_N��!�IO7�^�G�R���ݜF<#*D\G���mY�"��K�(J�䌸��ݶ����s)����4���6[�5�FZ~w��������*5�1U��f�0����I+��j�a(*�x��s�L`��0`��_45ڮ)`�PH�_�XG����8Uۊe"!So��A�w�)w���3Qe�G��2&R�z� "���q�� ��l�x�|�IL��3��3Ǘ���F}O��t���]u�w:"���ٖ�+�?mn^���e����?���v�!ϿrQ��:G���;�p`��I7l��׾��)�؝������,
0��a�-��0�x�s��I�sP�-�P�A��e�{��<t�����W��� ����O���``#쨃�^^����%���9�M�*��Ӄ r��s~��5�d�P�5��G��zs�E���x�?q�L�Ƙ�a.aJ�=�p�A �W�L��2�9���Z�$W����I|f?��M�]L7�z�C�1�@1�����u�F�!@�ݵ���0B�N7JSȍ�a�
�ު�4
L��Y�3���︍���O<-�ʬn\Sb�Cb��D�|� �{��[� `�:�h2WMlh`h[�J�y�z}��W�{27[��'��8�g�;/�rFMcI�SI����s����$P��4�Ԁ��}H��:*_��/ʥ+k�wiU��_ֵ8�Q�'��{¾R�s��:� 
��1�\���*�X�N'c�<:���MD��Tf�FQ��J���,kׯ����F��AS�/�d����J��#-�z��O�V�$����Uˬ�Xޤ45R/OͲ��[\�K��O�|��T��<�:�Cy��D�����/���M��W��㟰n�'�JFJQ=�>���n�dsyN�C�H9\&����^T���>��;e��%����#��'�D�*�RqF��H;5IUX�nm��Ӫ`���0�p��U�F��J��v�q��"EB�$&Áa-X���Xv8`Ȭ����f��܈8���1�T��%��L&�X�(Kpԣ�3^�a��+mSX�1��^�6�5EJLi#�\�A
�;u��4�1IO�K��Ɠ/��\7�+�G��T��R*ecs���s3��KW)[Wk9v�G�+s2�P&������Y�{��n������(p���	,���t�� 
��K沒)��gӹ�cӲ��5���g�7�×�c]G�M*z�������)�A�k{�����=л��ˈ��@�݋R�ߍ#�9�>����t�}V6*�z��B��  V�:U�C�.�%��:�z�u�'Q6�1V�r̰�16q)���*L8��SD��	��}��}�w��j�s�]0�=s͆	Ή0���k��|V(��)�߄��bn��G���ѹ��!
��F�阜<qD~���ВHmOT:��Iefe2"9�>� y��q�ư��YW1Y9��<�愑L�p���NS��(n�e��}|����)[�"���?��+M���)�1�C�6�>�B�Dz���Q�t���\]�[��"���\�_���L����)9{򴜿pY������0�0m^� V�D؆1���z�i���63;E$3��j(.]��H���DN����h@#��'��uY�xA=���Kj��r��y��K�<��2bZ]b�ȴ��#���Y��el������ ��$��P=g�MSق#�,�F�zuX4�_.��<���|�Cr���i4��o�+W�-_��פ8�Q%j2H�wP�w�l%��L�c�\�5�8-i�>�ӧOJ]����N9}��V���G�W/^&_A*���@ߛ,���y���Kț����l�vX'�� ��O�-�N��w��^�/��Ir�&�UBf���9�;u�]3�i�a1Y�g���Z�Z1|�1� |?@g� 晡7������%8JD�u�)I3��A&�Ƅ*�aO��D�N3�2�:�����L[@�#d~������#�D#t2)i�]��,����TT�}���:�~*/�w��M��&R(M�^����rH�H�X'���Q,��K@�T��� � z<��o�� �Z�D�+���E� H:&�]>_�^���n*��#�-��[&!�VSz�@����tܹ�K"��s�[�����o��}������\�r]����H>+�uA웎��"����G
�'l!&��>��F�`�{���L�ˁ�ʥ!�á��k4�ч��4� ���� t�`���%X~$)V2e���΁��Q�@u�z�2��S�N��ȣ�r�)� ��;��Ħ��{�ClC���l>Y��fa��Q�m�����b�z}���ӷH0@M:1�0��K@\_���œR."�����G.\\6F�3^�ı��1�a���9A͖�)����C=6��ĵ���!�\�ㅚ��@DB@�(��JY���r�=��}K�"x�A��?���/���^�O`����Cd[��E��#�����C�ӳ���Ү���Ԣ|��Rɗ���p�5�a/0s���({fz"�h�@�{��˚���=�F�T�ht���{�\���iĸ+U��NU���mJL���JZF����^���vIv��נR�G�� �>[�a����Q.�k�mO~��d��5�-�Z�Ψ7�Sc��$E5���#��9
S��:�F��������������u4T&�'�,�VC��&4҅{�L�<�U�tE��j�3�1e��b,��`V.2�\߸.�uV�ſ�i)��@	8�����%��]�԰d$+�SѕT~�QU<����-�2�S��zҧQ�>��m��"i��+V۠�p��t^�Ty�"���5�{] ��	��o93,(7 +���� ��M����	���u�&j��i �G�@,-�#g�Ր�G���?&@qj����$���(��z�h�ܮ�]�,_�c'����*>r%C�䑤P��������ӯF�KpҠg��ǏOsx�\�QQ� _6�:!Em�DyK���쒲���0 �T�S��q'��L����$0����������*�8�$��������L6">Ɛ#%�UkS��b�T�[��'f��䩋�seS*������Tf�5��,�p��xN^%\Gd�\ut��;���~J��}o�������?��� ��@�Q�9��5�$������1�kcx|����,�>�4:�����4Em���8�4ԨI�3��� ��L*�"�%�_�^���3 !����w8��9�|��3����Sߏ9�� �:Ѓ~GfTנ<���2g���Pu��=}��zu�'RYëOG*a��Bb�hߋ��k2<n���������E̖@�: #�9@��T����j� ��
���0#��P��bY�����c���o9#��{�䷟Q�7����G�rʁs±�h9��8&�w�ߔ��FC�'�!-l�� �z=v?3���,k��v,5:���dґ�_�����j@E��IQ���ƕuG�� C��B�#�	#�Ȫ�ۤ�y��s��'���#��c/��NC7�#[��;�H<�	�=bz��q��O��� �E�/dM�y�!;�;�`RRBO�^�Ç�g��K����˨��ޓ[5Z���y�p�EY~��T�q�m�Aw�2S,I�Z��mHQ���d�h��"�So�6�kU�%�,����;^O>��{���c�Y��W�;�x?̳/��X�,/\ؒ��>_1@:8*�TR�\�.���ߗ�����׮ɋ/^��:�W��ĉ�����U�Ɔ,m@������:[ ��8��=�qL�3�cU/ȸ�F��IFث�Mu܊����W��KKFU��Ϫqo�@�snf^n={Z֮^b�R�S�ӏ�C��^�ҫT*�a�����?6t��L�ivը��~ ��m�\��Ccl]w�����5�+����&%-�gubԀf�xhı=(2U����4�u)�BnﮱV�[[���9u�L�$��wV���ls��C�"i�>[t`�z���/�%��3���A��|��G-5��H�9��7�NsW|�C*B��̤ԉl�!� �{}5$i��Y����Q���/A�&	,݄�0�\�B�=ᙀ��?n�y��85��E�%@wҹꈲN=�Q������46l}��8Ϋ��nw�l��lt�ah���eoĞz�@7E< .�L�:�)�|Nv6��Mw}X�/�`@No����dCY蘡F��F/�ue���]��HvJ�EΠ��rL,�[��t1�*�I�����D4�V�N֜�"��@7�����ZA_�޻�`H�i�t �iC�δ����@<*66C2�Y�h5����8i4PMKF�tS�0�c��F�����!2p:���l�')Y\� ��Y�B&��T�8������5���B6L��l�}�ؑu�����O7�"n*�^`Fi��8����h�B�5�VO?�a$�����¹�Da/_[���CݘԲ�,�s�I=بL�!Y�f!b�L\#�xxT�ِ��x�N���c�w�(>��:
��4���������_���F�]��Ԅ��`��v�d`	7@��[�������3_�p��}������)�J�Qc�Q{<���6�9��E�0�H�

��]�4T)��_H=������ʔF;9�h���n^�i]�C�G�*�em�L�
���q���~J��oPH��<u�8��0��د]�l;Ƭ�ƙz5k��8T1���r��	y��w�����r��a�N��U����ʵͺ\��;��L�c�i5zz��֣Oʺ:|��*�BI�mZ�ǎ�\�P�Z��H��dB:��`G���w�5����!#t2{i$�P����lUa��Fo|�C*;�A���Á*W=��E����(�����ǜf(荍)�����=UJ����1+�%�2����Q;�GTf��@?���f�{�o�B"��kO�S�hY8�euN�SY�8X*.��O�����m���$�41T���F�qC��ړ��
>���tc|c�*ɧU�' ��eo��U��p��;�H~Sҵ��E^OQy��@�����DjTL)�6"}P�]5�I���ڨC`XZ�D18#�>�Lt�S�jh4�?��O�ƺ���u��aG{#K������ WHgi@'�̚1Fl�4�E6���I0i.�e��=P�Wg�?������]]��K�	�LZ��H�Y�A4r��#�����O���	��=�!�$��d2�RJF�L)��A*����?��s�ַ�/���Ge��9Iʐ�GA�{%��^O�{D6�q�N"�Z,��k#u�F�0�ͽm���|V�"b�fGRj���=I��8x$A���' �X�ڤ�ƾD)	�Vh3��&���r&ɨ���ڍ��:�� ��F����UNB*`7R���%�3	�b�u���P&W��Dt7��L�@��4(��E���� Ȋk� sw�0;l�m��l����?3A,�4�A��O���ʠg����0R�;aZ#4�l��?Mi� �t6Z�<��E�tC'Ab����ܤἶ�����E*X��|U~�;�!T�9�6�EHy��t�{��EYѫd�'ƈugp��D��e���L����T����s�h�d8�.��p�vo:Bu��A��B�/���P�z��C��������d�y9��$Nҕ��e�K��Dpã왬�j�U�duS�Q�ט����7\J}�ݔ��o�uu��PJ�7�zoU&�s����NA��&��F}p:��F�������� ���Up���ɳiA�'��Vr��s$��u���Ҳ:tD._�,�;{r�{��ڡ���V]�Ԭ����,��=���z<�%������4W�Fƙ�tZ��)p4���V(�R�D؂@g����rE�����徻�cG��׾����]�tqJ"�ʅ��gt2.W.�"G/h�֗��Qgc[��6��ظ���c��q��h�*�4A�.-�˚+��l�nW�M�L�Ө���52���E�;�/_�6te��R��ǔ����%��3����9�Ω���f��Q���JN��Q��Ag�i}dvW/��Q�Ʊ�~V�uҐ�4�MN�::;K����s��][�M����^O�è�er�KPi�f^��q��fK���=0̉�^���Cƈ�k���Q�����H�,H\eiΔcd�����C�>N��E»f�:c��j����y][%��ᾓ���
)����N����цb�:f���m0H�R�=Q٘�v�4��^\*3+7�O��&i�m���P��Sg�#�j�ݺ��oR��3�� `��5Bv���ct��(�j>3���\���e0-b��G���b:2�c����,J#E���i���+�AS�e�����-�Xg��K1��*@?j@�9��k��Ә*�� �:�XNp�����&�ð$�l 2f�]�dR�P��?|�5�}
Gy����5�6?=E�D�U�9�e��Cul�>��s�25��!2
�I����=@B��z���VE��	I{ o��T�5�6D_a�@�F�怈�H�H"f�6��HX�i�{B��4f"��Ģ�!zd73WQe$l	B��k�ݝ0���y��I�?}*N��	,r ����^q���� 0�MH�e3)�.��r��
^�c� .2�ɘ�`�2"�Q�Pp��fy���-�z�#���h[q���iٮoɸ�
)�Jb�!ҟ�'�m�F	���"2XD�vO�XJYW�j{�/|Aצ���95��Ր_�tA.�?�5�����ʞ�;�d_y�%�z��<�8!G���!:�JiC3k�=����{�T����*��� ��G��긨�V�w��c%9��4��GO�:?�V���;����.OL�36��3Tb뒣	�
����(����1�hZ�ƌ��+��Ǟ���=����o�F#�E���?���͟�t�:{�O�X��D�_x�%���4�5��ˆF5-u�p}s3�fn�?R����ٔI/�q�S��$�z|8��Bh7!� x��k�12�=0d<��1��g��e��K{���X.�3�u%�
/P�5q�� �5����:��=#��hFߚzl�k���C#����&�6��F~�q[F����!	�F��$�/²Z�0�r"zM`8���M��i�8��E�N5{�ͱ�qË�b� �5B����M�� Rܨ��@�۵5�\M�6��Ų����~��Re�F{�A�����t鰅Q(���W)�
�g����ݖ��>a��%��e����ʩN�^�7�;����i�G]�ބ���Ef�+�^C\u�8�C7R��qF�|�����3��:�D���+�umOڤN�6f���$2،�*Sވ��ޙV�D�Ρ��wd�q�k&'�G�@G�c��)ؓ�1��<q:зcC�R�mʜ:���,�5vUvיS�kң�H�yG���N:5i�~X�o��1iM-,v�!J
���&���uLdu��E��Ĺ��6�to.����g�W�i׶���9=���?ڝ�^��	��Ub�\�1�I7䧄�i�L"���T�Rk�esk�(�Fz��6��Q���P�ҏ�E|H򁉙��볛�ΙG�'��@�j�UR#� Fx��3��b�4��B0��)��5�J΂� ��n��Pi�!)��|U�j�*Sj�䨮���[�1�-�ia�� �2��B\_S�)2�.�f�;�L8�`<0�˗���[�������:Ou9qdANh�9�dwg�Be��*6�5� 9�|�$����Cr��1���{.���fԛF����d����u;}9��7K�7��k{�pxI:���:�N�|ٸ��r67#͚n�n�5�N���.��V�}�.4�	�)9��	B��Q};���A"��[$��DF�^[S�%-���Ajd�ȫ��˺F�KǊO�K ��^M����et���,��d��v2jˡ�ò����:�b<�y�ߝh
*���MF�4�A;�O��M�<�J��@^�0![���^_>��l�_%��X��l��ft�]��Ⳬ��T:���AGf�z���h�X�urFj�rᤪS�R�If�c�Nn��YFv,`:���CV��dql��>
� ���њ�>���yL�{Ɲ ���s�qv$b�t@-�4�u'j̆*R'���%@�:V�ᥤ��&��#3,���̠d�1�*�����k�ҩ�խE 3��Q�>�\2��y�bu�P��	�K���6[R��������0�Q�RխVW�_"��G�
`:����J�����"����k�\0�-��:Z6N"Έ�sE�0�� H�� �K']������,#a�D�"J0t~�s����
q�q��? �42���l��ܒ��!7L�Î�e��M�Đ�s�o'���M�z<�[�:2!�0"�C��]�g�����F�q�x����U\��z�l՚�Y�gC�"pX��5�&��X�Ȏ�.���L�>��|���ʠ���޽�7l�D��c��"�\Iz�0@�8@`F���F�%ӳSf3,�N�{���#�W�����ג[N/��̂\��%���H�W��U�� ���)p]�tI�6�j�gę����m
I#�!�J#: �A�Y�.�b;a-���-U�Mɨ0g�	�PՋ�K�M�'�G�D\�����E �r���.�K2�!5�$�U��)^-=!��Hq"l�P���M�4wt|���'��>�Q*��::�RV.��F��t|������r����a*z���(Sv>4��-2J;v��loo�9��!qn�������g�=�y��r�Yyꩧdf��rO�.I[��j_���e�Tic�����`I$�/r�YZ�2qD� :ZO�
m��af܇��?�"fd(L������7P�H��:5�L�ཱུ�-U��]��EY(��O�0���+R�8�0�ıw�2�P�hb[�w�6���|D�R.�[�L�õi�T9g�R�^0����b�س�(_���>��:�萳��m�033c�~�RÈ�b0��8|?�;��YL�{�V�!��?6����?J�N����:��U�ߐ}�����|[*�69í>WC�"$l�~�=.��4��@/~.����X�p�l�CK\1_�)u��h\0�#�+SEF���7a���cT�#��8�]���%[����z@F˥J���e��(r�c�WW�G����2��Fgi�$�v�-X�,��) �!�{��Q:È�s�$�uc�X=� ��5�Nl>�[LE���q�x�}�M=�+2	h���R}9�O�M����2���(S�:�E25�>,��XH�ۤ�L�lq������3�u_��y��Ŧ�ù��h��IMԹ���0#=O�-2ߴ�DI̩��܁N�=]��r�2�b���5֩�U��V�ۏ�@�nݑ:��P}��:���6(��s���t�7 �����y��Q;�k��7�A��������#0��g������D]�RE�T���G	�K�!�V��H��P�qSW�>$?��Zff���?��<��_Gg���r�ߓ��U�&����n��8u��|�	�h3�
��v�����Q�����r��	�sr���a<��e��V�ɨm��Qk�RT�;��R頶竁tS�4�Y݈j�@�	��*�ZM�`.%�rVϭ�"nӷ=�\\���� �8>R��L$Έ��8�i_�r�6v�]]��'[Uy��G���ޠ�J�
�iD;� S�`���U����� �3�~�Q_����#[3����a����˓��}��4ꟕյm�M�Ta�F�^��N4�	b�!�����ē*#��Be��JDg@H�Q$H�3�26��ov(����4b�2���P�/�2��-��Q��DN����g)�V}O*Ŵ�չ����ײr�%*���U���Q2�I��Ge],1(��ޮ���<=��G�~��D�5�3sgt�j�cB=`4���5�f��j��H�88��B���w�M`S��`��<��ఝ�-kdh�]�9Y}�0:��8����c�S �q�=q���n0�����0���ؑ��Lk�D6P�H_����粥��j+vl�I�z,�TtM�հ��{��f^�c�5�q6�n�08�(	�����d84���aH�������I�Cnp��J:��	Q�B�-K�\����� �r<=D�d���r�l�} �h$�hĢ��^y��L�A0�P�j�LJe"��q�,7`�!�4��VW��/<7���"���m��&��:VW��a�KbGG���te�CaZ������!�ͽ���QQ�f�O�uU1��X�}�������-��	F�-�C���F]	�t֌�ǑmA�v�*w�y�r��۫�T��������{�vQ?Gf����5QK�X���E��'MV� ���ܝ��5������o:����1�!�5 5�J��T�!;�P��( ��=�qZk3���G��\�P�A¤�����SC�����5��G�G��4뛒�����i��T(:�\��G�I��6��X{o$��/p��U2H1t5���3�:�\.���i��ڄ��fnN�)����ьq1�*R�xA8a(r���lnk��Q�VK�cK�.��YcX�aWsʹ��I��c:��n�eq*�����9@�8�.n.�fe�-���e�ޕ�?��5�f�\����
��n��G1�1b����m����e���u�����g������F������k����`ڟ�Q��C4�]J���[�K-I��������M������j�/�o������[J\*?�(�Hȳ�;>SϠpȑd��%�
|䙩x�����v� Y5���Se���}ղ�xA.��@ ���|��mm��2ylooq��3 ����� ��3=�`��3-l"��g�ǟ�g�n���ڥ4Z�tڌ�&i���
��X�a�x��� �^8G�P���<�C,�Y?37�]�l
΋�u�����g���:ɤ�_!.�n_��
�@���X���=�j�PC߭��X琙ͭ��@8��`v~��G?9j�p���7�H���^���a?�9(�ZpU}]�<Z\5���ga`|�#]��0���p�8܇k��	��fB�
�+wZ�#*DmE�lc/�{��y��429	��F
	�%z�rD�榛��>K���?��{~�٠>���-��w��N9#W�]6�����{F]��#'O���-��rY� �-����`��<���y/8���:e&d�Q���:ww�ȿ��d�~�=�5.���%����͍��h&���U}&5}��1�>��5o��� a���ܳж�jRg��L1�z�G�{|eu=��t{��7QǢU����/�,2�yu�Ǿk����}O�g9_���T���@�b��*I��5�(�Em �lx�Yt�1ӎ����ް���3+~���̚��,9n*�n٩��h�p`�X0�~��Y� h&���;��Lpv<#�0��	���#�5�2Nޗ�����ʑ�q��Q�d���*�J!-�D�`((D�@@�Q;/I��
O�?��Bꎆ\�>�Q��@�-�O��oR�z����C�P'���.R9�μ��x��iX ��*���;����_{\6v�ҡY��2��8���v��I`���K/:0s��,LƆ��}�qß�	�[�y�μ](ȡ���E�&��C�P:�=y��o�ߔR1��7Z���f�p�s�ؤ�W_���h�����������R?w��l1��P* )Rt�z�<e�JܫU���0���M}Bn��#G�Q`X�)����axH��1,n��8�Q��m� R��aM8����=�Cߗݨ�筧O��e5����S=�OTq�e���5��*kT�bi��\��ı�4(�N1t�9�9�q�W�\�#"4�55�[ja\�T�<�z�`�
�ŕ�Kjb���F/$Y���:�a]��!53�L�Q�	�zG*o���.�����HA�6�h1��d�? Jx.ulU�݁i�ZWC�>��h�T�+�@��������`c���K]�)�#��p_�cʚO:tZ@�:*[���t1��r��8��tZ�7�zv���zL��X��]Ү{�:(C�v�׮�m�����h�K "�Z'���0�qk��k$�E3�v��x\d �N�jc@K��Q� �&���%fېuA���FQ�7�����糰���N�Y�t6'���.�I�E�N-uH����Ⱦ$��s�5�N�c����3]�Ç�Y&�"2;�Z]�7�%����5]g=��ܴZ���h�����,���߮� 8k���5IRum��1�w�	�E:�C?�#���O��~U�x��1��	��15=�{F��`�����6��#�5DK[�%Pץ�&h�@Yp��i	�>��ſ589��SM��K|r�F4��?��'���/���fB'c����39�} ���	A4D�9U�_}����s�_�ܯE�
p7\��o��x�!�qӲ�:����?�n����}(���Ezz,��>,�}Ǜ�P?/�?���q�(��7��9t�t�Uy�/ɝw�%W�^�ӧnQKH�z]f��u�^�.�|R���q�v�~�J�u���MĤ	]f3bQ�<v*(�O���
��R�$�1����~��_x�\��T��0%}�?�S��^�o?�|��F/F�2=#ǎ�y�H׮�<s�V����n3���f2�n�J�(�K/������~PN�>-�h����F)��ɕ��\�v%=��w[��g��N��44�f�)�uɜ�~�Р�F�:n6��N�L��;����2ش>�ǉA�2ˈ�߯�E4��aЋ	�$P�%5^���->@�OĴVv�]��nm� %�{���p= wB�YSk>1�F��eA�~�gWG&iR�95�9B�)kgKwԐ�W�� �=M��&�[`�`{z�q��m��Q>��� ���[Ά<A^��+eR��⍁�m$�2�r�ja<�GJ\e�P���v�0i��N�̍Y5��:)pPȰf�ЀiX�J�I}.��M ^E��r��!7��Y��IT5�� �h�,��D����A�A���U������ӹG;�ʐ��9���99E� ���hԢӁ����e��j��LN��d?2Y���:�we��am�./��l5�T�5��0;�@�H8a��ׅ=���^�����Y3s'�k�H�V^�d��9��5�0���5{{5f$2�4�:`��P(eI���Q�z������d�L	�p8�*��323�<>��f�M�?i�1LE�#�X ���N�I�,���`���+�sD1JA����.�-ctJ4�a�jdBI��$9 ��;x��
�t�Fҙ����U)}s�,Y�\d�}�n�N�b��_����!$�� ���z*"�1�h ��ه�=ֳ��S�T�z�Wu���(�4�IK���
h!G��1�����[������zC�U�8}ÙnR�&�k�O����pq�,ǖf�=��y�pj�k�R����q�̔�Ȼ��=���+�M���o��}�sr�Ē*ݘ	���FP�_�����X��L�aB� ����$D��A�Mc��R�B:	Q����z��h }���m�Ǐ�$Rqw�u��@��=��
�ԇ4J�|�U��1c=�����知a��{�N�P��f7�iuA��dD�0l�fx�Kz?�k�p�<��E�M����[���:	�ܜ��s���P���AJ=f���m�X� �n�$��}z� ޚ [b��U!W&�#1��4	,`��G����յuH�C�2AFQ�Qͦr�D��s?'8C��h�9��5}��y5��k�b6���"f�c3C���D����K4~0��0��=w����&չmOv�) e�,�����N3M?@�F4��7��^+�cp|.��BcC������ٖ-�B�sA�c�,,�˽��K'S��{N���M�a��y�󔣪�=ZC����7@�%P϶�
�Q�vz~Ȃ�'���kQ�8���P�s������/B���B�H�8q7Ž�){(9��ŶO������sDYJ�G�Cg�N�ƨ�/}�KWW�� +��������<��wp͑�
KXò�`�k�{���t�|;L�\^�����_���]_��ao��AC;*���㼯_��_������_5�?������-��)�x =�^p���3�����?���,�������9��j�k�L!��ZB�ŭ�{��_�U�nbtp�-�k��_�2y�mH������������=����_�E>��_�`X��:s���o�[:��wkh}�8�*�$8�2��h���	���̀9�3È=a��бÖ�	���ĶNN<>���U΢���(���g<L ��P���CZ���c�������������C�a���>71"4rr#�6�QOJ:��1HF��S�2U�b.fR��F�.�k�F-�_��ۈ<\�~�lg����������Q�q�qrc����
�F��Tt�#�aʣG�d4�Q�倎��kD���0�����
��FUʋq����F&� /1@�Q	��c�+���=�1�u$�[Egk?`�"��I5�d O|�1�_W^�rޑ���*��e���;4JLi@3��^|��,�9�6Rـ�s��ɀ�+)��7�7�FwB�ţ%�g�f
�`g���d3�'���r�5a��'j4܌d5�ed���<�_��6)Ș r�8[�@�i�u��Fk�"HgF��k�l�8}jnZv5
j5�8	��P7g��Q������*�Q[�3�ˉ[�ȓY	c����TV>�я��t�\s��ƵC�����M�� ���}�|�#�b�����<�-Y
���ׯSi�0��I�>�؍�c?��r��Y*�H��E:3�ޓ'Oʳ�?'���'Y."�$0�������x���~� e�D��|��!��7?�H*���^{����|�G>̔8iU���X�>�-6���ߒ�~�����`T
����G~������*|Ԯ	����S������yF|�ot5ڿ��{�~�'#������ŝ$��W/J��g�<5�t�0��ݔ���@���������=q�����V��ɂs�J�?�7��{$d����7��(1 �c��W�Np)>G���i�Rj���y�;�M�d�ei�1q2f4�'�=q�׋g����fˢ:��� �z�'�h��������$��њ�Б����̂q<p: �!`2#���	6����0��z�{���[�@�x��=����ŋl��}�^ ��@���ג�����������z ;���Ʋt�\_�8_������	Ifm8�G���s���I�?����X�Y\����~��2�w�)Cs�V[��^�i�g~�������9n|��m���@:L�Ro
ޑFᓡ
Z,#�L��P�j��΋%M]�ݩ��7�L�Ŷ.� ��ށV��9�W
T5=T'�yL�-
l��fS%�87K$���3����Ӈ�E��`���z�|�A4/R��I���f�T�jZ�̀R����w'$�(���ݮJ�í#��zkպ,,.��%]ɋ;lI��S���7e~n�(�+W����5��nP�ַ���+<#��V5���Rlb( D��� b :���^��c��Jt0� @�p��P)���FS��9�g�R�="�7�dF7/�?�����}�~���1�T&L���_���`|Rl����ڐ�rAΞ:��pU�/O2���شF��Z�<}��hZ���({��6:5NGõ���z���Uj=�]3O�ߩ|.>��qc( E���:=��;ԩz�Fr�T�QJ�)U����8+��b�a�ĺ����g|��7�E9���k��R�1���W�Ա�˒>{F�`N@��w�˒��r�':	�r��ο���v�iT��!  ��
�������[oa;�P��5L��xXt��NV���� z��ˊ�J"�Μ�z>zLn��f�]/�;ԕ�cMrU�'4*[<tX���(d��; �[����gh�i�e�dK�9&��r^="�d�����8����t�R�4?KlM܍4Vפ���"2,s�Â��#�B��rƌ��#��i�q�3��o��k��y�|Q���:s�,Uk����� � ����� �J[����#E�?�x�-d! �E����qg�gb@���jn��#z�al�Y�p�0����l��{�'�M��a��?bFpd>��͌�Xt���SOs��2�èHv?�I�uK�"�M<�����j����:��-�n�t�(\e4�	�c�D�Q�
O���������^���m�P�r�nd�oK���b�e�bm|ֹiS��$'L��`|$����56�!���ԉ�d3��h�P�2Q����>�l^�w?)]� ��rb@��眽��!�R`|�P�_���>���eTB:kvaQ�kF{�Q���{lk�OCY��B����%��j$k��ז�œ��[��'�3��I*��Ǧ��iL��d�am/��Uq� H>a�?�g�o���و�۰+go?.���A��e:4�gd]��u�i�S�?&�[��9/Z"*�P�0��*�0N!q6�ҡ5wr��U���Z7mm���?��]��b�yn�U�F������W��k�����owe��ɜ*�V�����j�Q`#"K���K)*SF ��}#2;���+w����_��*(�����?�����vi��Y�cL�Y�R��>�k�c�{|��}�� ��rE�f�p8	���?�Lc�*�,�l�(e�ݵ�e9z꘭��X.�4�QtW�.E �z&�m��wЪ���j=���������s�K�#��;r}}��Y�A��ޭ׸�P��ݪ��5�̭�Is|'�%��KE����D����wJ���(8��ňU����Q>��/~I�V֙���Ըv�=C��2�~��r��l��J"y��%��^�}��˷�z�P��'��-������'U��S�7p��%���wy��){7����>%�f=2L��Nx�o�/��_6��0[�'�&}�� @���AȔ�f8�a����G�����̅�]0�6FF��̨�?�N���������&�G�Gt��n��U*eb0���	�%�������E�z��2_��Wd�5
8���a�	Y�;2HX7\J/0Xp�J�ٟ�������=���ق��}���pHj�`�D�ȷ�|��D�����	�՟Q����[�`�I�{S�4� �����<��7u}3Q��(�"{WC�ɘg��q��q:�ĩ��:1p���|�ЄY��-�Y�8�훼0��k�����������&^�B�������������/+ŉn%��v&�ϸ�!�j�@�P�{l���*���ݪL�$���lRt�Jc<`��K/HVU0�GOJ�%�r�0�$����~f���4�LT��ɿ��o�铧�F�_��G�	ŉ�pN�mu}�-+�ȐBn��2;wX��Y�v��܋���W.�&t8�hL�~�6�d1�ꄄ�(����$�P����z��++�3<�Hţ�9R;U�p6��t��uU�C50�2�A�s���#w���M=y���'~�W���ˬA�-U�+�7�!�z�'{��G_�@a�j��{���E�y�ӯ�����R����SN�<-�䟓�U���M*R__�B���"=�ʥX3���YF�)���ئ�?Γ�	0��Զ�A�Fꨡ�������y��E���;�g^VE�i�� ��
�����7#H��U�<U�]Fd��@Zݎ�����s�Ү\~�<ǚ�9(��k��O|�Q.� -m0؋j�_y�U�ԁ{�L���ȓ�}�/��ǟd���H4�#��0S��W�sj�C�<�ښ�~����f�T�p��Q�1@j�
�9Ծ!�iK�5F����%������Kb��J�9a��r
"�.��3�(BKU��3*_QG0���T��I�lD5@����"��J�k�e�P�H�����6f��8'�<�Y��0����e�zC�����/�3H]�38�9��&f3�o�
�,% ��g�g�K��l��"�'yf�*�Ԑ��'�O�哧�~��A��7�It)�S�	��h�ر�E4��q�3&=���a��a���qH)m�t\O'n��ٍ`�	y��W��I��Ϊl\����j��g�l��%m�/�O2��2����Y�
���6ֺ�)�Y�K�U0��� 7�)&i"��Ἳ;5^C��^�Ͽ�����(8I��\h�I�����:	��3�@D��Vh%D�nq~F�\���u���rh(��I�m����9��Ҹ�6ז���m�	bwHW&PP�zcێ�0�@r��|�@�v���0�F�=�5���-��۶�&(U̫���ە�rN��~�|����<� H��6 �C^���_���G��F?4��;Ҩ�Ǜ43�QgFD�I��PC��F}ԥ� ��Ac�;��vӌ=���<?��Ϟ|�'�'�-����9��^x�ɘ*�&{'A^��%b��V�PG����<(�7F��5q���S��l %��pN��CGٗ�*�|*'�3�f�N�z��������u���G; 
�\����������t^gJD	�2���#Oy���ԟ��^P��a.0 �N��`8	� V��Z{��І��?�3-L�v�1�4������x�\����ԶdKk��dv��-u�@6�Uc�nVՀ%��e!s��$2i����̼g �����O��dL�~L������KЅ�6�L��2�a��NI��,c���cf���ˠ��������&ih����WT��_��Ǥ��i�?!G5�� �%�$�"R��N���6#7C���Sވhx�v�d3�0R^壯Nܵ+�dxa���Ɇ� N�f_�;"�V����g�����U�v�#��Yg^�4����U�qQ;�k2_Ʊ�j�TA�}�a�����Ȇ��l���p�/O������ҥ�dJ[�P�NcY%��!S��� 5�� ��Y��Q����D>�����ڈ?eӬ�>�2.�@����1KKBl�Z�1].cVHRc��^�Sgm�����D�)��14ا�6��T��yc�9�%���t/�:p`@��il�9C6�9f��d �?��Ǵqa$*�Fi�I�����f����H&� 9\3C�����7<�+��Ĺx,l}}�T��@ TRg�@7BC��"]��!�(A�+e~C�8o�h�;p(�0{8�pNFHo�J�3�}v�*�X�f�ÿ�=/t>��	�`W��� �[R{糐K�íΰ���8`�c�a`K1�8ktJ�Y�s��6����2�~��c
�`����1ʾ��8fBMpCKZܢ�C仝!�s�'\���i�[���r��;�c?��z���:��V=�}n&�\��|�]�4�	hi��X'���>�:4y��8Ɔ�
S��pp$��.�$8�g`� � �j�
����kv�4=C�����L1�;�~�w ߊ�i�$s�q
g_=S5=2{��d�s�|]�jvJ
S�2���q�Y���iF�P����2�	F��w<���cj'>#�V�C��z�c��p�[�� ;���d������o=ɾspB�
�S�t�o��/�z���7�ȓ	k<qeO�[�'P�`c�4��!#���Ndf6O� O���r���J�<%'�5��9�o���R�r�-&F�r�g�܋d�I\~��ga�H���:�pz�6�+���Կ���4!ԣ�}[ƿ��Y�x�\���u]t*���]S�^a�L��=o�W�ʎ|����Ԭ���N��)�/_��� %��g��R�Dh��,���`"f���<��3� �%ձ��|;��F~�1��)~C�D�.« ��:ց���6m賄�q�t�dF�=��l����ro�=��a��A�j�{�����(%����L��#)��$���\O�2���$7$c`����S�F�x��6��I�^�O�2�=�Fӆ%�Б	�ƴ*s�졣������!��UHv�N��K�Yc�~"�&��7�����uD:�eȀ�Qx��Ģ�F�x��{~�T����R�?�4�B�%�k.��729�ΨAt����Y�7e�Pf�^��[�ސ�'�#@���;�-�bn�2g�����Ӝ߳�}cӯ�vM�[ܰ�����j8�t9L�Diэ�\�!3!�K��T�����.����wP�h����	������=���^K^N3�`>���=,�>o��'����2ͣ8嫗���'��z�ݘ�
jTT�&3�c`�Zd�5�Y9}��,_�,/�{� �(D�q'F"D��Q*�>1H���$*1HL�v�jP�kj`�L�����S���4��Q�^��J_ag�mc�tR2jT��4{���[�la C^JSKz�,�LbB�Ú�k9����Y�>MTH�����qc�JQ���#7v\����)ֈ:=o�֥���H#�P���gtC��i�u���Zc���2��bq?!�Ǵ�a���0
�(d���jT�Iii��4�F���QK��Ug�lQ�
�U��iT�Tul�@�t����x#�c�i��eG��V��amc.oL�z�����Z�NJ.�t���F�a�d �ψ2���}V���?�
8-��~�i`��Ȑ��{�
?w��>H���!�M�� ���P��i;�2$<�[�ChhC*� �b�:ch��:�Aּ��<���Ӑ�iT8 pCcvp��kzh��χ�>�7��������,���ν_N���gz��l΋] ����	.Ra@0I����,J,�UU.�U.�M�d["��e�*Q$RiI�DZ`�b�yw�N�����r���9������%)���.���p�s��=�G��S[*tF�Y��c��ʔR�y�	By�� �cT�ϒ7�ŜUKP6q�lV!�P�W��3������Xā8���4c�������W��m�K�c`�?�wn>�Np������hus�{4bF�J��C�\)*΋��u�ytF�ė��qw��� �>��F���u	�>�:)��8�g�7�A�lU/c�;\K�n���N���Z�ց�@��1J��wU~�0rQi�t~n+�����;�l$��[Y����#G�h�"ǫ�*0ݿ�59P֍
��IO���;r��#ER2˲dy7Q�Y����Y�`��t����G��b�B�֕�����LD/��M���!v']Dp�[�ی��*�*պ*���$F��u�3��������c��Or���%U��9��.![����нls+gm=��G��.7�S h3X�{�X]W%^u��2(#�(�C�T�kR�/X<Z��X�r��t[C)�WlNZþ����{2�]#�I��n�Ė��7
�#������Pi�gn9�x`)�RuA�1|w�g����я}���_��^>i@���W�?櫧���9�c�ա��R��j��Z���ٹY> 8u�vvV�^o���:o����;TA=r����Fز�-ITpY}l��yFV��w�8( �Ekw'�NLM�B�܍ͭ��ͅ3:���䶦�r�;%^�r�L�P���/{�xڑʌB�"P��]Ӻ	3�<ϔa1�#xyN�;�?c�O^y�����PaZ}��=7�s��� ��a�`66�2e���S"`\ܞ���j�~�xh<�0����uY3�1���[�����{@Sa�.��O&�� ��P9�����9�#��N�9�Tf�O����a�<\ۉ/gˌ�B���=79�Q��*���L��v�ӵ9���t���p�3��7p�^�������x�}�&Ix6]�8�c�q�Q�x�᎑��4�9*5#9BS+����US�Q6x��j� ���g��(���	h�ؑ{�l�P跤zt�r�ss`>�1�T9��'Tb�[ �R���������h��.ZaZ őCt�1�%pX�2q��4|���co	�F[)�I�.Zmm٬Uԧ&���������5��$�����~O�nK�gU�N�k/�B��蚬�����C�Q��ZY9��d�@I�*N�mL�ȓQL�H�F��Ԭ���m[��"�5����a��;�sm��*�=`��옔��	ʰߕT�U��t�Ols���8f�b�S�ZE��4\�;0M��X=�]��"�]�:t̀*����q�q����;�|EY[O������_�Bq����O�	�؛�9�U ��PW��
�B��8�[olc���3���'��p
�t޹x���`^A:b�J򳆰Ǻ�W뭷N�GnP�������Y�\��O�^2�
�N4L2�҅CK�YC�z�kTp�pT�<�o��G��ч���'h�P����,m
�J��^�R�PL�nj��:�2T̼��X�q�c����s��$A$��O��� L��kYD������p��m������Dft����Y�+��M���}�QK*�)�a�]���7�R�ǐ;�!r���}���0�A%�B��3��lv/Np�&��J@N��0 0.ȥS3��#��p�� r�?�q���y�_�:OT�\�4��PH��L�(���d�����s����)v�e�F���EcO?��i+a9V�y�s!�G�On3�W4"M3�\��5� ���R_�f�.��ć�ұ���X9�����1�@$M�02z�4�l�B��Y��f2�ps�Ⰹf��}��Ȅ~5[����9�3�d�C��T���ԯ��Y�Z���rQ��K9kJ o
q�y^�d�sҘ���z�έ��KV�b��^����yb�ȵB�0Z�m0� ����s�e%o�{�3�
5�:������u��%�V���o� Kb�A� ��W��Dź���CD,�6oi���n�¬	'p>cܰrKU7��	�U���6*l��F���0�XT$1a|���u�z�]y�λdF=g�yG�Drpeż|
e�6Qv2TA�d�E/� ��ݼ����&F��-�22 !�\W�E�\��>��4�{u7v*���ܼ�?Q��m)��n�So�)��v�gb%��!̈́6������B�S��Ao�����R �W���2T��|=�r���4���}�|��CE��_���Oء��+C�o^#<O荙��c$lg�V�G)Y��J�j��`w9g���[���k�v��!� �e�Y('�=�#޵�`��� 1�Shlqp�(�T1��ypX�j6'�.��{�=�� `2�L%�+�['���c"�OO�J�x"��}��9��-n9�L�d�$?&�4 �~�l��i �\�ad4|f`�0F�A�a,�Ξ���l��j�QJ#�k�Y^����o	�+dd�+��z&2����S��?\R*ۜi���s�~���X	�U���=m���C��ӑl�7M�5�u�V�<���S���9�I�-�rɱy��mXA� �!��8��4<��p@!X��������}��<܉��[VE1[����Mi�V沽�+�KR��;P��JP>�F����Mڮ.0I�Uڒn?��ٲ]�(�>4W�
E�n�M1//V��OZN���@�.l�����r R5�b,�X��Q� g#��)6��0��[R��S��i.����h:��T�$S�/n���PR�F@��*f���}{��6 "-q���|�;��}@Μ�ի7Ore�V����@��Dv{�֌&1�{d9���\bP�bޥ.``��EO�Χ�g{=�F�}�7�dak
����PhY���lo�w!`2/��ߘ������C@|���@���s��UkgO�����Ha�=KRB���
�=Bc��
���U+x�]�U���~��<�� �*Cӌ@�� {/�T�=Z�b�;��������������n���5r
�U*��hHa���F�Ti���I#�c�8���[�悩|Xϰ;�e,�V����iD�y�C�G��c�i8��ErH�K�Jcġ��l�8�T�q��U�1c�I�ivq�5�\�����B�1b���xR��Ã����E�~/"�e��)҄�<i��o���yK�=+��g�M��ʵW��8�]�E���1̓�r�f��ޒAV�K(cb�pM9�3P�n��-�hS#M�d��KJ��Wp�&���ɨi6�O6����[�%�P���憵�n
���Mф����|t��`i�f���[J��^�5�*���E���~�Z����_�o}�9�o�'�B�J06��M	�T���6�,;CY��6 m�+�BE�%
���5�v����iY�."�� V� K&�3��h\�.H�P�V����ۤb�D��Ҍ(�0$r-o1�j�B�����P+?W�_�� "�~&֚N��m81ZF4��.ɛe���\k��|���%����&pvv��w��%KV�:@�U��D[��CVSG�`a�z!�ڱb ᘀ���P�o��v '�1cV�hDz}�lw�7���������7âh��~�ރ��ϭ�P�'�5�)�3����z���k��$̧� ����{���|���v�|�~�A(0#����|��P�Y�._��N������C*8*k^�DGd_�,��s��q�4P,��e��H�0"z��C�J'�]1�9�$Fih|�ahgTE�cݛ� ��g�gRc>�
�J��?b�?�C�����85\C@ ���O�E�x�߻5G�<�3L��\��`q��	�+�r�g�#�i(�A����G\Ȟ[��Y�C��
z���p��:�����;�gJ<����=+_b:yk^���R���|���/��ݡ�B���U�xD��z��p�Aɫ��v��,<$���oX�^� �+�@��\�a�	s�y���P -=��#�M.ދ�����-�N��� ��âX@P�ֹgǕ���C��}����~�{䙯}Y�?!�y�qyꩧL�,iݵ���Tv�.9z����7�wL ��@D����m��_�s���c�Xv�jm���wJz��� �Ͷݗu�t�̬�n��܌����ES��G��5�t��yp��YƑ8B���fk��d�y�3=��g��Gt� +D)O���~����|�:�mpcW��N�� 5Dd`D��u��뚈�w����żE������Ȣ�>����;힅ہ���8f�D���ʄ4��x ��>;�j����=�ה{ཙ�Jf�#�?�!wS�w�9��@�(U{�6�]�@C氻� �@��e��t*
[�A��F���#6��0�$.��N�i"�	��w��T�0>G�"�Q
V�������F�
	%s�'S�ی�s&�ѣ���}R��{�8ǌ�7o���u(�L�G��̇l_"��q��H�W,T�4��=�p�}�9�ug40��8�u*q\�?W�(hq�[+Xgx����;�F�h��u.z)0�¨�[�ճ���3�`6��cpsZ	z]�7�(f���0;��k��RV����TA�����>�%}ܛk�g��?;�o  T�?�LxV�Ap-堉���\3��]�S�kX� N
I�RN)*x㣡��?t����W7��X�IUeY�{�A���d��mt<������f>Ώ\h�Ov0w���vsG�����Wda�*��������r��[2����Vs��0����ӂ-km'̓8ld��[�ǲ	���� �&Ka((ݦs&56hM������������@ ������֚�� �۶���dU��ԛ�$�>]�{��c���@������m5FvUٗ�������W�V��ǎˍ[�r��u9����;w���N��e֚�]-yjd.qTr������(��uF3xg�IC)�Mk5�Ph��d��R7�a�k��Q��l�N߃�FV������ڻj�����6�m�����lU�i����Cr.]aJ�9�%���|�wo�/SH�q���G���#�N)X�<9�V�׼?W�u�?��'��w8�˨zP�P���<���~����w�E��8�,�>�01��<���	 �N�
� ������\po�E�	���p](|�%xTdP��,����8'��6�щ��<`,��k0C\���ü������sڲ��3r�q~4���Pa�>qb������91׸k޻��i���h�H�0J�T�A��z�����g���q�5�P��4�זq��K�8�ɢ�Ly�8t#Dke�)����zB�� �cd-\���آ� X��ݞ����`(�=�gs��tFF��G�Ĭj�S�����_����yN��?�?���z�����vu�i)�G���J$�9t����V��-9qlQ��O��|�c��/mȯ����&�-!��8��wPf���vv�26���4vE뛝s��7j}8q��\-�UZU���:X�i�w�\���=��TnAU�1B�T���?�uB=�}=l�T<+,zz;h`�����/1�5ꎔ ���1*�+ES�C]�͝-Y8� ��Hz�m��zu����47'���-j����X�,7��c�c�{�d�tZgm�۾����O�����9(D ��q�E'H%"DT�G>vȀ_ps���9q�83�|��L�D-��5Z����{�$v9�� � �!�H�f)?��L[(J�!�5��?�&�EWo#.�} �'V�DZS�T]�_2�*U}��[�1��U9�9�k�-JM0v�{B�a���8S����P@���}F!�ô�+�P0R�^7� ǰ��4u5 Sba�?!��+?�{�x�帲�A�B�x�|Di�S���%^ 
M7��N)��g>礢�ر\�af�O�d���
�q@��9s���F�C�`L]����<if6�|�GɉK�}�Y%� ��Ð�EԼa��xc�h���z��s{��'��C�O�<?C�0p~4�!����SX�ESPs�NN:�[{����.pp�q���Բ�"7kk�v�x.<g�&L|��cu��m���>���r��[�60��^��-��u
��N� ��.�)a������O>�OX�����n�g϶��T\�8��u�����j���o�OF�<xom1�POMq$���*�R��������_tN�}O/�׾}�|���g�|c�y�&qD&��X8LR�>�w�2,�aY�,��S`�P�Л�o�CA�:���M���i�ʖ�>��*ەE���c���;��W�^��zȟ�E�G#|Y��j�r�}[̓�Т�^+[�+/?'ǎ��<�$�����벸�b�Y�֬$ncmS����Zb�7;��^��|d#!�V6��4�L���Y��b�A���3G;����������l�f,�O������x�alũS�0�` �^��34Ux!L	�����G/s�}���q��l���`�|�rL�����fp�I�G�ƱS:%���a3��L)P���<��`o�,��>�0���q�c����Xf��0��8�,�m��8�?����@o�a;>�k�[μ~Nz����B�E�¦1P��*#x(w�Ue C���<0}n0�� ���s �9�m���PZxG���P�P�̈��Z���fB�Gv�Q~�ܹ���,���ϱ,�:��s㚸w(���_��!G���3�'Y8��-��~�8y�W�����7����!�'X��5D�;�5����:����b��i����;��p=��P��qO�ÿyLub�`|�H��`Sg��`��"?��˽��+/���ȉ[��ads��QV�8G�n:���@*��*��o�9�~/���������Auh.�?�4���ht����둞��_��E�V1X��Ȭ~EM�4]��b�yl � �^8�1q����/��/�^o⚞V^ 7ظ�SG�2�ŵ;t��1���f�z�Nnv� e���[�;OB�-��H+�<?w�,P,HԚ#���@�?���ޘQ��� �}�LmӪq��ѿ|�j�A
>{x���P�'����~V>�׏��s"�����m4����-�}�pO��J�lFB���(tyb���>�(lqKR�����a-KcN�����uLWF��	��7���6n,T>K�@�G[-�z��oe[L�z�YzpţQN�Tp�*NbW���ؿ�\��+DN��P0���0F�k�1�s�b�=�!v�	�pL��l�CO���1	�c��-��o��Ҁ���SB"Sen{%����\!���Z � (�>~����Q`R��>"C��ѻ�"�_�*uz���?GX���rȔ@���Bc��B�R(>�<czo�_�x1��<�-@��_C��BQ=�M���g�yƼ�#G~�c�=j=��!�g}}MN�8����
�ǵ����e+\s<�8��w�a
��9M�\��aJcE�?x��W��n�}�L�y00J0������q_0<@J�*�}�#z�"-�~��{,]��
�,�q��18���lnp�h�`��k�Q8#���[[���bۏ�.���0��B�xv�υ��y{��D���[��	��L�Ҩ�A��4���}��ὺ*{~��Y~���v�X/�K����:I�� �X{[)��u���6�$�����=ܛ�N]��lK5�˯�.���)��8l�诽yM.��ZRmx�M�X�����秈o�f�qS:Bp��d9L @��@�M�ρ�d U����2r���}U��<Kl�sR�Ù�vX�irt��Ю���z������f�"���!͑NPMe=�gTQ�g��4��r��G���dgS��"?�c?&���>��=2e�/��Q�o%=0`R����Y�����+�\eBjarDC��7T�h`�p�;�9Rнv-Ǟ�O9�C
��7G���*�l8`]��Q?]��;��	(([�P��,D坒(D��%)�dA�>r�[�N\��r)gdC���*��FL�=���ʈwX���-�\�e9��<�DT�T��IUB��y)���tzP���5��ztQ�IflP	C(�C��݌�?�c,��O@��y]zu�����E�9��M&S�K�rx���eA��s���oy|��;Y
Ȝ>�b��a��%�{E�u\������5�}�ԩ,�=�8:�1�̒,�AQ��x�3"�	���7�{��PB���H�~� (K��
�ک[#�)i�8���X��^/� hĂP�4מ��w�R܃���`'z��� � Q�0<�9���� F�<!����(��s��������?��Q.���+no�e��d[��w;�����C���ý����u��M��b�\�U:���0[��ˡ#7�z�	Fol��El�7*�:Q;����'O�K\q>�+$��a|��N\m���+{7���ߩ�%��r�:8Y�`.2F:,��z{�u;����ؚ��|v�kQ͋��4w���E$88�o�����S*�O��lWu�����x�	��\�u��LD�
a��LE���1�Jsa(�e5:�Wߨ�K:���֎\�rK;$׮�<�ͯI�ݑw�'g�]��X9�����SO���s\i�SXH=���xc��s^��X�"˓�5��j(L� (����|��0�Pbg@�k��A���&�S�E#���	�'�|���� �2����d$�!!��T�*K����A�w.�8��|b?ɤg��p�c�'����C���+}����|)�$��u��9i!�Ja�=�GZӦ�p����Ut��Bŉ�Ы��� 
b�m&]��$x �v��{�=*�Q(!O!	M��g�*̩��Ya�J�9|~�ÿ�(A��p^��6���&��!{�3\ׅЏ������{��<���J-da<@��zo��f��1%�׃�&�:T�L�@�`�A9#���5�0Xp?���9��1l̺�m�H	>��$F
Xj��F�9�3y2´"��@����z#���ӹ6����D�J�S��Ч)~Ɣ��8�Z�Z����]Ȁ���&�Ɖ���)Y�p�_~��W���!_[Ppc�T# N�O��H<���W{�g����+:��a~�:օb�����!sH�qѾ�N�W덖ln� �H$�L�LP�� �a��G2So�66��A|�걗Uymln���RU����q<JM�Խ��ڧF�w���¹��$*�Q7軾��x��u�9n���
�g�<�M,r��J�Pq q=ꍭ<���i�Q�w?���_�ƾ��O}��6B0��̚�D�5Ԑ#�0_j���iu'���-]�	��H�Z��ܼl:V�
�b8{ތ4w���0[�~ÿ��/��Q�������E�p�������iтh:��%��Djڰ�綄F�J.�;-su9q�1��@����U�X�R��J��e�������N���	�ܱ�7���Vo =�#c����\[�D;"4Fo���{m�|D�)�X�� ������9��J,�H)W�ܤ���8�Zy]:.ɸ�����A�N�|���X�ј�
v��!�'�da�5����`.ǚ�����/�6烂4���=� g�M�YWN���.HY�{���@h���@�y)�)T�`���:� 5��'���7D�:�3��P�x�����Of
�!y*&�a3�
�P7�axx>��]� �c�� �%���ֵ�s@1cLpN�ډ���G��
�@T;R�0.��cn�7S�^g ��J�����W��Q�a�0₨ ���2ŹP
fs�N�38?0�qm*E�j���[[n��c�ݳ<ӭ�O3M�~I�J/����p6#F$������\q������1���Tr�9hܒp�=��������t��-WMPs�{��.�)��c�]��{>��m{rsv�5b���׽?Z���Գ��-�͎�dT�Ɋ��3�6��ą�?XI�.������4�P�*`K������
g�;�G�YG���H�-&P\Z�`�E ��U��P+¶h R,�2F��
_xL�(���1��u^r�#L�P���<x�1w�>���C���]y�7������~�R��dv~A.^9��T�g�R�3�v�)���A�J��(?˗�3�MA�-)3��@���Fȱ�@vϙ��m���_��k#Y�l���7��3T�\�����Ai�z��\�\��j��Y(��oK=W����zYn� Y�qQ�����w>�	y�#���Vs[~�w?'��:%۷n�f:�םU�搷(�˫0�n��"Sެ	�vw`hx���BU�˱,����Ǿk\~b@�mݬ��WChF������ł~�Ց\�j�����2T��?v!ʙFA�n���������O���>yJ���z��|���X���5I�ĕ��3t�Ci[����S����5`z���s�q������Uì���3k�<r�k�f�a��1��Y�P
�#�����wxd,�J����ʨFY-3��8&��>U+ރD�Jr�R�B��0)>��ҤT6C���c#˱x�=2�1]*�v �p�9�O���������f��M�/�} 7�^�P��N�����8|�4�m{�ӵ.FX������Ҳ�����בw�XBq�Z�͢N�E�=L@᠒Jφ���U�m�~��A�T�
XK�\�a��{������}ꤔ�M��k�eX��!�677t.]�3�;�)��E�#��PQ �B�R�5bp�&)9���n����EY�Y��8��O�Fbp���S�H @�s�0���=b<07�+x�� 0����8a�u��T��ft��2�t/�kU����F:vϸwC�#򥟝�[�s���w�5o�z9�����J�,"�����3�����y�t���.ȭ��K7"��
������Y���8���`�149f/1��#c}�|;�-�2����B���T녪5�(%�*�r[#;L�мd�n �� e�����j^a~���ӆ�Ycqa;�љU�C�N��2��W���l�zRUO���5+;+���vS7��*Т���{U��RQ�h��t��<�K��lmA����5i�Pn�!
�Z����hMQ��w���*� D�K�������ȑ'$��I�C��,J�[1�]8���Q.A;��S�yR����cD��C�p�<��o�cw��~��g�+���K�T�H��;��ݔr<��:,s�tO�vJ�َ<,�~�jƗșSg�Z��ֆT�M�b��B�rtE?s����R��~�ow�f(@hl��ei��f+��~���'�e�!�FKξ��������P罷�b=�W�|xإr"K�L|;�$� H��}NBvy����!�X��4�I�v����2�����^a.<<�Ax��� P�����Q�%]ɇ��#�r;�q/�s,��5B�6�9�X���k�0>��;=QWr�7ń��=x�[}�ֆ��=��H/�1?)k�G���n��'��µ��gX;NB8X.������x	(|(y6�q���"�<�l`������`9ڬ� �9�qm\�5�*x��x��%0��%7���8"/nߥ�~�H���Ü<���-�v¸w<�&8�Q�� c`qK6&>�A '�$�	�3a%~�����(����k�H ���/���&7�G�['��\��s	l>�w<n+��t��!�V�����7�� �C�P�yS����S+5�e��[F4&�v�^ɫ��z��#t�!z;-�r�C��@��� !<��@�Ò-UjE�0)�|U���	�J9L,�$Dk���{#]ܥ��&i�7��FIQYo�4#��2��^z�R�(�3�U-�<���B]�#P~6�<#kP&3+�Jb}��)�T��'���ڱUd��N�k�S��}�*��N�-�Įo17NQ��F�"��{�����PV/�E[*z�G�[�����Ͻ$s���)_Xt5�s��/��/��O�+��+'�WO�K����CG{��R�\='�hK��Ը�(_��l�U�]�������W_3��ٙ9}��\�|���jE.��"��:�^�C]��|��?,���ʗ�&�n\�JA7���#O�W^�󡑂Ͻu�a��GH�-�X�`��?�V�#�!���za�V�+n!I��;-L�</D	bx��J�`b}4� ���`ió�}/�%�	�T�̻���4���o���T88����(�#�����y�}߰�˗�y�� *�Ne��sϙB�w�o�8"���;�{��M�<��9��8�昳�\sl�@٪n����=�p,lm/|���O9`<`�Y�]�C���c��6����Y0?,A�Ƈ�f[O�-qJ���G�+d�M��%�|F�ٰd2̧��;����L&=�>K�9�#<��C�0bD����u��g��p�v�E>��k����}|ڌ�ng�g��E��3S�%����+�6S��?:+9rn�Q c��%u�N�{�q��y�4U"%X�i?[P��x�[�˰3���X	P�q��K��T��lB$'�䡸��q�Z����j�Ή�>�8��"�� �yN��E�����=��q�\� �ȩ��R[��+�8�,p�G�I�>z����<�a�ό���tw<B�yx�Y��ԧ3Ҭ[�g-��/�ܘ�͜N=���Y!��s���-�B��/���X�H�|��_lȻ�W��U����K/�n�#�ϼe�õ���e�\���5y��2_�ͿK>���M��� gwwK��g?#���R)��Va��z�*�Nˌ���e|��{���[���?��S��ٯ��|��U���y�)��
D��!W�V{C��<(��rA6���Lf+%Y��QocM~�s�#�+w�l�.���`�d�z���E�Fm��3#�ݜ)���3��&�O�y�$�t&�:c�G���!��[��VF\�n�`h�J� (zI:ahz}aI�! �3�F��Bz`8�'i
�6�eq��9.%��V_(�0��A֠#�:k|�4^G����	��@q��C��E �)�|�û��Y�5ur�\�����9��p=*c�f.�d4�?x�\���#�,5Vp\�k(�`!� �;tA��J�� "�&�`x>�~�����1\�WF+0�0�����x� 7Ǚʝ��S�ao����՞��l�;Ӎf++���gO�W��w<�W��V
y����ܯЍS,uݳ#���Sʒ*�qU�UKE�5ѐyȲ�%�<}SVo\�s�_�:$x��B<_�S�.ݞ�x�h^��lF����QЍ6X�ʜ9�XH󼁴����v�� �Q�[��V���*�C��Z�m�	L|���ts�n� u�Fz�q߱�a��q�X��{����F�jZx���q?����M�ۈhu�+�d�O��U>�"����r�0�P�mU~[�n�ڢ�Özl35�g�^[�K�ސ+���\�,���$�^y��r�p�n4��W�d;�輹Pܨז���n����o���3:�ݶ�r�Kr\�<�FT�Bة��ޒxؓ3o�,U�O>���6j�օ���\��
�A�s�@�i_�n]�͵jT<,C�~I����	�v�L�h�ڷh	�89_�'��q:�#��<��4Ԉg]�ʡ�y�U�237kq����
^��V�".�D�9Kt�?�w�-�(+yzy�d5�a��f�;��2��F��P-�.�&�~&6!���5l����)؉���ʱ�3@�1�L�}h�w���s�nq> �!��ozy7�'�2i�yH	K���R�@�#l�R7�h~���=(��9��V07��{�2'e0�|�(������\���N>�X��cT&4��P7��#��2��b�(K�²3�	�`�I�K{�S��F���>?��`�lp���V,T�D�2CE���	S��/@�vT�i�ׇ��{;oW�����Y��s� �������P����-�N�����[�]z݁Y�?��-���\�zQ�nݸ,��  �36�b���Yt�Z1&�))��H��؎�J�)h��� �����X:(�s�+�޾iHd ��;-U�=�Dq�B�q�*�ʌT�6V�o����r�En�Y�N�/�b��#؆�F�z�ǔ���V��v��lV��5j���%Q�掣+���>�y�U)�{��uCjey�}wɟ=󜜻�-qy޸`��#im��h'�g��4���Pc��Ӕ��M�Ƴ�q��[�_ԍ��E+آ�+� }��&,�Y���7en~Q��1�ml6��'�����bc��ߔ�뷿 ��cV��}������;^�>qDν���UIG˻z@����dk��ߦ��ob�BWƒ3�0�j$=���8v�r����c�R^c͐�sޑ�a�����Y�L�H.vFYu������&� "�J���5�$��N�|L{�3L�9��$#Cά)'g:���P*"���#u2�IZWd	�k��P&4F�~^#�(C���2���[�}XoMo�Fr٤��gIÉ\�$���ǵ	\A�TXd@cdF`��`��@, �*a� �����du��i��lq|�Ks�$E�Lq�8�0"I���Oc�� �lRCC1�Cb`������p0Hc�T�0���s�cx/���Vo���?�-�dh�ܩĜOW���o+�n��t*�ޮ��7���%U�瓦@M݀����|�&�ޔ/����+WA�
f~�.Uzj��˱��g/��䵳'-_;Q�>I=���ʎz��LT!SU� ُ/y����(�?��_�~�՘�f�G1���7wv����=�PO��Ң;~�*�eK/,��}�? �jCN�9/gu����T9�n��TUcA�S�s*P!|^����G�@>�a��Ȑ�dJ�a�0����V�oMS"c�C�8�a��ސ�9�mG��u�U��FF��w��ϜOԓo�e�PY�[�r㷤�ݖ�{  u���/�s�o~]���k7��g[5E��|H�U��+Wo�=�?,�����zT~�7G����W$�9_���UdW�w�J�� ۫7e��KC�[�}��7���	�ݸ&�jɌ��-��C�G��>�d�:�;d=C.c8�{��Z4��hJ[��	Bh��|B�z�,g3���6}�B��f�/�.�:��J�N�o�Y�([ ����t(;��SW����wqn*p�s�ܫ��(8Yn5���������K!���z�%|�c���&O�鼸��,Ã2t���,���,r�S!�k9 ���|z+h�I�O4uH(4;���U�2
a%z�6��ĉ,�{�7��u��.	q�Jcf&��k���C���I��$�g�=����\t��$�|�����s�_��G�W�Ϛ���-����Ψ-��k��-6��o����cv���W�NF�Z)esǨ63� ��$e�g�chD��o�����s聞��:U�ƾ��;r%2��$x�>�v�w�g��H��B�P���:k��zU-�ֶ)�beƔ�-�ԕ����aꗨ��Ku���2R~��,X�`�9���HonV�}����p�u
)l:Dn=u�uU����qy�{�����x��������*�'��J�нƬa)HgT��_yK����V����Jn��r1�ص�E�o'�]X8�9��4�R�C3�$
hB�f�2�2CE�Q�B����X��183l^5���nȍ�˲�v�Üܼv^f�E�?7�7e�,���̜�Q-֭�\R���¢���؝G���>�J�bU
���@�2�o\ݍ��^�g���_��ߗ��/����l���EF�]��m���;�~}��gU����@�nʫ�}U��^ԡ�n��5���*��ˋzщ^O=Q5�rŜ�w���E8 �Q�a�kr$�����Wz��l�OC��P��B!E+�������f'8E�g%	���mf���XW�=HeO��!e*y�.���0,�?=I晙K��$ʙ9g���d�Z'�����䅿�Yx��s$!��}�f?$����2�I��p_4&a`��d8�<tݰe+_�
�Q�Z��il���7�m�A�|Ή���%[��H��(A������s��k��!kV�L;�����F����z���i�P�����GX�{��gԁ
��4��G�)�Q�n�W5�[:���q4ʙSV*���Y�Y���Q����(��>�)t�|"˻�6r�Ϡ8��QFf\�"���m@ "�#�}��Nef阾�o��Mŕ��#Uȅ�
�z�C��4*r��q�i��PE>�6o��$Z��whiF�pna#<S�r)l�������=w�m��?��~�eW=�?��M�bx�!��9��˦��,#��lK�Y�۷.������rBڽ�*\�y5GPo^yj����+w�9Ƽ&�3h� ^{G�M�;S�«[�BhY^.Fmr�B}���hBR�p;hk�nޒ�lxpI=�vO����,�����o]�g�1�@������PWs}M~�~V�~�a���95�����a���������t�=I�/�lon�����Ɗzo��Õ�����m9zσr��w��J=W��Z�QT�d�%�����w�r��*�����U#�GV��WT7�Ofuy��e��ɸ��<�ם��9����T7�5�|O���fJ�!a�1JÐ^T��7z�,o
��aH�p�<Y�暌3E�s�{�F%C��A\�
K�.�5�NƜ4C���Bd;`����(�_4"p/�<�}�*(v�s�>���)�Z�g�wH{ �E����8{��y��G|��r�֢hjQy�
������-�Yf�b2�/��!�j��_/f�k�>��ԂGa��C�r���w!o�wd>u��I��C�2!��^�X��Bι��1�x�$�|fR钿���N	x�a�rU��e��¹�cj�F #_�шv������c�.?��O�o��祧�V[�5G�i)����(sIi�ı�c����F�؏���;\[�诰z�#��w1�����\����w��H��A�3�B��ZYz�1�P�P��d�
��w��x��\��Y]D�}ƞ���	\|��y8z�in���{�<�R!��E��~�ΎYY̺7=���g,U;-�9X�������ɋ��P]�D�o��oC�A�SχO��E�)I�X͹[���=�����SĮ��^�SťV/jr��gk*�c/�✑Q�����Ū�]u��rIVot�ˆ�P��_�@f���ާ�����K>�eks(���u�ּ~��������6�T�^���F������,�KS)�����tc����U�������93��� b}}��F(_ɍ��<��ou��,�jE֛h�qY�.W�j���q�F}0����#��\�!���R���S�G/�0�eT8!���8�ƅ b3������( �n�]�Bg�{p�'=�=�O]��N��#u�Q�4b��0eh�B�}�z��G�2z���`�u�_e�Ө��&��ŀ<��ؓ@��P~TP�qN�qF<��h�1tM�_�X�B4�" ����*ݞ�a��{�T�8���[���|;˹j����ѐ�sCP�I����R�K�g�b�1!�!��C�xs\�� ��i���z�',�.�0��脧�)�7�>��,����\����~��?�ӿ��h�.��o�w�F ��_����qxd��}o�v
=�┃�����^��(�C@���;�C�f,.A�JM��T67n�H'�v+���U��������ֲ�PQ�kgkU:M���y���%�?�L����¢-m�x@y_4.h�'��s�I.�rM�嗌�5�F�����:w鴼q�E[0��K?u��z����LE�������!t��E��y$�弃�s�ȕ�1O��G<˲�9�9����~�1r�CKW �@���$UA�oɡ�G��5U2zs�z�n�uH+�ci����4�uRd��@�w�e��-�y�Qi�Ʋ��1>te��%@�8ju�>��qO�"9���'� ����s��r}��A�����{Y&)��͞g���5�52���u�J�%C���Q*Cy��T*��1�eC��n5}_ꢌ����N���ԙN2�!M^o���\��FڥŃ�D�U�w�/8q>D�X�O?_�җ2-���Q"�q`����T 8��2�W�����ei\��x."���y��Ԏ�Α���
=W(w\�$.�<�v�C��Y���9��'Lb�Nr8XE�MC
�C��2�%f���4�6�/����\6ž�k��h'����ںZZ�?9~L^{�5���u�<��B@ex�S#�X(Lc8葇8&�L��rsP�`���a���c4*��1~�1�M�1���A���C?�C�`�������=���W���a���0�F!��kS�\�7����/�hW(s���7b�N��M���J̽�=��m�;W�?�C�*���gJ,�&��&���֖�j��w�RT+]��@��Z�)%�':�h(jC��*h';��$Z�n�by�	c�>&�$��b_�ܐ#w�b9g�o�0CG���3�|�	V(�o?�m�+�-���p��"k�kr�����ڞ2��N�+���j)�w���HOEAǴ��÷�T[�<��Dà/9��֪��@#��F7�N[=���أ}��n_��m)G95�&�ᶥWؔ�k��u�����S�&꥿���R��r���@�벺yM�db^�����v;�5�q�q��K��3H� aM�n�3�+�-5��%�
&���To��M�zl}��!�Ո�q��Q�А���aS�xjT ��5k_�ƤӖ�Cõ�E��7�hw�y�P��z�!��y�2%*�J^%�M�S����}��z���aiy����AO�A���������X��i<�#%d��,�:J��4c6=z"�CeAÂ����A���`��!���C��ׁBv�<��t����|���'���4�G�ǔ��13���A�!bB�o\��g�0崼�����~�03�*LaP��7wW�E~��G�5�����#d�c~�&Aq��9e%�a�u�;#��Ѿ)h.�Ƨ��ڴ���p���m������P%�yX��hd2u���5��y��͐�Ї>$�>����i�r��5�7�'�}���=Pk���V
=1-gu�����ֶc���9��O��G�K�� D?T��"��]��+�٧?)������'�����	|�y������,��Y.���!�+?�ą���`�[h���j���*4p�b]�l�u�����ѿ}2�r����N��JoN7���^G���W^�e�ؗV�KG�(�����QV�/Z	��`�R���_#�٧e-Y�=%�������3R��i.��,Yt���mZ.s(et�������kMYX:.�Ɯ��r�t��D����%��s#Y����p[;M�!D����y����{�%��ܬ�n�ʟ�ٗ�ܑ9�@G�=|�Ʒ����y�"��5�t��fTyW԰ʸ��5-)�R��JT*Ky�������!�$�����>%�K�
����>+'/\1%d8�&4o�G>�s�SG�R����z�y����^,�Ǻ>��c��|�~���(�_�N�R`�7�P�X�mP�dB�h
A��S��?�@%��!�ar*i��8��@G�OEF��%X�.�6s�O������ ������}�*���^����N'p���c�29<'�	��yK�bFTB�IE������t\�x�0���|�*��G*�p���4�m��0�p@�p}��CT7�����5]��~�QR[w	$z��̈a�c@�#�猵�{>"�Oh��}� 1��_�{b�` a}��:~�m����D4zèAt�'�W0��.���U�a����=�����>%�,���Q0:���<X{Nٕi�@��v
=M㼁��Req���k��s�q���o��DU-�r��!����uy����t�&�����{�Jd-��y�\�faW���*�M�!�]��$˫1\D!�r[�$����3��ɓ���=n��z�yBPPϿ��Y��v�����K�<'�.����bY�IN7;��,��U/B�D4H|�Y{l�igu@���e�(wZE|8x(�ή�]^�`��s���� ������d��a�:55:6%-�$U��ݑ�#G����*PG���	tEg@�ʹ*j4=�����8���qƣ�ys ��V�'04b(9Dc�`��O,�{>I�<#[��Y�
j�K���C����ɓ�'��_�Y5F�8q�J�H�@}A��.F���۸�FLo�/�A_=x�:s�f�
׌�f��Y}3���#�����P���(t�{�#��8�g�����2��\�����d<s�T��Ԩl�p��R1�:�4�b���(�k�C3S�P	���
���4 >��6"��]�J�cE�6�!�.s����c�0P�f2a�X*L�)Y�BC
������T���S�M�#0L�0�l�p�ib�0�A%GE�9cI!=��`��j�����a�y?2�ke��4<x�ҩ�H��1�c���z�xF�G�)����%vP��l��'S�HH�Cb�#)��~��3aF^���Խ�(��8p�i�wR�!�?���i��z�cI�|D��T걤Q�K;��NIEƄ�W�Vf:�j���-k1
�	��&p�@)�eU>;}�S����u"�L��W�/�@�����&����9rx�� .�ZTk�&��,�Ϝ�J�&���ߒ�9���H���tP���+�+���?`B!Q�N]�yF�R*�j���8�{j;�� ̛��7nN�+q<|������Y��xS�f�� �aGC�X�e��
�B�d����U��ڐ箜�F4�ӯ�*��3�.���#2б,�Rm뇋�_.!D=�c��ʧ~�c�<W���/�"�p��llޔ��9}�����lC��*�R%U+��Q����J5��)�|�'+�|蘔�٪p�����!����B��ݦ�G:�U4����+r���~����kWl�;q�lo�µ5�&rg{˺�A��$�):0K=��ɖ�5�:� ��3�mn���is+'RC�LelPLP��hO��gzCc����d(��DH
�� ���$#����zC��!�~��4 <jz����r5���<�#�D0���s�<9P��!���;�6�>�m�è@�� #Q��O��i���FWX�@ϓs��kY�g.��@��c �}X.����Ȩ���4�8��*d��y\a��r�����{`�k�F���uF]�+ehdq�p�3Lð���߬�`؞�<�ǚ��d2���ݨ|���0�>pm���^}�+f$�|�>����ڟʴ����V
�i!S�0t��^��K���s�q佼�Y�� <b�{$�����ò�ޔ���/�͛�J�����ݲ\_ݒ5
͝��wU���V��B5A>�Y�Q�y .1��{ �(��ԪG�3`)6��j�����X}��/���4Ԟw�=�z�iн�x���k��d��w�X��B����.�G�ʅ��Rj,JO��ܵj�r���;z�9�d6�X҈�v?2�`
��%>�c���\X�q�X�u:NQ/�uc��VP��TÅK���LY^y����~Tʺ^�5�f�?�qy��3r��We�R�
f���-�6����iE~�COIww"o�|S���dyiA���+RH��ܲ�|�!6�{�:~i�3��5�Pdiy�,| p,4��V~�1nv ݗ+�2;��q��t��R���_�/����G�ӱ_��_M�<��zS.]X����{Nnn5%_�ˏ��G��o��%���䭓��3�U���c�n�wy���&�w*2�Co�lMᾱ�����>?�a�V���}�|'�A���8~���9ư&��bH�����5���d2��H�,�\���J�X����I�A$6=?z���e�r��W(i|
<9Koy��!�yn�9���V��`�V�76i�ܱ���AC�V�1�5�ѱi����R[��=蘻u�8o�3v���-����R1��k�)��/;�Qo�D묘fф�k��@�K�V(;�;Y4�L~{㍨�����z,W�X9�Ů݋3�J�H�1	>�9k����sQ�$DXE��*w<�(0�h2b��+;��t�N���}z/�s�뜿|-34.��n+:���ྡྷ$��:}�Do��m��(�N�B2J"�؀P�b�r^�L\Ո�!�Z�H�T�:��v��><��b�93;�3U�8g]�_����Ηͻϡ�]�7.T���2�p@���{ݖ�S���GV2�h 3��R�UU��f��? UG�Otc��I�{��%�ڒ���,��U��,�ɭ�X6o������ؖ�����z�'`gkH<(ʰ�Jsԑ�Cw�9Q&56�WS�]����2��H�:�xb}���Nlñ���������QRS���w�z�đw�f���f@��+����7�ȓ��r�.y��9���_~�_��������37ըiɂ*�B�(�����Jg(2��w{K�'�F�(��=�\cIn^ZU�eF���:����T�����|�'>!7nm���W�ݏ=)�.\��j�i�L��e9r�N�LH�gG�Ks�,�8ƻ��ſ+_���B����ܐ��ȏ���}��q*KwGǪ�X��R�ycF��@䓟����?>i�R�b��z	u�-���U�_�z�<�K�����K���ڪ=S������/:�q2[ב�D6h�J�:,;�WCjXE�7ڮm�#
��k0�u��ǁ�%���ʒ��ng��ַS��I� ?TI��g�L�
cC�a�p甏�Ϲ���\�A�EGEb�� �(����,*S*%�e c���$�����u����+z�T�@a��Q
��أ����`�]�p�>�qA����XNw}�ke��Փ�j��SO=�N�-}�U{n�Ռ7Nы,�(�R��9Y�`N�����S��L�ݱ��)��aGH��gǚ�gd�"�Ô�"i�팕|Z��B�"�R�8�5gg���ow0�rf��Y�0:���[��_}P6�½����4Fi��h$~�1����aDíO�/cӽ�:2ā�R���"�Vu�:�o�q{)�<$$^�xzQ����na��r�9�_���ueF*�`�/-�ZS��#WG�?ri�j�i{�¥V��L,���Q:��s��Uf���,�����lB���S����=E��«�"�`~An���P!�W��N����Gx��5Z�/�ح>c=�.ؚ*�@u���C�H:� &����(]3� ywz��Ã�?b[`x���~����4Q#*��6vk9X�^��B�V�[����Iʹ�����s?�I)��3k��/���J��ll놕�zFGe��:������7���]�^M��}K֯_U8���«�;�U����e�5������wk�
\����YTT��fB����/�'�W_}M^x��|��/HefQ�������9����O����_�e����Ͽ�]�;r�<������3��������qD�ܸ!�g�ٳW������/�"���)tx�Ǐ�Ȩ�6��,̡zE�-�j��hGe��]�{�G�5D�%+��4�yrT��sS��`m;�F"��IS���瞖,V�Ҳ�M27J�6��C>q��\Y��C�WLϔyNzS��{����;��x}F�X
Eb*~����=*e^3�0� HC$?��HnX&�g�k�Ջte�����Ò:�o��P��ر���K3�"��7RCx&(B����ds#ҭ�D�J�팛$�aą���q�ݦD��\4��!�4��3��R3�r8�ZJ�zpsN}��'A����V��G��,�!S�e����f�#���ĚV����{��m�Ї�=I�x:��V4]l�cچ�u�P0���H�
[��`R��a�B��!x,���-��dai��ES��(����hB�W%]�E=Ra�Eg0,��ղ�	O,/oV,�$���H=�~Z��W�T�5�ׅ\�]�!B_XX��Ջ+�ݞq�����Z�}����2+�us"_����{���g��gO<>ò}��pƌS�bﹺ|����Qj���ac㠆��\I<q�sz�q��p�4Cbnv�ʺ��y,/�䍓g�s����?�����z\V����U��_����w�'��}TΨw���s�籾Ց_��o�bY�G�}��������YYTo~aaN"�`.ݸ�J��Y���5�^�-����h���#wHO���"Wol���u�+�����~�V�Z�����؃�ʋo������<����8(���[��3�uc[������^|E�:/��Y����ߐ��&O�}��d�Q�ϏeN7�Ճj���m�Ns͔��S��~��2*�p�����6�I�H��܄B&$
��Z��F=���*�(�6^#�&���v�Fa8�S �/�����gX&GϞaV~��	4��2g T���� �iHX3E�c톀+������g隠 �OE��?@�|����$�CF	��p�q��ѻ��jQ;O�K� ������O]�t�����7D$q>v���/����9~(r��	Z�A���N&C_^Ȟ#T���yB�5�k8�a�?����זK��2����/���D�c�p�X��@H�Ź��0�0?�ޭ�S2�j�N.v{�=���S�o?�t�W�J�O�O&��/��,�~��� ��ys����rQn� ���N�zŨ3F�>��<�ć:��k2b����[��eZ��mȱ}��<,Rx����峒td�º_��(����_����
�JUnm^�J��JX�8a�5t�`�ZX�Oݸ�q��f_�I�<�4Q�W��:�BQ�;r(���;�U���/ب~��[⊤�pu��9"�SOx���Q��Br.L�(as(���	���t�-���:V\6/���U����|I�����|�ߒo�y�]O��k��ȏ˱{��j@��\۔^sG��|�����릟��j�U��U������EN���k�T��+W�����&2<}I�7��*�r����}�.����m�X,>l5�(7;x����ɋrqu]v�H\P�=I�2��ʫ'O��ѣ�������▼�k�%G/�xؑře�����ֆE��AGV�g�{�g�����!�s�3����:C�,�
k��-�>|��S�-��8C�Q�!���)���a�R&���(��qPq���=��Q!g|h��`�*`
�0���h��L�z�q�cZ�%y��{"Ush�г�ӆ|N^�
s�}X]@�W6�V�� Ri3=A*_$��ox߷t}2�l�1������)�*y�i�А��*��܅8�5�q�wh�G�Ǘs�REIf|p��>�|�D�+�n��a8�f��@!��k��aF�؍C�_cS+[W���7�������GEn+����l�"2�Á��=s�����Q#�[Χ*\��w=*���W��5��׾�@e�� ���0O]>�U�W0�&
�[kb^i�y�����Ps[jZ�>z��{���hh	����8�]��*e����-����*�+���z���h����̡��t�SW0HP��h�g�������Tu
6.6�z�9�k�AI�%X�����K1������Pq�\�z�=z�~{�G_�x�V1��.��¢�^�^\:���<�ݗM�� �_8 ����v�/s�Ey����zk����(�e��%��HTg�׬?��\M�r �Wd��Br�!7�GqK�˥Ʀ����4��Q"K�N��K�1�R����f%��޼���iI��A�i����,��#�S9��몜rx�yJ3K��ܕ�g�y��1]�}}����[�h�0 QŇ?�!������w��^x�¢��ԛ�R x�FT(N�_����r�̽��'
ܐ����;����"zI.G�τ&iLI C!Ǽ+	z��wo�[Z�����?�9�ܹ�Tݚ�J�b�
�`��-hFE��	��V�M�ml�ډ0(("*(��EQ5Q㭺ù��y���߻���o�ϩ���t�q��>���7��]�r��
�Xk^��s��n%��ސg1�]�E��If��8,G�#��`������ñ(�-ޫ{�>�xt�J-]��u6 AIU���PP|ifl���ƜG
�](t����7y̑&�c^}\��re�k�8N����3/b�`�5���$766�q̕g1���M����e�iyh��a��q���7pp�04=���;�{ѐ����r"_� ��ge����:f��}?��ף]�E4��5U�kW����=N�a9ƸG�X�r���h�k�ic�nm.�ɓ����C��
�����c�=.k�]�x#�o�(\�؅Ҳ8���@��	���/8t�
J�D�}��T��k��#Ʊ�abQ ���{�1�Jf(�]�XUa��ϼG���'��V���|�o�,}�����R�0"ʽT�IM��� ��VER�@�j  ��OLp�g�
߬�@$�!�yzы/�LP��-0>e�X�ঀFVOyر�h�8����$�9��r� �յ�9pP�̳7��g���.��G��ӏJ���jX��9���'ͱi���j�|��lH��~<�x|ĺ�A��(�s\�P�C����M�djfRM��ue���z7=(f�D��xB&'fU���8�d��4�ŋ�eciK�W�g8���ʅs�lӊ�<\�/�D}\�׷%�bx�4�u�S���w<!�����������ʓO��gr��r��i�UG��� @����]I=��Ɓ^�0wZUz8��)�(;gQQ[�u*����p���"6ç���q�^�{�N.�^�߫�����xn���¸��=?�����"A�?�{�.C|l<�o��0^����W�\�߯[TfD�olQ쯎�^d�rs�s��A��H�y��.L1`��B����K� |�<��q�p/��E�^����tD1R��XY�s���M����2H��؉�:/�.��ދk�g��^�Yd(t���#`��aJv}���Cu�{��G����<̟�h�����@�#N��]ѓ��������7!Q�����%�ӓSrp?�r����G�����\h""K[:���;�1�q �p³Fa���i��&,I6)��/]L��>!Gx
kvT�ɱ�l�-���3��c�O��������yTz�z���^vg@�elb��+ڄ�\F�Z�|��J�;���C��}U��ǣ�l�J(9�+9�(L�]K�d���$
�X��0�������,�����a�٭��g���O�v�� TGȣ^y�Pq]Ω�LUI�O����sv�	晫���'�й�H�(�ŭet���Ͷ,,�Qe:-s����gXLm�l�̯�d���Wy7�������� ����W�`�齏��RmD���`aK�������F	����� ��X���MVIT�PXYl����@�&��;�����jԓ�W�K��o��j��ڑ� l�75tC.���ρڥ"�<�r̞t/c��n x�ׁ@ED��z]���.�����u?�{�8��T�p+��?33������J�W��¸��?���"�X��;��Q�E�����>o����d��9o�" aqϴ�GDre�
���M1��>!��cRF������w�M�T�~N�=`��F��.d��"�{��n�C1�쯹'�a{�@�X����r��c;�;���X������o��^��eyn�9z�s�<�O�R�5�<#{>p��0�K�����v����B�P��ڣ�a�ۅ-�'q����%L��3�`�q�F�۔oet2�ΰh{���_�/�m��m�裏���E���,�5M��םl&vtl��B]aJ�U��9���0m1�T� ���Ar�v�n��Zƀڗ>J��LWorm�'���[�����ٔ����X�6 �G�Z6�O5� �%CC�e	ƴA[�V7��IJI�ʦ3 �@�8�QR
�-n.����ĉ�l��0e��xB�N!EbM�wL��Qg��ڐ��s���C*[���r*�t����k�(m�ducU�Ty.m��2o��D]�k\�ԓ>sw�{�,=�>x�tt�-��ޜ��B�}L(��v����*��C�,YiNα
@D��"���P�"G|B���⒜b]���?++�.JoM�$����o�B�T�>� 5ָ.�]��+�s�/��̄�P��A���^:/��{��N����6+P3?�u2�5� ���ҋ��yу�lA���5����b�����8/:zA(:�w �{�`���)=��u�N+�ݿ�
��Mε��ߍW
Eo܍�̈)(�b��"0�=�"j�,� �����@/���c�,�N���pC��������}�*���Jw��F�3�qSDi���(���{�G.k��}m����b�`o���'��+F��)W�������`νϼ���9�u�mu�i���������G�2���jw��{��n'{�"�����h���#�����ƙ2��g��?GZ��G����4Ԋ�d�6!k�-vA+��-exS2<>�>{]0���Ui�u��r�m_�@��6���i	eV�iI�	�<g�ڨ�9�B�y�)��*\���&�B�q)(�;�C,
$@��Ӭ�F�P���O�t����8�`��P&J���k�H-�F�f�g�{�Rc�ʅ�d�����7�e���,a����aA����p ``B&�Ee�����#�	���6_��a jF��X���C���&�0��,V�����@�/������r���W����NcJ6{��(Y��G��;t@���YS}fἴ��-HU����!g�^ 5� �+�����I,,�.�B��(xL	=�R�$}�����`���O���/�^���[����j$���CM8(d����>� �/�U�=G��#YYG_�2�/��8���Й�:pX��1��dr�<��W%��r`Q�[��+�Pq��ȱ3?m��b(�o�Q88����l�v�֫�y^�B�Cp�n�ő�k[9?��*��t��AbV5�(lQ�����Ѭ��C̑\�x����y���m�[�Z#�Y3N,�õ��� 7`��U�j熘�w��C�<��6�r`b_�u��*���7�B\�={�B�灡���^��Qo���N�륈��1t/�Ah�p���g�QTv�!��9�/_�C ��U$�
k��t1҂��r��2�&�ÍO�5_��R�w���� qO���8o���{)7b�5.�G������p���M%��,Å%34T���.�2�ȥ+f�t�v�A�C���
Rl#]8�{�'�~��&)�j7Di_AU�f�k��Rң�� �`��wV�nx�X��,)��+McW$�?N��~wD#z�Q,�� o� 6"@!m	VVBE�#Jl*b���@^�J��g �	b�j��U��٨�Z��z4T�@/m�k����}������₴[���oy������E^�����{ Qg$Z��L���'V�O�V�N�{g��(���4�L8�B�M��7����e�@b��O���u� �/��\S��r�5ϕ���4�21>��ū�g�C�NZ:�Kg�ek��,/m���<�י�������9���:�_B����z&f�����I�j��ͩB`�t����ȁ�t.����k^U�E��aW֗�n8!o���j ��~��djr�����N��ܼ��*�ğ|RT�<QnJk�z�B-�z�k[k2����Ǥ��+�URe��\�s�����'�k�k���ԃ �Ɂ��U���׻�y�N/��V�.���)6�`�m�_�u��=�^0 8Ax9�禍�<ʔ �����i��A�)��V#�S�1�z��+Q�������Nh!��TWnΊ�J�ñE���:����y],�J�4C�=k�����C�P�<O7P�lxd��al�6��ͯ�s���ϽiJ1/�!�"=��{ӗ"[��1�Ɓ�x<U��������{9���'<4_��`�|��n�Pn����(\8�����O���XG�����{0�p~�o�)Ϯ2R��|��:��S����d�y�P����ޅi󫋗&ݝF<�G�*��6�.��SRR!ߌ��TxE!��S�|`�z�m�y��G���S����z�VWnw*8(v��%i?�s!��R�w%��z)�A�_(v�cr����7z(u�w]QO0V/��R� �uy�5iT����ũ?"�*�`C=�~{M�-�nV�V��c= �Ճ2��k��i��/�#��mOQ;ohL-��:��3�p|��9/B�_Q���z�Bc5��6��I&�jT��jD�*ֱ��D&k��OU�;���d{g�h��6�<��Wdv���K=U�ωZI�*<�y�Y��6�Y7�t�]��0'��i��0i[� �Yt�J������C�fM?V5U���Z���M�p�9<)��U�WDV�wdr-VՋ��䑇� o���sea�aU�+2=yP���IWZk�szB�C,�뗘kGh>f���Z�%]�b\�k��uB�{��=L/CBn	A�@���N��%BPHŲ�e^&�Q�$S�.���Á�A@ȹ����������k��DU˼!z�(Mr#�S¹h���π�J��kg�&|��c�Y�Ӻu�FCz�xV{~C�Ë����<���F�ZX�^�0S�n� �ޯ+$W|S�+�#�K�\	S�+N�o�VGY����V��?:�|D5�w)Z_?9��v<����!��J)M%3� p��[��=|�%p�����8rE��ׁ{��ׄE�������>�G:���jr��#/����YL�!�W!89�2"w��r
���aF"� L�B]}��E��
��Z�x<�m-�@��#M	��%����u:���?3Q.�j�R�T%	���Q�q28w�R4��Q4��|���t�F3�Ի��X<5Y�&/m,GC�\��U�Ywvz���u���!j�ި
W�GVo<���9d��hJ�#�1�q �@��
=�#�R�1��(qT�2��øo�����+U�T7 ��WRz���\IZ1`�TT��7'7<�.�{��`mrEFy��96�H�Zb�j����j�ڇr�ퟗ�3�Y��ݗ�3K�Q-�!���իF8(*U��G�T���=��C^ �	K�҇�9���
�-�A7b�ϡ���5=oc��~�rJ� ֗���d�L�
���*ן������{�=���[H7|�.۫r��URkJC���am~jFV�6�a
v<��A���§	�#q����B�`2p���UWC����!}��C�riAf&�����*��|�M�ikc�FۄzzK��X۾��³?���ԫ�m�@�R�֎�\�H����>�
G�����)�kH{ԫ�LA����A��M��u=����4xY��Zv�e�޷:�B�8/~�X(�Z]�p���e���.����k�V��wՀw�[�=�<��w�(���7����zq��1~0@ �9h�d]�C�˯pnS@ә+����u�^��d{nߍ#�`���3�ge�1������pI�sB�9���źq&ż�߃Gf�)r0�+{��\zD�H��qnx`�<�eda�{/��Q����=uRLx䢘)����Ϗ�A�?�3��g:���"WX?�p;k#��	V���:ZT�W�B��r�E�NG�OI�M���M���v[����F}�k��U�cC���(�!K�iX�!3"G��{U��I�7w��=;��������^{_���	������u�m�H'1�Te���0`"ƨ��z�.*�垪݈�-�S��4 #��؈���%/w��A 0�5\�z���B/ð�&� ��(�Z�k��������䃍��cd�`y��xF�l]�Z�Ѝ<h�x!B�ҡl//�+�?�禛,6�|�J2�B�)J�XG_&n /e�m2p]�cB����i@�y0�H5�����Vé��}�)���Ŏя��\��}Ӫ�k������7JMixb[�r痾�M���6��XE��Z�u�t�1i��i��҅���c�!N�c8��yoaU��R'�Yuv<���Ғ�zI�XI�̏�sĲ��IIW��%��g����}��_��!c��EJ����@i8�[�Miw!��r��IV$DC�����YC�!r�H=���4�M&)"]H���B�������IM%�D8"�j�Ig��܏zxm]�h�[�f�A�Bh;Ry>��=��M��^�<Ȕ���)4�=(nx:�����y�{9���zワR؍�r2%5�ʾ,u`���9(|g=s�W���{���U�{v�;~��"�vp י!p�V�x�<ރ�Dۼ\���6�����ZW�n�I~<��J�z�[x�ָV�vo��O���E,����#U��ѡ����%�Q{�`[�*eB�7g�s� ~zY�q��gQ�b#W�n(a<��k��uo����SO'���e�t#�=sD��\^�� R�z$�s���8O�PY�	��b_u?/@�n(���)LJ�p�LC���U���[j3T��OSٚ.��3g�Ձy����[t�N�O�t(�����	q^-U���(}ťKKw������?��?�[]����Ss��	�����W�C��X�:Yu�4T#i��2��*�u������H�^�d'^2���,4!a&6b]2�>]h{Z
)hz�Qb 	�,��^m�'�HWC�g9G��#�ߓp��X���]+��zA���a䩤�dGKѐ".1�r�6H�ԛ}(��Z���u����HgsGJjL��N5�~(x�X��Л�q>�R�q�Sy������ok�[�f�<0V#��f�9�Ǻ.qUN�*p{U�-��6dnfRZ���W%�0��G�?'���Y���3i*����?=5!��y�>vJ�<|@�^Z��ￃu���iY:N�g��-�� i��[�1FX��HF�6ij�S2���7ƽ���4)�@���A#������:hzwV�Wɥᖼ�%/��z�	�z��G(0���[��7U�[]1���'���m�GFG��˟;�_VT9=�ȣj��JmlJ�z�j�5*`�Q�F cC!�
ͅ���<#�IF�NCVP^W$��k�7�\�"�o�uϩoomgF�^� ��|���-\��������s
8ɽݩu�B�Χ�@:7N����w5 $���Q�l[�}���V8��Vίn!�Q��\ā�'&ǲ6��u�u7�U��=j�s�
И��,�����Ȁcn�`�9AMƳhE���xs�kY�+<΍s�SW�.��y�Y#O�x�q��q�:p��u�` <��üW¾�������t��wߝ�݈s��tT�ü���� s�2��u�T���W��:�Ѡ،,(tth[Z�d5�u]�*��#��eFZJZoɉ>���_Z��>������_�{4Ln�=�
5.���n�`�o&<��y4���G_���!U�zS��NdS�r��ÜHtD"%�
�a!|��+����Y���:IJ�4�i��j�B#�q�Gi�Qc���P�q�$�{�}�&rZG�3�nVw��߱q�[�;��#*�N{�!w����þ��Cg1TX���R��[���� ����F�w��R�^_�ז��,�}��Ժ���>�4X�T���T��t���ڐ�Ld^���A sj�%��"gTU�vB=�I՟�** \T���lo^T���ϮC���ϼ���|��a��p�y^t[8w�B1e{�1I��d��C2=��ų��,��lS�THo��xק�9�ip�Q���2+b��g��l�r��?A=ÀJ0�!�,˄�_(RPĪ�]��9:7.[k�277+o}�-r��Q9~�J6��h2�2=3�e211%�.���������[�ron(k�[rq�9r%����!�87\uL��Ve����G��ʠ�#�a�%�媅�Ϝ}B/-gJ�ޏz~'O��uU�~����k����V�44N��R^���0q7� ��C�@�"8�
4�	lĆn_�� 8�i8d���~����<�n!����:3
B����%�Kz�G8��n��f���E��p��e�-��gtĵ�bO�:%�~��3T�<��4*�Ν�9����|�7�\}��y�ZyW���0��=��#w�q�.e�
��`�ܯ+:XKS`~p_�җ8��T���qg�����$�43d�����T����x���z�[�"ǎ���D3��$���7~�7�q���Ǐ����v��޴C�G=��W~�W8��v�^4�;��N�+G�܍F��w�ō����}��t��C���gʻ���P���������o{��2P�K�{�G�GY�D��ds5R���|�����h��q�
����i�%zj����4y�;sK��N�����Ǆ�{�-��xpt:����B�&U�����U �T�O0��o���ty���Y���7S�VJ̳�'B~xo\p��N6L�3�6d-vh���Ήӛ�n�FQ�R����м�l>P��V��Y)5Բ�B����]���q����e��U�5��[;%�U��4����Vx�)�|+�K��L%:VP�%���u�Y�o}��X삦�� �4���Th%4�c�:��{ý��a3�� �:��>OW�Y���©]U���m�𞞗�N=[N�����~��*9�����1�ssR�����
����B�:y���r���IU��ɱ�4'З{Y&j����c2b�[��<eZ��rI���}Z�C���5u���1FF�2�uz\��ι����U��+��]o�#G��SW���՘���6ט_{�K_�Ȋ�wZr��S2P��z:g�8M����nW�`^ϋ�8��e�t��2UW�G�X�O{��J�M���>�9�S�s������0���j���6���iS �[�%���ۼ�~�^(-��Q���~�_H_P�E��^��ڔC� 0�2����=T��;poJ���Y����h�A��D�����y��Gآ�.�eV^Q	�ȏ�����y����,�E��w����3��Ͼ򕯔_��_`TG��۽,���#r���`��G#k������-�"�z׏�x�g^�{����L蓟���uǝvu��(��o�E^��W˦�Ihr��tNa��u��:f�z�����Q��LB.����7��^���s��t-S�Q�����W�bu��v�<����^Fc���wޢ��O�� �����ȃ>ȲF���<5V��=�y��n"�l��nߺ�sn�����?0"�몯f8
�$��\}�ƚ��-2)|?qk:� o������Uم���zֳ���~Y^]a�
�x`�g8��xu�5��b�� �Ĕ�g�<R+��_�W�(�e21`���t�Z�y���QKߟ�+�8��	%j#���	���O>C��#�����ۈ�(If#͛�<�pҮot�6
��^������ظ|�Q�8����:Ґ�-���Ӟ���ek�4:1"��*��9E!O���6�*��N©�*6Tϫ�YN�csk$α�F8=����z���j!���f3ĩ[�"��Pxb��NX���!��ў1�W��M39�*���P�H)X�C0 �AISd�2^��A}nP,G��z5c��-#g<
y|D$Z�yZ�BIv���^�B��'�cc�.֐�A3T	 �%=�P�5l�Ko���$�>S�h�M
��s�r�+_.�z����
�F3x-�,�鵟'N�`�g����&Ir`xm��X�)���o���P����R�}2�
,x���.��1ѕ��;��:�m���Κ����C��-���?J����GU����u_YZkK�t7dL���_�y�k��<��U��9z&EJ��ّ��5�WC�P�zpsS*<��^�^������gے�G�ȹ��R�����u�2M�616��&�^s�xn�/3j�P����,y��@�������3��N^������"���A����?�C�}6�pF3�>�k��L#g�+�&�p���Զ�~�]��V�u���I_y��.n�vt�N�gU�9V!��IȔ��5���FҸ���7Vj�4���Ս��@��g��<���{�P~���\3�+�{�W���˪ ��j�Pq�pj��ӏ��xϽ$g�����D־�ϫ��bcx�0�����1zx��a��!�JI��P��>����� ���^���Pc�d��%���;��0�`�yn���fy��Sǭ�y�8��i����3� ~:Ҝ)-��#�)��{����&�:O��t8�#pD�׿���屇fo�^ې�ztf7�7�LtO�ļ��C���|�>$��s�#md�� �BE��ڪ�[䵘�1XYYf��\�z�������ю>�T�ų��r��~��HV[�UU�� �¡���կ1
٬�)#G}D&��ن� ���K�O��b�l��x���u��Y��%����%����?q�����K�ݡ^�y�c�yC�<qF��rq�T0D����s=�A��O�B_^^�8�p!�V���L�[��<�$�9;@K/:;��.��k:�FN�GO8�t@��6@qq�3��CƱ{0�A��/#6�ӂ'pFz��=GN����A�����
X��aA6Y��
���=��`�ݢ���x�B#�о��`S��Jk{��;�a��4�'th�Ȑ���		`��B�5�S�Z� �`V��G��˺=a�����C5U�c�)��U v��+�7�Bn��7��Uy�?is��oxQ���J �q=�pI}�1y�G���(G�?���Ի���Y��c98=.g�<���+�21���6-U�o����_zL��Ⱦ�}�+��7T)_���7�^����HE�W��"�'��=�9�=��I5(vZJ�!��_�,���P�m��1��l�Ѕ'	/!�;�S��)+����WO��0q��	���?o�*������i9��9��W��n�l�`��_��,'���Jv�1��*���^��y��'D����J	�n|��-�>���˙b8�}�{��>�O��	���b�$P"�E.�����w�}�#�o��dm}�Q/����@	�L�z(~�_��2������{��#e�g$Ld�������<�������� �����˿�G?Cz�� 	�s�Y������������@=��(�\Tcl]=S������8�?���( �4�J��{�-����ϝs����ٳ�����۾�C�W
��0�ʋ�z�+:���1][˗t��70�ʈ���4,�P
�?� ",Lp!�BD:���[��H��Q�Ȱ4�Ȁ�@�#����jo=5�;��&&'�v��и��#�<���W]�3`5�%(Ws�*��"�p{�f�4���c���ӏ?ɵ��v�� ��Qʇt��z3@|Z�����׾�55(O�<�Ci�>�F����3��b��7f��uLi��t\��$Wʘ5����!F���U�:��5���~Zz�Ӊ;�N�6�+�����ʇK��K�%&�N�w�3��Q+ge��!�R��Bd�x�y�(������f��w,@,����Sn�uԂ+%v{�߯��%��C<���BOn}��:G�~��[^1׽FI1����1MC��4c�����P��D��}�&V` Eu�Ȣ��kE^xn�!����,���TX�~�Z_���|���I���k��� �JQ�_#�~��u�1(&o� ��J�VO��z���(���OS���m������,���p/,���Ӳ��#�k#ٷ��Jz�
���p�nV����NU��\ghxnnB.�;'��������T��$�u���;4<��a����H���{ks���@<I@)#��	�
9E�����~�>����(v|~jr��SW��>�W,���I]�S*�,�ܖ�3D��jk�ʽb5֘K����hy��?���(ez�q�hRD��nxA34^�'qiqI�����YU�[�I��2�8z��3�� �uc�D��J�x�a�9��w�#� �;���7^�w\g>�L9�V�x}emM�\����9��mD�h�Z)��yuDF��J�7�At�¥�\CŒ) aP����W���Zj���!��M�4m��qx��2�c���Q���!k�11�E�N?y6�W�Zߐ�y��s]6[;F��Փ�5C�7��iI/����� �HS�K�z��(:�!���X���Z�������uY\^�_#� �p�M�ΝCO���� p��6YKo�i9���Z.�U�71?PZ*�Ѿ�e�%���L�� '�!a\`ȌP92й�9C��x��I�(`�"�x^b �f� Պ�L�@b��u�P��V(�Ú�}l���.x@���I4���!����V;����R*��0�յ O}[�aM�`}��P��� �Cj��ԅ�-i���Q1�<$BJN��F����B��Ӫ�+�F�1�H@M�����rlPTR�u��#Z7������шE�dG��i�j�73�\\�w����|:ʕ������w�CuKe�݅��!B��\AI��������a���~��s{.GO?q���:�S ��j��НP�����n��a�A}`M��o
=��ɷ�Û����r�����꜏�GU��(G^�a/	�5�f��f�.��7���Ex�bEX��'ev� Ü��M��n��2=�_F�W�?�Ct���㏝�����lI7�yZ�/~����{����7�HP67T᩻�h�h���\l}�e��z��rP��@Hri�����p�����j�C�0$B�-���)�����4��SW��z��KK�D�{�����h�&��[Y��AB�G#B�y6���1d�B�4� T��	�״�11<�e��LF�(6�a��{Mh[�]G�XL�����]W��"24�����Π��>"���c4������A(�9���a�uU��NYT��|�����*)��,��v����ň.\=��a2������[ɓ92(j�T���t~z��.��T=���q��y�>���gg�aX���w@f	���y�� ��=z�P����0�2��j��#a����h!49����|�#1�Sv-4C%��J��`�AHK5sC��vw%;1ah��z�;-�ܢ%%��gc*o0 ���@� a�.�y��+�����B���P�'*��n��]đ�%�z>�Lƹ1^����6I W+�
{J�N��=�B�}���)���_�$�s�a�GzRQ����i���#i�-���4$ ~��yхQ?�vN�{@��I��9�\7�U
^��^���|#�k��<��*�d ,��$��?�]�#�]�4
�b����R�&0_���΍�<��B����ޅ�u�39b/Fv_Gq�U����k9�K(A����8�F�;���xB�߁T�U	%`�H���y��z;*���W��n��dY�^hG�..���������[�.^�ݴӬ=/��Nӧ>G>��CJ����PW~n&����,D:�{���7�T��b��J�D�kSR/˺z4���+r��U�����ΜWoeBΟR��O�?&���������Vy��S�(U	I)x�)�H�*%�,ꂔ�x��V��#�3�g��0��)4�л�zիdrb���Kz�������h�$1�~�1
�����
�Z#��Ԝ!�'f�����7�U: i�)�K�Dhu��W�(R���Paưg1�<qTz�W��� u�U2�Xfi <�a�$�ı@ G����34������[��^
�-~#�*"ނ������F9'�$�̥*�/^*�k# ����B��w�<��ܐn��OC>��a��(�S��X�2��0��V��[b,ߛ��F�fJQ`�[��賣�R�l�S��U��u�ٿ���:�g�/�^h04\"K^B�oct��ֺ3,����B�#�q�հJC���N;��ԋs�*���}�TM���W׹��[�ю��4P�"R1Ji�C^�`��s6�WT�bS��˫������A�{C���!��en� �G���ٮas�Yj�;�׎� �>V�x�D�6?Ñ�aAnc߂��$*cB٣9c w��
kvR�����GHSV٭Jg��<���(SK�+�$�>`��|�Z.�sp&�fu����]��M�����J�!�<�<
5��,$E��
��U^N1>f��-��jXq�"�=����`�4����F3�`���Xk��.%ði\ѧ��w�\��5W̱�S���o�ߤ/�r⛢�a��n/�lpd�d9I �M��-`��p�``�u��E�ޒ�*��*�Q%�3D�no�HK��_�*y�[�,c*�W�V�ء�l,��Jlfj��noڠ�������{&W��mԪ�H���Pm\�.ɝ��-'�<"O�='#��z��L�g~xnL.^\�����w˱+�b�9��}�j��m�x�<��A���!��������Ol���>�U@S.�ݾ����2/6��½�c�ޓ1�u��馛�ڧ��/�'���m��vNkY�T�O���x�u<C�'x	��P��򏥒�YW�W�v��@ �r1�(�����	J3���ݯ.���yN_S$6*��IOK��� �0+���f��	Ld�����P���� <��)V� %�6�cǹ����^,��R�V��6���-=}>���|�����[F���0�a�X�_��|q��4�x6�!r�� ���Dx��y��+�!�
��4rt�s�q�$p� �x1T�n������ቹ٬֛8���r���(Wq�ץ�Q-�R?��'��0��N�00ּ9Ͼ�s�N����]���#(��ZT�ĭq�0���-.��� �aprP��)�[�3I��aP�!d�a��d��L�AX��#�����e_�X6����$��8���x}W�"ރa�(��Ç�`�b��[�`1"4Äi�f}Lr${�l�x;j�C�N+k�� z��ޭ�)�i8T��,1F){��%;'��w����>����B����[��a	Xd������Un�R��G��G�ye(�7�	@��Wٸ�������\��"�z
}�/��� u�%}�OfB��}讖0
��ـv1�爍�%�u�C�u�CMz����5a����A�H��j���ͯ�Y���oW�!e^9zw#l:;=�0��G�Xz�W�cY|�(v6={�N��6;3�B�*~��ǟx���y�	�x��J2?Ӕ��z���ޯ�k{S�f�c���>����zy�5Wɹ�ge��	ݐUY�tI�*��N:�(��7q ���D*��"Ж�.w�B��9�����2L�us�����t�}_�������BS�^�ߕ�<�c��[�8�ÉI�Q�� �F�B��	z�`Cԁ�̵�� V�
���W~0ʞ���	�C����zn��FV{l)/���s���3�Ye��zmL=u�"d�O�$���
qD���Zb��s�F�a֬�T��8��{#g_;Ŕ;&���)S�'���+���Ag�'�M�-ˑ�f����d����p��S:*kF��٩���b�� �\z�pp�;��{pP��|82)�3����~���F`W�V��c�c�{��Դ6���0���ؤ�X��<{�N6>t:"��4��e�`9|�k^�u���|^���IY$4�o����ە,�&�jF�ʩ������ʾR6}�|�am�gʲ>�1��;$<o���y`t��������u.�z�x�b�n��eH�����1��Ėi����T�@�����0s��j(TqV��?"��@ǡ� �7\����[V-s�f�؄Iu���&K���m;��MN?M
=���!f@a����F���	�{���@�kD�
ҁhN���w��m�{\���S߭`���F��+���LRŐ�������p��\X=k�Je^�����ƚ���T����ѕL1����W
$:D�Xݺ�]����<���|Cx4)�q5Y[�^Gn��j��x�4�%��'������衣�(���ϝ�W,��gv����t^=P�3g���Ǐ�[C~��cW���M��XUa�kO��u�D֗/���j	����]/���W��]N���v�Cp}��k��գN����6�5��r�d�B�G����GH�@q/-�X��H�.����3��0 m�y���	5bΐ���L�H%�m�����[�]~�gV��'>.���2e d���2TÚ������LF�b��@�����`J�6��O�>��͖��5!qjZ�����Qk}M�W�meu��7<cA,�n��Y_�����	b�2E���dc���7qJ|�� �!h<B)���Y�e(Q(�}���ב��)�*��Be�4U�XI��6vA�B�Ye:�B�"=%Mʐ���J��"	wP��{îa0\��S�{����Rh|��F��]�2䫆	�ph �Nh'���<���؋������{6��!��[P��.��H������գDmD�  ��IDAT�e�(�7�X�Ȉ�b���V��A�j��w�����{)��*[��$2*�z;{44Y�[.�o{W_�z.���F�q$AZ���>�0ti���^�ӓR��W]��`m�K�8�:F�ށl�z�O�p�E�O�} cAW�^���*�D��2ə�4�;RR͉q�o�e]dl�p@cF��f�g|bJ���z�K֤>u`�zZ�(���t�Y�Bbi:B�ّ�@3z�~��Y+<ω8 /��P�i�!ȎRx}����~�����5/2�C3�#؛�v#ď��`�ʻ.��ċ�q�"�������E�����һ���S
o�� @����4z���]zވ���myZ��4 �z�V�U�+I�*����o�^��hr㱫U��|C�b��"՚u*(f��s�P6r�7刐0}��Rh0�!Rh,O��8���e�x˼P��ēg�!�4�p����2;D�t۝��pI8�5��G��?~�[)P6�79�%d��,c����<�J����?��4�k��V�>BF*0[!��eY�M���u�ygC����_���P���Q��l��Q���+u���krc}�!�Z���1�j���<=����F~���*+ˋ���!�%l�T_Z7���КΚbB;~�b�x���0o�~펟՚5�`�M������rͅ�Y�W��-q�Qq�<��r7�"�F�ᠪ%RU� +�_ (n ��y#��x�h�2#��V u/bJ{kkC�:y���G^�X��7-7�����c�W��E��lR�s����������?# �mm뚏"k֢�E��ʧb�
@��ir��,L��:�#��6�����^O��C���bր?�����)�d�0�+U���P|B%IC�b)6`���� �[��G7�m��Y�R6YKi�ȝEt$�K�[[[␾LF��B�� յ;|_F;�<uH'"��(ň�-#'Dc�(��1�"d�����2���U)+�� �,�Q����}���5�	ekXǵ��%����84�ĦБ�	�،�G�* 5�*��鍤\�/���ld#�y6��W�D�����eg\c!��'yz��$Cb���ʛi�~��`��]9��~��W�^��*�w}Ə(�vAI�{C���fJ`7Y�^O��:��u�o{�`�|���qN����z����Ŏ�H-��UQ"�;
��S����rxC+��b�֒&*6;a/�u�vU!w���ݕ[^��r�s����e.��-7<����$� �촹Xz�!� �E��Çs�ͨP�L>�� �M�Oe�y����i>3�F14E9y�z\gX�c�w�%���Srõ��ӟ��Ǟ�f#�y�ur�5�S9�5�����kD7���2�_I��h�އz��r������Eb �}�7}���Mo�"��9>��q ?���*~���8����f%����Uqą������4Aw(��P%��3�.ʁ���W�ec��P6X�>c��$+��r�6�,70'��IF��r�8T�D.l�{-�4:�(b(�$���~@5��ރi�PO��$����|�$h�����)/D�kM"�=�?6>-�(��.�h)���>H�Z���ȡC2�lp�n��:����`�����ߒ����i[��֠"�X ��Ѝ��� 1A�����}�=,�^�>4��ABS�c�Q�0	�b�xL�k���"�V"���g�.��4T�����=�i��`i��Ȟ-��#�B&��,[j��H��P�q&�����k�y&B���;*��pfK�#���3�)�~�I32�H(��q��l�B�������ϜJ���vq6F�E���8ʝL2�\wzB�-(��YIq�4A��4ס�ES|	�@��a�.�OIz�˼��� ����Ss�r����}~�k�M�撁�lbM�=�H�=r�[�\Eao�<W�ç$�Õ���9q������
ݍ�R�u�e�P�È!)(�`y~��+��R�٘݁sṉĳ���y���:MU8��}ߧBN����~�7���},z��!D��^��.r���/��\���.Ꭱ`	U�i�a'0�w�r�)w����?��mZ�gΞg���+d{g��\;��w���r��(+�l�ǻ�q�am����9�veM�12��К#��jy�z�`���.�z����9h:i*TN8����%�e����<p�(E����s���\��bww����a>����}�}���'y�n����˪>��~��L�k���s��
�l@T��e���4~Cz*����H�4I Ñ����ӀOI虐�R��J#(�4(p��(�q�3?�P�6j�:�Li�1���(�Q/��d�%xa(����f�es+ԭ7dqiE�=&���^���j@�ҔMu4j��P�$һ��4�,�7G/1�w����N�M>�P�*�V��c�u�J������fQ�����r%����O�"�u�s%T�6Fyԓ��ؔ8���"*IG���D�n�W\��w�8�s)�3�a׶獃�`��֬6.��8���F�hWf��e�Do6Y�3lo���6'���Ӳ��0>5��vDG �s���ڧZ�_$�)v��!���@`qz)�1��V]Y;H��H(�G�8��¤�yE컬���W��{=�����y�^�܉j�x�����:���Сx؟82PH�	j*ۯ��pˆQ ��a�d�����	{��dB�'�C�@r����W�Ln��Y�p�����u[��#��B�x �pP�Ǐ�=����n�ǎ�-pPC�M�b��n��An�V4Ta�Ըb5�cr���~�G_���0�}�~�d�k�ʴr���Ry�7���ƾ�@q[�yr����̠8�����������>�;JJp-4w@c�sx�>����O�u�nǹQ�����c�Q�5�r6pX#��|�%35�G6��u�X������S�6�J?!��;�A~�[�(�c��*�B��E��IlL$V�Vn��o�[S"��r�w�v��p�Æ����� b���3��4�l^��Q�%��,~�2 �-��`���/[k�j�u�y/x�<��rם�˱�7J���wS����5��]h��)��vO�8>�a$+j =��?���=®���E�O�β1˵�����vL/r�Ǽa�蔳ȇ�!���"N���-���e��ę7�]�˗ot<UY�UP�YOuD½}��_��3*��!�_�ΗGy�]ϖy�������^+�WK�nCd׍�BT�h�܉+*���tk`��e��H�b<����.Zp>��8��9��T���������Ңk[-�������iS��L�6����kSZ�޺O������26;"n n��z��Z�4��*��Y�{��[�Q��sߛ'/���nn���)���:��׈���g3�=��d]����n ���F$�(�Y���`S����3dg��a��`@��߶�e4�H���B�x 
�t(�H��9N���]��I��Sʳ��.z�~��U��(k�����g�������R�!�3V!���<��<|�^���5��;2� s�s3�R��df�&�}�?�J�Bu;;���ú�@���U2e�uua���q �~�u�ˋ�����(S9��ƽBa�gZ��!U�h0����X�x?Ix2>�͌����\sJ���/����ij�k�u=2/��K���5Ը����VO�}�y��>��J�u��{����!C�ۺt�w�y����h`����4��k�$�X�_NY���o^z����I�����<L�|�MZ��AS)�	P�K�9.Ͽ����	�zdZN?qVZ;�����n��km|f�����V�7����e��������qAc�D#q�S�]�[� ��N�q�C����09�4(S�G4BT���)q>Eٴ+��
�_pE���`�]����}�|9���GN�b��aS&Oq���8��}�9H"�f�A/|�����z��<�T$�
9x���p��Z�D��`��ϙqG�?e�T��w�[}�#����bцy@t�iQ�@�(̴{�y�bNca��!���5(�"���;6�{��yv���9��%T�g�W�� ���H��ʽ��	�aw?�*u��-�������+t�/u����F��,|]���I��Ld}B�� �9.bx��xd��6�"�g���#�:��z(��3��?�w������1�@�e]�^��h�C]j o��c���޾�����ۣ����	p �C-9�=5ݔ�͋�� :W�ap��$^�v�<�ֆѭ�����W��w�����k?}�4;ݡ���7�͝z����RqlUžѬ�����~��	*D00��4'���>���!��Y)�,z�[�Q\�� [)��9X��^GD�6`��SI�y|��LB~;�U~�\�Ey��cI3-R����n�޼��0({���}l�?Q4v��F�� �?����xS*�I���A>��}3r�_"Ǯ�R���̻�_��������(�z�UדLLaS�3���c������e�B�(��f� ��<�+��/#ʢ�D�ॖ\&d"��3�F�{B��"{.7^~A��;*�QR��£�]��E�o�W��3�8!�޿�=Yڅ.��q�^���a��X3��M�C��O��e�)�k	����n�M�P���S�x�4OEѨ�!���+u2&�dC�T�6�R8��Es��x�r�Y�s����մet!,(�P��X
Y�\�|	k�iYW��@M���9��fD�n�|!�@�<�d� �.8����e�w�������w9�n'2\ 濈��k���,��B9�}�cEN���{�P�Hc�a���ވ�\�����O����r�"'Q��(�i������"ؠ���0��Xz�!�|��(��E��ɼ�	y��_N��*�W�@�#���9�� #[�L�b`(ָ6��������w�T��̲{X�{��5�#�9�V�-�@Ͳ��JP�����tQ��{�+G����7ȍ7>��͇CT�w*��c#(
���������O�����	y�k_ˆ!@�����4)�w�����%����`h8Y~������ �0Q>7=џHI \�0<�z e�K[	�S5��{�B����X{�Ϟ ���l��Y�yn��Ƭ�_/w�}G.��v��詊�=3���J>��s!-��X�H`hD�y]��/|Y�&�)�:���v뒜?�(��~����-U����;��Ӂ�l����K����| ��ĕB�w���a���xg�l@\��K�s��<Ȭh��@w4���7m��R��~9�}��\�o��X�w�Ã�/����c5�)SD�"ɰ;f)[��/����W�d?��B�%�]�/���QpJ0w%ȡQbys�����V���7�n��'a̔��*3*
kr�gyg�-��n�e��v-_�-4Oa�Nh���`o�Xwo��e�ݓl�i8�C�G��¥B>w�Q��0e�+Eo�b}7�����7eem�̃ۍ�ϯsy_��Qw��v��bw�b�����^;X���}���ɮ���8��p�z�F�W�X#�P:��/烂p��2.��y��2=��X3��2��s��-|��s_SeyT=�ɩq_��
{ߣ�>�Mw�'���}��l%�#��FIr��X����r�7�|���o�;��z��z�$���Y�nD�L	"�bx˸&>��g���Ggc{(������r���=*�ᨯF������_}���w��򒗼��=�=�Ǿ��>������9y�|�`?�o�������я~�D1�V���~�_��#��S�4lpO���`�J��3J<�'>�'�T�+� "k�����*k�Ƕ}U�z �*����
�^�>SR��j�#�D�Qm�ni����G�U˽G�z�k���_o_fGe���\��|lj�n Y���ky	e�3R��O*V�>��Qw�H�7�e�oeU���V�����e��(�+�����:�	]�\vI��ՠ�O1�g����nY����R��*o�I�?_u���)��
/��J&3�@���*��\�B���h��]�O�.J%w��\�J`cp�.�Сt�f��Ġ�q�q�Q���^�iH=�ЖX%Uxd{j��S�dN%Ajq�|DN �f��B�)K	�u]c�,��	I����&AG>��y�;/Y�0�ճ��	%�C]�U]��Z�yB��"8O+(��W��z(nȜ�{s>�^F�:�',#�� ��"�ۥ�C���Q�c�nh�p�n<(��Q3��s��F�cSH~}���{cA(W3JA�g�õ��Hp���>�|Ǳ8�P,�ݍ�8h��
��몴�P��QOu��] ��� �kie��v�l��7R���}V�M�T)ص�2����ޖ�����z[��UC	��}�������̍CA	ó�½�λ����#��?����Ǩ����w��k�&�_-{}�ٟ}�m8ݓǜ�m)�	�:�����=(���Sr�W�g������h9�ȵ'�-�@���ɴO@��*5�\ߔw��;پ��~�b�;���,���?&�S����9z�q������o&�U������ߗ�}����T�gnf�z.5KI�S��1_�+��3��U$X����!��3f�!M���BN@�^�E�.M{����
�)��Q��8��U�4�C�hSY�eF"���څ��Mz,�@�uV�G%y����*�j졼���Hs���}�R��'h��
[���#W2Ú�JvE+R��ݠK�ˊ�"u�a���rv�N�Xc��r�X�����'Ǥ3PȎ:V�k�15EY�M|�c��7�5�]���<�ʁU�قj������#D�X(YE�@L��.���7�4,�ɑ����ی�Kt�-轌z�O��?�(VF)5��dO���2��:�;�)�r'��1�v�ݘKB�c����kX�����ب��8�F��ӁT֨<���^����\��vo��\��H?�"\���reJe�S�Ӌ*�6/-I�f�dyeI׻H[�W9�i��ñ��9C�`�J�5��++�?j�)''��eK�Ą�Wڌ��@���Fq�F�~�R�A�&�vUJ�j��gc8�IT�U��~oT�\?��&ɾ����P�S��OlRL>{���D�: ��<i	a��+��C�ޓ�jN�⹒�ao��"���v[�~mϱ{I���~׶�Z9S��p�������.�r�-��ލ�������Yω�B��^7 �����{����l��pIZ�G6��'�n_�*x��������&�8,�o����nB�冒�A�
��<�z����_�b����]�Ї>$���F^����>0F%�wQx����N?��G>���|�w7&��a�ܴ����)�*l���Cz������z�!c�ld=��lH�t�#�с�������9>�яQq����-z�W�|�����|�S�����|F��;��	�����{��^�N�0��ϟ�q��z����0�iD�����E���Z&����.Ԯ������l<��(�@�
2�A|�����3�K�.	�RB��^i�����>�šo(k����G���0��>���g��F�d�(������*bX������s���; ˽ 	��q
��~d�K��G�wm#�~bP(x�iI�_�o�jv����v��CУ_��u`� t��Q���*
�Z[�X��������6�����8���S�h��(�d��uw�i�(����'��ۺ����Ao%��m��2��=�O<ř�Q[^;5��P:%y*��^Өi$�7�qԐlԍl���UP���j �x�}A&�I�}: �s���Aw��}sD~��=je�/�3���/���M:,pd _�D�C��>Ay�Td�>��4����x9b$�ɽ�I��Ȝ�X��<�Уr�����)��kRN#�9;��`�1�v���Z�vzb���x�|ffz����Kj�V�7w�ll���]�o�\=L�����\ks�� �[����ؘ����z�%���z�üS��"׹{�,ي+��ny�ݺ;a��K;tK˕{b�s�F��I��!u��;���ƽF&��8�B��C�c��fy���Q\��@S�{���2n�?�0� ����i�l�&0��+������KuZ�i�������~�{�����z:RE�$_����y��S>��O�W�W>��RI����3r��a5(V�~��~�x���W����;��c����촜;{�
��Pk+�2��.6U��T|�2*_�0�$���٬�,J%K�ӆ�p������?�c?�h����|�\��T�(/��1V���ɟ��P~E�:˼z����>���ϰ��NV��.s���I %���u�q9������4�@3_���Rn�V�������r��ޣhd���k���؉`��g����2BC��Uٻz�́�@c)�v.z�~�!�o?f%uR������Ha���w�ʰq,�0{�F�(	��p~0w��H̐gʦ���>�l�c��Q�\�S[�j�
��$M�O0�,	�G���L����<��c�\�u��#�R��]oRb��2�vފ�TøX+����t� Z��EN�:)�X���uxH�4�/�[!řq����iX�ev���*$W���0c�9�<�^�G�����j���`7?bC"�i�L��cU� H��A����ẂR���5W[ۛr�ú��yO��Q0$@�����򦨍U0Oe"v3��yk�?43jxھ5����۷_&&cYZ@{���\{ݼ|�ß������מ�-.]hWdt���q��#�����/}��k�;����o������qG���;w�}���{��Z��r['�f'&.��13�������(��iQ�%��˅���]�����'&�=碇^��Ñ����*x���<-c�2��Z��E�=�~΂���O���n@���s��EN�/U* H5�u������6�֞8x�q���|&�f�@OP.��PP��ox;��^�~za�5<���Oʖ�FȜ��:>�=���ൾ��7�Y�zD�C(�����!��۽D��q���/�u��a�	�(���y�t�a1���h�^�r�w���������/�����#��Zq'3�\�y~��~��1��@�zǹ[;]iN6e��y
8�3�����uzdt��\ϻ@b6)<U0���*�dh�����ߜ�f�N�~�*�I�P�P�h�^";R�����D�(A$����T����S�oKQ�^������/����$�w�WfFg�5�Q�Qؗc�m��1W�O�쵚�z�� ��Z�l]�f��{��p��ַ��c�Q��7��|P�ۭ�	���K2��%�mF��<��̙�Ja�����e)���t� V�w�����-F����(��#����R��s?���ر+dg��2L�MI�\h��d+)��uH��6d^�L+b��!\�?̝F�
�������@c��y����*�Qf��pRU���;�l���^D���5���Q�h�=&1{�������bP�Q�" R���������<瞙�+���������.�;s��s�9o{���gzei?����9ە�1���6
!S�H{�*J��??�ǂ�K�JyޖFS�� ���NSYΖ�8��3��+�86��fH?ׅ2�ɤ����CW�c����m�������HpUS}˿��g��'_|��+�9����"�;��<9||m��o���}��E-:3���^P���$uN�
DY^ �u�c��}Y�~p+U��/ho/��~Yv-k̭wEs�����w�w���(��!�p�(˘��h"w�`G�Y��G�Nj�)3��fd�2N*���uE ����m`�C�{�&��FY'��w�����!R���T�ÏZTl2Dz2%�c�D(Ny�o��q�s���<v0҄X��H2!8V^�_]�1<��5��{�aF5odT�ޅ�	"l���z*�G������T����wS�nG�.�m���{n` `lpM��JX�������5��e��qb��Y�ދ�K�1���������7ȥ�^�{�ܹs�Y�׀��Ȓ%K䡇b�B+���I�2e�L�i"��!���=�l�6��_w���ׯXg;y죑�3'�Ζ]7�	f:��Y��`�,(j����P���]3FS<k��	�����{�P��n�B5E#��!"��F��'�r�o;��t�}��'���Y�9� �;A��cG��=d����>󬥩ى�M�1K�;pP�o�~�6��E�l���oz<S�nAL��9R���mj뵴8ڊv�H�w�;e[]=�Щk�q�\�C�k���f�;�)[���!� G	�__� ~��d"C�j �x�ײqs-�YkK#�+Y��8�B4ȹA���3[���4F�!h�#
�c��F�9�d¼OǼG�� Z<�R�����UU�|��Gs�1Pz�u���J�t�A��׏�)S����&�OoZ4M��JrW��� '����(ZH�����3Y�|G��-��kʩ<Oܟ�@�>��dWR*��ƭ��p-(.�`gOwlu2�x��Î����n���c�z�r噵/ϝ��3�������D����x�� Ȍ��C�5]�X�(b���j��6��56�w���0w}�]�vG�'����- c�)��t�M�Z���5��m�ܦg݀���]{9N�@�1�}������2�P����GT�f���q��v����¸�6�H�F|����HY!-�I'žǜύ~�M��p������f
�kuc|�ĝ�����M�>�)y���/�����B�5j�o��PGG�,j�Օ9��m�i6����?��R3�q,M�+�Ʒ�sMO��T��^y��7Ec`�D) Q�'�|B����?��Y<gd"�M�F@��ŋY*@K�	���W^�E���='q�8��#�h��#�N����!B"��Uv�d��Sk�|g�ĺ���RD���7u�!ӝ�����P,E�A2�m��� 7j��5��KRgC�	���A�<PY4�$��q��{��7ѺΚ4B=�|$nk�gJ�q��e���k �w���JP��@�9�ȴ���5e#k�?0�-�M,����WL��y�L�	^[VV.����<�=oX�LEe��Y�Z�ӆ4;6�`D����7p0��6q��6иϛ��9F��5kW����׀�`w".Qt/��`)�aԌ��I�`���A����p!҂{͆��)q��Q�����P�ZL ׏�d�Rо@��c�O�������R�(k2�-�"�3j�E����`;nIۍM�f��C�5�0���Ca�N���$j�V�Ђ7�É�y��R+�ejT��(���eD��@�N5Ȑf`�3@��x�΍b>{&�6�QL�3�}yذa�H���>�D ���ֱm�s���[������O<��wf���F�8N>���O?ݴ�����y_��d�%���u�<8��t�=;(B�(��1��I��:������n�5l�����
��{M��#ye�}���m��5��,1��,���ޤB�9�\*�Re��~��|C���Ddz��}}T�q�y���eAn�<wT����(�d��^��!�X��g���8��E��L#�H���jY�WN�z���ܘ����b!�~�~�Ǻd�ҥ�4��~���=w�M�8��������� ��_|QN:�DF�˖-sdQ���Fԋ��~��G�:r4;Q5^���<�ߛ�}�����c���]����Q�&Q�<�q@�8j����]C��g�#���~����/�����6dp�p\�o �Ps���dժU�h� َ:0�V��f���q<(�!�ȹݷ�Օrwpj���1�N�ּ�k��P�͝�3S���46������|Gۙ�凙6*��[��۝H2\��(�*�s?ѝ&���ȃ�L-V����h���f��#��b$ww��dSD%FN�=p"�>�0)�u � �W�I_x�yn��<�"����~ �<E���'�p�:���p8$'q�444�A �PTL@��}���A��Oj��l�u�K3_�ٳ�e�6��dO���H3ݞN���WJ�Ф�7��(p ��.��!&�z���aJ��'�K�l2:X�����g�����T�G�geK��d�d��BǍ�(�u�.�8>��]B�Z�d�I{�Qꬾ��:5:�]r�����s��M��X�:���9s��*5��jTO?�4R@/^���G��Eg����-�=;�R��t��I9�Ѓeo5�H�?�χ�����^{�i?=����D�S�^��HA	�#�����Aiy�\r�E�~���_KH��w�t�+*��K.�A���K/�"o��&��(#���JIqAGsS�7�M����_��;��_�g/��^~b鷛jҾ�O��2i�O���P� ��ߔiI�Q���N���es�I_YR7`Τ�3��tw��w�@ݠ9���8lZ�����2s/�\�o�m�â$y>ooD��=��֟��P�u��I��v��;;���[�[2��B��`<��4N�]����О&Z7�"씩��:��q4�K7J�y0ض�m�V~h�FB4�.d+6#Բ��׿ʸqc�SN��"˃:�F�e�ugx�V\7P� �-_��c:|�p֜�7���ΐ�7��5Z]qL�θQ{��Q�Fo�qp|N� )�C9�����ϟ1���0�scs�9�x�n(Gq��k���Q�	'����t�Mt ��{����g߽پ��h��J���jK/6��g��<+>���Wۢ�Xu�,�ii4���&�ʴ����#�a���t����	
2��%Fˆ��:�2���x����f
IZ� �G�IF��#��g����2��@Yq֏���L
>k�`����u�g�,yA3v��}�����d9�bB#t<���Gn��^u00kr���ԩS�=��b�
:�(�`�G�q�Yg�/� �Ǎ�;�C`Q��\��o+߬^��}�F}�=v�_��W�O#���63V$��,��|	����"�͛ku�Hn���s!� �y�9:.`�k�FNx������6o��V� L���
| �e<:>�@�`�i�CA��=�\I����Za*# �uBD��>�c��~�I?��;D>xo����J��C�u�<��R��� �̣s���j�J'#듩g�Ό˪��y�M�60����ڥK��S�#I�{�[v�u5���n{�*>�w9��g2�q�ͷ�Q^�v��1�gRT\.��9K�f}���(��(����7��Z�y����X/'�x��=���%˖r͏9�����-(�q��D��ee����y+��yY���O?�햿?�p�֦�k�;F�BE� p}���'���M�-��Bp�EYpؖ�n<��^F�n�8,2آ���ꋜ��M�ߘ����%T�Yd^
zt�h^7
�$$� 5�Q6oGT��,��i"�|h[�l��M㽈H-> 瀗�סvĥ�'��6�i��稬*g�mkS�zK��VP'�F��/���`���L����'@�ZUD����a���d+R���[��\y�U�v�j�0�����4_EE�n�7�{G�Q-�:�Y�����{Na�<|����,!Rq0�@���x�!��o4\�ͪ��n�SD�UUe\�o���V�{�1�8�AX3���F�6�G}�}� ġ, ����gn�����>�ʊ~L���KxVpl���r5�8�7߬���Ngr�E��>�p�V�,i��aN�n8��ύD��&p��5F�1hw9F�q��+���߫� ����&F���.�'��a����jX�4j=)� L1Kd~c(~#&����c�ñ`fy�:n��u9���lX�zj��P�A��R}�����GR���R���(��`�����Jy�Ǹ.>�h`G��L��?��ر�%Eq� ������Snh�&��yMft|�J��t�by���%����ك��/Ȧ�[�QXX�(�-��u�ḷ����W�������:��ӎ�7�(>R��v3���9\\JU3� ��)UԜG��}E,>�Gp���][l	++�S�1�6�?�Rџ��g����ߤ�"�`��~���''q���dʞ��)?>Y�}g�|�Q9z�̟'�j���:�{����GT������g�^x�))�}N�{�Nξr�o~-������0^�y�)��OO#aU[s��{�Y���,�������0��q�9�H�C:գF׵��|�������䕗_���"Y��r�4eO�����䣏e��N�'�z�m�Ao�	��dbۄq�ޟ:���/GqP��_.��a��}t<�<A�_/=�`�]�i��3��;��}�(�w
�,e�����A7��>�y�p;n�������He�t�pG{6K`k�6�����;Z�)n����38ȫ�ˣD�sݶ�uI��)Oc�}����`�3�u���D6l�) j�����Ė�!���>��V<h�.��*��¢���2%�T4�@��8�?jԹ�6�����˘j��.8x��^{-#pm�n�>v�x�����1A{��
���3�#D�0�����u[d�����`�lOlMM�l�:��s��j�8"0���Qܩ����9��&M�Dc���������yٌ�<�����s`C����#�WFT��=�}��NI�<��`^!��t�1�H^�C��3�����io���q�<�X�\6o�N�bFf��E���:��ϗ0,i�!{�x�(cy�A1�sPS�L�I��4q�qyĽ92N �����۴��n���SF��hƤ�A����F!�}>T�#�9D�܏X�c���_H�l�(R�S��[^y�5)�(��O����D�
�Q���������5n��y����ϡV���ur�I'��aͺE
A� �q3��m�y�|+4��y��Y$7�w߽e�K��;>P��Ka��M��r��_�Ҕ@CG��2�!��1R��1�Р��s��z8IԽ���~�QN��?K��B����C�`i��Ur���bu|�Z�lC�X�l	�H���gvذ!t0�x��d������d�ɓ���JiE)3r�z4j8/!k��*�*������s=��#Ҫc8t�H�z�2>#�'���+4@�Z�Mj�FN���(���:l���\�g^p��/#��@��Jć}[�+0��D�'�eʔ=ֿ�����:�=���;��fk[}swv�e�7���#P��<4�a�J[���/���u&M>B��;�n{�=ӞekP�g�û���w\�K�;w_��,ؾ`w��ll��Ѱ���d�:�헵�u֦�t�ub��`V�S�wv�lK`~6���"7�� �[<�d~���?�,2����hJm���o�J�~ՒUG��Ġ�a�,��'� �`2D�0hwݕ���_~5ǐgk �!��ܮ�O������e�FW0��^ >��]�δ�i�׹`�B��f,S����_r=#��>�\��{:_}����H�����6m�H�xL_��˶���
޿r��n� �x�4�����eox?.:az80\x1�]�3Y�4�!P�n$]B�.(�A�0}���KƩ�2AM6�I� ��Hv3�2�E��r6h�LѱX6o![�R����S��t*j�ޤ���ӛ&��,F�H����Ey��,��jQ#sY�D��սN ��o3�:/��JwW:�h
�SҭNlee�\z��dR1�`+|��j�r�����W�x��5��P�T�����������u^D�$I*)�����:)(,!Cc��L
����SN�7gϒ�3^������f3�|��iU�_��`�ԑ%���AM{�]<��Sq��F&�������(Xe.�ZC��s���S���en������;�wu��t�p�2�$�>:���  �߲I~��.���uk���=<��c2{�O���U߮f��7b�h�m�It�}��d�g����4��G�W��M2N���j���m-<�`�ڜ<e�a�+��m �N:D�v�=F>��3�w��|hЁ�2�����R��{oh�H��H*���o�s�=W���ղb�jihjֹ�d;�#���n �e�Sb�_>Ə��ђU��m�5�ն�����e�K~'zu���!9�4K������6Rw��w���ջ��F��~���]���on��܎�=_����^�m��=�0&8�2f�3ȯ�< @� ��t�_B$������V eI#�� Zu'�h=�|yH�"��p²m�:2b�t�4X4y�nR��~�D
�^�9<6AD�@�"rE䉯��Wҹ�<<w��i�
��~�? ��x�hma�s�p��fC��ŏ��	�Ø3R.5��Yǹ���G���_�\��>�1c���re[� �[(�3ܘ��;�<�C��#�F�������d���D50�o0��i���Z����΢�~#L���dL�:�gY���>8r襵] ��:�=Y#B�v�|S���x���De�F3ǟ|#D� A�`�?�T���y^����<ב2���]x�&�'�5�m։��+�;��ϫ��=F2�s��9/�e�="���� ]lUB{��ԣS1�b:�~��ߩ#i�|18^%�5o�6`k|Ai�q�jD_P\"�׬%6��O~r�̜��,[�B�ԍ�9���wߕ�|z  ��d�a2j�N�֬���k����/��Z��[	!���7Z�`H�lR㺷5T>�;D�=��0�he)n� �cF�g��b�א�Ę��L�6<Y�h�@2�k.��G��Q2��o�喪�<)/�bMz��`�kkm��!�d�ر�TH�!K$�g�l�:����I��Z��-��-�>��K/����{���YM�]*����I���&�Ю�hE�Ԫ�~�a�H\�C*�����m�q;�B*�r��p�`�v�m���[��،�e�{u���k�d�ٳ6ok�:u�{t��(k����-�r�����O>)S��SV�����J*�y�a"�;]ـ'�+���-�壨�<�?������Զ��g����l&���w����Ţ�-W�=�;�a{��^��m  ���a{=ݹk��Ht���)b��B��_�g<���]
�����10�V�ގ���|�~�9�c������X���!�<'��=*��я9�.v�;P{G��x@u�<����XWs#��;rϑr�E�4� �F�FF�/R�4Pj a��h��D
Q�'`��(��e�z�0F��N�����@E;_���?�����S�;린Nߋq�
h�ɑ	YD:Ə�s�����N�/^�{�{p�_����`<�T��@���'�X��c�6\v��Ӕ�
�����#e���L)j�ꔅ<�S&��0Q�C?�F��7�e���fS�e�z�Pg���� ��m[�_�*�醋3(�A����P��3��<����e�!iqk��z�Q�K;�#.3��ݢ'��I�ߙ�j�65\��A�5"�3�<m�o�h�DAuN*);k��l5���'�l�s��r�Yg��~w#Y��~�u�ɲ�v�,X�D�U ���7ˑ��� 3u��y���PuF7ޓa����g������+5:}��b,"��p��pcMG���:���~wgB
u����d�\�٣�ڴ�9�D'fO;,~0� <f�A��f��	1N�7'}k!~���:�yO������üGA<o�4�C��wd���v�qG�ĉ��rx�:�'�gV郏?��{�+Gq��3^�Y2i�޲r����'�ʚ�d��˄]v��3gJ��T2-�:6q)��O~3�:���2A��ig�%>��t�ar�ԓ䡇���C��ig�%���X^z�Y�Ӯr��˟�i_�Q>��Ǝ�X�!��_Sb�D�K��C���IGo��A-*��7Ȍ���/�?���3[u/Ž�1�=e�����������	�_�����9��/�c�^�G>��]�eF�i��6R�a�]�#`��"��uTr���$�(�]˷��{}����m���͊�X��;%������n?��o�u|G�5�u�->�� !�p��0�Hkz4�J�t��Y�g?�"q��vl�|Μ9��.;�>�x�R2<�������k�a��#����!���u��aL����N�4��~o��Z�c4�������` W�g?�C�G]h{���t�4f �[�Q.ڕ�O�}?��q�����e��8/6�~��Y� �[n��-!RsK���1�/�pD>���\��&�dc���hQ�]���<�@��u}��~^�g��st��� ��ѧ��7�|:F��.�r���ҋ���� y�!ioh��+�FmP��ńk�>3����7uZJSfM�7m벮��m�3�����'��>,��2�)�kЉ쇣�3�p @j�,-�����۪��F���@$H��X&�'����䱧�P��Vv�i�<�ȳ�ƛ�į�q^��Q��&uJd��gdU��#�;~�<�䳼���5̺@F�=��#G��A���C2���Ǟ1������dOt��p������
�hi"W�E$~a9���XL�L�0,QP�+��A}|т��P'�f������gV�4�d�@F�bU+Y��O� �B �s	����
����E3���o�5W_&{N):@2t�P>j�\z��D����l9���[5��n�Cv�8Z^|�m�􋅲�Y��"�^p��W�>p� ��?2}�<H�j���_�s(g�;U��?�����䅗^��3����Y��s�a��b�p�\Tc�k�չ]��ٖ�9�G���D��\t��RRX�iv�eWȵӮ��/Δr
���ѕqh���J3��w��9����N���L8n>�42$b��0b�~l�s6E���%����82+l����?wj��Y�KI����i}�z����o����ǗE.�,�;�&����5�M��>x7m���Fȍ��5���9C�`X��T���̳a}m/����H�R���)�oo!�um��p�M��avg-
�V�δ� :�"-� "CD:H7��O�rcD��r�� b���Ĥ����4�����Qȳ�/2�f����m:�F��{�_h��^;z���5�[��1ئ�o����
������q�k����1+$c�(E�8K�sG�M�[:R(u�e�Z 1�c����2g�t6F�+��<�ׁ��js ���L7�l*ìC�^�9����%��	P��w��}��ܸ^���,�d�N��4;ڰz�H���������A����p�����϶7�ko�Hک��6覮����a�S	�Y�4�����kE�'�����l�5�|��'e���щ�����E((���z�*����e��5�ڈ<��S�XZ&��w���$��Q.����K�:�⺤��J�X�X���6Ss����)�g�,G�6��~^�e�2��Q�I�BEM9A��	s���$��cM�5Z�~����-~3��<6�k�:Ĵ5z@�N���>�6i��5ۑ�ɚ׿��9Rӯ��s��w���T���V:y��U���r�]������5�s1j�F�	�3Y���5k��,[�u;j�8٢s��76���:��OV#����3^�%O����̮���2�gSՙ+���|T,�n��o���S�d��I �ο��-R�b ,eղas�:t>=~g���O�W��5At��յ��F���=%�:lm�_<��M��Tw$�����eAP�= ��z(�X�3j��������L�s*�
Ez���9�Ծ��}��F��k�!�iM{n��|JߠqI�M��T����M%	>
�/�C��jg�̆M�P�R�>c�#ܔ�� M�_n�k�=ش��A��r�iKJ�1,)*aj�9Dψ��Vg���t��
_FE�n�0���k7��{�v��G��������nFJE��c��ދ�������;묟˼O?c�������mns����ugk`4PR�:�t�|[���ϕ`,� �	-&��f�ѩpZ� �Av��#�#�<BN8�x�ݼQJ��dS����g�L��!�����aÆ���w:��y� i��p��c Pph ��V �ׇ��}��_�{�}�\`⬧��]��Q��v&��Doih&�ϳ���c�r�r9��C��	V�u�n�~ wZ[�e$GS�F_1@Y/�����w}^Ņ�8G������p fL�!_H|�����R/k�X�Q���l�T'!m�V�R��A!�>�gӽN��R�2����8�h���9�]'�!F��;ׇΝ"�`��D��J�U�,�ڢ�
)W����Cb])))��0*1���-�d��+�N�}(��k��ӅT��`kS�dѽ���[�}�E}Eң����l��:�k���j�rk�nS��QL�Ԕ&�C݅����6SR,��ǽu��-&��(�Ad��g q�0�>�bg����4��=�a�T�(�XW��uO�gL�I����f�\�L�XKII�0��MZb�rϟ��6A��U�W��hW<�k�;��?�E�:�!]���|���7��{~��_ym�<��'���+-.Rܦ�q�<���'�V����ț��ҁ�=�N�X?���ʇ���';��{�P�u����(=�c:���	i4�ч���s?�bu���ZL�0� �2l�,]�B-�Z��0f@6�ޮ봰 ꋵ��[���H��ǶƦ�Tw���,�����]#�p2����⒩���6�8w&��uc�}�U��QJ2)S�)9C�Hf^����q.�_[Ͽ���G���&h����t�������|Q��RE��gb��&k^f(����@���w��$�s��F0@%�y嶼3�/`6�iT<9� j�	����&����g�KӒ%���1�:O:�M��s:N�X"������@��F�=���w��r�M7Ё@��A$�׼��V��2n�ŵ���GMu���	�ȵ���\v��2�� ~_n@r1�[EH��@$D+��.FUW^uk�Ӯ���E-���Cf�H�d��kzG��.���zW]�O>��C�喛Hn��3O��7L�U�|+a5J%e�l�����QMU�J�v%���V�^bl2Pm�*�� �R[{��M ����&�Yj7����"{O�K��e�����
J	7��������!�hK�p���V��'k�]��fWAXо�̛�@Juc� J���*����`�C�"��x�����:з�}"�*7>�7����[n���֩�+�Ts��'K�*\L:�GBVB��$�Z']�M�����Wrcg�6T(]��!77�m��6�Y�4�lXK�H��*�FL�ާΪ��y}N@��HR����Ji�Z�N���U�q��UT�k���a�:,@:��y��������AC���4�ެsy�n��<�F�&T����DJ*�u!�Lu.�H���W�]*]:;!���ް���F�^uN�:�A�B���a�aR�7�]g���+L��'e�����`�c*ݫߓ	f�,��$=�i���_"q��H���`(̮	��?�$�0C�3�,K�d�@:����HޓH�$��9ZQN	��U���<Bb���tJ��\��T�h����)�p��aXub�0�*�d�<a�:�%���C#��v��{}i��_#�f���q��o���9t�@��G�eL�qay��}ku��	S�����,J���i�9ZQg�OHAG�*I�}����z�Q�0��uL�d����ߟ����ҁ�>�x����/��W����x<U$���B7���j[ScT��gړB��pn�N�g{�ړS����Fޗ��}�5����4}���!nɥ��!���>�Xʛk/�.2<dl�ԩsn��=����Ms���I���r�3�w�fS3�[�g"S�5��A?��b�ͩk��0��0L�mm7�<X��K
"�,{s��3�=�4iw���M���k�q�T���n��~�pc�Q�b��v���/��?��n�~8��x7����6����Q�*��csGE���)źm�V�s�8V|��4a������g͈��!�ȫ�����7\�|���<Ƕz�U@d�g��*��6��u�xQLڔJԘ��q��򫯘�?��|o�,]Pg9� �H��E�e�77.�<�j��zG��c�<k�3��NP�u�޻P�XDiPv"S�I�2`F;���d���������<��}Wu�tc��hT�1��T6�tc���w��d�}'��]���E_O�ܸY�@f�Ջ��w��9��sM�w�m�^�~3i�����cB��$�@��2k��e����ܡ�m�9ɔ�lА���~�}�Ο�[��ya,��pO�I'4�nVgF�+�!�Ǎ3)��8|${�A~��c��e�.�����tT���1���t��x�P�z�"u(p:�������ac�n}o�f˲���aj�8��^��?`���7$\Ee%zݭRVZ��^�*թqد��.R47�k��^bS��-�i�|�T�q/�}�C0%� `PhFHB�#e1e �hPn� �G\I�|�u��d��<��b5����螨΅W�2��Uj�;���s��SZZ&�j��!/ "�'�_�$�jТ-,e@��
�6��S��3�W���vqY)� ��fu�%m�N#�{ZZ?#Z��K���BRX�D�!C{iHK�w���Á����$�@��7�j~�˕�N�c��/.�|ؚ�������=Ǟ��H��v�A�����ꐈ��ir˛�1I�^ui���l����K��?o伮׺��v~�?�S���~xm���0�J\�59IB�׸m=���a�n��칿�qX�T˰�@.u]\���L�� T����C�5��Ajq�34b���$�F�t!�魠0*w�u��0��;�s;�H�b�������;��3�z���Q{���Y��Ѯ���vҸ��5ꨙ�v�T���j���b��㏍�;i(I0��O V4��x�ٌO
�Y��|?7D^y�5fUn��zy�ɧ��{�,3_|Y*�cǵcOu�["4���E�PpD�5۷P6�J�05jta��cwb���$������@jӶV���a�s�ϑ��Q�+Ug�w{��t�I$6��8f�8:[����UG ��N?�
��!��zo�9_�]A�!�´i���:嫯1�P6���Lz~5� 2N����y+�c�;T.<�XHx�?~N���5iڰM1!*�:'�A��\�2If�Y�ȕ��P�z��ws�� ��S�<��:�h�J���J�0v�P,�W�ʇ�&O<7C/>���1��*kI���5``�x��hO:�x�y®,u���aj�L9	z̾ӣ�Z�4�q�lH[T���vҫ�������1����d1�z:w7��͋��,�������9�ੜn�2RH�wBd$���F�muL]CڴA8X�CZZ�!�^*R��a ������	�3j�S�ެwO���� ��Ҡ#��28=��(/����t��B���%���5y(���`D␡��za^0t&�y�D'�3�[}}�-����'��\�p&���֘^O��tk��6����2] ԣc◵�7K�S��qTG�M�YF�"ץ�lS����h������0&�r4�d:hpˁ!��::e-�-?z�ٗ����_�7�\]��[�Е����1�t9y�D���C'v:���&��HFr��֘�������pw�ǭ���澵w����Àz~�h������fzޥ����{���]
�9-�m���?�k�[ ����k�"���l��a#l����9f��\��^�"���?��N��),�҈����r�6u��h`�R�5@1lr�u��hc��P����͵�L��������U� 5	(P�"a�ڍ�6|��	�d�(�5]��Ef��fs�@7�
�ՓO>E��+��R.��9考����&�#2����B�"�XOeE5��[cc)x���d Ep��1�e�^�e��q�W��g��>��B⢍S�7�i!�id5���KiE%3 ���������F�|���2d��+�(�l@���;t�(!u�T�~@e�!�ٺy���ګ��D�6��U'�U~�!8d�� E�Fp|�t�AX]
#A�k�z�M��Ň���	r�1����NU��Y��[���H�˩��]��dK;<h���s|ǘ�����r����6ȴ0���H@��f;��̘����n��w�]�=�T�G��ᇟF���'���1���H�:��=v���ote��FαO�"G}��t��u��!Q�� �	�5"RE$��u�H���
��%���1K���k���2��1G���1\L���5cbk<���D�$�Hd�]���}��F<l�^c�����ioC�3�C�<x�re���DB�AJ2K�:�@L�L���FH��z�NzW[�lٴ�%=p෴4IY)�Y����Y7Q�?��)�>�0J�,�~
���tQ���,i��>Z̐� �$)0{��802�E�Υ��'���V�GeĞ�d�׫���Fj��K@�=����x�m�eYS��ծ����M�:C݉�^A�+���Ay���ɵG�����w�|z�j����B����������+Wm8^<	�:e�̘�K���2�q���ԫ�,#�=_� ��q^�<,D)Ӄ�uX�
[_c�נ������美������w~ z�<��� �Au6r��m��~�}����}���/ڟ+M��)��a���� Q�-g�-	�ϴ��G���c�9�BD�g�CR��G#���"����p@|��������������mT�B*�]�cC�F<�NA�q�[P$ q[�n��R�`Q�Q9��{�t��5�)O3�O�('�"�u�@�8H�F?�a��nnj�̫*kx�/�-��n���h����(e	n���Υ!nkk!��"ؓ�$� asJ�����r�A�y �}�ݹ��(��;ٔ��\�!#2��P�B6��.��.���w��/��-����)'
���=gӋ�zO(�f��q�P:0��q��GcY�;n�Ӧ�&�￿�p�-��ϔ3�<C��R5r���E���K�j�tᒐD}Q��dIz�t�w��_)�v���o,7��������6�媒R�[��7��-��ʃQ�
 b�$�h�,e02~�^�$v�ʫ.�%�i4X$����:2~�yP��a��)����C g}��K�?�X))ʥ�\M���a���QƏ-/3�+d�T����,RԨ!g3I�+tޡ.��x$`R�pH�pH ��x�L�8I���[x�[���3L6�m���o:��ĵ��ɡ��X~�����I�zD�uj��|�̚��t��*,*��z�>G07���})��ك4���|�,'�L�oдa���m���Yٸz�v��RӯB�����>�ꈩ�k�fLV�]/ ��3����t�Z(���65���dۖ�g�+�����lm����%7l��A�H�۝0��X�h0"�Muk����S�d��ǝ"G}�\x��v�*�OejWBL��Q�¥:�e�ҙ��+��d��2f�p9�ܳ���:�P^������u�*�����3�����{W����w_}������X�fMɿ�|9��O��U]K׮�ҪP{k���L6&���e�����"m>���F�g2�����s����v�(}�����������j��k����=�\�8l����@��{��v_��c��3Ϧ��ÞF�cJ�F�V_�ԥ	�x7��"�H��L};ө���2�E��؈.�XG;�)lL 4j���U������.�D�;�By��Y2��9�l�R��.��(j����k{��݃j�;����pz��"�� ��a�� x{q�슏(Z���Q9��tD�Y� �qM�̍z}7�!��ҫ��s�f��W�.��Ņ�t�W4�(!j_�l	j�� �ъ��c�J�����{
<�S{��L�8X���p�(�ذi#�۪��1���l��:x�˼�>�xD˫�B���tvh���>��,���h ʂ�p�1G2}�`8��Y!���"�q�o��#O��kx�ϫQV�;A�fW,#���3�^#�쿛v��5�9g�+K�Y#��rn�i���9� ��v�5�s�ؾD��s�H�kHsg�D^ � y��]�s�B$"�sL�e�\IL_(��W��4��pB�	Ή��J}n�673�2����ޓ�cF�#�!kV��x���q��˥K��h�fT��2"�x8F
htuL��9k��[(O�g�r�6��a۳Y��9�~FJ��Y�;���FN?���/._~�\>�;[~��h�&]~ٹ2r����0ՎdT�

#�
���..��ɍu�a�B�CJ"�j�#�SC�D���m��e�Ʀ�r����GM��r�a��]w�)�-���y{�IGKcK\V�� y;�X]]���e���i�r^_?�Wj�[�.F�)�1�'ʽ��Y�*�󌬵ٳ�d�fҤCt�g���P�t�v�1ҿ�P]��IsG�:7_��M[uN�\��/����QDo��qc巿�J�;�h9��c孷>�/-��O<Q.��t����e͚-:��R�Rw�[���}��<�l�[~��K��v��ɞ< ���_���+s��r��omj�#�/*�����g��Qv̤5������A���^s�5~�W�;�w��4��kͷ�	���ðf��݌l�3⽍��k��w�ϻ��~_��\�?��F@O�F�a��F�5��S�n�so�7�N��1w4�}�S�N�r�"��׸2�l���ς����y�� �ٿ,�O/�c-�qx� m�P�]�n�w�������#�:R�9�x5�ˤ��AV�:�bAd�i:Q=7�����R���|K�	�z�2��UTVр(��m�t
�ԓL1� SZq�ڲ
�)��
m�p(J��HKo@D���v�-����+�����r{�9Y���Amk��	�S� <��=R�h}A]�[���;8�;:�R� 90�Ct�l�H3��z�Nv����o�>ZW�U��֛�innQ�grΙ�#2j�XA���wfK�:��j�'z2N�\�@xi\|>��Q�ɾz��S�~=�ۿf�,ђJwf3F9��RP�xtw�1t�~�P����4�E��ݦ}H����s��j.�dy'5:@i�M4�#��Ȗ�"���з65��S�gҝ,��b(h�+�{��G��W_!=�VÈV�0��,6tш����Qg�X��'*��~��{��?��'��C��g,5��jK��]Ft����3�:�7G��O��1#�u��� �7��Z��Qr����b��@ƴ��5J@!�)g������E�\�Z�Z.��|��������E#�29b�q�/�g_�.67HiY��sԔ6Ժg= ,��v]�]M�wD ��O$Z�שQ���!)�,q8)^p ���d9��)r�Mw���o�]w�!o���\w��e�̗��-++�a�Z'���}�ↆ������ٳ�˯{���\>��_�9�+KV����}�ϡ�x��:;[��.�w��3�0㒯VPuؠf��kl����O��^?���e�ރV5�XKcF�d���c���/̖k�����9��=���/���H0��X')��԰�t��ٳ��_������K&Oܭe�qU}���MM��Vm,_�aS�?�|�����in�(�(L$��ޖ�gXb��`�a�Ű��tu�L�h�u7�o쮏��h����}d2���������c��1��qX�5��G�����@��{�3c���s�ϸ�� 2��r��֐GA��z�Z"sq�!�8#}����X��I����e�Dп�lX�Vs�����bil�~�ÌADq�[�Q���3�i��d?������2J�"�wL����* }��4�θ�������_�!��`/+��ȕ�kd��huK�9���}�(���m�m�ۍ�)��W��Z3ރ�s��e�[���u-_�F|[�K���8dN:�D����P�ՀD�YR )X���M�p:���+Vɶ���=�Q�$]2����EJ[7)�q ؁`�ҥˤV?ϲM�k̀�,�P@-����F�����5�>�赵��$���755t���h�����i���|9���X"��L�LB��^{��E�T�L���H� k ����nv7�n�L������rן�ū։'\�g����{���j�T)g��3)��j��d��E푔Fd�F�E�R��$H@�L�{�	z�!��t�b	�K��N�? -mq��+ق���\l�p�BDpW�HA�_�O�.�&�bl��$3��9_��HJ�[j�jpÑBӹ�y��)�tO���Fq�KUE��B��w���Y- %0�4�~_n�2����à���sM�F7��02�m�<`��w���Tb�TW���l�ߢ�S#����Ր0ayD���=��C�C�2S����Liy3��3ձ\�i�i����1��t�}����n���y���=Ŀ��O�(�ܤ��[@���;���OZ���ҿ��<������w��R��nkj�A#�ȓ�=!�xx'��cwH7��󪩮��ƭ�裏�W�?��n�A����y�5r�QǨ���y�9⏖KW: ���i�*Z�ٰy�<t�Zu�u� �M��fpS�^��q;����ֹ�֥���
y��.]�q���\1��z�Wݵx���+�+���L�����?<�Ӗm{5��jk�E�w$2��h��t��� ���s_�ǌO*ѕ�=�%��ٙ�z���9�)�HUj��0^0r�h�����X�j�[�����E����~x֛/�e��n6j8����|���>��5�}�#�~����~�V�|��i�ʈ&��NQ�V�\����*P�F�Cp����_)K��3�^���.�;�%ػ�fXX\&��z����<����0����"U�'R��W��W�n�7W�i�y�GK�+�xܻ�ѝaz��~�&9j%G�I0��E��Tk�6�Ö- ����: �d+(5[4�ӓ�S� x1:
d��'���v���!����V�C;B��gyeګ���2�Ϻ�/Y�T�"0=��x���nrؑ��m�a�`D�g���,⽁��X�f*Y�9� �b�1c�R�%�r5@p>[�Ht\+uch��<gf�2��/ם`vd����8M���ܰU�<X�PO���,��Q��|��ZO*!��r�-������|"�x�r�ŗ�7�N����Ԡs0צ�&2����LR�|�R֮Z!�^r����ʲ�d�{���S��H�}6�E��Tw�B7:0��V�ㄝv��v��-#l��_S%(��k�.8�A�}Q��T���"Z�� ľ���ǰP�<���`؆�!�«���yQx�P�B�܂�L�G$�U�aLן=��b�Zt�RY1��՛���Ȭ�rF�)�$#F�o��I`I���i��/�C?��W,�$�\x��Z�H��m��X�5��LO9�Y�.���&���Q�@�cLKK
�ԟ�z���b]�1�z�)(��ԉ���}�����n`�ұ����d�	;�:"+�/����u��A��{�I[�r�CO��v��j���l���m�>��jy��g�e�9������ff�P��frX�2^a5��@@:�E�4���ά����urۭ7��g^�ʹK6l�L@`�Cv%#�.�R#�?d耷ضq��3k��Gȯ~�k�,+��?��Oiu��t^�=L���"�;�{�� �^�Ok����	�w¦m�D]��v��e1q�=V��.E��|ePD=ި`	]�ttI \�9ոU׵:*_�\�Au6���&�j���Q��0�*g�`��l}��������wk�ܿ�����:��6�>G�k��Cirw��cw]�ޟ�����������o��\�i1-��H�z�����9����n��k 1Hq�)L�=�/����Q���7N�и-�|�X��wyeY���i��g�̙\��]v�E^�m�4i�L��������'��<5V�<XI]۪�b�[0X�|��_z�7o!��&5v�h4��g�;�- ~It4�a��ZN�h���l�?k��z�Fy��eب1r�	'�W5�MuuR���Qb����u$�m���=F������`�;5*7\�I:�p0��O��13v�,_�D���IjlF3�Ƹxv�OFm���=�`��:"��fPk6�S'=?j�1���n�s.:_V�q���"�@Ɠ�����KJE)B��'�s����a����Oe��2�W��O�g�ȿ^�7����f�e��1c��0��^T���xT^|�i9����0u�N:�9�cd櫟�SjP�a�u�3����w=��^�=�\�tm�SN:R���o�w�}��#Ͼ(EU��K B//�t@�#�PX,�J"���򯿔�;TN>�h��_�I��!�AY0��;��K���d��!��k��=`�=e�I�3õ�NQ���ҁ�[P��~�>��A 2`��Zͦp�2=Z��� �.@N�"��T������n�C���Jy���ү�I�+&;M#�B�fS��z�=�Y�O�Iz�%)����)�<:D#����i�r�nX���j5|�h���W�|�Vc��98f �F���se�.��k��C��v�,�?_&W\�K�펛�gg+C�up��Yc�a� ۮ�.Y0�ίn	�-l���dcL��{��C��,JWV��Rz�.�LY1�1�`���f�\z��r�yg���XZڌ2��:!iC��G�N2/�\\P(o�����_���lfA�lPǤ�4 �=�tj����7�z� i��J4\�2;R~��Չ���J����x��u�1Y��C7�R�e-��8dcR�uJP=��߳��$��š8������� #hR������0R��D�>���o}�������ݨz{���o�a��{#��� �o}��a�k���'_G����c(p�}�o��IH�|�U�#��3M�0��7qP���j��:b�pL���:�h������@�7��9���5�H7��Θ��lި�V>21 ���xD,H�o�ۦ�y��mk��'�#������2߲�N<�H�<��kD�f�f.8�%1ѷ;�a��+��3��.=OH��"���}�5k����Ԯ�,d��uD�(����n����g4�@�1B7�V)/���F�v���$���}�eF5-�q9INfœ �f�~P�쁄"�@�+ꘁ�c�7��85b-e9cӦZ�F�q�r��u�RV^)uu����Dm8��4���n:�� #���5���ۘ2 ��O�<["��]ό_�w(��$�I����ݲM�|�q����R�v���Ug�2���D&�YR�vkT�y�U?)�g�%;��R�*uV�@��c?�7(�@���Q}^���@��X�ke�rӭw�;���ͽH�K*īs-�����G ��ϛ!���A��_�*�w&���^�Z|�aR�z�%k�^7X� ϊuFF�1cx��/5U��nͷ����W�_@4y���Ys?a�'�\��Aڒ�y��6뇻�G�|��ȴl7��d��\$��{�K(;�~�m��̱2j�u����V���_,���^�+ģJvR�4�O'ۤP�7�S~���Qd���nm�3-:����A��C/�C�{�:����ȴko�/睨�OJr�:����r�M��ܖ`v1֩ν:���Jt'�xA��l2���dN��f����Qޘ6[�RZݟ�BQ�A�gt�ĖJ��Ȱa���kW/��2BAyZ�u���jt<$����
�~"�3j<�6m�K/�X����Q#FJKs��q�z��x@�\�D6�3�1Q
�#�5ƳDu�} P̽��7錋�$�te���#U��h������}S��*� <�2d�����aЁ����.�eI�'�o�=��-7<s������ީ��������}{G��5��pk���XT�14?|^Y�����n=t�盱�������ҭ�,qTF���!�[��$��3�y�������j�D��LZZ�L� ��l� ��j�I�c3F��q��(84j�Q���?�L���c�c�$7n���F1��O�I2�N�Y�
K�B���t�SO�י��l�)�8��`F�����s�ˆ)�^赇L���"��D�d��H�������/(�5j�l�n5d9@�|˔�7X���_#?��k���f>r��!��cM @翮ydY
�N� �<3��VVQ��v�hQ���X�f�����8OjD��}���\����CEҦ�<L	WC����#��8QG�#9��_�Pl^���1U,��!� =����|�ei'I
�dwF�v߃�y�:��tzH~r�2k���駟q�� �IN���_ʔ���)g��c9����X6l����>#�|��4�w�s�P�C7�}q�u�N�����r�����!N��]w�CN8�ly�/��s�K���1�,��>���Q,�_$<�9p���O��Gy��{��Q��	[��*�}])Y��e�F6L��_^y��y����5��D;EŐ��U�%�HTRh�J9�9I��MZ�
���tւ��/83>�ҝ�ĳI�:�[�#���#֮��ߛ#�6���Pv�4Y.��26j���JmC�4�Ʃ���RZ֩��^p��TU����6�j'L�(SϾPv�m����d�ڍRPV�`)�Ư�(��cz�"�jo!a���j���Ŵ��Ev�yg~��իu,
��;N�C��[�F��f�$:h���L�n����R}MF�/�/�����{��u�8�nP~B�-���G}F�8�julq̘�U��
p̏� z�Q��1O}��֭�2|@��v.����!�g�M�]�N��s�=�~Tf���TT&�	�/�[�k3�W�P!�cy�	C�ut4��� �%��P���1��:O��xGAг03\�wH���� ��)N��;��Zk$=J<�ԋ�q�Ɯ��u�^Qzv�in��n6��=�62��{��Aw;�����`Q� _ذQ��렸�< ��R��"�p�Hio����e�﹧'��%NF�l`�Z����X�(��̀�6a$�/�4�C�ש*AM����d巌~�w#z���&:n�>iU���{U�.�j'�����^cbt�=,1`J���F5ZN��D"e�*�&�����!�&�3��$"�mP#R��
Ԙ����y_J@Ƕ���=���x��ESC�F�U���W��L7G�\2!)���������b޾4ٯP/�wc���Q҆ �S�A�Z��p}C����V���wu��h+ּ�n�0xH��is-��l�(����q�,�z���O0�v:9�Cؓ�e�;����(+"�9��1���~�uｘ!@�\���O��V��@tƤ��\�Z0O�=��445�O�IJD#㎮����U��(�|j9	a�	��m[�Y-jc2v��2L�����'����,&@ 9�����]p�v�.�eS�p�9��)���r��wȦm-9�^���� �Bz}��!R��s5X�ȸ���[�~뭠4���G�;��r�Xe�gt.�6}$��:�� ;;Hy��愠���O�m��D׺G�o�"5�`$6��Wǌ%�\p�vԑ2d��o�����%�J��R�K�e�q�7oS�i�-�Ǐ������?2pp?�L�<�ԫ\g���I�:5��0�۶�J<Ѯƿ���FY�x�L�{����r�����M���Y�b��RI4�j�TF����vu*�!�V����9�����qC�G������X�vC�:$��|����=�-+˫�g�����M��a��ME�+�J�%��
Xb��Dc�-Ŏ=��2�m�a(S�~{?�^��?k��ܹL4�'���~s3̝{��������������~AP01x@��Y��ejz����������ٲ���:��n�CA~��Sİ�ZvjV���Ž]ҮA��'�Uo�ZV�R��ݹy��޽W���A���g�
|ZfA�=U�)��}h���eH{@�COE�i��7w�e�ېϚY�}����~��}��ȼc�g;ʣ�\��K/�J]���{��	Z�&��}�����[���^��J �v��~�s�~��0K�+����kx����x�`t��a�2C�އ�i��e�s�����,T�s�9[ct,�{'��<���k���d�E�,���G����jtP.ë�/NF3��?f�@��j�!eu�F�kh��b�+�i�ϯJz�IC��ea�x�0��P"E��P0�e8.�f�pR��x�Р-�쑂���J]z;�$��k�vH�PLR]!�;�̱.E���}T*��ahk�Y�L�ky����Yf��pd].�fN��1�%���|��H��_�ś� %�rs�����Z�r�Cۤ��O3��T��zY�>�C4�D&���Y�?�أj�o�����.�R��h1����	�bdϚ��r��l�@��ǚ:�<9�As����;v��1����7?��*5���c�cr�-����~�;�J��5>��~���?)cSCҳd�f��R�(0�Y�ci���ƺ����Ay��W�k^�z����L.{��d�д���4� u�����ΏC��޾��/K6�RY�t�|�3?�7]�&�W����O��ߧAD]�	�5 j2�D���33S̾��>y���V������y���XըkG$ݵ�Ak�Tc���>�S�+r�i���XhU�L�'&P�Z���u�r�J����2Z�:9{�)���a������>�E)� ��3�����._��w��e��6���+k����0�{+ɫ/�BυC����t7����JMpO{\�KCo��s�//��B9���ˢ�(�o}��o��|Q�_H"Ѡ̎����|�6�N\+('�;^^���ȱk�����
��>��O��'�HUncL����^q 4G�G%��oɱk�u��D�?�,��:�#2:V�k��7��V�A!Bx)E��{����%{���+$�z����s�=Ζ��;�T�{xD>�����Ij��ճB�3�8>����3�%�4���c�'H�7�@���0Dof�b+���
�!0�zqbl����e�.���s��5�p}��|!�����!H��o���;�h�39����|�<���� 7����|��M�}�u������^Xz_����>caв0�^(���g�d�-�JC0� z��p����_�\Q�#Y�c�Fa�PQ�* �F
�H����v�9{�H������y`S�$<
Kd���d֌�A$�BT�VM��ll%8f���<0+Nǎu��1;��-�mJ������1d&�3k�:�>^�ňa�^	o�`$K��l�M�^s�Lg��̰���2�NUul@@��,�EpdS5Kÿ�.Hp6(s��H/A�@��=c� d �/|�Er֙g�?��2�C��.��~~��y�]�QV%�N	
�<t��h��L3H��_��W��>�Yy�{��5�#�t�<��	�XGZ�bUL��c�wM۬
�}��ByR��f�$W\�f��jY����2S������爂��2g�ޫ_�Jyr����w�Sx�!����Ȼ�{�|���˻��!J�Y�:���2�byNz��7\&?��]?��p��Ne��u�Uo�}��Ρ/��,:P�vڹ�ʥ��X���o�	C�s�/{���۞P�n���Ԁ�F`�Q��f���{I�������3����L�N�=��#��l���Tgؤ�@��=�h=�$��=�k���	�
�������9��L�1lK���]/����ꨛ��/� =x�|冯�I�#m1ubU���f�`|K�ҙB�o|���]���[~'�_{����_x1�	���sE=���Y���#Q���3��y'�U��B�>�d�e�O~�s��x�����%z�)-��Р4���i��]s����?��
##Cr�'�5�|��Z�،|�;_�����X.���Р �L>�`���k3��xԴ�|�_�;�zd4P}Z>���˛�~���~	��zFqu�uj�t$���Z�`��LH��e��/|R����z�c�w�E�{����TƆ�8��x�
�.�LH�UG��#�`�UXu+gK��N�1mN<F� 6\36�x|M��:d�Yj4ս�W.���'��w��s2� ���u�%e#?jؕ���� ��g�,W�q���B���/ۣF�k��6������=�Ѻ�g����-��oe�[���}/+3u���&��sT��e;*@y& �H5(p�6�n�F�߇�H8�4�����#��o�_�G����P�Z߶�.$�F�c���:���!u��0����F=�zON����
R�U��&��į�¯8���q����dY���ׅ A �FY���XF�����w�Ú��M����!/RFY�@R"�1��6Y�<��$Si��O�W(0��}���K�{8��C��GӖh*��,�k�BPp|>O:�6Ԯ��w�S/�B�a�Ȃ��5�Q���vu��$7��U�n�:3�U�Z�u�l�*���cc8�E C!�������n���my��K����G�N����$�:H�smm���l��͕p<$�xT����,���l��3N���ۡ��I�u�����[���&�6�i�����2M$eŪ��tYD�y�eϾ�jD��s.|��tu��I��P�Ҭ�T���}rpD5���_g�w��~.��앓6=O.~�k�:JШי���a��D��K^�b��7$_����7�7�q�|��_������oO�mA#k�k�(�P?z H�@H�O>!7���{�5�˯�T�xӥr��>+7��^���i��a^�^� �"���}�d��ٔ86.?O�9�l'�uc�-�XE��|�$A(��DY��}�a��������K�3+A��D����!u�Q�g�fY�b����D9�쳨�p�i�j:!�rA��	�Kx���B1�o3S\�2�+k�+���d]�ڪ5ꉰ�WV��D��!S?f�:�� �IO�th����s��[�([~PN޴�}j�� X��6�O�3� H"w���s�fYw�J�t�2Y�|���%/c����4��Y=�:L��0�X,V�M�3*`3�r�o���#�7n��.��=v���T�����8$�qIϾ��7櫱�'Y�Q��f�`������
!�M��-H����@���zn�{oy�{o�ˋ6NὟ�X;��9�P�²h�ay�L�����-'�J�kt^�h,��L=yw^��d�~��
%Pf��&ǅ��f�ft�^f�9W8^��A\36Bt�c��~d�#�j.��0gYj��y�wA��5�L���O'N�@��?�C	sdʌ�'�'X��� 4Q�1#�i oAF�$�����+�1�&7�@��c�1 ����&2+A�Y+]�l�\��a)�B�I����CA����fzԩ�l�J��d,��a�P����&�����h(��X0t5<U)/z�ºN�~ͩ�A�鵁��3��e
kj0A����g�]'&���G���&�Olod�7�Q�=O�"�]�c2�����'�KP��?��!��ՊQ���Lhm�6rD��r5��D���(K~(w�@����3�)T,C����1�l�]<�F�o{"�T]��a	ֵ	�`H�*D=��i��M?�����o0�N�YÚ�����`zM�N/h����d��M����5�:�ǟ��;�I{W?���u?��>�F��m�!Vr��r��Tc�{�l�t��Ǐ-��G�Ε��_���n�_޵U�z�j4��z��W��%1��◉&���R�r����#i������Vg@���S����a��_���7~C����y���˞#�I�w��^2�(����J��%K�J{O���n���æS�'q=<��K�!}v�NǞ䉽�tIa������e�_I��˖ˎ]ٳ�����v������?�Ϩg@*��tw�Psd@��_m���b�h;�*��)�y��Wݑ&Z",�j�{�w�}�r��_��W���N����e�<OS'�g߰2S�Vu���������<�W�w�_k@�H.y���#Ǭ�������R6o�&��)R肘�X��l��R��d��7!���
9m�:y�;�$�y�t-t�J"�=�L��W�!�Հ&I���!y��'e��������e�[�Δ��|���O��Ndp�"'��Q�mR���̄��g T���c��N�$�?��f��˲E�r�K.�+��Y�o˘���\�J���-��:�]�*t���F7��ζ��ʵ��,����;C.{�%���n���;��=�����yҳ��@�_�u����d6g롽�,�ғE��4 0�Pw��4��	]� ����tC�j��w��c��K�Z�i9��X�\��B�F��2�g��ZYZ+�m	��q$sq��R\B�����HY8��W�������6�P��*���[Yd�ɶ@
��!j#뫃�ĝ�9���XLiU�k����m�A6y��g��~�jb�W�w@5D�~�� g]�� #n!��([��g���=04��=}�R��(���f4=�k��F</��J�Q�Ԝ�P�\:���w��M�l>fي\ �01d?�����Ĳё�sf�r�ө�1��ב�g!uh� u��y=V
�5%qh�7kޣ�Lߘ�!�k�B ����}]D���4��	��ͩZ��Ox�.�%e)��A%��L��K߂ʊ�~���p�ʡ�S�g5�JCȯ�"G1�vL���SSb���C"��VD�s2ҙ���i� x-���}�k �� �m���p�r讽 ��k��c@ ��o_�A����-[)U��뺀��.�P �`�7�\��Z��^���5/�0��k^�*��O�A_@���������ȃ�wH$������V�l���8˹�m�O~��R!s��U+�7�z?p�X�B6'A `u=���8pH��K?U�A�+ң�nJ�1k������gd Ѯ`S�[����hWH*�<��S������k�3���:��b��ړ�/�Owj�Pa�Կ�b��p-�*��-[��y�|�_�b.�{�*���I�{Xn�կI������8P�p_$VRüb�J�����={�����<��6f�0�tK�]}��L�YAkP�^��Q�5��5I�k�LFz�3SSQ�<h�'��i�� �e�Zٷ�����H\mƙ�#���J��?\Gs�����><�~�GU���ȸ��IIh xx�3���Hn��6��|��W���y�,_}�|��?����2�Q�V�LƣiIh�Z�3[����7��?"����̳N�^�����%�zϻ���:�'4�J�Y�%��K6gD��]��9|x�|�[ߓ�����q�)�~�:9�s�s_��<�mP>�o_��xFi�>�3�x$��^�d���F9/������[o��k��+_�J��=W�k.�J�y����и�Gs^a7��g0Q����3�%�H���<�����[�cW��'�,W��r9����){�~���mVDqMV�c���#@a'�@R�6Az��g[��i>��+����@��f~�����?X���z.z@X������.!�z ���V���6j;;Rj<��֞�n5�292�Pd~�[8t��͟�[�g.��V���
�[1��.g��2��UIЭzx?�:2���UzG����]�|�mT��Ba.�at�M�.�h�K�Q���p�����G���V��B�ОV���(m�6�K�%����Y�|�P���z������/{힗��nv�����Lw�~����;��ۭ�W#��@0��V)��(B��e�N���1Nf�.���Hc)��~�M��]3U=����ဖ���KUF�Fi��yZ��XA�9���Sf2����fƾD���-P.�X��4�f�w���kQ�K
s��c���:���d)83�rh���R4��A�Ro��� �Uil1�8�\p��iF�J���~��2��)[Mob�s�M���d��R*r�tu�F�-���\F���fR%I�c��\� +��"���;���*���FCz=����˙ua��,���lP���]�HRy�LՉD�횅���PNt�����/
ֿ�|�oIR���'�~���ч�d�Nt�	r��-�{ծ0���x{ǀL�L�m��!���f�ǣF�S���|�c��w[%ܩ�-��j��l�]������Uk�I5�W��mrꆓ�=�!?�����m�ID?��>���9����L5tm�\�z��5=��	��~^^�ru^+��R�����������C˖�h|��:�8�w}�Bi։��|�7�o7o��-\g�MN04Ț%��Jp�>�v N�`�mO��cC ��^k{w;{ݹ�q����z�Y+����E���Lh �(�r��w���S��t�.�`9���� ���#eu4PL�͌KGO���vȜ:�ى��}�LIiv=��VjJ��i�1��LNO�#	�e�x����5 ��|�ߕ/�Fy�^&�_q�:�~^��lrF��J��e��6���A/��,.��7�l���s�Ҭ���_.�W��{�f*2�)H]�˒�%��۷KVϣ��J�ջ���9�y۝r�ͷȆMgȺSNeF��N�U�wB�ܩ���	sm���jc�D��Q��}�ɝ�'Vs�o���H6�'�.Ce� �)��Yk85�ٞm�`J۴>�W�?���T�Z���V�}�׿���������\8�`���)��o�^G�P�h�B�V^k9*����GOO�kfff����5r���a��'�����
 ^ߚB�����[�*12���q�e�Ey�z�a�lkArd�l���s�_�.�q�k��G[Zf�����׵������8f�=�7|�������SB�P�)s]���'4ˏ��Ԭ�$��h$����ؿhq�O��}����s���7�@��_<ԋN?>��_����|��w<�����]��kn֮F��(6�#���Is
�5�n�![�z*1�6�P��S5�/ȊeKdjlL�GG䜳6�ʵ��S��~9�K�IaV"~G����p�{��-8�	���5�A����R�Ԁ�����ב��$9�MP�"�<�y�ȹ瞫k;'O<��d��԰��E�De ��H�B������<�4���<Aщ�=;�U��Gnf�=�p�-��(�ց���e%��x?ѳ����O��folw�G��4f����LN� ȋ�lA�
�&�@Z�#�*j�5�������z	�q���)h�L0Y�J�(?���}���}��e@g�:������"C�0��i1iVj��ެ��Yq�L����5NOM��}��n���ưPa�\?�G na|=�n��5��%�mٺu++���z6��(����߃J���C�WCR���mFqQ~��[d�c���!H�VD��]R�3�ٞ�|��ɉZ���J���pǧ�9Eejr�6+��8�Ȱ��1�-Z*�bU�VW�� ����-I�����T��.kLhd�'���m�~ݫ[6�̀�Mp� ���v�;�:�I,�_.��f��4p	���*�ɨ��KU2��B^�B:Ej�|#+=KW��TF�NH2���= � 4�1ud�HX�mLϙ�\V�{:�L��F\a��m�r�t�/6�Q��ҩ�C^��S�O�:�F�B�X:"�D��{����η������?�F�����T���~�9�Hi���\�ṫ�����ڭ��*yL)Db�=<����CO ���㣲l�"�鍏��i���I*�Ԟ��������Ͳ��=Pw�h�!��ZB�?F�P��9E�%�)FU���}�Y{|�����o�}��ع����>��h R�J�_�v��`���_.��"b[#�Y}hO�ڭ�1�1~s�2�z�Өnx�q��,���W�>/>��e�f@@0�k$7Mn�c�N�&�R[p�V����큮Z_G���lW�1q@�G�c�h��y�z^��p�#���0�AGC��\3�7"�O�B}���in�cZD3(~����=�Nr횵��C�ý���^��w|��W_:�?y�o���	��~�����o���G����狕v��P���p����fU�g{���09�$�2�YGT��qǮ���	��K2�+�}��:Q5Bp�w�~�:��^sj�؁L��W,O�ð��12����A�W�D'#��Lu��=к���j���򖷼�@�A5씡�IY�j������N ��wi���G%��c�k� ԉ ��aHhd�~;h��Lu�5XFJ��'��3ڞ� �5@m��u ��ef	T��� G�o��������G�� �o����-� Z�p����Y�t�^�/��k��'��Ma�r�.�x�Y+Z(N�$��6�t��w�Yl�8��~�٧�����;�l�hR�B�f�"�]M3�D4('�=I�8u#��s��2�T[���>,w?�����$���:���U�5���3r���{-鿫aT'cH�r,�-Z.���/�Su���*%i�<�T��wȚ5'H,`�c��!���j�����L�3��96�V�Ҟ4��Q5�ͪ_��p���B�%�ީ�N,�v��Kr�@�4��)����6��ȺC��K��!T�4X���\Vci�~A�v<K�2��D	P���1��.ӳ��n}o̊C�`btJN<~��u��
zjGl)d3�[�r�>�}��ݩ�.}_�R��=թ�<
+�/���,G��ռ�i �}<33$I�j�6ɔ�	��1��MJA<��A�����[Ȍ���������qR �t�23b����h������)f������0�סvU�R/e�#�J�.3���u�L���&��ߧg<;1&�T�D�qR��Cz���ptO��}�j��\ӽ�T�_l�L�S��
�wN�S��B�c���3e.[\.�U����J���
w�xZ,��v��S��w�����e�8���s��	��W�h���j������x}!��h� �' H������\�
F왃&�Q�� *�+������v=�a�M;�r`���@��#Jۭl�ԥ�S��\�1��=%81���Q#u�w����QD��'h��o�ڀP���1^-��x%k�mF¦&��g���R��4� ����H5X��V��GЌ ����Ittw����L,|�}�]�?v��ƍK�޻}Ǿ�n�H��hG{[���Y�EK �"�x;�r��������l�K5��+W�3����fx�r�ϓS7n�=;w���c�x�4�5f�L�q��)���N4m�R}j�-�O�t4E�nx3��v�
�9������7���ttvʹ/�@6�z�|��ҀhX6�v��.5 ~���}hPӬ<`�,h@xh)D4���7�=�QU�OY^��=j3�l�K�"�Gv(bH&�YnoMz8h�W�U���y5��� '�����+9�8�s�R`�H��dD���o�5~�:H�;�72*�,Fu��i�~�/�����k�,�CIS�z�(���Q��o?$mm>R�"ϩ�@���G�v���Ȉ~��iW����:�h�����Mj��m���\I�3�֬grZ�4��$N�'��n��5�Kk S:;7������7.7h� ��x~�/?0 �k�#oJ�r�7~!���m�RxDs]7K6�t�\�޿RG��A&�fG�aU3I0����?��ȁ}��9j�0)pʶ��Wɫ^y�P�����x�vfs"�n~H��߿Js97+��mb�~�(f��rl#��z�ઋ�:i���,�n�W�JW����sp�f��ට�d��a����[�u�IY��k6����#���g4 ��Q���XW�����=�����ጓ�A�	�<�s����6ѣ$�l���ޮ�;������ȹ�%O<��,_�/'�p��ݪt�w�	;���H3�q��;��sRӽ�H�ٺ������W��Ç��K�~	��$��w��q�=26>e�.A�(���l����sx&��2���Jcf.'����>9�������*���P;���)����t�
���+t���p��/Y��M��iӵ��#�?%?��{)H�j����9x�G�>�H�B�UL� �j�Y��L9t�q�����������zN�_u���s�UC�,���j��W3Yy�d�M�B��j�]�UC���-O�d
���F,���?Iu�ݔ���VL�vϝai�g��EtLÛ��PX�I8�d:E�����F�A��1f՚C�#��p�(�pf|Ao{LZ��<�p5���P:$ 	U����z�u�ޯc@���s��Y���8��2����X��K)�@D�����k@~l�n�II&�@�5�����\t�_������|�y'g�|�M�~�?}�:ցH$v\�<x��՚P5�����YL`���twvHv�*+�-��N���/��|	.�����{el�0g��D�Z�\7����l8d����%�r7,��^[ khF���V*s24��U���=ݙ�w��]239�k�8��'�������5� z ������ه�Gﻢ��^�%S�i�N:���+��C��x� "�x���Q�cuK�3*AȌ[���6�G�9"����i])��[)c�����c�>�=���׭YT6������o�WfY����6	8&Geﮧ��c�r�AiP�ux����-ۦ�iE�5�NQ����eyu���<%�''l$4���=���A��ֿh	����9�Am-�NLiM��2z횁����He�� :5f4ܝf�:�9�d�d�^b�g\�'��IqvJ
SU���ɩ�g��XA+�mF	J���k�ǯ೛��\�������p��: Q�e��%t��j���]�e1�{	d+z~5 �=�X�e&>�8i _�T�<8��!�)�4��slODY��Sܹ�1ڿ_b᤾wNv?������yJv��E��Z\3ђ�8G+$��*�Kp����$�̂w���Q�}��M��R�ը���E����]��#��kvD6o�/;v< 1P��=�J�YR�sTF����
eV��������I�B2W�˗���	 K�"��-�k��`_�jS��ǥ���z���9i]b%o��&y�: �����Xi�֔��/#��Q[���eU����k����\}΁PK&K�HC;15-�W,�v�fL	����޻��J�36M�+d0T��9�Qx��S��N�A0��ɶ%�s�v��3`����^��+/X?�����¡Wl;���-�0�n�&4���q|��D�\5��:O�\�4m۪�W��t��5��\n����/���]����̽fph򲮞EI<��V9�F��ȴS&G��"��8�	�����nLd���V�Z�
�0��B� ��F�P��{Y ��Ȫ��' Ã�V t�!㇙T��}`�W���<K�5�����1�����e�����~V�"�'�x��Y�j�� �[�w�o`\߳Z�2pX�j�^�IT�ڼ�
T�u�f3��U+���w��W>�G?�_y��oy�O�<�팙�ɞX�����B�#gpxx(��b����0��,8�����[�~�>([�W3���K3
<���q�����F����}�Op^�^����Q�\`EL&0�v:�>@`��޳g�L��pA�F�b�$W��r�=j(מ�����%���,�����8�Z!;'��0��tϠ��j;Z>0���q����QDbt�h݈��{��Q�z|�0���[' `���<)N�H�R�i�@!�+��`h��l)�2*@m]D�>�3宻7���H��g�^=[���ɇ?�y��ߥ��I*_y:��>f�q�;�-n��R�%���9aI�u�/~�9��iyۛ���9 ����������E��Ï�/n��c��|0�&�����?~\^�ȚK�:@A�=�͏1�A5�۶?�Ye���~� 5�;�=$7~���ҋ/�!���PĈ���x4�@tFm���e���9͐��c+�1������'�����{﹋������A���?��ϥ�QT�0�,�#hp�G�e�&H�s�R��z�C�%݆`@m�ڑ��t/7e�޳�Z���:���6=G��<��ݞ����!(hV��^�/�w"i65��`	x��ܔ ���ig�����4��d�3���R�@��a��w�i� n�����?�Zm]���f�P�t�$;W�tT��@�k@�ogV��8"���X�"��e�8*��u�Q1������ʌ���i�^����{d����9��/�g�_n��f
1��g�aO'��܌��.9��>�U���>#���<��b�U��L���M�Г#Piz�E����eqt�ҩ6��=U(�H#<
�5}�|%�cQW������3����CWc��v�m����4���^�c[�f�ϻ`�ٴ�����O=����Z.~ı�C��矟=�E/�ӭt�G?��=�F�陊��"25>"v�>���rhh����-3��M�Q p�O������s����`�
��'��i4�#QC��erE= � �7����M�ddrz�\�@���`�_��W�r=�F�Ոv�� F�s�1Df���jF�������h�Zf���;n��3�5�>9.%������� �+}����T(Đ�g�p80}�yg�j���S����d��-��-�X9�-D|~C��������z��*l3DX>eS�է"+"@AÁ����>���wo�g��"(�5��4�@S=͔�1�~������_z4�������$,�)D ю�Cc�g�yu�j,���ܷe+���ӧ��U�>�f犎D�!V!�ecd��w�<�����0�@ R+f��ҽ��>DP�K�����{�U����C���G�n-.�R�8��:c1���OV�Z˟?|��4�^��:ŧ�,ZL�$@�U���쾎�}�9�V�">x�f�z]�HZ�	"�)�m��Ի4{��/|�s��]J�<p�p}�l<����;�0�����,$2�P�0ރ���η���7d������p�&3�G�j�3TS�p��~-w� U���FxT�L~V=�4�w�sN��rwW�:���{@>��/ K�	�Em�1U�|�8�~��06���ej�/��W4�s]�D�<����&Q<!�j_�+�I����q~�4��"@�49���4�Rm/GMsN1ɡ���,��M�OnF�>�����D�Hŉ��uG��v��ٲ��Mi������>�+���{�M����]�xG�-Cfd�@��1��A�=א�M ��˨C��{g����Ms��;>5Ɋ"�`��[�L�%$7��v�aa*���\�
9/ٲ�V��7��"�c���k	����J��O��!(mԁkH�yZ�5�w8��w����U��'"����F! �`HQ]�Y�+��\����hj@Pid���S���Cff�����3	M�YY���o�A�9���N%6�m���L��-�D�����������w��9�r���A	�;������ޭ�Gr�^��ԧ����O4F&2�oxN�ƌ>���N���S7+�fb��/�Z3�׌����p�O��'����r���s#�5�D��[-ӳ�<���(���D����x�܀y=,Ȝ �I��P�*�}l�R�x�i�p�Z5�yRY���fr���i�[�%"9�nho�[��C �-��%R$�l��Y~V��pJ��"�~Mn��f�Zń�n�B�,�h�����'oX��������VN.Z<045�Ӡ��-21a}���3,l�JѲ�åc׃�U?�8�lْ��L�Nr�#���;:�\��֡��b2�G��g�+�#�f��TI�9�.^���W�^�:ͪ���8˄�
zjc�*�� @/+���7\�����U������CY#�F��V��&���s^U�8�����^��J^�!0+�qk6h�2#d�#�%$$�� ���>�ѡ}�pN�d[:IU�٩:Ƕ�~���[�� y%�G�`S���1c�&h"���3�D�Z3E�G�5�dh�R�������q�Ų�q�݂^{2Р H�]��@@B��l����t����iF�-����Z�������{�^r�bf0��`�2*#�77��5�#*�d��U�U"+Ya�jXS����5K<,���v֔�]#��W-[L;r���' WНׅ��8�, �C���2�5��o�>u��� "@ݿQ�� g�Qf��2�έQՀI�`��'���F6[aI�!@�T��z��\�Hv?�Cz�5H���3�Q�SF�鷼�[��f��)��P�jp`F�0p#b+� �D9z������K���-�����5�9��:�G��525v���lU4{_�|1�~�9�03�<��cW0������y@�2�QO}�(l��� ��R�3v�[�RE�%ݓc#��j�2�l�F�`XP�E�(��MCM�h�c©\��d��Z � ���-<ô~&���S"d&�L��.��t��>GRЗ�Ź�]�J�^?�����=�H8���_�j�����7K3���������4�?��ωC�C����C�p4Y%�-��͙Ќ�*���k"�p$Ѷ?�$�}Ao{t��s�(Jo�6�Z�{3�%KԀ�����235�Q� �=p�>͎M��Dx��Ű���F�gmׄ:��J������ɍ������4f��xf�a٧�@,
��J��:���ذ������ݲs�^�	w�������+�C�TչP#]��(I3t�zm�D*:����+�'|��|y��o���ᑇ^�j
�?y��w8n���f[t��R��Խ}��t$V���h���"���m�S6�|��o[���O�hd^�� �X�l0��8oI��R	J3�D\ʠ�uM��Enu�5(�#3i���[ڻ����X�T�r%u�]2�ې�&=}�hT�պ��G`�`,����a�Wᰇ���U��0}Aq����|N��fh��1�W���8 8xd�LP�����C�L{��3�,�y`�
��2d�~d��Q#�fz��>s�/ƁA������5sI�C=��YuE<�(��j�qMM2��T�n��zo��Z��53L��N���l�3F �
dr�hf2n"X�eW�EL���&��.���b!�A�NTw��5�hNY>�k��2�<�|�,�Oؠ�{��I��z�E��g�V��?�#Ȁf�-�B����p���i���#Q'g��g\�u\/���N�jf�S ��!���?�lnI�%[!ص*K�]��%vm��:~ 12آ:nq3�͍J ��l���m���q���)�ϢB��N��|� :�� �\͙*��L��P�X�њ5+d��ܛ;{��(���Ӡ�Z�%}��Y)��S�8a�瀟���i�-����ol�5�M�	�����3���5x��P�y�q�u/OIo{T�bR�kG���z�
�G��Q[�����	��3�̳#�G���)PݡZS�= �/���ݖ�qHl��G�aIj���w�}��׬ߑD[Lf����aY�jEC�����ж��,��e�}���\r���R���C�c_�������V�a��"VeD��c���趿Iz.d���Mo7�,C��$f�+���v��}X���/_��Y#fAqZ*�x�ºP��j��e�YpM����� t�a# O���epdJ>��$oz��ҥYÖ{�aFE2�E~�df��^)���=��F���-[��=*�ӳ���%�D��:��Uu�Q�*� ��?��a9��k�B�?:�:����=��bŝ|1�Ӯwx<jӀMc�M��4Kܹ�i9��Mt��EX�-� L;'�.��|&D  "|2���NL��p4� ����-���a\�b˽(��w�;X��e����p>%yV|6��k�ʕ2N�%��R��f�ad�(�7 ����ei1`{U��� ����m!��Iww�������p�83�^ՠ���$hYձf=�	\_�_���kWk�=�ٸe�Y4��gg�� p�{v?���

�o��V�
��gw�h#��O��~v��$���-��<36Z�rŰ'R�R�{:��z���m���76�ۄg$���*��$��\2Y=SadVP���ءH�@V3m�h�ķ�pĸ�|\O�'��|6�Vf?�J%��2����f���Uk�Œ��q��'G8��rԺh1�N�'���8�`p�G�%��s�~�#E�����>���4�jr���d�J��FG�$��XNY�ˢ�@�~5| �M�q3�h�:�;U�Q�j�8P�@`��c��z=$Du�f1֩�+˖V���FI�]2�B`�nB��f�~h�g&�l7�"���>�S ��C�F��E0]���h�?z(m#q�&�Ys��*xNj�ʅ��kT�Ùf����@���v�;�|�	��чGN~�\��4�^ `�8�K�(�j���
������L����|�2o�*�sj;��rĳ�g�:k��d�$0��d[�ڼ��fF3z�O����e/��w���3�[�g�Ёx�����{�p�����!3
d���N��l�� M��l��m_�4�� �Hw�GZ3�s#j�}�(�90�6!ܻc8]��1��lSJu��){�t��r#�O���q�r�ò��{�(�"�������=� h`Q,���E����286+�v��{eي�z�U�L>��
=�Y^��T�H�REY�r��ϊD,����pE���(CE��"J����E�@� �[k����4Ȼ�쑍''6�"�<x�|`2���{���Z���E<C�8O���=_����՛5�8��mr�O:�961��:ʉ�����,�\���S6n�g��5Ǭ�� ��|�2��P�i�"�IХ��6ԝ��!� k[��*����+ 2���L�(i�w�jvaP���k1$/��C���[Kn��8�
Ȅ���ۦ�������K��Pe{�T20_\�+�GA<�<ᕒ:ހ���edpAz`/����pݒ����mUCZ:�!�Ly``@��R�e��ic�g�%5K�����me�SC����.���Ү�S��*�m�`@�jޔ@m�M�S	��MtU�T�k��@P�A�B �c�c �M�p�z���{�e�Գ��#�<��8J��Q���sM0��n�������O��;"����ظ��[B�,�� U�u�/��O����>V?�ѿ'����@*��$��=�_��<�HP�� ��jU0c -�P��cFF����3M�j�2�?[̐�ε�V���M�Yrk�á�NaRE�D�Tg|��F6%���Q��#� ɯ�qߕ9)dƨw��7*V�8��r�s����s�(�{�D��ޣz�p�z����|پ}�<��A� ���3plpʦ&�R�^��w<ժieU-�QQw7{�>��i�T�BS=�=�sss���Z>7��w�p=�B^b��#͊���b>�oT���؇?p�����9s���:rY��+�('� �.S�s�&�mv�̆�jٲ��:������T���iJ�\�+��@F���P�0>�@a�n���4�FI
�Τ7�fѝgx���v}�ޅ����xr7��,_��i�7nxlu�0����Ⱦ#�}�nu�����	�<	�*Ah@�Tא(�=�d�i@J��ڶkܣ���/��z�Ơ7<E7���9���zY,��+�n�6��q`�����u���Er���h���3kf�8`-yЖ�j�lG��Q��ǚ�h_�U�<�?LG<�䓬`䧣�KV�Y)/|�E�R���
��
`�����[&���d~���Q�"�m�Y������>�Egg� B���UA�!�12��()��f�/�#�Tu�$3�b~Όm�W��X$x���w��] �A�d��C\��HF35��6�P�rs{C߷Q ����1.�R��߇"9 l��I��98IЭ�r�R;� <�����G��X��V���Y<�GC������333�iqbZ�����:��m�������iNOMG�h�I����Wj'ׄ�_բ��3zz�dx�tu��x8(�#�����}f+���V�=[^s���d ��Bx�Q�=|������Y�T��^�j9��U�˗�8�{�&�,Oת��/�k�5H�Y���zY������.�!��gC����0�c��*����7
A�A=;hS�t:t�I�O&:uπ��	��(}wv�o�"�v ��`������`��f�!�Y�����沙y�E���W�kp�5i0�������-E�a�������UǌjŶ���sf�2uj9�����ho�����l[�{��j}P�V�>;o306�$a�G[��$��H�4)LI� =��^p��p�����r�U�ں��9�6"����SK�8k��ϐ�@���̈́�7�Z�a�<��F�Py(2�Q i��0�]ҍ
[��㩰n��LLN�r̶�`�A�L��òH�A�Sgi�Ԑ�(� adb�����&�f)�5���G�\@���iZejz��dR3_�:�I:+��]ʒ�l�����r��=�S>�����5�z�0��]� �,G�9SJ���/�#O5���>?zu���w��Y�T֬\F���]����$��0\���V&�^�M[� R;�)�7��ke[��)�F�c�z-�N8�`�2�c֬�%���sNZ
�,�Ho_��zU#�h�b90:3���L�F�*u#�rf��¶1�t�>�w�����ׂ�s�S��C	��V�c*R��8�lY�����q �� ֭��
�P�؇p���dB���� ��������@���,�`�ld,�k�W���-���*�4��!/�u�uO�>Cv�c�?*(y9U���h���F��" (�&S⟙5׈��1AsP���K�����$�g�*�~���cC�� ")�`�X�Vu���a�C�>�\'��6Y5q�T���j��M�����0���������A���D	Lz^ Fd����/'��G�i�� �M܏:{�ޗr��sD��L���g�Y�3��1X�_�Zn�<�� ��H:���cT��Q��πO1�Ӧk��U@`�R8�u*B��pzlF:�| �A(��;��2tx�k4����-�S�Rտ�Y�(�J��o�v��}-��4P,�1}�Oݻ�R��pȨ�e.�JJ�%�vJ�[�m3��V�Z-��w>��3�ʓ��V}�| �Ǽx��~�SѶþ��jfx���=]����&G���6{.+j�֢����_���_|�s����r�%��a���1�kt�^%��A�\UL	���>7�PP~ئ?mf$9�A��2��?�,�Y�n�ٹ��^m	�}���"��2c���d�2��z#�e�~θf
��@)W`�����	��v�F����B�
���X��j���=�gȦN1�
ʌ�S&�Aӓ(m�T�1��j�����?�3��<�6>1�F\�a�畽M����I��9�L�B��=*���A���q�}[e�ꕲ���8i��\ۛo�� z��;����lt��62�JX~��*N���F��A���j_-�?\oWW���՗���w�~f�����Փ���uvuI��
�!C�C-�:�0��(��U� ��z�➄�6 >0���k�
R`/�v�|1�*�M�����j��8
d||��#dD��p�k���EeLv�i�,�Y�&D:X`D@#l�M;(o<C���r��	�J�b����|K���3JS��f�$��AO�XY�(�/����O�<.�ep+dڪН$���3�S7�{�E�]� ;����3g�gkη�id���˲M�={�+PvE��{\�K��H�r�	F�NӫL� ��0z����N�c�'����f`F�I�z�uP޳k�\}�r����vC�JM� �3�X1�U˖�7hODҟ���h�7jM26�y�>��B�����2�F�0���`�O���8�g�@o
���W�T̕�v��?⡑ab`rz%;@R"���"h�W*��灙q�'���|��B��M 3P�qM�S/�&��蔯[�^�ٻW�S�?����p܎��&���O`SM���z<����9<k�;����w�d�����a3��K�ϒ�Ez�r�Sz%W!P�]����#\�c�ퟕC�3�HLG�U=�aI��>�,D�O�"v,��!ؿ?�Ǿ�L�T =˞��"d�ao3�{��L�X7nؔ��� �L�kG��FfThèG� ��piI,�5�M������q`��0@��Kv�xJ��(S"��J�����&	�CoԵ̨F��1n�p(n�k����ڲirr�q���g�oס������v*:�-���cpG�d�A�>��,��
���;)Q��F��HB�'f�[7�@6m�(����r=�}4 E��%Rj�%�t��$S!����!�+�k尲Q�}0:6�4 Z3M�f�c����SO>���&��g�%h��tjP6=9#%͆#�)�'&u�Pb������P.H'��Ѭ�-!�7/��J�e
?���t�f`� �Lk�Gl� O���[$��� q�L��I<�4�����3����O�u@P��|@c�cr�guf�&��'p�9���#�^�ا��W|���h�pL� �4�|�`K�˒Lǌ���CF�U�{�p���NQOC�p2�O�7�K��c��1�x�,3����~��=5侮�x�-�4UQ����6���i� ;��h�m`Yp�1��V2��`l�{���:��0�Ha:m��빍�wH"q����O����&���Y7�Xh{�/)�;��0�'DR�y���p�9�����V[���E�	Ѵ_]v�_]/�Ϡ{���JeĴ��`��>�� 57�QP��[g`� A9�&y��/de�<��8F��j��r�/"�6J@�4 �@jр�U�,p#?����R�g�����Y�T������Ԍ&)�GKv%d�0%ղ���zF�͞����v�:���ú����v Vh��$W�+���3�3	���q=�#ȗ$�N=�vkj2���&���ko��:^��.��<t����J�X%]<a��,���Vm��O	x�2��V?Հ[}�g9/�pKԔ�4���0��t�ht2��r�"�C6f�%~dZ���1�k���-Q�@�23>1�,�=�4���l�t��^w�Z��u�p���n���2P!ZmSӳnݼy����?�Y<⺁�~�3kʵf�f��p�O"K�|�[=bl��D[�{F'�Yn	�=j�J=��e�3�YR��	f �Y(�t_�����?�l����p�s5�t���!���]�"U��q)8��<y�g3���T��^}����F���7��E`���E�F��V#95;!�]��Y�ȷ�@��J�0�C/H �Ys056A�MiQo�,@�� ��Y���;���X|���(��^�bk���dG��^deh5��`�[d5���{j�`��4�!1`O�*-��h8���u��/|3mbF3]� �������n��@�GJ�$�����%U+��Z
�G��uM�6��ڂ#��ǽq� �	��3Z�a*IM��ϴF`'v�������E���D�ۦ�B�!o�����4��<H	�:&(w�#�<�ѤFき�ƽ>�� �Dm*��"�a�zr��ip�*�)�7=��$�*b5�r�;�UpO"�
�:��@;K���6��o8uTxLo��}?޳����OEL�c�6�{��������1Y�h�<��J�jۀQ�1�g��#�7����hx��4���7�˞�hz{���i���<R>������]f�'�ĉ蘪��[<�U�Vi���@k������T⾠��@�������?C���9�82�@啄�l�+P'�\�5�EF�>��JgM�e&�-{�<�&+FϨ�r�	����P�>n_ ��^��ay��#�m3U��M�yalh��F�M������i	�v�+F��`���c4�{�ɴ�,kȃ�o
���D��b�ƲS�禟���]�&�w��k�%^O����m�R���Z��O����ie�VaY�ϵ�F9{�.˯���� �`���"e-S1�D���F)�����k��hc�ǄɁ��4�c�?[Sҕ�#A+DF�c������6H"�i ��ACԿl/����^�b$:c�ijd�b�:]V��G_����\�b�#P���fpM5_D��9�]��::Q��@��OO��<�U�˘ٻ�b1���k4�BA0�ՉՈFS��QfN]ρ~���������y~�����B��G�� �f ��"�ֆz	�0��%�j���f=����; ��)7d�2?��0x-6?S�=��������\���'ۢ^�w�';̊�w=��_x~-2���ۼ�2�{�h���8hF���8�{؉��wo9��W���`��4�ES��5
�&���d-oT��Z��}b�9��r�����y������
8o�0��F�+0_�ka7Z#-Nj�L���2.�L�@�M>����YJs��W��;����Q�=ͅj���f�D76&!�k�T+�`>k<>������s� �_�䌑���2�^`b�7�xd,�	-q]#څ�f����16J��gK9�V��+�Sh�R󜸧���b^]=�Ʒ��џ�C?E��{>?2�Q,J��ɠ��X�o";�B�s��5����w���N6�Hzs��|�����R���g\���7���;��Q�o���"?CXo62���1� g<����mo�ú j	�3z�b���::I�0=5McM�%�d���1�@+C�+*M4�=���y?�喇w��?vRoo��,n���o}�篝�ɞ$�D���IG2-��[!C��p���q[��`�7F��;��-gi��f%0�A��`$o� ��`���2�L��}�G��G��Y:/�G&��;��y����`%S���l&7,��q�1����N}��Ġȁq��?�jn\wa���Yb��
�7 �4�y  �a�0����P��aR��`�1�-۪�3T�,z�3#����I�
�A��=dZqސC�L}j���f��N��t�|鈽^y�7hX���Ϋ��8�"�_s�Qۦ��5��fm3��2�x��{bμ��;�֫�P�~ƿOͱu}����2��ubWZcKGz�G��/�F �i"�~Akm�#BC���=�z��	
Iy��R�C����m��چ�i.��7�@A�l�q��	dI�������� � B�˫�w��eq�G,�'i�Yj�䴪%f$�9_Yl=�VF��2��-�����u�d;p��n�;��簆ã�\O�t�Y73���wQ���AA+0�{�L��O��h�����y㐭g���jd���GkOL�3����//�����I��{�������t�{����e�)#�!	q "	�l� ȋ Yd�mVFVYd ��_p IȰ��%�4dZ����{���U����7��νU= �V�YS�U��>��;��w.��@+�Z�9�!��z��}��?yQ�s���F�4�D L�Gy�(t�\��I[�37�j}1W��^�a�5�B���Wt��z�m�����eg5�����|C$R��=]��u�q{ȱ��0���ذ@$�� ���/�fy����176Ӎ뢟�O-J����j�m��ͦn����5����G����_~y��g~W������~��|���k��V<�J���D�4)請���8f����Nc,�5����{b]�����PsF�Ň���>BȽS���;����S���k�Ũgf#(�*U,��#T�c'!�2=�~2�ڤ�$��P�V���*�?��Z��!�[��K/<mB�j�?���\}G6��^�:�7�AO�~F;B@����Gf �/�#��΂>��!l]l$��������el.����HJk |����h��'���~�����4׋я>��P�] �
7J9�]�j��w�n%~~!��V�x����m�Q~�иe����Wb9��D;����^xT6�=�?�%�N!ǋ�@�'��1����)ok)-�|x��:����W~��At�ҥ+�be��N{-y~���3��N(��ܢ�����ӽ��;�
��-����G�k�	�r)�~A��1C������Ç����6��h�;�s{�ɼX�I!�1�� �Sx��є�2S�GKcH��ȯ�ޠ$Б]�dݢ���� �b���[<�����9�an�0��@pc�1S�AA�e�
��hL%�����J�R��t���!���=E ��O!��k�� H�jzU�a������T�<�9�)M6VV�[���?y�a����2/�x� �z���;��F���4��͕6�lz::��,K��y��1gf4��CK�S�ױ���GP�f5�F	���|4��3Ft�M�<,ʳ���Ăa;���O��"8�K�.��O��N%S�1���_<�K�?"�F�,��7���V.�������?X���џ����������������>������o�u�?����Ooݹ����~!���pcSm�L0�(B��\�\(&"����.k�Q
��<��M�ya���ϯ���U�KA�	�,�"�f54�_Q�̨M�2"�:�b�Vd<���K� �6m���(�[���J�r8��0Έq�76��pm��F<u_���
��`DT]c"�e������V���`AIS-s�~ﹼ����o�3H7�� (36-��>ڰjHR)X��2ͭ��,ЃY�@�g��	s�@ǣT�$�Ȕ3�ʥ�T�Ƥ�q��![
\��S�%�2��%-jX�s}w�?�a���HG��i͝ks���S�a�<Ϟ��/"f)�!`S�9]��޸�R��Q�S��t^70&��}�	��r�	h{�-p
�+C�3�5.y��GT�0Z�/G�䤡�D�������ηJ�L�4G����}�ôr�0�Б,~�s�e�y��x�@�7X��H�
���Tʚf���R*E���5�-R\�ݼi^}�؇�Y,�M�cF,x�Xw)J�q�>���'���RONN�	���9A*�M�c��I�Rx�>��=m�(�i�pzm�������Y2���aSY�l$�fKs}��,�,w��٬3���L)t�������(f3�@N�2��e1[���1��n@3�u���������38�&c]��Yb��F�lEa���,Z��=��p�B甇�x�#� `���2GŎR��瞰iY:K��}2=��1�<�+�N޼T�̝]���-J�Ξ1�jl�������^9�N�?��ᵓ���߼�������֍���魭I�e͠,��~[�T��o޾����/���k�w^�y~�{;@�)+��2�q-��0Z
F��(��!Xc�H{ã%&�h�Bׂ�'��V��>�S�πT�^ ��/0�a�{ay�^uk��hO�C㽠�s=z���-����g.���l�`�u��G4��xU�s��X�a��$T˂��W���ޡ�X�pvTV �a�s0z���z����u�X�+�Q�W/_��@l�h�	���O��Rh�:�P��aO�"0P�A
OB�굑�{�6�{p�b�m��u��� �=2��`�(�{��������T�Cr|��
�L)������A5 ���05(���Gg�)���bp+cg��خ2c���'O��a����E����@�4��;��q���@v|tBs��u��~,�&6k������Q��؟�ۤ���~��) ��Q׌�w2����R`'��b)�:=S!�&���q?>�gv|p����~��:�|(��ۯ���W�w����|�p�@�ޥw��V�M�5c~JY�趇�$[.��@j%��_D�'"#"�~N��?z��T�o���_�q���H����?:Z�UH�,��Tr!#2M+Pf�� :F��LӢ�H����F�2����>�ː~+:�,�r1V8F"�P���s�51.0��H({�� ���X�Oc>��R�8z��2�0�T7�F�XY���b|W��\� �s];�GDrb���0F�Z��3�~�d;6���.hT�4M��.� OY~8���#�ki�0��n�N����,R�����D��o����:[)H)� ����#�� P�R���J�Ճ�ն6�7N操���l���w޻u��[w�VW�綨rq�'�v�d:�vpx��l6�6�UD	.lf�gX��R��̼��ǅ�1cP�Az!���Y������D�1K�����wt�V�Xk��㸑sz�H=(P� cWΨK����J��5pJا�JV?I\2��ަ�:jh�{"����DWMGl�H�,�m>��C�By�����|�W�+/?g��#S�?2�G���\cM-�?��!�@�g�������k75��F��0gyW�`�j�ԭMY�t����+��A�̎;`)���޽O���ի��3ϳ�(���ԵsfJ��[�,��T`�Lw���{$��`	�z�4
��b/�tԓ �P��]?:rŗTV��3k�e�r���7+�y%��m_o�s�
 �����G��H�qO�;7��[���_��ٰ����6���AX.h�����C	Dz�2�z9�<֮��K*̜�t6��X���׎El�鍖Ϊo��e57�������7�nU��Dp5�3�0���*�@�O]}�e��UP��h�`��@�ٝ�����%dؔ�o;��Y�?��jdH�
��D��uK��a��������y�o��v�k"���a���@Jf���	{v��9,�+Ox[gϛ���_׽*r��;w�o��Dh�Xy�� ���vP c��H#��k�x0f�Ps�J!�ZĐ0�#w�_��ԋ��� Ym.�ucuC�:D����n���!�Oy|���^zq���m�/ԇ�`��l�������G��
��Z^x�=�V<?�^gAa�L�)�<��(Hx,�;N*JO���c�f�M>�L���� �.~&�u��np�ˮ�����s�EE�����=@jM�@�{t��ؼ��{�;�3��evEo�L�ۀ��f=�v]�s}R|Ɇ��^�!+d�����u�/[��gu;i��J�=��<=n��x�s-1`QZ�u��K�q�@n�3�2�9��2��f�r.��/�WaH�K��5O���4���_�8��;-�,Q����f1��^����!��s�[@�B@ �E��m({U*"Xv̠74� =1��,durL��≐%k� �&j���ͽ��'"h6.�CY�"�̹�W�_�B5g���Vb	�����	qШdg�\Y[eר��y��3qUh5P��j�#���Kf�W^}V��C2x}����xy���g X;��Jc ��V��3��f+(��q�&�xe0��2ocD �e[O��}�Øc�tEOA�D��9��@e�j���#ݗX��R�xag�:�7%b�e�@�8�0Gc5���k�BG�t�P�d���J�%X"�5t;a�����h��"C�������i���nP�.�概Y�'��Ne����|�K����u*!T�t�|{��.[�UD
0H� %�W����_���Ǐ?6��C�GT�T".^�j�����&�(O���8�tD-pb��Ν_g�eH��W��	87BX�b=`��D�U40���ߥ�x�)�֢�Hg��*���M�p�cͧj! ����ɺ�:w�l�='sv��h�!kֱ�.����`�eo>z���w*���d�贩̙�-Yk��U1�/��d>������-RPon�3�8Kc1\/?u�T��<�~D*c�U �=�	y}1.IX$�� ��G=b�6y��_0o��[4� ��w��
Hݽb%�TE���)��g�7���o���Wo����>hm����D��.�!�b��	`fl� r�e�!'�ō�yf�Sð8�z�	)���3��5�r3��}��fi�ŰB�
�3$�>��Q�(��C�Í�	rgm|,k��EHc1I���v��2�{֧�_ϐn�!Z�
 Iu����zz��x�Q�痵���gOb�]�"�4$�l�9���њT�|:
�R��Q�R��F���%�z}��4�N����@.�e�JdRW�FhJ\]^��g$�V�L��1���|C���Z<���J/ê�����ks*�;>���jϔ~?:5��j����3ċ�:e����ɑYo�yr�ɃL�V^���ѫ��\og�H�،�L+&D���LP_l{2>E�3��#�:�+�|~�z�����d��� Gxfz�P����`a�=�����S
P����>=¡F^Ę1)}˒D#����^+�ˢ� \#GAD�ó�Y�9��l���/P���S.�N"2as&����# �H���p��sd|���)_�/�tZ�����(�]�Φ�h���J ��;NSvVyP0����ɨc����2��&��W�j0�*��/�O�:��_bm<�tG )�_�F�O��f�v�'�
B��#�&
z(78787��d��#��/���j��9t�D��\�:>8�*
^����@����g9ǵ3s����Y���8<s�g�]4�/\fEɵ�o�jֈA�F֭�1*���,M!�{(�����c����sb %`R�l�S�n�k��d́����e� �˯�b�,�m��g���T����)��������{�������Fv�ˢV�va�C5[JI��B����*X�����(�9Ȭ�U]xU`cg2��}B7��H�4�ZE=<�[j�b"c��S�����1���?�3��#�z���P��A���3܉�9�l_�C>��"R8�����T�@O�1� z��M�#GH��D�9��m�8�����b)�b�q`�?�:��=�6M�"�5"�`)R�����b�ī�z:���,U:x�hQ �Vh��B�}\�p���ජ���*Rp��_�pb
z\���pa6�����`�<��-]��#��"�SΉ�c ��p�a��h��_j� ^����x�)��ը�[�^� OD#�Y/�l^f�NU�Ε?g�d�}ԁ�� cG"�0�5�C�l�$��xU�,º˩D"+���v�����4�gh�9Mo�\������8S)CM�L��]�Β, ��q����А_x
a�+W�q�c	��+[��0�N�0 +գC�#W��.`�i9pC�@������w��="����E��o�������@�SN��O5�ʆ�%��c([�q���QE=	��H��,�����n�1i�˲l�]��S9n�C	-�@�g�r�yI@�L�qC�@AeS�'�����Mt<� K�y"�(<�3{���|&LΟ��\t,��a���#���|������,�խ�4 �k�fgw�e��(f4���|m��q��`����ڤ������)���}���Y��@\��Uo��<=M���{���|��������)t_��������ћo�����U�7d�lT~��Bl�5&^Hȕ���:���FVT-�r�*�Q#�m�;��S������m��܎�3lg�l� +������% E�A���V�3��@Q�z%�qrǢ�z2"B;�Ŝ\^���_�9y2��6�YR�[܄����� %�]��f��*9l�ޠ/��XZ�`��)ߐMl[�	�[$x��ޤ  	@IDAT�kĨ��;D-�.���F�6���w�^ФE����p&� ؘ�P;@�A!b��[/�wD탋����~5�����|�Em���s �z��hƹ�]���̻ 
\�rM�2.Wnu4���Z���S2�2�NlA����GͼGj9�Br��d�����)#"����$�:&]�&��z���d̻�7*��.l�(ā�n�+<���&��X��>��=3�j�o��"WL�"�	\�v[dD���
}��~a����}P9�s��(�`�������:��<hi��[�JbO�u1�b ��cyB��Z:|ޫa>�J���t0&��W�Nl�5�P�����ıo��^�ڼܫ`����[׶�&GhG,r(�A����������/2��(���^*A��"�[z�aQ��"�i���=�Q��	V�:������K.��zGOF���G/]?k��\oQ����(Ѣ]�GN�Yb���~��a��>4nauiDN�"v�m�� �U|��t���5�S�kȽ�t�j^��\�|b�O<>v(d�:eΪE7F�7ZI������ǻZe�{�q�l�A{t�9��+RG���i? ��=*ox�0*h̰��.��΁���qɀ����U3}��>z���?~���?������+�����g�����^x��Y=>WM&��|�Y�\��V�d" f]�9�E-���,Tsm����BCcWtxm��E��6�
Y4���'�8�����}-���%�����a��E&"ʉ����񆑀���):�u5"�-)�Tt7��d� ��
�{�)���l,%�[�*��Z.�+6N��],~�d׈�e��d�����k�/E?�z��܀�~���+㉛��`'�ߠ�E�3�ᚎH����@�����uy�&�Q���v��=�(P��)�Wx@�6�u
h�]�Z�u4h��v袁�?Kِ0�>��a��n�;`��
N;��d��<:��i�؄�,�Z;hڮ�[�9*'����s4=�������@e��ڰ4u3+&�G�,rQ$a6i��"o��=�M.B��ۼ��MS�\��!P�"w��$�cG�dM3�ɂ�I�^k� ��,"�"!��/+���]jP?��^�"�s1.���V��;y޲����3yz)M�,�K|���(�:�qA� �Qs��.�j���]�.�r�FYqp��e�<���7��!�u�O'�mi�K���k��M�@��o���>/]S�e'Ƹ���!vŚx�Ӣ�6?<�ӓI)K�'
|JtVM{uUm�����uSȸ���a���G�F��\�'`���u�� ��^�P��xu�(]�Zy^�{��@�7��}��͉�rB���� �Uv�5��iЈ9+6�@[���-���D�Dޅݶ05�%@�ṧ�P �BRa�4֑:��eU!ZD/$� %B�!Z�̶���v�<������=5xRt�]�8R��
�-JR#�ȑ g� ���h]���J�\�jRd��rB�R<^`���@�4$��+�R -$�l��H�@������?��Ё-���XW��`K&������nQ���_��o�濹m~N�gV���uk1����������]�.���K;��;�	��s�U��9S�����{"��}�؝��p�-��4P��K�����p.�	�~�]�r03�3Sd��4_2tG?'b���'ڜ{t�������1%�����e{�=�U/�e�>�x��fw�Y�����Q�r6ݳۃ��0��ɇ�Y���U78س���G߬W�������L�Y�=q����=~��ѡ�x�t���~{{`�?�����࠴x�������μp�WX?�!l�^�*�f�n�B�V�A��L�F�U'k��u�1�a�N����,7�w3g��ySTkE�r ���t�+�Z����d����I~47G���$�vu��V�<Ԧ*��>X*31�ꐣ�Y)�e6�d�'������7�h�3��e�O��GS�c�������'py�s���Y��1b�&+:Q�aj���ć�S��5ѸM�f��du	}�ս��mC{U���]9�ۺ�Qq�L^
<�x��s9�Z�t#�5����Cl����Q�Y�.��@��(be8ۿb�1�2�c��m'�nK�F#�滁B��a�E	
�{_�Q'#$> �O�z���Yy>��-� ��8H�5����p�H! M0>9�����Mf��r�=0n0xD�0�I.��\F������x<�r���K�ݹ[���JN'Pృ�U3F-�idjq���pKK>�G�w�_�_y�W���7�Z���� �Dʄ��    IEND�B`�PK   %�X��%� V� /   images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngD�eL\��qw������;�ݵ��݋K��www��Nq�b�nv��Μd29�I���L2��r�H�H�
�Қ�{�^��<��9�]���r�53�g�
�ھ&����$�O[g�����]1			c	S����##��/��!Cj�pNȈ//��#PJ@B�qr�Lp��-~AJ��h��g��ֲ?���+��5���9:d9{��#��.�>j��&`�cbϩvac��]��o>+B�Վ���	C�0�����E0U	��1.*3��u/z�a ���ߪZC��{��c�/�C��/���U����,�x�.4V� �|��a��Hbd�|'G ^��*���w�~~5܏q^�7ޙ��uF���{z��Ls-�7��g�����n�5����M@�����ǥ�b|��N$+�MO�����7�ਓ�Cd�-ϐk&�{������D����AUBC)����7�&D5"��GeG�˖��O��W\�����e������1}���>L�v8G��([�D���(������#O�BZ�C0@��Cd�I�z&�je��q�/>��ە�[1�,��(��dxc���y�*b5{��8�:���)0�zGUj3N���yb��A6}�ϭ��&�Q��XveH����ʈ{��`h�(���c˸����e����Vg�wm�j9�E�����=�o0f��	-� ����~T�"���XӴM8&/��~���X�O��T꽴B��>�����<D�ՇS��K �������M��!x>����2�qb�2�;CD�=F���ڀ��įTr�����*F1�Z���͒f�?q:��kk!E���j#�>�x�Vmջ�f�%e:<PK����5�NsⲂ�Ж�t2�2߂8����D/��+�3��r?yE�� ��B6y�Ő{:߈������ ���X;��D]��\��,B�r�|н+�g�_��$z�'�*D�O]��9���a����83~�C� �j�j�;5���r�a��Ë��E��O�H,�2N��BF�x�B�0_!��_فU��7�����'0P<ɘ��1�J�&�>��A�X0_�9Fb��Z{H��c������a�����D`�i1�\����(������#+f�*L[��f�-��K;Ǘ�)���ys�	F�L��f�.�Hs���������f#"��fc�G���E����Avt_���;(�f�G�j�I7�*�E�՜��M>݀q�f��\8G�h�P2�(�Jr��nB�]ƐL3��Fuj�]�&b������P�t���+��R��Hu�?Q�UT̀6P�7���H�%�n�*�����9a|�%��
�h�WCI�#�5g��&�;R�a�$��*�؀FSSs����l֨�����TRR�]��������S���� d7�BVa�8�/�Q��ࢆ�!n �7rЙ��&��\V:i�E'g��:NΕ9�L��+w�0�j��@]9��|����Ka���A���+�&�P��S�h�3��*c]���ꊯ0�PR�Isר� �w(^u��ׂ�=���G�K*4I�\H�B3�o^r��)䦋	/	�}�/��7P�@�r3$�h�����g�TX��,L�׭.���rf��7@"'qa���-�B*y+�E��Of�Ks{�US9�xzG@2�Κ(<}���b���)��Fv*�^ w�eHyV�7
��)���h������_�cI�L���'8�g��8`k`��O�X��/kA�͌��fT1�o[}z������*�kE�/Z�����W���@�W1t9�5�s>m?~e'�U��n6�C�����I)��xN��1R,��Գp�����7�u᧰�{��y�������e� 'RC��)��F��]�sᄰ�����؜�؂i�Bb��FFѼӛ��厎�2�`T.g(\FR�#?UR�2"0�V,%��^���P�ZňNQ�0�ҿ�5��x�&�Z�1�1�_�N�X޿Q��5��E���f��ce�#�Ki!�~aW�tZ"���"��3���>ڡ�3��{�K�&WϨ��Ց*)�\=�?�;����:�=�� �[����v�
[� ����gfe�N���+q
	G�`�����n��]6�]�hCh�d{k���8Kp&?��m��*P���1�01e����xH��h�]ۤQ�	��x1mjoz�����)����:���W�J0�Z�^��h�ؑ��"�|� ���2xY��n�l>h?���!�d�=���B+l�i=��N�C�&��o��,����38W�-((���/��y�x�FP=�e")1J�~�/��>i�P�9�s9���z|.ypL�@=��܀1���( ���>ӏ*A�5�5�ogrQX/���>ܰl]#�aّ��<���̼DOG/6u���^�濜����̿���u8{�����\�o# 1-Am�',o��Ao�|��ifUX3���t�
󏼔�lL����\5�'dk̫�o���	�H[��btM���u"(���������W����QoF����>�D��GC�MJN��F�ki��+y��k��>@ڇ��~8|�gNʶ�r$�E[Y|d�2�P�2b2��b_��ԓr^8a�M��vchn���8ܼ"�á�_��{p�_\�\mwǻ���uqG�vƦ5j�=u����Wh��/UBL��ocE��N�������H��x�$>��tgñ��*طZ�_g��DA�4���}��t���gG2a|R��?����UB�eb�_�SB�f*�{��]-P�JÈ��e���y�|#]b���j��1F�b�,r��;Y.+ �#Yh����kH���{_:���F���.�"�Ɨ�иfӱ���o���QǑ>�w��bZ}�Kk�T�J2�l-��Y�����Uի�L��w]���s		��}+��ӓ�>��>zv��L9��Ug��V�*B���d	�+�ڂ�� �E��f~A�?�Z��"I���_�[0��GFk.����X��&��R��Ieƭ7�{��lI�F�ǜ�3LM�X�;�)�>���{�V�9ԓC��w�s��,��ڸ�]z�5TiaR�9�*�%�b� y�-��1r3�?�A�!$�jC!�����"�
�����m�ϋ���	��x˫~�5@��W>�P�꤅�Ռ�*�d�eW0Y@����`t��T���/=������|��u)���\��
cl���/�_�C)��y^~I)�:�\��>�f=q!@��O-
��*�/��PZ-�ݢ?T_j`�`�<�u���)�x����r±n��x��t}��{�c8]�9�2 ��c.S�S5 �ĨS�x��,��Q�΄��?���e~g|�<{�9��$4��/!��~�����������,��4��W�vh�hf4�Wb�8EO�1��<�������c�G���CHM%Vgrl�BQ��P��^}��WP�����Ы����`P+��~�r�ŐR
N���2�`]���@��B#O�Ex�*c�vv��#��a����=��/Nu�N|N�}�~^ �ԫ�qp�|�V�,<ĕC"��Y�|Æcv=\!,
�w�e�	n�����-�5B��8����5������C��*�!����ZZ����,����H3!�9X%�w��f<~���U��Ʀ��0h:����y��ף�s�"\2U�]��{zP?��#I*s��L<�̾T.�r�=܅8g3��E�����>�k�x=\v>�B�;S�3����q̵>M�]����X�>>>�#�9��1x��#�m<�!*i�j�/.�D�����B@�%	AM}V����1	vl읾X�E�
^^I3�<t��wN���JgR�1����Kb��0�^�ܠ��(=R�=���M@��wt�r��ʅ�Q;yd#(T&%��/������b�׈si��1495r�����I�_t���)M)O).U�,���k�A�� <�և��^��� ����C��#�L�[��f�+Ð�<��'c�7bڸ�&�^=99�����E���H=O͵�>���e\Q{u��l&f��Zwc0�an�&b�P��U�X.|F�"��'Qb	u�^Ԉ^�'<q������������J�?��ʗ�	�Ȁ��OlP�z��2��_��Iۀv˒��2"\��g��.�	K<KS�_�hG���wn9���y�������B�²�9����-��N��dR֘Mw���JR�`K)����K 1������}���9H�G=3�MzsT�U6S�_�h){�>��l��͋j��{�\Cv+vVA^�+n7���H� �#�t�h�������ŕ�2q�$�P2�h~~�\xZ�����p	��t	�(q��%�&��d�߻�iW�.x���^�<�V��2ֿ�8�`[���mc�3��e�e��o���⹾�#�v��"Nrjj���b��`� �� �q�2�+��F��1NNrk�L^��;v�@l��o�0��~Y�����96�2�B��������ﮬ��/$80r����-P���N0��\�큪���^�bM�T�P�﮻�yv^I���r��%-�}jj����.��`�Gx�@n�aM�зg8'�5����(L���࠸����?<[���
A�GCd���W�?�p7��X��T�`D�~�D5�#*3�������](Ϯ֑c�A6��]Sc�����W�������(Bÿ-ѧ��m55ˠ �<V�\2�^��+�����ڴ� �hZ�%�0�1����o�$=āҾ�yA��>c����K��9��۟q"�:�NZ����< B	�4n���Bػ�^��z?�Voj?K{CnoyU;���}�LJV��卒m�5Ӟ��	�-������J�z�G�,!-�����l�W�(~h��JO̭<�19�S���.Ȯb�6���Ijy��'�
�0�^N�"�䜖�إ)�IL4��`� q�D��[g���1��,���Q��	*�E2����������9�2�V���g�`��nn�c�R9q�ɦL���P��c�R���;RQ3mˆ�.��D��"gKd�F�>}�+��	}q������zf�]���@���GDR�̟}����Nf�,��vl|E�MS��U(��3���}���
�G�����f_�"�ʔ�h��>LM�����#�fNF�Hp_Yu"���<��2��`eU
�`c�&���584�Q<�\��N���heov(jR�L�B��@]�'�<SW#��7,�������n3��sJ5h
G�be6�����O��]�XJM�5j�	�hh��jeU�֫;��*@�9�ޕ@�I�e%̩E���i-U�N��XZ��򔯑��v��S􍄆Нi"Ź�0[q�VԅJ\���:�ߤ��*�PNV+�� �4�K38�!fJ��iI'�$I���D5
x�x��������;��@�ǌJ�N g6�f0UӮ��<�!��O��j)�[M
8yN/�ҋv���Jlm���_�9�� ���lg��A��������#�O�&?�I#Sl�� �.�_/�!l����|�LӴ��6�ֶ�e����^I5/./c=�~qr��(�o/֑�'��ɢ� ����?��h�㬈d�GTǝ�,�������M� ��['=���}p]H<H��'~L�{����U�_M|\����y�����>������L$�Y�����\������6��|���ꦒVi��� Geu���^�����jvmfjwV	���@�s��.y,HbE��[��K5���T�J��c�!�{=�=�G �c������@7��>g`�]�J;f��X��X5u{��Jd��jo�����VJ�!����)����]����G��b����Şq��yx��Ơ<k?�j�e��+���g?�\i>���e�X�m�O��y7��0�"��cFɨ��v^󰦜�r��a.Z�'bUYjSfP���.&�̢̲��r�`�O�Y��d�eY��V)�q�	S��}��Tkf�����wE��k�_�u��Da��=�v���Z��P�k�w��ޣ��nf�^��ز1*�dM��#ʃ�,X����WO�.�O��
�%�'d���kq}��Ԯ�,���kV�\��v��iN�
fE�ld�\0�gY��,JJC�t�U�����P�y�~�m3!�>!�N�j̬d��jH!*J��C$Y�Y�~ւ����=�,(ɡ;j8�z3�T���F�� �����ìKO�-Mb��L����w�+�-��L:�9E<2"賨��"�[���!v��@��,0�;D��d	(�3�qF���k%�7��8Lg���R0�HE���������a&�}66�a� �f��sq%tEϮ~�;�H��$�1��*��%�����i�k[P�� �:�ˢ��	�p�̟�<�]���ћ��F�R�#�,�!4��Ѕg#nکgB�Ǆ�1��6�k��JU��g��+P���6U��`#�& !�,'L���M(�H?�&y�o� �_��S�,�t�#�kJ9Ws�2a2J���ڵ�eE�igC=+`t̃�|���l��P����2��$c�9B������D��� ���j8EʽU�7��G� d�E�Ţ<�5��7��&Sb�^���y��9�V����˽��������Vx�'x�|\�߫h�����0�����෰L���*�?�~s}�}=�哽�|��E|E5�u,s�����-},��������kr�;�vT�h��(!=S-�>0��#�gll�沽�g֨$4B���9p���+�$<�n#��&@b�Cր�7��}nl�i���ML??[�`��5�{>��>�%�P�ƯԬ7/ ��ó��y8�,`�J!�'����lj\�c�����p�z���Kc�ˊ�LU� �S��}�l����9q7Y����I��i~'@�B*it�j�N`jÑ�;�}�7$Pѽۆ7I:���a6�e�g`C���Aqإw�!H���ƺ52~G.L;?�*
�m�v�
�1*�{}������HK¨���D$E��Ϸ�HB��̩IIH��%D��v ��.�iό�1#�9ڍ�)�h�r|�	��6��0��+��|#�o����"��}o�=��j��@Rs�T[Nm!�R(d�Ij3s���7�6أ�ekbB�'�d���pLJ��d���ϳ7���q 2?$��rx�+�f_b�ߔ��)���0c�w�Q�6s8�tOsj�Ec���Li�<9w�yf%���k"�C�[$����-)�rr���|����:��r> �{x�O��L����8�)�=�z4������l���݉�AOҢ��]eM�&ޏm|| �|���r�hj�r�?)0�NOn��G�
2���W�$���G�%Z����>cO�f�{t�.P�­�+����p4Ϙ=�� �ue����Ҍ������|�ɂn0mlO�}
�X�dx�%��9�,� �_ð��f��\R���lKl���dǑ��+n��L��x]�3�A�Jxr����@��BN����@B|wM^D�-����ѥk	JU���ؐ��<�ѳ�&��y�kp*��M�i���tt��T���M.����������i!` N
�tj��NP?ص�{��?/0��0�8�o�]��W˼��������'f":��/Q~u,��u�|"�s��8{��Pm�I2�w,��?��L/�p�����n$((b�]�޿��gLx����~�3y�ܠ?��A'�	'�7;�q9a�C쎉���kaÈW�9���-���z9A9���;�l��_aa�����t�� #p*0QS��*X���Fc� w��CJ&)
]���f�
���W9T���7G�K��7���G�/L�>?lU�|�<Y�[�a/eC�U2Y���D[�+�&t�O�r�/^�:�)��o����_9g��̆b���b�����������l�b�2 |�'����
��F�J�� �=��%3,*�������$��Y|�oҮ�n��[�D }��\��h��yC��և�IF�����{?�**Ȥک�M�o�"^�k8.3Ӗ~���`T��O�u;zGێ���?�0%����a�t��:�̜sp:��O�$��	���j��
��栌�T��3Œ�>�~���W~���n� 0����Z��Q)���ݣ-�rY�ɵfR���=����|��/��~r��<�S1��V`����r�����R@H�����vls<OB��Q�f*:JZ|m_��zo~��I5W�A��1kXm�M��W0m��M��Ps jB1Ϛ����O�Հ]J��_��uuS��)�Q�l)_4���ccj+%"nm��з���D72u�R����tol�RPBty8+�k����ā6�V0H][1�!����M��[�&��OD?o,Ǔ��	���cV���U�t�3㝼��Ҫ豙I'��U�^����6-;�S:�ݴ�n���g�ͽGN�,�C���(��>oUƲ�����eU�/�~8���<l�םVNl8�P�r��v�J�AY9C��NZ�m+�=0u�!�ɕ�zp��!*����mXh�*W{YB�م�k�#�;}�q����t�T�2ad���������'���Aݣ�Ĉ_[��S�y��+����ý�7���I���{Re8�s/�����,kq1�{�GO����pa�Rfq�����K}�^��4�Hu���r�qb	�o��#�c2&�_ç9����.�18���鈌��ʔ�X��0ڳ�u~8���i�5Ҽ�k�It�3¢�M�qJ]R�L�9��P饣������qE�Է��ӫ�q%!{]3[23�FB�F
�;<��	J�@��E�c�)�(�d߀b=�^�"e���QfX��j&���!S��ݾ:�\��|?Q���^�3�UhzIA+��3�1�9t���ϞǛ���p?��o�D�;�:�_	�.��記0���:���aeej���g���&F)���#��A[
J{m�	��]���I�e��b�45%=�|�	�<�?e>>�-	�V>>V%�L�
������9��A��~B�Ɛ�Ϣ]����3X@³�g�M���`#�*|�/[��c��pG��6�ϑQ^��������?h67�	[4M稢M/N��qgϮ$K�h���=�η���\��\���	�v�#|xݚcm�w�P��b�Ȫȃ�zS�3�NW��1�|����b����}�*�u�;����d��3��H�|�SD�j$&ng^t�5V=&Z�����0���1B��*'�S9)��AmF]�k�W0C�x�,�Bb�a	�e��U���F}~4ZFtQ�K�Q�Q���i'��"�T>o�3�m+k�=,UJ[f/Hz���W
��-M�����fA��K�Hiȱ"�i��`�>�qr��X;��Yː9W.�u�mA��7ޜ�%[��ዟ��қ<�/c��?�G�,���^T��&C��g���e��:�ݾu#�����ꅫ<Ui��,��'
�������
�%~��^�qM��v���cj�9lJ��,'t���d�N���U# >΋�p�p]Vk�Т�#;M?�b�OH4:�BM�X�T�\��S�ŞZ�;�51|D�_�L{B�\�tQ�K��������ڱ�K�1��Դ«�[*���e�f�����B_�����&L|�7���@���7`������FiD���~,Sd�L��@
J;�?U�q(w�V�G���q�-c[qlL!�jJ�17�3������019L(�^h@AXq<�%���$8O9�����>��1>����PE�1���	"���>��3��B�r���0*�ə�T3��a��(O
AƆ���Ba)l%�Z�Y���lp![�Y^T���:+Ꙙ��r�l"ٛ��Ԟ�,�uH�,�q��{+�����i�Kd�qBDU��.�k��- �"~�y�5����Sۇ��,]��(�����~H�l�}�M ����fB *6�#1)I�]�n��[��?�{kS�z;,���w����F�����5�ǹ2��\�XE�Z����j^��F�N�6^�d�����"L�r� S~���-F�kj�[��M� !�Ďr���߷�F�9�Q�+��-�hq�Q�u�8^#�zE������Vʜ�}@�cB���Lr���p8��a�(VIhV�#7�z���q���E�ۃ{��,���P���Q�T����K��e�A+��4��y�����B{�,l�S�7�����?ڰJ=��M�C^��f��ԙH���w�z��n�5TҾ���z!1?2N��?4ax�$�ə7`V���҇]��ȍ�8��"57(�%�CT�����L3yka��%�7p/�/JA�X?�}=$���H[y���9ƴbU�ۡ�§�RE,�y/~<���㔜j�����1�
��f%�C��*v�
[�$�j��>N]WGc�{�*���Z��c˕c
�3�K��j͒��=�l���M����x��f=2F�0�$w[<S��$��E�T�(t��X������f�"��a*��x������X���tK$n|�=��@<�.������l���q�|�W�;�)Js��:#ԅ��c��'�|���'&֎ am�-���@N�6s�IN��2�r\�i�T�A�lӜ�~�>U�A��)�����c61S��,��(��h�u�d駂�MY<A��\�9�R�
7s���F��x��M,���2.��Ur��x�.�5���w-3���8�ܿ�E�+$��e��q�c��F���2W�@�۷e��s��/Yq'�x�wq-�1��ҵĖ�����(e�|�έK��{uH��l�|(sQ�������k�΀
ve��=r[c[��A�5��#[]c',ׄ����qg����T)�3�f�t`Ѥ�ɝ����Bب#��zcٚ��дޕ�K"����Xɚ��@'���.��G�����0{DzI�����Q��TF����;��.���H2'~F��Ӷ�O���Ϛ��Hx����b�oOc�/��W����ӄ�fv/���ڨ8�\�X=/3�
ϵ<���&� ތ�:o����:�o6(H��=�(\�e�&��\GEb�Wݬ�ܯEg�+���?�����QP�����@��!��P��M��c��g��e����Q��y�*�
�S2�ր%)tT��ǔ+��J�����+2��4��م�q]X�0Z�ݿ�'�}�	��~��	*�`�x�4��W�o��~��+~�:Je���] ��i�:��*߃�Wܽ��L���1h��:osO�`����ʴ�T��;Qx��(�.d�W������6�P:��eWСν`ҏ�(L���#�8v �ˀ��`���{&�+���Z������ ������׏ذ��аu�R��U}���JD+7+w�@k�U#n�x�A��xL�;F�V�g!a��0��XWۻ۫�� �;}�|�	N��s<\����8�7�@UqP�_��H�]�g%���;^�)�3�����_����=���ٝ��Fh�3���|���2J�{Z��H^��0��^�o���H���S0��L�8����Љ(��ɲ��	���+��m5E!R�(�\�dp��'����t�)�4��H��v����G^{�x�㿭N�'1�i�����E��D��B�X�(�G�s�e��t�ԣ�*Mg$pL���N��۳JC��͛���ᤸ)�L�R	Q)��2��p+�<4{-�S�j�Ɐ2FN���^g��;���b$6�NO'�G�`E���Gth���ac6w�1\�\��5��ZY�S��y���r�o���G��*Ŵ�e��%�9 �W�:x�����vq������m:pwQ�=.�L;5��,��q�&%�?L��W�w<EL���'�$z���
��ԷS���O�S�nC)�:�Q�#mR�P���L�5z��Sn(u���o����5���>���<O���R���L;m�rt!~�c��Ś͏�4�7���S�;F���1f	M^��uw������(K-�������.���,Ew�YWY(�Ǣ�d�	oЃ�
��\%��z{�=^T괃{� �DƬn̪���n�?�ڀ7��c��{��"�p��J���O1Wf 1R8F
�m��9����Wp��\R�uJ����ӣ[�P�soh踠P
2�38ԗ�����(	���{5M�eK�O4�̟ņ���O�Cq�YԴ��SS!O�U)>6��l���O��rϝiR�-2$�*�p串0��a�za��{�wN�q���j�2��<���L�&�}z�`��>�}z>o�N��m?V���8��}?���`a�H�ɸo�|nxEN�������O)ge9)h����Ǽ��)�����͌ZR��g�o���K�k�P;�̸�$Ƅ�U��τ��8P�l�f�;�S�RV���]7��Tl���XZ8 �,}b�|��|��7�~�w����+�n��]���ˍ��W��=�U��Ǩ?$@\a��.��4��`K�Cl#�7a>��mn�<���r�j��A��ck@�������0OR���Y{A�xS3a4֮:,^�?i�3���.S�T��~��S����Z!��mB}lM��F҃���l��$8Pn���2�rQ�)�J:�ȯ�t�K�q�>g��)�)�(�|=7�Y��XExI��s�	C���J:B���a�>1N�P��d���}Q��s�(�i���Xˌ�4#���T�? c=�|��stǬ���}ڏ㮵Ӷ�o��Wɇ��I{�<��X'޽`Tׂ8Xӏ.�~��J]�����e�S��0�ۅZ�����E��w�k���&��m�&g� 6gr �zQ�y�\�L�3�Y� $iMo�,iP���
�������e�DgӨ=IX�8%�5T⢂�gП{�Pr4��T4bd�P-�}�Z_Z!�j��"���s��B���^�>=[�����hY�{f�̈�ĝ��W,�G`�������j�z�� ��=�'�����PR�������Z���S�8㫵;al����%�zJ,O�3v|w���du�M�M		-վF+��|��Av޴
���]��V*)��>n����l�Έ�/z'z_���z��.l��_j�wIp|9�|��B�F/���p�{�[���h�Ϊ�J|�/�� �����[B�Ed(���D��ߝQB��p�]��&�'̲Ѭ��*��C~Ǆzf���4ヱ�&̒z |��G�9�Oj?�^;��e%^�}o�[EE6ޅ��.������4r��h#��f��t~�n�}�|��;�"vq�w&�������ǜ�N�3�V��>�����F�L��<�n�|r.�7
��9^�8�S��^����ґ�O� �4�sO*PZ�2qA�lY~�߉�\���F�j�B�����D�ѷ�H.ʤ2�!��ųI�]/�9J'd�$�Gz�;�K�W$�KIj�ņ]ȝ���/��hH�P��x IF)�~���6~�6B)q�G�<��j����'%a��
͒���^��<�3��9%�]����S����%`�z*��Ӹ|9E�����Bk��YNJr��nu�7����|%~5�<	Nxâ\C� \em�rw&�g\'��$���-_<c�ωuA$���;�KƲ|��n�Jh�5����
��# T�i�#����>��l��/'K"�� �) (+R	5{ -l�#�[���}f�퉊^ <0>^/�[76s1p�=�j�9	)�-7��M*����+���?��-��%6�~E����o�F�}`��H�_�����~��N ���>�'6���itNI�KB6���3�<k>ʖ��/�1��R-ͯ�-���^L�ӎ���v��4����5;x���'FV�t�ySR��!e�"�5%����U�M�r�3��$�g��3Z�p񄿮('4[+����y�%ڞ������fv��_傭X���Ҹ9�Ӛ�����jE��a������8x���B|����n�O�Q���E� m�r��sc25���a� �d�	��@e@�
��D`R֖3�{�F�Q��@��3T��E�r]р2.���$���BX����9�еM��!�/4ƫ��I��#�IG�X�x-��H�0f��_J�K9���L�Fv�	e���#%v�ǹ%�������Sw�r_\z���g�EU"�EJA?�|Nx�s��qq��!m�������ϴ����=W������y�BR��ZG����196+���L�{kR��_��/！ίpW������o��ޏkI8aN$����i�f�#�Cت���𵄣3?�0h�%��Jq����5
]��0@Ɩc��(��}��%"E�o���&ι�D)�m���M��1q�[�A�Sl,��lݡ竵 \�:��p����C;�7�0�3;���F�o\���~I�����q��6�,����$��ٙ����흷���Z��~[gI�=�*fJ��� �"�J ��5a�rU�M>�ϗ�#����Ŕ��`~����og�~j-fg����)Yz��JϢ�2�=%���{�k��$�W:�4�f)V̫k�
1�Z��%ª��,xs�H�o#�qZc�G*#�z�~���*Bf�TZ�:��5����5I6�U�/�|
H�me�9і�G@��N�gџ�|+�7�}�&���C���<Ӿ3��*�yd2���lD8R,=6��Q+EM������q��=��a�b�MƊ��06@.C�o!��t�����N_v���Vs�#Vťw2	z' "�tꥏ}��%]}F� ������#��ڨW �*���
}%h&�JP���s��0I�Vtж��nKDjG�lc���x0麟��:4obd4|�L�;O��QG��*%S'o����Ǜ��e�+R~ ؏�8�=�|��6��5����ڝ��߬J�Q��R�� ['����p����G���E��a놢����Ze����l�~U,�f�3�P�|��3�F&�  ��9<��Oj��W�e?#��Ty�<�	�]���%�y^��pgc�U-LO2,M*�h����\{s���\G�]�����qٖi�����X����{S�"&�^�i�PNsIޛ� ��x^�@��k���[e�g9��I6��N��Wo��3N���_ⶢ��K��`U�$��TV�� �v[8^w�_8���u��F�rَ��~���6e��;,���nv��?��bFF�o���s����!��}��e������D|W�ӥ�m���d�Ad�d�p�L/:P�	I�_���vs>)���j�.�!��OX������,����g�ca|��ct��ac��%�|�K�&G�Wr>ߟ�+���`�8�H����j<�D0�ť��rq�7�O����v��4���(����u���9���ﲁ�~��kA�s�b@)�qE]:`�5��܎,�gDZ}�5����.Ѩm>;��,�G79�Qr6(O�fR��/Rp�_���r
�PC&�r��^P:F&*l��XF6����+�L,8F�G�>�"
SO�gw���7�[��
eFy�<�l^����>�3j(w�Y�x&���X�%���N�r�!!��6�"y̝���zt ���6{u�V���@�)�Y����;�z�b+�w��ͱj1O�ߘ��[�Κ�)5=~%��OJ7c��sE�l�>�j#���\Y��"�F�^K8�z3~S
~fnr�c��V��in��%B����m��{�M��cگ��֫��ߧ��}h��J�VO�!��ۗ��� ��Eְݵ�f9z��V�w7����"v��8V�������Tר�6�ϙ�%3<�>���Z]�O����B�h�_��\єm�.���|��<G��`�2��ő'q�,�d6z������FVo��UXc2���dۣe���IN�LK�V�ʹ�6إ����KU�xA�6J�m�CY&�|x��"������R�4�>4\��ԥ1�]�GVhhAo�Ԙ� �Af�T�6��c<����tU3����g�7��SQ��oF�&����PԵ��l��4���F2^G���g��K�Er�/z�a�u!q�M�"<��z)q}4�ť�Z+��37
qf	}��a��\��c��n��谨^��	�;�fu8��h�b�x�Rc�~��I�I��#�L�VX�g��m�p@����K4�MC��Eb���:�,@ӿ6�u� ���`Z�):������"�H݋���H^ 9q��Q�	&��`�5�bcc�{o�p}~���53�ݫv^�FA�o>���W����y�o)��r ��ǐ�|-�Ģn}�UZ���{xse�Z$'x��x��Zm���Z��	�i�ݳ)�p�����2�;e0V�F��.�d����.
f��㣉e+:Fj,e��eoIҳ�t�������=ɝNNt�N1U'S��9��>p��3<z���?����|�ҭ���}��?����p;�3�q{��"�����ȫ�p�晆F���A��շ���;Xi��w;8:ڋ��D��h_k{)�
��S�17$�1�3b.��r�0~K��J��<��|w�x���k��s��{�Ê�k����d���Jϖ��p�o$�P0�@��M�N��u�i�����%��e�P���JfW q���',�)6��V_�Yƿ��o�fg
��s�:A���*+� i�ű�]q\�JCͦeS�F�&�.��~�+��U�0�§l��%����	s�K�Aڐ�,:�� R$Cʜ��d�a�/�H!�6ġ2?3�R�E�[�?�N� O�^��?�����ߘ_d�1&Ƅe+)7@��ZM��P|w4Jc�͓#l���������_}�oߥO���}|������&��h�^�an��k7�ƭ;����Q�����ӏ����.^�����}���QES��HD}Cʽ�s<\��|��c6�1�L���/}��V�������x�⩈�H-��;2���M�#IQII�(���Y_��DM/��ɝ۷�0=/sh{G@��OޗyN�����7�ǾU�R�#�l��Mq"�9J�q.ݾ�\������4;����������O�;�P}�� ��L�lVAmJѱ��M�UQ�.b��1
)�W��Pc��p��%J�.��mafV@�^!CDF�E�et�뒖����"o{	��rIE��AP])���I�?�@��"�T��8��z���E�.�Y+��f%,SbG+6ݠ#^�D"�k�QmT11?-%v�����Y��&���q�3.�T���6�HS�/��3�	(k���HM��JEk�Y.H &+qcq��X�X����[�Q��|g�����Z��;�0�'��8j�#�?0hy!��x��]|ia��&�O���'x��!�J�f�)�d<�V��Y��;s�R�m��s���[R �'}���Яܑ�eٌ���ʓ7PxE~���� kTi巽�/[}�mnIYgbJ_�Ru����zUz�����V�O?�ç�0�8����x������|��w�x{���&���U��ʗ$=+��Ə |��Vg��������b�����/��`wGr����9j�^U
٨�s�5��7*�WD!)��b2�ڹ;��᱈�nݺ���x���BG���~�����%HF�c.u�b^������Ө�dcoWG|��¥]m.Eg�r7��{U�u�-A�)�D�
�Y�J�%�X#;��]���y�Xlt�[���>�v�1�w����n>�.�x�F�/�gLu-�g.H.�z��@���Ѫ��(T�X�3#��#Q��z،�]�8�B{����� ��Phl�z��M1�e#3�u�(���0��)��^�|�o�ۢe�f�1&��#���kbCQ�*W�B��R�s�
��a�`W@x��������krk�;����P��&*F�~��ﾆ�_�^�vY�����)���q����^��o��V&��9"��I��i9�8($�l{=}���S$A��K����+7o���ma,=����=��e��jbnv�SowDXEG�����4�,õ�=�v���'�$�s���"n^����i)k����ǟ}��}�ؙi��"�T�������"r�(������X������Ա���Wp��u���%b��'���h��4��� ;�ڝ�2�E+ eo�Bp1����iE���ʨ�a��s�ٝ�ݷb�0+=��73>)LA��c	¼�إ7s�E�wLU�X���2.�sG���*�d�9����/Q�")Z��Nҹ�V�./�u�:a�XJ*4r�9Yj%&�'�bn8ϥ.��ĴKa�{���X����,��W�yݯK����J��R�K��2��BO����Y���Q:���+����_�[�m�FA�{��ş<{�_��ޡ�>�KH�R�@h�Qb1�EX�����k��ʊ䋲�1�~~k��j���Q�F��EU�҃�eY���s�w����d�����l�|؅�r#�(a�y�(�/	̉��/��zc����_v���|�5����1,,-�Jz���(�
�5���q��S���Gx��48x�7p��=T�g��Ώ��G[/��;B?*�y������կ!sudai��@c"� |s�&�77������S��D&s�|p�Q�����"���0�i�]�:A��0�v����%gn߹��[74��>��O?�/>�f>�)˖���	��Q\nsǎWe�i�+����M�%">O�^�Ad1�(KC#⡂�*���� ���Q)�O#�F"t2H�1G�41��߸��}�_�\��t4ċ'�� �Za�N��"Q7ǎ`,��p��iI�P)�o��G�p�\)]��z���I��NGup���Y_�n�zP5M��$N�gFãL��)��(da>�����ƥMcbs�..��7���w^����w%��3<|���?�v~'���0GUk�1=>�v�^�.���xnǌH�E>�N��rw�,í[w�ͯ~�����o\���w�}���p0�ݗ�T�V~�/㛯��W�]���?}����\��wn��xCꚛT~e$z,wR��v������&>{�[g=T'�1=�,����n,ߔ���/�����|�����Ot����;�o���5TÊ�27yi�����:���c<�B��OO����5̎�HZa}}M�����H{B������,�Z W��]'�D��C)���x��)�x������������>~����?�Ѡ'�R�����ƨ��+K�R��*���>�'aJ��]E�Ϲ�K�7�'���Z|��wt��YO���F����t�ũ.�0�h��DU�.�K����.M"�n!�.��e�t�*�Q.�_>�B�#_�u���G���a��YJ�ؖ�cnn퉎�_F�q��TE@�u+��c��v�m��T���wc�%�R�{�s:\��>2�,��*��Ca8N�4�JDc�Ǉ���r���^�� ��ߙ��������?�y��&��ȉyʪ���&�6��=���������Ǉx��'8����̔�?�dG'YP�V�fi�A�/��i�ab���v��C6�Nz��
��b�@�>7�	���J[��h4[�+�n����_�\Uc������
)�8=>������_}k�{���#|����/}I@�Uq�;·�]�_{�ճbÀ�	A�Q*"�!u��Ғl�Ψ6�RV�'��	��u�y�c8�X�?�	=�\rzA�f�T�2��� 3�qܽuoܻ�z�"*c{'��@[��e��۷�`��u�[�{x��g�����vѥ��%dk��격�l���w���h��r��[��"�&���*�"���Ar����t���I���9�*ǖbh߉�F9t?�m��\�����rkY������;[�/o��cY�_���s~�s�ꜧ{�gv�R䊂iB�HÐ2$Ң(C@����+ئeS /ŰK���ι����bW�^��8����K�6�U��zu߽���s>'���&��.#zflP$�"��!�6�"�L��u��j�O�Kt&��h:��K�es�Z+�.-	+%I��<��ӧ�Q�͝��M �	���� R�r���E���¹�8s��{��O��l����U��'?Lgk����2��'�	Q2%���_n�Z���2�ss ;���<��s�"|���;s^���{;���WX;�A�Z�S�}!�WO�U�D9�ƣ�����������8���qD�d�r%�A��U9U$D���B�����&�w���t� �;��edd���'�����󧂌9-1�fx`gO����,N�$y�7V�ƽ������m��nbsw��2C�`};��X�i��c�^L�(dt=��BFA��Ē}[�&Q�����k���:59#�H,���[���-��P�dh�	�_��]3!M���m�7�AL]S��ߍ<ኚ�N�t�ku�M#���ʲ�+�aC
�QS�!Q�ϓ��0���lh���#���֎X�6~�JM���][;�7�OS�L���Ҩo�1+���zk�C!s�C���ֶ�w��E���y���8qb�DDA|������җ[$M:��:��Dc�Fԇ�'f��\w����+�0}�e�䒪�侪��W����&�jvwD���Ӊ���y�����Ww�_��k����j7]e��:���khu�s�.7E4���1=8�S���K��I���"�v��79wht��#
�%ȋώ�'a|,�v\�XkT�n��iw����3��o��EN9:5	�_ ,8�A��6X��_���I�t�B:�b��R���w;W�_�#��t��C实XX��'��"��m.�u.�2�[����������fL�*�4�ov�wֻ��<�	_X���R�wo�ŋg
�p�!&B�B��P�d���c(�f���A�`�$pSn5q�����8J�9Ұ��q`;}�;����+�V�bp�A��ӱ;Er�G����Bh�d���R�,x�2�0=���_K�df�y2Y�ƎٰO�3L� '�b��KZe�)]ˮ=:�`$!��\~��E1��������T�����"Ѱ��:�CG2�~켻�%1>:�X$����+j45]7jU�\��͇�����6窀;fD_P��B���qŊA�%a4j	��F���LV����!��N�<��'`��ID"9A���l��ǟ�X��F��� F��Ba��7٣$%c2���[�*��70`d/�Q�юɉi\9}W.��BO����s��m#K�%��M���Ϝ�;'Oc����#᧋pp���A�s�,�F�eցvC�8C�o8�9��͹�G�>NiҶ�h�#�皍���Óh����Wx����Y�#� �Ο8���Y��^��%���'$�$$V�ɖH�\�\�rUu��à�J�8���=,��� ã��#*М�ɂ����M�)�))Y!y�Huۇ��e������/���.���s]W p��r���D�{���ޚ�y��Lk¢D3$i�š�/i]B���? �\6+�U!�G&�F�J�AB�\��0Ƀ�Y_��u����;_Ci�q�=�"��ςd~h��A譜m��ș�e�,k�[3Cuh�T<ɴ�y#�]u�~�L��u�s��ldx}�=��'��8�/��p�AᗫW�����&q������R ̀�r���h�o�C㕴�i2���C��V����V˫+X��p cã2�3�3~����^��w������g~�Qs� �X�(~n��yh9�M5O�����$�F�џ��R�a��sl���C��͉�9N
"n��P��:8����ߓD"���E�[���%x��ۤY��M���M�i����&঱��`H���ju�k����1���o�!���b��ۇ@$��?�cs�H���/>C0���y���#�0��w����ldS(��"�IX&!$���a�}����9�E�^|x�
./,`,�@�p�����z��ƣ	��c~|3��z�����lEӮR����l���#<{�
�٬����D;�C�|p�_`��l{GP=�G��0���`�+���0e�*ʘ+82
I��Ml�Y��40+B�&=�����{�IL��oeKdf�h�l�	��.��q�ǯ��!�=��l�����g�H�>�����`�l;�rP7^��Q�4d�879���1M"�Bmժ���i
#�6궝�ϰ��N;��6*|J�.�~���L������Ôdv��_����~�I^������^�����66���F077���i�xѓA�}?2��_oয়�DIJ|Nȩ`H
�\ȝF<y?'���8b ���-�l���{ldO��Ջ��5�I���74)��M�4~����qe�$��QH�����{x[{k89?��ΟW&Q�.�������C�6�ҕ2�D�B!4�Ad�Մ����I�k�מ��ۚT�~���&��"񇥇���n�,����(I��a��}�u��&����T."�:���m&{�k0�s�͸��P�(b$�xz�
���B^v�l��>���C(���f;��Bٸ�p���O=�ܦ���F�b�\^(`�V�n�T���9��"������i��w�8���KX^^F�莟{Ә^�����[Y��&q�E�"kYzZ��l1����B�,�q>Z�o�WƮي'�&ӷ!h�N3	�D�>�&�k}pp��i�B�:��O�8���7�#�����sq�I�Vʨm	]%:����	8�HH�P���$�	��O�e5��dz���QN��:V�^ck�)b���ȟ��ƌ?��-�����ɻ�k�t#���{��'�%у�Z��y!xஶP�ˠ����8..�cvr�p �\�˯���9r�i��O�bz|B�vn�"��#u0��}�'���с�UC�^�$,Iu�F�e�	$}�A�٩�W3�mf��	��n�����XY]��������S�0����x��)H��o ��U{��t���?��X��g����9�gw�Ƴ�+X�$�",���6Yd ��b��&�^h��� �6�.>�t	�0�L"{��;wo�ٳ������1>0��pjz�������I��b��d�q����=<_]�Q�����}�ҟ*d�ŭ�����J��2��-i��lm,��h�lHÿM���ے�y�s�w��z݀�����z�r̴*I���룍�Q���#�C3iX���wg����ʼֹ�a���0��+��}eVW�����E���SSS�����+��!����4�Ƈuؒ_�]p��Ӫ��'>�o�ږ��N�����|A�Ʊyk5�b߯,�as{G��p�_'���: �.�;�4_�l������=C�*���!��"S�`}k_}���"����h��%�;1:������)�`! "Rn5`�zU��u�{]�����sp�8��Γ���w2i���r}�(>8wg�1C8����{7q���X{�����˗U���gS�<��ӻ���歋Z���l�<6'Z� Z6��8��$z��D-����'q��-��F�E����L��!%���{D�D���ޤ��T>��l�`�pDB�É5����{��Hd
S�؆�f���֚�W,`,��.�h��$w�$��s?;9��xRF���
}���Ѵ�P*DCl�X�Y���U�U��d�U���%ɈiWl�H d�4��y��Ǧ�>_73�9���'?�	n޼�X"�P$"�!:��$�,3����h2H���lk��oMÆt��,����4,5��G	�$_��=��V�nH��U��eul��8>J����X_ٌ�ę3�;�C"U�������U���l~]���J�g$B�5Wc[���g�j�ᇃj_4���=�	@�� �o>���kZG�Y�����=�o�\'���f���/~g9w��͚7G�Ntv��n�զ��M�d
���͟�œs87=�T��c��"�ص��9���̌���LV0;���A�%��MD�:Ъs\��S���6hdnP�V$'Bj�4��v�t�B���1���x��	�8F�Ş��j(�JXz��K	�P�q�"����:�(�g#�rav��B_߿��/�a�pu&��\�G�a��$�D��JeGeh�w��2��A\;y�9�ف>�l���;x��)\~�:װ/$����w0;2�����&%"D�~8|.��up�}�{�    IDAT(ʘ���k�ULLN�l�����1n?��[�+1�جi��̆�Fv1	
|�5�������єOPÇȰ���a��Ci˄���%1�tBS��H#LZq{��2�M��L����m����b$����~��������q��+'�m��&���Q�:���Y8&FF�)�V+��(�e3���D���}6zf�d�I�[��6��\_��bm}�;j����Յ������I ��(Ei��Ζ^�4D��{51u��n���"[�akg_|���,�n�X�V_@��;|f]�*��x�{x$�]�ْ�_*�G�����8�����_WN���.n=}��4��y��l�z�1|��%\���XO/Y��q�ܸ�6��qrfJ����B���<���6e<.�ЩZ��խ-l��b/W@��؈��N�>���q��,�,���GX|��}�$��&�QJ���E�ɏ�j�Fn��P ��"WW��qx���2���u-��������F���+��h!�W������u�=Ṣ尡Ԭ�P�
�f�8�cJ�(�@�P��ξ��'��Hz�v��6:l�>��Ľ59���DdDRe�8:��ޮ\�(��j�
�T*��C��v�
K&����#|��������3��(�F:�%I��_K,s3�����-�٘b߆����W��V�v���X��7֘&J(�����Y�0�~�3��*	���k�C}r8;J��!I��gV@�S�U;��NN��:��^������g��ܔ̍מ�M�\���-�$�+���������
V77�p�0:2������w��s.���(������;�����7ocG T��Fz��Pi��B#S@�P�ɉq|p��?��|�/��au�%��>JI�l�	Ny��p� �r��Z���D���H�#���h��M��:��n7�s�o0r	����	C�:����r�;�XZYų�/�G��A,���p��5u���O���a�3p�K�'����N�{�ȕr����ѯ��e�첣D�:3�U���ՀqHP1����lq��<��Ϟ��� R{[�{��>{"ؐ���7�]��3�G��Jl.�'H&���<���n{âps��&��14:�p$����<����a�\@�ӐIm
��ܖ���ʌ{sɦS:�nG�0�j�	_Qr��I:E�=�-�=mHF�.�F�I�v��0%YѦY�����F�;�FKE���$~��{2�	���g�H��$"�I�x?���A��LI��ɂ�!�ߏ��AL�%�pr/K�C3Mt�<R������X����s ��0N������HA�x�xB�C�3I^����{�jU����t����`o���y �b��2v�v�駟jj�K8=��7��gWr�c���#�bp`;[x���RAQ��BV����Q\?w������	y������%�ڐHW��.^���Y����u�n��
�k/prv�/��﹓T]���4LIht�Q�T�cWc�x��v��v�%19=��/bzv.�/V����GXz�LM��P��$���196#��p�/��O��u��\�� �"�v��~!"s����B6����Yl4c`�S,�X0�=8In��yҔC$<�M�q7u�k�B<>��Ԡ&���d���/-8W!|_�7�i��u��,2$���Y�K��Ѓ 
h�LBٳϱwt�ׯg��B��X,iB2><��x_P��'?�_}�b�p47�]3���DM����Q�f��G���5���o,)�9�=Z�5%[EX�im�ߵ�0�iC�f�y(E)eȔ���eQl�������~I%�T�~�ѝ����P��!G�����sC��J�"�bq�	^�|!�U���"�e��jM�	ዄ��olmaswG����؏G���/��s�����G�Ϟ?�'/�F�w�?��X Z0m�F���(!���kWqfa�\Nę�WK8::���R�G�u=K53g$���[�$���� �b���岌�q4��4��c�pfWLU9;�bg�f�6�+2��S�������\��&���M����M�x�.�������s��$�M������^�r��˶z�ʶ�v柒hd�o2���fː�0d[Y�v�!��U�����S���s�����ܻ�i�ߛ�� a�J'��0?>%�jfQo��i:�5�P���:���R��R�NΟ���(��R�n=���O�a��U^+�Q��b�!��6��5=8ڷ���,dS�[���V�,��?�C2;P�l�?o��v�F���%k2�ŀ���`,��!f&����D)և�cS���?�X$
w����Ed�S(V�Fl^���b�����%��u�X�����F���-nw�h7ʰs�ީˍL��lN�~�ƥ�[mJ%2�*�$f9�>ll����k������%���4]�ϟ��sg�JF$�dF����0�"��4����d�����O�Sk�Fc�&�9sJ����Ɔ�}o��GK+˸}��`�|��\���kbl�.���>����Ζ��$f�k�\v%����х+�0;��d�v�������`kw'f���3��w�]Ly�q�����q�S|�g�˸�dK[ȔF{p��i\��N�>-r%u�O�<�J��9����L���v�܋�I��S�t��6p\(��M��b����*�Ʀ�R�X[��������z�1D�>%Gѿ��?�=j�L�����u�<{�3�k����c ֣�.'a6{t�Q��$5�d8g����T����Tc�{��)Mx�a��<�e�C=k�Pv�Kś�!��C}CH��j�y_��/p��MaN�(� CC�OR���{{�U^���5Q,Cl�U~�`}����l��_U�ߞ�%%2�_�Φ�4�&�_&���Y���p1�O��'���O�ŷP�%��rjV�ŢS�9�s�����ava^H��۷��|Qk*!ᰮ5�
>�ܭ��H�?��
H�N	(���������Ͻ��_�n�/�����o4��,HJi���0�@��U�p��2��~������
�^.-by�!t�?���1|67
ق.2!5��z35�<n���'��&\�v�U˩�y�F j�� �ł�>��F��R��r�%;�T:�6�Ǒ8�C���L��X^]!��AxL
.�[�ھD��877��7�l%����s<�X����Ƞy�������e������I{�B�f�9�/���-��Í۷���C#0�p��[����	�ZTR�CG'�ب��DPnV��z+�;8�eQ��EV;s�;��������-ls��9�$�Jt{�n�.4���/�/����[�HN�v�|���7�td����<_��X�,o���ьx�K�a32������U;��F�}�09��~�=�&zhv������!2�,r�V�@�і�s�oP��I
��k6>6���D"Y�v[�kEc�kմv����@�Nc����Q������˕�7��-m��?�'�����ށ�#|B]����-@�Z�6>0���1�\�"����v�j�o���/������wo�������!�Fs%
������/�D��@�^G�P�nkhh����+V�N�?��s<_]Vf����~����b8W�ݻ�q��g079��'ψ��~�!~ 3�:��<������e<^z���jp�}"^�zUr)�)��/���x���"� ���0���a$�I��)��#�<W)�ZU�������+�tOr �O���Șo�jU���{��\�:=FOx&�X���|�7���N��k,�ϟ� ��A<;1������f���D ��{��'�l3i�$ucq�s2<8���ii�I����v��d�H6/wڌ��Y$b�ߏf<sj��͗����ۚ�XP�AŌ"e<^/k����5��_��T3X�[F�%Q����͎����{b�����l}=��K,q:����kptt�t6���u���z��Y���Þy�햌6����(�%� ��H$O�(���!l�7qm�5 ���������!�+y���~�C�E�$N����P��߿����G�G�n,��J.�[���/�"�8�f~�#�>����@_ ��x"La(�@&s��Ϟb��K�xvs�k�:r��n�T�BA�4|��z����r��$�C����QP�����0�/N�v7j�2ԡ�/-ߺ��+�]؝�g�4H L!�Ӈx$�K7�j���1��)q{�z�C=I������9D\>���7_ai{��c�m]T�v4��*"�H2AMRc;�M:��3m�+�7��kW��$<�ߧ"������Lĥ�k;TxǓ�ҟ���y��Ʃ��J��"�}0}��mH6q��Ua®��Cܸ{�<���j5�K]n��ňr��ED�R��`��q��p�Q�����wr�1��9�')����T+
MWѴ�>�)9VV4�K)�"��$[PZTi�}ft�|�L�{G���p�>�� ]����6�嚈V�N�VՃ�&����FF��ᠳQ��lE�8(��nWQ�=&_���嶡�"��*�8<~ll�J��i8�#���(�Սu�ri�)�	�&��̟w��3��*�n�"�FkF��R^r���/�w��6}���J�N.�Pq���C�r�K��/WW���&�������v�2.���߇T!����%��z���`8*�h�^�>=1��c�����je��bztT?=8���`x���� �G��٨�:x���ŕel�����H�Եk�p��E��o�ʺ�E8_������<��&�z	D���e�)�'"�
B?.�4	S�OM�Q&#k��g�bfrJ|��i=x��mBg���W$�WK��i��D�
���bT�X_�a>/�jafN�������
���G��e3r��^�֢����zi��F_O�ٴ)	Z6f�Y)8�Pq�%�J��*Y�$��P����/dB��b	�!UPo����)c�M��i3؆g��"jL��N���oEZ�ۅ�"|��!�$.��e�dV�`3e��<[Ԉ��*��oM�d~����%
�4&}ZhR2��a��&�+i�M)[���ZU�ao:&�8�#�
�*���+^��di�����.�����ɑ��<�?�������?\�����wVs��>hԂ��y��;b��^�"��@0��Ӄ��^���	������G�AH��D��q*�|� Ȁ</r�N�_#K��5,�h��B�a��N(͌Φ�>C��B��.ػ��j����:#.���e�`����y}��$z����P�Ţ"|��y������4���!L��|�ݾ���]��(2���5�dS�jNu**�y��c�(S3�.�����û��`$��7��!���"Ls���a�Ē8<���z�än�Q����,����:v��||�LN�#��`?��� ��ZI���ܝU	]Ɋ���dx�&Z3���.>�7���a$��{��Ƈ��?o��(43���X�t������Z#��)�~���j=� z�𽹓�k�g�Y��R�zIh��ڶ&t�����va�O;���!�%�#���<N���֑F�eX����@���_zw���wn���+&�;wp|Rnd+���T�!9D8���gu�q��%132��!��mM����BN���Ѿ�:$g�SGr�����DB�n�L6�o�0��,�/����E_��N���2}~�&�6V���l\6_$O^�]�I"
���ʟ<{��O�a�� cC�<����1$i+��XIb��I���6�����t�%�R���8��=�<N�8%�eusU:�G���=<w�,�G5;��È���Cއ�L�븘A�ZUZ���M짏�&q��E��=!|�Z*h5�� ��#Rb]^xY���њ�l]i��ż&�ͣ}s��j���<�&�U������sMY�^���=��t*�f�&��Y,,����FzdT�a&s��g�/�noc-S���d�H�-�r�χ�ׇF��b�(8<O��c�5��V�4r�����2eYK�,ãڒ'};�ϷIjշ��*�oO�1�*�Մl�߆��asʳ@pt./v4w�2	Qf���MDѤ�P���v�iD�f��i�A���#^F��!��P��z8!�C~��kM��Z�����WR2��k�zݲÁ�h3c�"��ϛ���������/����F5 BZ�+�"d��}��� �_�?��9 �N�ѽ�x����u@�͒�_S����A����1�RBH��6����J�4���{�<Fi��$v�>tG!w�Z�Z�jS�,u�1v��BpҎ�{z���1nt�r�Ih�T�E��|dbJ���7�\��?���2�HUJ�;-yG)W��C��nC;L���-Fk"�m�ۇ�����K����=>7���{�%��C��Ņ�S�!{/j�^(Y
@0�G�)-̎m7�����`��+4;N������?�����G�#�yx7Ʉ����>�?�ǩƄ����"QV�}�?���ɜ7!�4$�����݀��+v"&O������:kN�
<��c8�ڰS%�U�Bf��Ű$��O���D���l��O�c2E.T�9lnn`ms���ꠏ���K�{bG�*ƲQ�I�#C裵�����#H�$nd��t���Λ�o��p'�j�Q�6��t͚ҥ2�������� �}�jA��Ӆ�^6���zg&5����b89:���!�N����D�Mds9��~���-1g3�c��xo���B�d���N��BN�`w8G8�@"
_8�h"��d?�N��i���~�[G�ȓ��v���~���IYV�Gb��0f�������踈Y�Q<*_hR6��(&Z�<��*<Y~���{�����$1�7���q�G�++�߻wG׊�߅�Y��z�IEGf%�C
|�m��V[�dJ��޻$����*�g�N�MM�"�mȡ�$��X��	*��@.�����)}�a6-��y�i�[���C ��mKĂ�^����%٩҅�rBJ_tޑ?�A�c��,�bE���ǵ�0Y�<W���������mvD�I$�o(+����8��7��;Ϻ�I>��H���?[8��מ�N5��lM�yGlM��d����ǀ�͆̈́�y]eHM:�:3������m�χP$�t*��,�m�6�V�1o�	���!�V&(��X��A�?��9��'O5lp�~���1��<� ���S�f����X����=�ǏoU��?���?z�<;�����R�h�hb"�����IH� lscvp�p~n��
��ܺ�;�n�L�?94��gW�&{��5PoT��Ã�7�bn���ؼ��v>�V��3!R�y�-�N�z�AJ�BL�͗H$�`JJ0.Ȑ�Y`.�$/�7�VN��!�bzxc�/��,���}�3(4��,3��i>M�2ʙ��_�<b�*��{D�����xC��� �g��K&��n|�"L���y�V�����1�?*������Y㱳~��7�<«�רԻG�x��u�N� ���p���`3�C�e�m>�.��}�B��N�g�P�M�i�A(�+�n�G�)��oMhe��P��a�A��Ņ��܍����%��yO�}%�$H�}�K�eآ&�p}jc��v'��^�����g�8�F6_����P ,΁�h՚�u}4A	e��K!���|p�lm�ݔ��)��q`�O;�9�3��v�X�
aa�{�і�\�\�Z�9L$��E����F� !0:W�G� �J]V��6g�,�m�ۘ+݅H�r�K��>ؓN�Z,I'�{L��<d;]�P�E�{��]<���x�h�X5���.��>��|��SGx����Ҕ��4ߎ�׏���0:�~A�]��K�/�ʧ�1��w�P".���=�&�MN�V/L;��dK8��d��8��Fџ액NN�˯����C=�JI��p��$J�`L�J�(Ґ^?=߹.a�J{L�)R]�$L���N�]��9�PY��X�w    IDATe
�ˮ�+�D$
'�T���S�Tnl�^�T>�Uw���BVN��a~n (@׿�dGg�x��9�,>U3�g��ף��Z����ƁȊr�U�:�Jq�i��95��~a1aa�Z�k6�|�����W��9ck��oC<�T��*��8M[�Ħg;ˍ`,sj4s�TK�dA��$lV6y�LH��/[{�ad�s�.�\�X�˿�v��:�|Ǚ,�3]�-��9�}m$`��pre����F��+D<�X��qa1�$��Ŝ�R���g���,L/jE<Bp����݈���SM�J�͐��s��i�w�\��|S�~�۵W���������[-�m��Y���6��Lm���0�^Gb=��k873��d�l
����[7�ɥ��ux=�Vjڏ�qI'a���c�\��EǢ`���`'��V��q��fsz̬Hڳ�M�+��d>�n0��A?��z�t����FW��|$�����%�L��/����3)�ɝx���\���ǅ��pH����@�TA�����n$�e��PwH�Oǁ�'������S3�	zQ.�����D�	�H� �ϝ.�U�+�֦��s��7"�u��,����}d�U�f޻�Μ:���^T�e�����/�z�B���v5d�6y�9�	�X��d`�]���e2m���uho�C�74;GP�����4&֒��&Ꭾ	2*�V4�v��@�&P�#�`:փ�S'0� �t���)��ы'���\���T(j����!D�^E9_�^3�rc(�@2B�D$���lʫvR7ܨ
�Q��I6S�If�����P,W���\��Ad��s�N7��(�i�>�h��)������X;�:���LLa�!��n�����|���}�JIP1�D��Pw�!�]��g>Z�0��B�\B�������%�?�}Úy����.��2�*�ӂ���I|��u���J@	���Wx��6������c��xA�q�ȵ���>Q����6vw��I	��?u�N�Rq%q)�e�aoO�>��7�֎��"���ф�0�I��T��Kb�渎�M�P%7�s�SE�Ĭ�'Y�m������C�d9J�_��o0ɤ%��QJĴ�G�qI��fu���nY�Z-�?}gO���̂(n޽��o��Q>k�k�vI�t��0u�JW##������LS�}�3�{}�O<O*�l)�E�E�5��X�*ƙٛ��NXh�`d���0�6�L��T�kHy�}%Y��S�M=���aak�U��[;e� [�^����<�-��۟k��2@30��H�&&���L���l��߇hB����h/٬��s�FM�`A�����k*.H��s���'-b�d+V�|���ѾZ�R���c]�.?�G&~836�?~����C��"|��;������;��[.����CW�6�u�ޢ��HQ�����Q9֓D�Z���.��7�h�7���|������M眢�Uu��{+�o:H��Z�N�<d\r�2v�
wr����ś��D�n�D�X0,GBq:�Db���4��)��)á�:���nv�ÒӕK����/?�����j�x��z<����5�����ر�	Ӂ�%N�v橺���_�.�͡/�G9��N���(V+�$��ŉ�)�Ebހ�	��ʭ�ih�$L����k,2���(�
\n?>��Ν;���A��e�}|�ݹ�M��v����:�	���F����7�d<n�DMX�q�{q��
��e��4����O�I�>����u�V�P��3�j��f��,��dJ�,� �ͮv��'gD���9L��;�ȧS��_n� S)
�b�r�RG�f����͉�S���,�Q�7��2���0hA]71����Y��XX����(r*�J�:�����x����N�#��"����M� I4�y��EL�K���4&��亡CIDCƑΥ���c�p|��!¸:���V�(�#W=t�b�@�~>�	��`���3�|�
X:{���l`��I��ך�����)}(F��
^�z��+�d��K�c���pX��M"Bʀ5���:�QY6�$7ɺ�V��)�ӂţ��2�Y�X�5���_���f��A��'g1�7�kC���t;���m%��GOa�ze�P�U�/_��+�/��1f������v�l��L�x0�����`93JqhlT|50U-G�ITtq��y\8{ss�ܾs_޾�c|p�ⲩi���\�q*��S-,��΋�d q�ǐ��㺡]k�[vl�0�&�4%�x�����+�H��>����|��I`!!���lk0����)O;k�8���Gk�k�n���'�tɲ
.?�ϟVV�C�q&�ķ����l�m���V�ъtd���h��DX�G��YR��A67&���F�afq�5�>�ү3�Fk63��e�[,��\�L�^7��Qv��afd�?Ώ���`����w*¿�����^<����Rq.�� -�ݍF�-�W�������&��1�����&w�6�6k��?7{s��7>�܋��")X&C׃�4�խ�4�1庲�Z�c�{�3�~�E��6_0("�f��Y����t��ɋ:d��|�L��_����>�S<�XA�\B�;��XDi4�G6���x��
�G#����R��������~�+'N�/@!��g_}�[woiZ
z���%㜓���#��&7�	��8p��{|����39�J����裏ELB�^T���=l��ȵڡ�����qN���PTr�r��L�]�<E�^��E�xD�""�Y�#舐������v�FJY�41���!���f��|P�~v��azZ�����PW�f0��G��B�� �+�9�C�rtQ�]~9W�m%��*M3�94K%�I�k����m6���-���>\MJ4��Å�
��ˍV݆��kMEr��q�inS��/Cbp�^���`�-#�P>��L�b��$���c�o ~�!̗��a�e��,�������0��F�Eu��3��Ǝ�lF]��NE�-��`7�B�Y��=�i3�`��y>��r�^-ac+;�88N	a�5�'W?�j�Ұv���W�X]_ū�5I�Bv7����"���-�kj8H�a��4��6ﴔ�M�ǁ�a��.`jh����Ą2����cܼ{K�n�dG_�|M+N� ��>�.�K����|��Y�5�uDc=�����{�pU�g��z����O�N��N���+W�U/WQ-��(����V�^.��ƪ<����!���K�t�"�g�Q����R����z�[�
��1:9S�B��55R�$�rFo���,��l���Pn05��kp&&��"��Qa�M[+�x(��#
i��t���UEWiA��3`V~}+܁EXE���ZE���ZRC����M�o�`��͝�_G�=[��E����a�p�"��a���H٦/���A��"��D�:�ﳽ�Z�.K]�V&드 N���e�b�7���&ǅ���X�;�;L�,�e��0=8��������w��NE����_�ꓽ���.�N��**9%$���p����۰!�������	���5Az���4&3��T˿����C�_��{���MKH�Lh�oՍ9�p+�Q������o*�ӄC<^�������`W��Z�1#VōՄ])_`n�!�0� ����m���<{��t�m�^��IL��`btD;�j���lI:e�a���bm�3����ۿ�Kx��	�C�e�d���Ay�W�:v�I��:fd^��)aw�1!��˻���XB�c�/�'}�KW.�-&SʘfT���&�$�uZ�:3��N]�f�r2���]�w�����i��D�7!M*={	�ӭ��J���T�aa�zyĚ1�
I�d�Hq2<c	��U����AN���Cb�Ë�P�&�1��C��B��˯���>D���k����c�J%6l$2�)��
y4+e�p��%*Y��g^��%�9A�K[��H�ǖ�jN4���U#�����
L����� ڛD05���\�pG�\BYx��E�855+�O��K�ｉ 8l�U�X\z��8�t��By|z6Ԕ�e40�G��C�HĦ�Sa����������q|��{*�4�aC����r�
���g��<���1����v��$�{k�.�B4��KUI�����h$��*udD�lZv;�ՊtԴ�É�i���}&˝���ܾ�#�7�
��N��KWpn��
S(��
�|�k���.>��s�G�j��~|��G����ܹ\F�)?�����Z�eO/Ν:�3'O)�JhI����a��M��q��?y�LnYl�������2��ܼ<��?z���
}`��Uj�B�U��|mCҧ_���4Hh3&`��l�9����څ� S��p)�2�����O,�$�Y)b�|y��H��a��\j�=ɲ[P����5�J^h��&^Yd0�g{��ec�w뾵��U�4	�jMB���1y=���EC�R��5�0�y&�ĈB4v�W�|ތ���]�{�Bx�q�5�ҁj#����gW �����Y����Z` ���_F'~��h4��Ѡ|��{�������m�Ŏ��ڎfӰsw]Jb<_����.���8=9W���dy���҅��h�@�Y�˔ŏR��H��~���iɚ��b%,��];�t�}�:3ʝj4:7e1̓�r�Q 4�lxCқ�؃�#�J�5&г���X7��:�����?���{�6�8,�Q�^7Qv/j>�|N��X��?vy�"���EM�	�D�*}�)��sS0(%!��K�����a�|MCk ퟩ�#$���b+��A��|��P����\d;������8(�P��<J[Gp4�FX��0��Q�Ԓ���  �X�Vw�P����O�5����4 "�UH<�t�l`�0pU��c��Ώ�3�%�c�J["�R�i�я���T�H�|'q}��⽈�](��jm[rc3�ßMC�Bc|C��b��
=��T�Y�\v�aȤf����v�|n��i��F����>��:�tt$i���
�$�!�"�ܑ��M"��q�ݔ4�³�pz�i990������5��2�GGm$ݭ��@*���;r�fZx�X(��ĹPDE��� �f���ua��=�C���%ˡjucU��ԁ�����P,�c G�pe����]��m#ߪ(��Nf>���k,<��&#��\Q���H��{U�v�$����yL����p���`i�9��u��7u��N�����NϞ�=�:>���jT�Kv���%ܸsW�*0X,9	S��޵w�[�g�"�}�ӿ�ͧҪ<nɌ�7fx� �f[H�������6��VT�	��U='�.]����%U�A�����s��a�ATK� s2�	Ul4I65�s$��Ź��-w��/�{��IH���H ,8����%����Ȃ��x̵#������v��#����XE���3R�E�Z���#�v���lM�V���1���p��;��h6�f)S�Ôܩ8鲉��c�o8�ڠ8(�ɽL�2�+��|���LT""��|��aq��)�%4���*s���w6������z`hP��,ĩ�c����(׻�c�?:���������;ۿ�:��j�f�;TF��G�뀫�F����Sg�хK�8=!���S��rV���F[!�,�
q�/�
ܑ4�&����إ���b p"Q!6S8X�Œ3�3��Go�A`W�}a!������WU�s)��3"rm�Y�)��Cwpt���!S�i�\���q�,-f�٢$��m��b@����jf�%i�L��6�9�$|ea^E�\���/���|-b��X�0���u���K�&�xvd��u����vSY�+-�z�����ŋ�10<���~z��xtG܏:�:eX��$J<|mH�6�_��_KP''B\�ܻ��F]�C�,�<p�X�0���U�n\=���p�%��d6�?��k��_5X�>��\�Ȋ�5��1N���<&"I$�^�JE��-�5���`O����[�jؘ�C��;���1rGG����H{1�����E���aA���;J�IA31��a���a$��M��K:�L��IȺ7���>ɱx�0�!J��k�u�m��o��L)��K�G��l���>lPy��ǚ~���R����d2"+ٺ��&z1�;�O��@�?�a��
�Sک�>'s����Ѥ��4m!\����M�|v5�$.Ҥ�h��M3�d���q>W4�B^�" �ɯ����t5�3�3Ss�E�A��vv��=}��ɃM�S8�,�G&՜�����ޤ
&�S�<Ք�_<�����^���r1�Q����s�@/�#�^�,қ��f1|������%�}�H�q�#<SX��\���s:;��x�;�i�R_�4�T�'�KX��u�H�H@b�<Y�x�$T�2��|]\V(��Y7��}AT�5A4�%%�"�,��b%!}[�y�򹳊0��6S���`r8��(
b!��IR��"l�����k�'n��ZßM�-��3�����bN��J;b̽�x?"R��x��5�	5�n�Q���dR�H��x�2zac���q��.�u�s��ZC2?��h".N8&<q�Qȕ��􇃉�?|wd�[k��0�~�I�'�����[�|#w�n�Ӓ3TU:1c����~�D:N��p
�=��'O;]��V�>!�z��5�+P�VC�)���E�4Ӡ����C�alH��^4ª���Bl	��}o��J"����euy�E%[!{TZ���I����C���E�׋��1���
U���<X\_������J��kgG�)�{(2u9��X\�t��GV���pin�QƮ���W?ŗ7��*IXAB�}�����t&ep�>̈́j���n�erX�����]�����ǿ�ӧ΢o�{�����U��K�]v�����d!e��:`�S�3L�a�*�"�l0n<���;(v�.�Sz]�X�Z.��`:oq�ַ�0��$A��<GSJj(	!���7��֛m��-��q\[�T�I�UK�K`?�B�UW:���LCm��c��ݝj���Fl`�����
�R�J��&7vϼ�x�1Ӕ.qDX��jZ�Os"M(���Ԝ����G��ӭ�W�D� ��<x�hL)��zY;,�i�%�l�b}�.Pi9o��P;��e5q��CT��U��˘����ب]t��tJ����T�����`��s�����u�=��3ҁ�7�#�涺���[X�]G���z	�6�-Ʉܡ�n�����C!eLy����*ַ�`102��!��OM�`~t!;�J�8:>ĽG�p����i����?�~��pB�U�YA.��K� ��/����?�'@3�t��P�����<���Y�n}�
�>l��)����+X��Wc�=2ܚhKJ�BN�7���7�d�j��W�j/|jnA���Ǹu�.^������i�^��k�����#�����|ٍ�-Y�
����-�6��:Di�"�~��N5W�=��6�N�;bL��$�{�g%�o��b��$Zu��i2��-����A?�A����-k�2c\��.���F(���%��v�a�	S���HY$U�vt,�cG!�.8�ߢ��~Š�th`@M����.qL�$��V_ڽk�wkh�3ĉ�X���� s����r(U���w#��ui��N�_���|�to���gS�st���?m�Ȥ��%U"�o��8���	|x�<�=u
�j	�r�J^)Itw"���"lZJ�Fv'�$a�h��W%R��&���Mk˺�Ī־����n��@�!��t��%]���1�-��V�����PO�)�Suj��&#�D���Y9���9l�-Қp�W_���
��4��� u�M�I�G)! o���FWy�����f��Q-೯�/���|���8]�alY�(�JSx��Y�]+�/�4�r�"�rkÓ��G�����	o�ᳯ�"�[ʣ�.���[���CKRd�F�,��w�)��pic��<��yݜ$gթۣe%��1��Xl�h�9Y�4�l�_���Jx�p:�.��]x�%"ְ7��͟�
�*o    IDATL�_�'�f�jU2�6���`��$c�a��E�R#W@�({��b!�)���+���#�L	3t�����t�+�;i9I>#[��T�!���HD?�$&tgl5� �5��t����&E�"feCE�ו��ˍe�ln�(��M%s�iSɤ$��e��UQ�}YF8cҊ��&�*�I �ۏx(��� >~�}�d����ʨP�S��	�#�	��c:�֗�����\�O���x�i�5���K%d�%���q��3X�Tɸ��.�"#6��J`a|
'ǧp��9<���W���=5N^{_E�7��r�cL`ux�������cx#A�1�n���㓏>VLa.����
>��΀׏��5LOL���8���3�^��|���y�fÝ��q��#5*�rA����%���I��ݻ�bͤ5�.�&*��Z���0�@�O]A_���"��\�/y6Rnǟ��l^��ݨ�p���r�d@��Ģ��������Lm�i����pb�&׷W'��^���J��CW6���]��o���?��|+�ؘ����=_��������5X� q��c��谆�x"&��b�w�Np�ͦ�h���^C����gQ���F"2Ҹ�^�70��&#�.��2�ޱ�ٳݑ����!�����"���~#s�;~|�I���ዝ���9�^����E���eC�ޅ�넳֖����i|r�.,��V-���+��m*�ّ6��J��Z��cq���I��)�R�اƔ��;�F��ZS�6�ʕ\��0F�E��{�H�$Q�W(Q���UB>���,�ˬ��l!�(8p�~�����PmTD��!��q�h�v��|�j����vUx���g��]M'�o���I���;�MeUe�,�}w��ތ0 �K͒�\,�%�����}�.A�+�(B/z�YJ A� ��i�m��.o�\Vf���s~y{��^�0lDǠ��dݼ��}���i�W�w>�'��FgS=2�8�ݾ���/akkCl��C��in��%�Ѯ��$�G3Y�<�����Y�@4K���}#�=<�"��ނ��Y�u\�wk�$�t��^Q�p�^%�2%`.��/����fu�l`dʝ\<���)�#?��0��q$JX_G�*�\�02Ȃk�\ZS �,*V�����5t:#�3���Q��F����5AIɸ'罐,g�y�ǆ�M��$�<��_F2��B*��;�;"��@�`�w@>�DL���-���Zu8q��R$g�X��C�6P���:�y�4m�r���5� ��fe����bU^/vb	wv�uM���c�4��}���y�E#B#<Լ��
���6Ԉ�P�� tOc�}�뽴���%�l��.:kB���Y8)Qډ*'�Q}��+��F����&�6f�N�ɳ'X�XB}sBM-���ҽ����ڊ�Y �U~xh�C�i��ױ������S���`���{�w�V��"g������[k�8�� �ޏj��a��1����@_�����,�<}��/_���b)��s���O?����w�фɿ�rY��T"F�1&���ǘ���z�t�A��r� ~���h6����3���n����Ҍx�Y�?�65<�/�)p~��)˫�tG�k�k+~��7���no��O��<2�<d�Ƥ&	��#�����IU��j��L�Gb'�?Wc�c�Ĭ�������LϦК�p��cl�I\i*x���P��f�i`�wV����oѬ�$�Y������'��\Y	K���,-x�H��#@Cc�d���W&��;�2��Z��ZW������O���j��2��
	��.S2��"�#.1�nq;�4�W��o��s==߾N��U���b&>�,��DYĻ��_��HC[��_<|Gv�������x���槐/�e�(�V������� v�q��T@%/��&2���0��J�!��=����.C�1M�5�Z�BWO'����&�5sy�-1�N?�\����v�y�qh���+�]�'\D(X�d*��3S�g�H�XO�0��JlKE�@;~,��s��괹PH����}�!��Ewk3��$�޺��/)�	'JiF:{�V]�I��d�V2R%c�FI���*��$��A�k������������$|��m|y�:V�	�]� |�]7w���Я��T�������V�$��u�(��� u�pE꠆�PN�K[F��g��gқZPw�$��d���,Iif`S$��r�j����݇p�w�M�
�s) ���"rB3J�hd��p���T@�1�y��w��3s���)�S̢`sʤ!PU�F�R;>��B��$#���^�K�����9ְ!��mmi��يBlx��S��,R\����������m�[*�'��0^��ֺѾ�H&I	4�	�ֈ���"�c��C�
����6V_�j��ih��Ϋ`m���5�	m�c�g�=0�û�ʿ�Ex��ܾw�?Bm�mݝ��R�G�Sj��!{�6��LN�3��zxۛ��nDWk;B�������յ��-�����!���v]�v4��#ˠ�͠>X��()����􃞞�����N
�ĎX��!>�$L�d;�7o&��_��B������Fs�Z�u�0�Ю��ZF����	��?����s� ���c��A��'t����_he��Bcs��:��`�Y����|rf���%�r(��t�g���!��ʬl�Z���/N�SS3�wq��������
q��$�O�
���NZՂ���Z���ϭ�xX_˚�9	[֘�ױ>��ޑg�cQ��X;ʦ1��0Wz6�ET" �F��af����w��	v���ʋ�ë*�lny�)�02E>mEi|�".�e��$�o$�V����Q��{T�P�Xq��Bl����zo�g�D��������m���l������뿾�rm�/�"k�X�3("c�}u�t��ܰ�:=��7���á�!�q�x� �����M'ڄ	�pRp��R�P�ޔ��������	��/�;Im�m�$��P�u8Q��b�7�dJIv�݃��!��5c���8�r���h�����N.�9a�-��aڧ�����.�jMDp��=��c$�y���X�cɸ&q�l(��^ټ����N�c9��j�{~������%dp��������B}�hW/�j�h�W�X�2wMO2�(��Rī���oh��S8|�7i���:n޻�"���Q�^�E�Xj"�0��irJ�ǳ�K�P���V�06'j>[�G��ݾ�]�3&2D�A�'�r�t���������g[ŞE�X�~���|"�������>��wA@�zO�;f��4��Z�{���/�I)Pڸ��nC.�B>�BA�C�4x�l�mm���ַw�=Ї��N�ܷQ�K�biqQ��'���A��C�82�����5�1�0I��嵍'v0?�|a�4H��?������*�t�ٷG�^�mM�Kd�W'�*��I���-]�5�	����'�JX\X�y��Iaav��B�At�7��O�O�
��-\�qEZ����Z,rgvptT{���AyG�ݿ��7�bbn
�Z��w���f4u���fd����.M?k������9�C��^0P��@C�}��.|#����9�r����I�_KMH��ɍ8jk��hC�e��<{����DCk3�ڟSj������y�&�hb?��/�@���*^�����Cq��L�((Q����޺!k��yJ�_�����,�/�kmn66�Du\��Q%��YliC( �q��$	����z�Ɗ�f�$�Ɩ�3�w����炎��㝕l�FI�Йd2m���
�1��M�u�깤Y�e\Qi�Ɋ4��}_��3YN����� �߳ɔi�;�,�C�^�0U%JR�Pz_�0����!|���+���v`cc3s�X^^��м&;"[[���|��I�����`�_D��<��5
m T���Lź�&��A�*�RI.]���Y�U~@}cÕ���?�N���oRO���͊���������0Y;���H�"����9��n ����E��#GppxȦ�z|O����k�>��eH�h�i��<�+"e�@t��i�}*/��ܬ"��Q\��Ig�+�d"�n���;4��F��g�(z���<�b�RV_W�`u@�;��	�&�y
lgRX�Dp��S톺 ~�{���&���._��o^j:ɹl2�H1�d[W&<��t��E��
�b"O���ۻ��9߸sUE�7�5�ܗ�VQO�:����y9gqJ#��e�zWcq$��H;w5�Fp��1��Fxk7��¥;71� CV�s��0_�Յk�$�IC��b��I6!t�����e�W���,u���eqbQh��A�L�lZF�**L�!�~�2�0�8N�>����$�I$��tf�Q�;tGw�Q��ӗ海�_\@6_�ٳg1�;���F��{����9m��f�)����{��k\�{�H��C�5*�bN��TRi`/_����I�tu���C����Z�}��%1�z�=��_Q/ʟwl쉮'���aM�<�_����#y��KI�Ǳ��2�XZ��L����=�5�R�}�bȍ����T���-bmy�^�3ہ���~���jAl��ܐk����$/d�ٻN�Ɓ��j�޼�k7����Ե4�+A2[cKzG��>�$0a�a<܂�Ɲ�ρ&�(�0���OӤ��F,��Ҭ�0�#F�-�Σ��#�}�e�z��B�|*�<�)z�f�[Ե4cms��r�c�x���m��,�������0hˉ��eO_:��QW�D����MAx���ǃO�^��U��ӭ(���V�<3��LoiiBs�IIW|؈J%@�?��Jx=_;�}q`�&�7ߑ�7�J6�a��DKX�9�Q
)F*�˗��ڵkF#� ���'��J^�/�k2�"�ZE��U�M�66�V~gl8�n6��76�F�oκw��{9�jB*���]F�P�RI�<��Ta�GC���?��
����������4����s��]N�2��gC#�[;��֮a��$��,�o"Il"
��dTzH�Y�����Ư��Æٕe̬,bm{MM͗;:���;-�E�?|���re���׏f�L�h ܗP��/���E�9���?�����Q8���Wc�w�&ތ�Qɮ8T۬,͎�v]���-��ÈF��@�;}N{X>��}���>����d�0/�Nn�a�f"��a�o@T��eu�G����VW��� �A}CP����);�L�l���]C<�7S�*������wT�c�|��_`l�)ޮ, ﴡ�q#+b�u7f�B{M#0EEEXl_�v¿��G`��h� �����ʗ����*�-�Z�,�9]��$�9#D�z'��R$�7+��L���Y��	�;{{��b#��kwoૻ7��#��p��&a��<pޱ�y#��D��YYv�4��Ή���Մ�"?�0�y�r'Z�T��I^dYw57����L[�m,��be}M�?�6���M���c�˽~�Qc��39�����Gpj�4������꛷nau}U�O>������0�9%+�tO�@���b�_� �����FD��C�ȡ�z/���q��<:���y��=�3g��ȡChmn�K�$d>܃����ž�0f�,��k�n�Hq
c�������ך��C>�g�8��kx��^�v*.��������שqY�XG�,��,������TL���x���¿����wqm��a���,-�9⾔������߽��"xp��}Ϧ^���]�=X�l�d�|��|(�ɚ]�<h	�S�KXPNM+�jO�{�e�J��3
Y�]j��=A{�Y�-���[wY��,�1Mv���E4��bm{[E�D������3�����W�����O��ӻ���#����ӧh;�թ�Hl�m�\��8�M({�Bo���w<��/�f���WV���k�)���	o�g���&�F%��
Ɍ��	��!�ǲ7tQ*�f�C�VrXT.]���W��\�i�d:���9U��i@�,p���YŖ��w��~a5���sXE�TS���l��a�[E��iYlhc>���+s�����n,�F��F�p������3�����Uli�4;;�fju�!�fsJ�"B
5���C�����˗0�8�!���FA���U1f�����J�p(:m����m���~���oη��)J|������Ĭ���^�$�"L֦�y�Z��[��z�OE��8::
g>�������}�̾�^�����[���^�	I�b����ے.�݇�~�����z��5u�|C�$�q��ʦŪd���)�ɠ��I�e����p��)M�4`����B��rϢ��2���tYN�>B����!t���}�5u��#��?��O�0D��Y�ܱ���tv�n���h�b�fFoځ:��s����[Q.fT�/_�Z�!z��>�������o�о��8������ە5,mn#O���ԉ3�p���c�yS���U��XW�-8Zt
�S�>�?@�Xsh�Zf�_��~..*1?F�F���w{�&	6Y�w�b��R�B~�٬�3��1(�Nd[��҈�u�@��f�"t�Ke'����v����8�:��0��5ݻ���5�Q#�u���@��4��oU�31�zp6M��ܥ{w�卫��S2j8��0>8~�K΍[70��gg��=|��GO�a�V\�l6If��j,��Ng��"�.߽�l�(��ĉ����<}�B�luC�w�)a�F�6�f��ܧ��7;��ɤ~v>#,z�E�!���1<73���Z��Ceg��7;����!B�$}t���9*����7p��5��y���.�4�u0�ʇBI��V��� O�S��*��0��nG��^;���^x�.��Q�ќ��d������sT����
�.9ȕ2B(_>y�B�0�Am]�G�D�jo�ƹs�p��1�UT�'^����sl��ERTw��~�A��h�A�@&�֮1�u��6�;u�#��N����{hH����e���7!?���]`���l)����ѡ����&�I�/,(7ziuE׎�3md�>��0tSS˻"�B��W_�ʕ+j���-��U(�/���W���d2{�"gY�0W1�C��^�
���hm�������L����U�0�����X�9l����ȳ�?�-�t���h@�D���Z��F:gHb��i�&��#���=�KkH�˗/+&�r+"d"��7��*���*P���6����`��LH��󶣽��]���L���MQ�E�O_�����,����kg飒�qZ��lQi��9}8�?��O����! ��ċ�>���ya���=������]"//aB-ܵ�c����/e7�_�{����E�䏕��dV��7��� �̿��;u�؇��&����	kj�o۱muQ�(����]lk+��5)���I��g"�ƕ_���1L.��q*�r�r�"��a�I:�y����儇$�x�7~x��>����J��q�2.]����%�׸���7`\�<>Y��h�M8�����1����Vװ���H,��
'����s&�!UL�����1�i�h�|*�$�)Ɉ��^X�XA�"+�4,/4��&����I�D(hlA���M�<��Ł]{��S��(_u'��|8��o'�|�\�b$P�P�|�{�F�߯�-hzi��ܑ�p訂B^?��۷���3u�]"޵�Z1<0(a:jo+��`r��p*�Ć��7�����؊%���wX��˩����������##J�RCGS��!��#\m�����#���10�����'N
����i#I
�;*εȦA4� �M	_{&���ʊ:vA����
�
@novY��a���n�6>�H�*v��+��\��[#E8{���ŉ����S�߇c�|��i
�W�Đ���2��4��p:�a�or<���QSP��N��}]=r��c��4�d3i�Y���L�P����z�~z2�Rtg/_����"���	:�    IDATܸV�6�������=u'�FCm-�-LL��/��\��a�0�M��FƼƴ�d��fӈ� D@��*��[�f*��a��Z�C���R��}eu��&R�t����tV^��HT4clX����ʤ'���������c�/�o|ml��9���>�`2�Y�	E߼ySn|"R���6��pMƿg��ݚ���ʓ,�NH�&�o�U|�~�/�m����mlg��c�%"�Ju`^�
�<��@��庆��Z��Q�ْ�ΜDgw<^��.�6����ׇdW[)Q,�l����hm�R���;�n� Ygk�����PUS+�sW��{Ss�[Z�������֞��7l.�o��7�	���O�=/�xzc�c�M'�^����m��[2��J�x�0�3>,���'�0��!��}da�و���G$/v)�H�ry��Oeae�ʯ~�+1 �f9z��U�0�0/��$'h�@7�6��B:�����#���C8���/��X	���d��l�\u���uj�ƽ&��?���G[}��|}�<z�XK��m��.U�J�@�(�KM�ׂli���pUف\��sGa���l
Wo|���\��FX;�Pu5N�=���.4Q�O���,�M��r*f�'����6"q��=uF��辽�Ғ@�O�o��"L�'�0eg2�O��t�F^ci���f�-�Ĥ��׉�DN��]�5�)��Cسk�",�v���;����ثqL,�c#�c�O#��tŇ�t�v�w0���#�x�8z��0�d�n���5�k��f&�n��O�jkk3|U���`�afs�x8��3�"ۭ�oi?t��1\<A�fv���ܽ�ɉ7h��oatx�=��L\�k�"�Ѫ��a�߹U�K%0���{o_˻���ǙӧQ��J=1���}��pfmg��!���D*e`~:�2�����bi��p�Ю�b�ǆB0[��C���C�lʲ���y!�"R�a��h�I�2���>,��
�z�4#�@J�8ue%'��hnihe�C#��!�C��,���9m҆�f0mM͒��m�b��[�KE%��PNt�0�9�׉,H�J+���jyu+kX\Y����4斸��m�C���P�I���~��߫{mt�wb�޽��)��\ES�]�;���&m.�,����%llG�{q��q���`����&��$x��%�8dg��!��ؓ���UC�g������1E�M�@�Ը�$�^]M��4U��1���5d(c~cbEm�w��m���?�ZEٜ[�a�����tK2�#�\-�8���p��C������CYMV� ���7�M�^l�H04�m��&npx �u��n9ʏ�
izS�|�Ue3�u�������ud}�TM���
ei�YCFGGU���&�ʯ����9T˴������������OQ������'�s�qr}��wJE$Jyd���εÖc�!��M� �tt��#�e_�L/��	*d������V����G7G���@�l#c��KcC�ҼQ9	��z���s؈D���Юau@��yA���WI�N3��67�����Jxe�o�j�`A%bymi��/�I���Y�0&21@��>��4�"��杫����`T�ܚ�yM�f�H��ts�	ji[x�p.%�غ\8������A>����_a3������āÊ3�km��0o`�V.~/� ^NO���x>9���(�Ξ8�ChמQ�w���{��f%��b�������T�������Y�|mv�S�鋼@�!���勨a�����Ÿ3Ԃ�#�51��`��;���h&�7�s
��\^D4�R�eWt�W��ع��3��gƅ������g�p��5���aF8�,�]�Â��{;��E(Ԡ�0�H�0"t� �G/�c~cSz�h<���~�s�=�ɞ���7�x�x
���I���!�d�I���6j��#�@�	L�󳘋lb)��f:!���|_�/|�l\� #�v�ك��$
)�Dkx����g��/�XZ!��,���{�*+?:�����,�mL-2�|N��D�λ\�4�����^D��PW�Y6������A˙�2���g���W � �̜.�ux�~*�a�Vl���✰��>��<���k��_�����qqJgr2�߈�ى���W���E������EOG�����I���?��҂�ǎ:"�����<K2P��Y2"�q�T!��]��a�>t��m>�SoU<�5~�>{}�-2�ȧ��U?mQ������U�`��F��0av�v��u5uj���}[S����B<��U}_����(�40.�aB��=ճ^�|5�����ZM��C��D����������5 �\h�J���e��7y�1�4�6E5�D��s',0y4J���]�34�\�"��� �f(�%96��ť����^6�6�{��%�$��r�*��*'Ps]�L^�:̂�#�5�-�-m��������Q�o�������vc�wX��(�o��|��C����l�� FۻT���= Ǭ�gO���-,�� W������FOG��O^d^`�&��I��#{���������)L߻of�W������HtK�#@^���&5bB�#C�8z�jj"l-�̩@+�I3���'1ԼHx��
�`=���Rsح���#���#�LT��=�=N$JE��-��W�q��GX4������D5�)�c���]���ϱ���*��M�8�� ��z��ܦC��'!hn�([i*���<z���Laay�9q椙���ٍt>�n���;�_D���$bѦ����aȨ��$��	��Cb	��(f( �IX^�����X�m��[��ZW�\,���j�]C衵#�|N$��tR��)��a$��(� q��@�!�<��
L`�j��ǹ��q��1t�7`r�aNq��!Xx��(����Ѧ���)�#	Bl�b��EH<��"O{T�1�7��{HOK-9���[7���C,//���Jpd]u����#�GC�ΐ@�ەڥ�.�ى&���Mx��6��%�ƃ�{�[T2��c� �W�w�>x<~,����o�WK�V�H��H�:(��,�r�%Џ�aB�"Y!ꐌ�#2U�j/B�T�]���J�����p���O����p�{�2r�=���sC9��n
���s���2�������V,���L�N�S�	�ρ�`��P���m+W��U\v� ������;q�mE���SL����V>s�z;;�����~�˿�=&FFr/M�~>G���ic����{�`�Λ9ů�0���x6+)��ٯ��՛Wx;=�k@H�丵�����TȐ�l��HP3q�^���=b&s�e��N�ѡtdsV,}�]��Jƴ�욄)W$��������wE�E��6��"��l�}H�(�Ŧ���(�[0�!���m�D�v�֚�}��OM�"6a4�\޻��9X���"��	�2a.�y�P����EzP��u�6�`v��Bz�x��$ƨ�b*bi�E�U̡�R�7]��9]���

v���x�g�ݍ�P��]�m��ӎ����6�����͟~^�󩍕�zW���CG"���9��2BN/v�wⓣ'��TN�1���&ṙ)�s��^��5���W�� 	
�Wf���?�׫l̛�o`��b�(�*5Y�PU[�n�Kv?���x
�,E�)��N�����CsKH��m�D������Ң&�x>GU5���Ξ��������	��;�N�q���~t��&�g�,E���.FX�p�)�D�9	�%Թ����8sp?v�t�V���_�����zv[�$+����$�?$+���:�n	���^X_���"&f���)M���ELٻw�]����L��g�.��,�0��k-xɚ�Ⱦ���������Ʉ�(5aes��A������kT�}X�[c��������
�Pʉ�@8takM�Ӌ�X߉"C?�bI��E�6q|����m5��p�>8z��A�}9�[7�ʯ���.���]����{!@r�����$���v*&�#c�$��m���Á]�p��Y1��"�v�1�nz5�Uf�t���Z!�A�OG�<�
��/�];]�:��+�:| v?�8v��k�~$cQ<���d�T���z�u�V�]�(H^�t,h:]M�dcr4K�`LB��0�iK�X%[�k�V�aH%���:�2��l��W�Y
�I5�L�k$l˃Բ-�ME aA�c�:`X��&X�)�1Qr,">�GX�z�]���ڂ�S�q~�8��]��s�(����q��S���Vi�L�2�_\���
�k���S>{�z������7���/~���U]G�R�^q�a�͟Ŗ/�'[P���d3�A��d����CM�t�����3�n0b�?����5�'�UQ�-�7�8"܋
���hg�������4���Z&C�*�u^�S�v�Tlk�����7A#,�*z0E�@�f�7�͎�:��]�
yew�f/O�zSFޗ3�4M�I����w;��I�$�ɚ(w��0�%�IaN���4
a��p�}��G`�B��\�0��J226��̭"L�d��Ы��<#c+�n�٥�՜SP���9�K.hD��l>��5��i���O�����"��o���g��1���q�\�N9oRw�\�Þ/Ù����n����;�N��}�1�t�9ݻ�����2�z�����S�`˃�7z��Z�������a�<|�Ϟ�mgh��� 6�#Z��ͩ��UFJ�Ig��'u�yM-�=xh?z{���_ZX�Mh�"���EAM�	�x�I�!ɔ�[)������w�?xx�����"� w��Ln�@��o��é�JvѠd��Fw~��EM»��h6�"����X".ؑ;��`=��*�^M��x�r��UV��$��Lbyc��M��v�9~Ο3<�I�ڽ�`~1� b�^j�+9�d�Z0'wN�z@��\y`y8���i�u�8q����B���+/�|2���y�]3�����n�5�i��*�O+�tRrja��֕��Aw�|A��T��	���T�?<v���}�wn������H&�����	��=����+��H<����v��S9E���䤢��&�����v����]Ѝ[����C�}�Z�z�<h,������$x���r�v�0������3kh�/X��WMIG��-<�}_I-�*?N�?k���@��B���["����9/%q�3݆�&��]tb��vE߭ưM�ɬ�FؕL�=�yr��d�?��t�5w�p�쏮c�9;�*P<�,8R����1[�No�,R��E!�	9�S�*���i�XS%���,��b-���2�Ns&w�^t�d-�lŉ(�����Сk��4��r#�����
ghkiF"���So���_b���TF�+2������ڜ���ĕ[���!�>`�M&��=��.����jf�=��w1�l�cld-d��+W0��2�{�ŗ��7!J{PQ��RR�_&/i��e7��#d*{�|^g&�K�>��]���eɀ�"l�o�H���=洊�?��3��)�j���\.�N)a}���DkMgvas^�BBr��ʲ�.F"i|�}UպO
�R��̚��:P^���@Uu�dsl@3i���������0I���!*��1$2DJ��sJfT)�\��2�6/:�������;���"�W7r����"��;�������(��|�];a��6��;�E�ًB"���Oq����L��E8�؎��Fݐ\��-�}.�B�e"�pǘ���<~@r�"�GF૮Ѣ|ym�^X��=Ŷw���#Q�7�So�f������my����CA�י�99�PS�ڂ"��@����ى��?I%�I��û�y�6��y��Ӵ�E�D�U���C���� ����R!�������s�l<`�v�T2�)NwV��/M�:�Fh�@�E٫�sX���N�_8w^�p*�1�ʽ�x���d1�۫"N��Œ��R�lX�9!��Q�t�,�l���gَ}�C��7�j���M�hl�������)bVwW'Bu5�ȋ$��~>|������-�z�FA
of��������\����|��I���`v��޽-ol�GL�i5c�P�l�Ŵ�d׫��lS~�j\�$�Q�So���]��:�T�i�@�3٬�n]�[ڛ7�!��;�!���Ԡ��qfh�0�)T��Vj�g�M&��zޖf�kj$�9�� �}�lF���CLL�B���A�67*��!�ds����Y�i�b#�儔HI3KdB뙴$��}^xU2��5[a2��愬)��MŦ��DP,W yÂ��ŝ���<��	��!["�lvφ�c�étF�]	B�TR�KJ�b�&UX��Vc��Q1̹��A�I���k��7���̤Y�vPb��"�aJ�l�TFp9B��s�،}����3�D�jij��z�5~���a9�$ȝ�?�(d��:�����GJ��Ћ;<~1�H*��/��~�3�����2�+7�+�:_�km��#jX��ӳT`����n5��^����eFx�S��'��"gJ6Y���-��2ai�	�!B������4El&U�	&PQ�`����L����Ǭ�m�����[6�|���_ϸ2I���S�e`銓��
rc�d�=ͯA䍱�K+�������d\(w�%�O�1V�)$]&^DT������St�8F�5�{�㱸�|��#�9���üb6]F�a��BR|U �ߙ-�����pW��n��?	���OϽ\Y�˩��3	I�����C���]'\�"j�N�56�'����ǣ{�{wocq~V��e�`5v�J¢��ފݻw�#����@'���?�s/_��]I�/
'a^Tv5\�3R�E��<������zd�]W_+X"��ޤ��I6x$5����zt!����5}��o��D(�O��G��Q�̓��q��<�x��ێ��������l&�o¤]�f�k�N8VD��Q>{� F�:��&4	�կ5u��$�g�C8N�!&��@(�N,���KJ��Lf�ϟ:�I�6o�|J��wnbbeEE���+¼y�;уZ�ue�u�!͇�d�b��*��L^.L��ط_L���l����Ǖ\��]��}���Ӄ��l���#D6ԙ��܉�c����}�+�m�Ƣ(8\�0��@���Ȏ>q
���X��Q�~�lL�04<8����Vf�4���<j 9�ӷ���e\�{ӫa�ӈ�p���}���E�C�|�2�ܻ#^���!?z�v�Q�rz�'a.�<c�^%E,��fV��z�-f«�3���
���ᩳyk�؉bl�)<~�'���k��Cu���V�a2���=_V�+����̞e�TJ��	WךL�Ps�D��5&d'=x� �B��_Sl%ҒS�BH�v����-D77�O&u�Ry c�e#��
�u_fsy�3�����3�a+{l���/�jq��a&{�9�{qykE���L�ij77���.=�D�h�� ��-�$MF3h�El;�C����Ο��3g��X�x4�Wo_��?�bxI�2	֡�)$}�v����.�lǃ�P(���l�"��������a?&���JNe|�X$�Ӭ��Y��r��>�$�]N��s2%������6Cs��&��%i	[��}@Mkc�Vrʜ~��������a�-�˰���h��x?���H���+��w�s�o��ZP�;*�JV��7{�Jm�Y�77����4^�l�p�Ďfַ���a�Y,	��~׸�e��P=5Ȑ1�a�h�t����v!��w��0df��fP�}t��!^Iq�����$]�����?�����;�/����?��^;��YD����9	�p�����F|��\8|�dϟ<ă{w�^�S�� �;Yd��	�Ji7<00����v�\V�'-N��5ී�zhH��UWIwL(�Ł�Ir��'�'��n��o$:k�5���sBBө$�v�{{����~\X\���jiş�����n�&�ѓǸz�:��G�e�0�K�a�KJ3�T¤bM�%Ih�D�e�>�p��;;�����k_��_K*����0����ѮQzW�u¨��    IDAT$�0H!���S7����E�7^\<y�Ξ����(�s����y�<4�Y8]-��i�gcE�o%T���(u���t���pܛ5x8�� ����d4��%R[Qd&��7:e�r��>H/a ��`;���ך�T�ZZ����x�������9]ȱc/�D <u� ><u��i\���{7q��5=0�������?"����4٧
��Ц�{�go�����ѽ�����"�|}��޿+^��}{qx�>����F�`�_�N�s�h�L
�TJ��s�K�\]�Ld.��u�(׷���T
o&���gx1�K�M2�hj@SW;��Q{�/�����Xd[��0k¶�����֊��VIo�������V�`F|G��U��6@��(Õ,���N��C�k�1y�D?�H,���E���H�,�:.x��K���x��9pMM�: g�sx��%r�2�^�X�K�a!$Z��XDKc�B8³�}9���(рr�S~Ylڋ������h� �bb�������ʢ��E�-h#B�ޮ��&�3�HmĐ�Č����?����N,�gϜס�t�%�޺���x6]I��RԺ���e�#}z2-r�f�9�}���>��),$��
j��H�}f�4�H���I�M��$P�tF�ZX5�2	�BW��Y��B�~�>F�Ε��!��	�Rl-=0���[���ኑ��8%�P��O+X�c�^�Y�lxiV��2��aB��D}�~8��Y0+`��I�Ne�$Fv�e{)�2�+Zf*{�w�bNh��5'fʣؼ2Տ�8%����˃]]�����o���W���K�9�8�r@!��x`���*���(;��Ј�9��E��ŋ'����==D�	WUaqi����H)omm���d���it��d׼�����5�������;�N��H@��ɥi�7K"�@uM��@+P�J����Y���s���$�ˍ��z%Z�1�����ֆ?�W�=݂��=0E���]vdx3x�(p���XE�0�e��"�i�/�W��|��'�c���DT����5��bg_H�p�e�?:�[$���u���y�����a�7n��L�\Ю�ܙS2*aD�Ͽ���"�4x�ގ2'�]��Z{6*�Ɇ��(R�	��.�m��8}�:j���`{uMc�"��*�j���10Їֶ&�3)D�;��)ѿٯɍ8w@��r�
��)���+�2����p���55`ei7n_ǥ�W�1��0�Q��5 E�H0?\�S.k|hY�ޒ����q���Q�6:����D�$�pxW�_�N��zǎݻDګ&���Pf��hv��l
�b����x�8����:�p��I�L|�[^)�Տ޾B�1��֐���>�MbHr�~�ˈ�@�h�j��x�[Z���ݍ����%�[�����9��ő�CT,򊾔�SJ�*��wN��t`W�<r���16*D�����[��3[��e�l�T�s%�4qz=�� N<,8�d��o�x�9\�>�kHr��ē:��]W[���ҟ���xp㶚^��`�~ʡ({���EA�\y�Ķ�v�~��ϰ��h��ː+RGOBm�פ|���l-� ��͂�_>@,r6�����Q9i��<{5���ob���D�4�|nleVK�Eͪ��LV1�t6��ˁD{nJ��$��"y����c�!��J�Y�YE�9�4�7j}�B��"\��,��j�̴k$F�^�2ڰ��ռZE�fDYK�l�Sd>����B�F�h	
eyR���H��j�@m@�?�E���	[p4/��>���pT��VW�!Ǿ��٘(����B�s��˝:v^G!EJ�*�Jl�:"�!�1D��	9G̿����`uu�\�M_vw���g��߾Y�_|���//�x*�~:��.�c:b_�����W�p=>�p���ݍ�E��QBD��VL+h�@��߉E�H E��,�l�ɸ�C6����2��hf`�wt�P�v\�ë� ��whO�ݯ����4�1 IP�iBF����������M6wcO�+�hl|E���I8S!f��b��q�y�(尣��by>\8qg����A�	ܺuWn\�o�t2-���`�6��c��4���o��YXT�- �N"�����8s�ܯ����[��������u�����ܤ
4H��(��.pZ%ZIJ����$\������H{'F;{0�ցB4��u�����*)!iim�����G�UScP�o4Ss����9�~���d�I���4n=}�gӓ��&<��./��هs'N����+K��]���������'80�W�Ry��/8=&H�{0���ڒQ˃�/0����:m��Hp4�Y��M���/�ե��^��G�{dXE���Ȧ���E>��
��3�1I�\�Y�E�Jj��o#�͡��߿��kC��|-n����K\��Ȣ�������ܑ�S�w �)�i{c�<�rPb�4}pɱ���0>Mc�i�b�`�NEX��l�X"w�HX��鐮|�[jù�;e���3��p)�G��憊0����>���]�7�^�������ʇ�Ls���>���g�T��T���|��;�4qz��?�B�a�Gl�TŦ��ӈ67������~��?��������&4������≔y�˫��m ���M#O���P.�l�����}_��	�����%��ڂ��^x^CӥS���1"Q$2匧�b-5��1w¥\��FS���	u!!��;坔X�|?ؤXE�d�А�3ް���_5b.�Zf��
xPz�9O5�W^��Ѵ�Ϻ_*llM���Ng���y��ׁ�4�{�m+P0}�-�&گr������q��g��ou�P!Bʔsq]�b��o��ѫ���m<W�|�VL����ϐ��k�&���9�<�.L
��@WO�|ݩ_�x9�`m�/�;z�����_��'��|��N>[^��ɍ�w�f'�Ҙt;Kv�sExv��e�@�����s8u�(�����s�Xʼ(��X��&��DM���M����<[S�m���$����	��D��Q��u��&muq+ka}.��#�!k����]˥��f�`�i�0j@��:�\Q�?S sﮮn����+��yܻSټO^���"-i�et�"�R���$Ex�Y���l+YDΝ<���w�\����k�v�
���C�7����t�Q�iT��D4k�������"2X2����N��A2�Qƭ7���+�ZY�������_�a���A��́�+j\	��!dT"wN��-��-��m��ӇV��
HD"2E���"��G&w����^��]ax��
���wL,���"�����>~��/_`�&���)�q��\8u
�!�����ۊ�#<G���=ؤ�<r�k"���i�u��e\�K�����a|fZ�q._��Ƒ=������v���|��)6����ߋPC�r���T�QΑ��5֒"��$���Ƈ��g�����a�^ۨ"�Y�$����&�Ø�Z���El�2H��HR�������Gqs��5D�7�����pC#��Bb�S�G���$zy)�~��O[I�(C8�I��3&���&dh�H�b�V.''4�ˣ�,��$;ҳ�����<��:���K�1��EF�R���UN7���ؾ��58�d�������눗r�
5���M�%y��.b���c����$R���U,Nϡ�ʣ��_+*�O�8�ǎH��f���4~��/0���	�������kK&�t0T>���D$�B<g��:5zz��ɛUӣ���G����! O^<���w%w����vz}�(�@�hU��G�UI0?'3�'Z��L�(�>3�E�����<����9�L�ϕ�^xߑx�g�8�DZ���4�����"lHa��F�mp]	}���:�Wh{�kU�+5 Yk��?g<��ͦ�Q���ڊP$���|��w�A��X�u���k�H�#'��vtYtre�{�e�d,�,���V�Wx���0͊өk�3��2�g8�ҷ]�"�j26.p���Ő�����@�?��v�٧�m|�E���c��?~����N��4����c�L�F� W�W� _�.��'����#���x�Ϟ<VYdhR���7hmC<�*�3�5� �QrY����®�ף9Ԡ�-�Laiф@���ͭ�X2�h���bjwm���b�$�/� lzCt(QII,��
�
���T���,��?�$l�4aZ��P�.$琣���2��pÝ*�gs����8{����	��_����������ޡ�����䋗�R�Ix����� ��	�!���_^�'���GU�i2��w��M|}�2f�����1��Y��h#H�''d�����0���\^Ը��	����C-m��؝���XZXD4������E׍�Ԕ�q�ǉtieI>��TB�:�0���9gM��T��>{"3�|���hCU-N:,N�ˋ����&a������k뀷���U�e+��I�$v-�0X��y��U���S+�x;?']kk�YS�����e��8� �,ڧ�w���.Oݱ����v�8����4B��n>�a�cy��௯G�m�b"���Zu����,p]^[���2��I���X�$���x���6�3E�b��0����"��w�����]��9��1��+*в��$�9u(���U�7v��TX�b�����,O�|�|�`e!�o�Mr��T6�NYa����˙)̭�be;�C�p���C�݁]�8�� ���a�~�6V�[@���.��kM����%5c�6'�R��anr�X
�U5A+�Z�q��a�>ym--�1s�'_�+[:؛�;D
��ƹ��{)c\o�TH�;��kkj��K<WZϿO?����'z�<{�k�n�I/Y�)���e�ݰ͹[�����ޝ
Fv�$�BX(�UX������钉���������m���F��IP*�n�be0�3S��p�o��)éSA����W_�:YN��	�aZ�Yk���`�J��g��Z�'���誙�}�7����0�����[L�Z]5CA�M�U`�պVD]��՚z����!�i7*ZT�k3�Ͱ�]��<Wˀ�>�&2��l6�U#/������c���WÈlms"���P���G�l~�E������+���������I��@�xz�"����ޢC�,?l�W���9�=~T��ZxY��AH���g��<�����Z���Nq�ABC.��5ux;�U~�ѓ�fw �JH�`+�n����y,��1�?{���a�dS�?ӛ�E� oB�*^������������ |~�B���?Q"��g���)�P!'{6$��4�?d��bc@�R�ݔ]� �9v珝���{`+eq��u\��?�N����ݧ����w�2�7Y]}����RQ�����$L]�����ԙ�8r��`�[�o)���f_�i2
��nN�=ѭlzfF6�4e��:X��˫Ԣ������A�����5�B��f�9=0^WZ��3mn���Kk+rBc<d:�ԡ�i�gx���������x�j\��LAE���g�é����+L����|���,��������87<�8���y���+��l͝��][JI5�,����;��p��ܿ�ETW�1�ׇ�{�H���F.��^��6��~*��/_h¶W�li��&���0�c;h
��Ӌ�9B��Ǜ�����B|�[�v��
���#O+�`{eM�!`�hy�t��cxh@0t=a;5�f/G�)1W+�O�R�I��\��ؤB�l%��L@�"n+�oC��]�Ȝn�i�@�a6�g�S��4(�]]���[%�-�����C֯M֭��G�Z��*����k���%�*�S=zw�BϮ!�l��)�"D�qyIG�H1�`CG]�\ks����+�ܩ3hj�G�֡3��/~�D>���:{{���N���ѝ�H8����fd�uWK�,<_=}���w�ݏ>�G~�"���c\�}/&_��fCϳEV���8*�e%�q�d���X�"QWDM��E;���p��H��Q�,�-"�Շˣ��l,K�Y`�P�Cu��BHdRȽ��Ҙ�XEXT%t��O�7�r�����+�W�AŠ�EX���>I�V�0��	�����~�1�M)w��ц3�b�&�02?��"��$s���@���8|���@/i����KgRx��&''uO�֯���ԕo�zQæ�k~�@�/%�T�-5%U�\gzA�@xo�.-�������w��lt4����饡�jy�(��ܫ�V�7�Q?�9M-͸x�4�;{��,5��$���,\����fZ�9�FW�P � ��'���N�X��[fxٌ�>�Yc"�tf?҄@��re��ԍ�r�r��g1��>�|�7~��������D� ����ܾ����)��]��ȶ8i�)�L��2y��|�m��\�=~��ޭ��ֵ����W�C�����BC�-�'&Q���ݭ���Z~Չt��Z�5���ؑ؝7֡�Gp��	���gܼs��^����,
����{�ؕ�Wb����9�Yd1gv�n�;��W��a0l��<h��_��o���7�X,�4��G���f��3+�㩓��ֿ7�#��.��������[�
�����X��;:U�g��p�M[��=ɋ�����]��&`W:���6�'�q:���(H��.=yّ����uDKg�v�k��[\P���Ɔآ��vw!�ڂ���x93��3��U(�7E���]��&&�ceiO_<ŗ���Ozw7w���]��<����҇��i��0|��<�;;�ux���EM/����Ə>��P@��_��w�>���"�	=��g1���ө�Og$$6ylΨ%�ZYF������x9;�l���d#~�G�����W�&����kL�/���(�� 
�2N�22�(g�jB����֌��l�cW0`&)�ek�"L��u���F��E�M�Z��Kl\������2EV<�'Y�lb���2�`�H�2�W��+��7/el���+Y�|ܐÍCg��B6u���)����q�K+������]C�p�8arm),׌���Y���k�đ�����,��)ܾr���'�2dc�������+����Ds38\� JN Ms�bA+	jp����\dD��%d��������mܺyS���1�<}���9I2�@KS�TcqCZc���1-FvѤ��'C�m=.�M^י���3� �!�M]ɗq����T
�hܘ��|*���U����i�(*I8]r���[b���k%��n>�4L�2�Qئ ��T������[[j<X���"�D��'Zm�3�$ˉ�Œ����:a�U-��PNʴ	=7j�1|\YlZ����r�&�4O������//��(�/���	s�bɄQ.r5@B�K1��)����c,ml���8�}����Կ�OΝ;����������ѿV�Ȕ�D��YwR,�ܑt46�0����:��T�B���t��^Hn&t{ក�{��*���m�#k�%�K���Z��q��$���NM�k½�)�M��>vU���{�9;C�"�J�gj=��qӿs��-�1���o�>��ׯt�V�C��e�&I��<��=�*�1��KYC����uܸx燇E����]|��/%�hmk�~z���I��Ʀ�C�u@[���Q��'�H��+�q��+�/�֭[�t�"�������+,n����9�&2Yz;NLb��f�L&��20�T�X��}���D��#��7W�G/�=�Ծek���y�pY�@6���7w�hǲ��cX���gf1��ۇ���Hv����^��`lnN�v�qw���!��;׮!�aqiϞ=�����T(֡y�oX�p/��3�;������9,/,cue�B	��m8�f���l��?��4�������������\]A,҄fh�g�(~��nfj
飔i=nL..biw��fDP�yu�0��?��O���"��7/���#�Z��92rd�8�^d�4�Ul!�Y�A���i"oki��5�6�/�    IDATƼBdcG��eާ,X\eЬ��3v��%�W�K�a�^��FI�3+M�:�h�X�.�׃�J���>�drs���=.r
�}��g����/���x�Wp��WIaGF�ʘ (@׿����G��{3t�
znJ"��O(��1Sfj�Cg�9�J���s�������m����,�xIMR���;����ג�P�Sw�ԄhcR\Ƃf���8#�-f�g�P��p}8��S����׮\�ّ�bOON���ӧx���I����Tc{i�Nu�J>G-*M:8��=c�Z����Ζ<�9rG�b�B9������r�����g���f����`¬j��.s�hj��֔� Kl3���� �� ���k�]��)�\b�����/{*VP�`���;�OH&c�c���?�Ή#DH�g�qEHF�zl8�&j�k��q�m���O~"R$������rq�S�h�	ܐ�"������ǐ{�ۣ�P�o� b��6͆=ӫ�o.�:�;9�k+x��o0��w�5��߿y�~��7���-��o���I�7 w9n��A����H�������>��w�Zu2��á�Txjؤ1#�D����At�C�|��7��b��]ݏ�՛ǡ���]";�
;h��I{դw� ��މh��UQ��Af7kUgސ�X鷻st���,,-�F)+�<	��~U7��0NP{�e��c��}�n^�"B�_y����'���d˄���u5�'i��%�}�LB>����P��ffG����+�s�6.������op1���z����:e�z�i���*��~&-���o.v�-��j�BW�^�I�ӈW�����ԇ�B1����9u�|�Y��b�$��7$%E`xF�T�!������A��r��F<x�K��^^��Y1W���AoS>�qw�]7ExaO�<��_�"��;��#8���J���5�<ډ�w������:��Puz�7<��ǇÓ���Y�G����JLZ]_�w�ػ7ؠ�q!��.`C�N�X�E�����%T�.L//cyu����(��o=�5fg'~�'?U���ӗ/p��}<{g8�t.�/�a������������N���G�i!Ad�VʺΉ�0zj�azixTL�v*�U�3�Q�edh��|5����v�5��$�
�7�ߒ��+W����"���t���]X�l'E����ɽ��]=�:2���gP+�87�Ͼ�{;"�9B~1��D��@�ʓZM�59%��]s �tk@� g�� �3��8��c"p�51򹣞]^�(�r��8<���a5Q���F�L�>[��0�$)K���w��M�"+�O���G����S�Ex���w�G�|�������}8'F:�)`fc�p(����uMlI�DN��r������x,� 2�iw��_ �&჏)Jt���ơ��;M�>��X��1���-Q��
��Y��I�Jh2��ba)Tj��rQ����B�"�3���~�l)��,�$@�
�jYX���?��8;:��&}����ff�ͥ�8lNTT9�U��B"Ԓ��� �sp(.
L�~l�Y��Y˯ҼV2�miԍ�-L.����"e�������ůc'���y5��?L�,��	C��/�(X����HE���Zs��H;:�_?@�%*�*%Dw	�Pv-Vj�,�a\��w�Q;� R�I	Pԕ�o��'w�"�Ԍ)/j٫��>�jAʢ�[N=|�Yl��$�m���c�`��<��r�rSSl���=vE��X|�F&c�;`�c��ګ�]*��+Kx;F	̊
%�7�+�p��yM6�ܻ��~��U�#5�X���}��F2N�P\��J��� ���l�`�d5��ś���܇]9#y���߈y�"|X.��v O�K�������~6�,Sp���ђl���&���$�Ɲ��O���	y2+��7��R򴾾�"�)���Y���¼� �d���h�삷.��=��a�4e�e�B]�:��2˯�@] ���9<~����R!����_f�a_g7�Z[��ݲ�0����5lm�bmmC�3�����k����A�l�~�?�;��������ԛWҜ��������*�蒤D;���GO������%�o�'�d�ut�'��7U�=�`�/|����W�$�Ǩ�|p��x���EH(��GwW��X�Ȱ�*?ɉ$��S����
w�4�Q�N8�|���C����eCfVCN��&��\��rA7$F�J�P��\�k����M(���يh�*<H��^�� 1���\��)���ζ���k�4H	 	��s
�֘�0�E�!� %^|��KS��Z�F�љ�@51��H�i�r�}}&_@U���R���&��X���4ծ D6r0���!5(U�{I6�4b��n�>|�g/�J�S_�@oO~��Ǹxn�r�"�WRz������^��7�w�������G�7��X�X�y�s�L�r��|<����?���c8b�(�����
Z��4Y���&a�i}������z�
���Fey�����xlx�Hs�g&r�����|lonij�'p�|�E�S.Qe���������������)T��3s�	M�|+Q�"%�qgN�kw�,n��D@=yl�u䘴��S�h��.5�\��"�*�#4�Y�����y���9���_�����/�]z���?�/�L8�TWn���&���e�)�2	xd�ν!�"�������):��8��H�}&�W}4�������/�J��bF;Aj�����|L��՛�EX �L�x"�6���;.+�]�v�4����2���^O&E���M�+E�]n-��]�(ז����sr/Lw�|��<��+UL�L���g���c���֩��폔������_����bgG�a/��x�X���rA��\�?قI(��<I6Ų�y�^>?�k�.���K(�ڿ��.^-���p7����+�t�pIY�����.�2|${�èK$�[� ��Ó-�}���$��=�20�S����R$��Q
kۛbV���D{gfHD��Vǻ��&�^�Ѐ`��L
o�~|�=�^�:5M�j������7o!��annZ~�_{�<]�<�d��h
��W*)��tJ��rف��Il��{` �PP��=z,g�����[���P(����K�{���q�lobxp?��S�w��ZSGǂ�Mx6�Oލ��1�(���ܼLIz�:�?�M�|�:����o�ᠴ��	�^��*���7ݻ\���7��#_�q��h����ZA�퓯5�=�C� 
����7�Q�}�B���uŰ�H��m&a�9�A;^S2r�C��$&R�HJB��T���ɩi,�.+G;g6
�.�9�O._�پS�<2� ���l�h�Sq�4+a�Q�b�D�t�0;8��t}PRƵ5�<�8��S�+�ij�pH���!]-(%��H=y�����vB�E^N�,�z��K�J%�x��}��&�	�����k0�8�_�$�T*-���z>Z��w��K�c�f�vb\����x�*..���hT��z�����3���?��\�h��7���f&�&op��lC�6b�^����!x/o��K��]��d&٠~�C纃2*����$ςȉ�!;D8�ز��YId���G���|�v� �ݩ�~�������[�Z�����ذ�y���X4	U�n�3i�̽0��T�Ј�����T��N� �ld~u2i��O�s,��j�ȗ��88���������������K�����^�.�O������p���wӕ��{�-*=�F���5Z��a;?�V�!o�0w��l����2�:3N�071a����S\�s��2^Bvʁ��}��G��ܵ���nE�}�A��B�e^��k}���F����d;������وq����xW�ɚ])'>���E<y��>�N���G�n���[�t�<��#=��'���-���<x]&B���o�B�/c�.���y��̡��A"��*���x��}}/fg��QxPP�'��ok�]�L�S&�	)ҘD4Q'x�!o��:��r�|��,�q��0Nw������`@QbL����������zA�5�D�P='��wS)��2����!��
eM@���m�������ɍ�����ܻO����&���D��xvԄ��jH6$�H�E �n�1ь����1bu8)��Iaum]7%ؿ�[?F���6����=y���$�b���ę�a�ҁS����k���A�����ށ/E �q1��O�!�+f�'?�M�������_����_������ '�aE���b��:��Ԉ��Q����DLV������Y.+�룦��B�XTҋ��5K�
~��Ѱ�:jz�e�(�kg����AO���H�G�?fs�k�\�f����+,���)�9��*pa�4n�^���A$}Ax5's���{��V�V�n�?6��6���!,����ӱy>�|2���)�ϰ����*�F�)i7�(��u.󗔮D$��ɟa\{���S�_>�W_�����1�Ώ�E{S��s�K.YD_N�SJP�O$E��%b�l��`f~�++:�t�L"w���ɺ:$�q�h���>���Klo�2�-A��b3Y��c�����C��=�b��-�v4HO~�umM���[�,Ҝ^�|�xs���.Ml������c��dz�ϓ�$�̒��,�j�Ô#��d�?��KW����M� t����I��Mf>#߷��F�[��ʅ�ۿ�;������=��:�*c@�v((�u��li�:�S���2�:�f������[��f���G/������3ã�8w�������.2�#��+��	/v��~ͮ�:C������Q�~�7��B�,��(��c,�D�	�˩��Y��/.��dEs�L�w��GF�B�ө�"L��.Sb���4Ic*�V���:P�P`�2���s��t��%+�U�T~�����a��j�M������C��E	�xSܠ���+�|��=�g�+!O/�B��\���.��%��L�+�p��`"�HơĊN,<%	9(�4����{��<|�F&����U%�UCu�$�:fN�*�ᎆkI�AJ$��:��C�,L�J��Σ��`sz[��F&�7�'�y����K�snhH2M�V�d�Bx��>_����R�X<�E�ZF��;�E5�p���\��O��D2���2�=���}���#Ч��k�%�5�C�����2֗�T��O�@�]^E����4�OR�H�s�~�?Q` ���_~�Ǐ`nj��z4�r�I�b:�JL3*��><>F]}��v�N�����*䱸���s�XMuȇ{����V��4�Ѱ��X�Y�|��h�o@?m^��0�
%6P%M\����	j�]d�ל�	'�Q5��y�o��bmw[;a'5�t"��)�C�k�=>˘�a^��4�b���G,�T%��9�E��7���B�''T�e�Hß4	Gnv���鳸6z�@P�/��E�--�0-;���J)��>�\ˌՐ��#�C���<g*����*����2�}��ـ9-Jjh��I8Er����0/τrM;o�*X.R�VRQ�.��/_���_���FC"���j�j%_����u	�CE�Ɋ�O&B���j�����r�Ҍ��V���)}�уﰻ�o���;=&�Jf1��1֛J���>��R�,�g�5�|`���_��!���`�[��s�/�K��?��qiK!O~���9qV><Й���n�dI2�����&1��F�I�.Y��X�v�&���Sm<NIS���&밗��������|~!f[͂�Rx���'��ެ�pw�PCE"���=]�/�_��`�����O��������7�����{�#�/`��Y6t����槑#����9:�P��=��'?�j���E��C�P69�nȰf�t��TS�F��Ho�
���4v��s��N��r����A̴�b�l���w��d~�ߖ�%�f]p�_��,��[z8���%����!�t"rr���B�|�.��� ���!����W���7X#����+�p��%�xa���N��%3�%�.�T�I�{�(;68
'��4lS�����$%��~��Q���gO�v�Qq��!����B;f��9�[�ڐ�X �xD��(��9]��^�S�Y�"Ru�>1��=ݤ�U�K�����ކ��aߘ�K?ev�iN����������}�dOdTA6#}����!ݕh��^�oܸ��hD�ݗ�^೻�&��uu�������A�k���WJJ����ց��vh��݃�ww���!�5�u����}�V~�K9s��Uߐ����o5֑F�B�N�J)O	0�������U֓�o侯�����*�4b��5�1�jWGy^�^/��:�i>�Ќ��$�D٬V���M�\�jc�A�<#�h�AS�&�D�d]\;;� 0�{��d%;����|�|��ъa������6N&#�5��{=5��}�k��C:!�]�
Q����&����E�da�i
%���נ|��;�+�{!�$p���9�4Ҝ���s��E�PC���r ���8��keT<�gT��U�������F�����18Ѳ�}��Ξh')BU:��Y�e���ЬF�X,K�����n~v|/��`�$�`sg[�1���7� q�ǂu������[�똛��F�`�P�_4S�b���b��K��f��|�`cO�z-�,h��Ōc�����+���,ȿldP2#����5^rg��b��cw���َ�e*m&�"ɱt¢�C ���9��9�R�����?�M���I4f$���8��B8(�0��,3>o7 �O�8����σb�$n �'N���<N/����������1	�՛��y7�'뻻gΌ����i��8վz��}���m3NR�6DͰ }N��J��`����N������S/�P1I:�]4���mb�����z�C����P�([sog_$$y,�õ<���b&�ޜ$0�NP�U�ν�%	JD�LF=;d^$bZ;$^�f���Ȭ��м��فI.2�ښ[$�~����յ5M:���F�O춮]���-�=���`�O�����K�iX�Msai8����f*M��������e���bbzJA�Ufor���b�_$O4K<.��6egڲ�>~ޙ��K?J��[}"��8�hЁ������Nt�4��q S.c�����3'���û�	,omamy�U��p��C7W��\EOc;>�v?�����^�|!v�����0ї��^���"D��;�"<�{K`�����W��o�#���.����������~�c�$��������o�ݣXYY�!��>R�R��]�!b��v�^��̞�}���m�l��|��bzq1N����M�2�#{9��w�L�PE����N�+JKI�[:hQڗ/�%:�k�\ N{JS*�#-%)�a!�mr���ڡl��}̤.�4)Qf#��H�`H(�H ��'�w��<��n&,�+c�D��JM�NN�t�FS�Ijkh���:N�r���ߋH2�Xs�ѐ�T��UP*���h�^#��ȗPe�{6�ƈ2 �	�1T��}�7�f(�P}��P���oK�rުCʏ*}��6��O��ZQ1��o�'ĂaE�� ��K�/$󷬘��ѱL8I�eO-+}�noIA��G$
~�Y(�hѢ��ś��R��C�X�����|f�U�Ȧ��mm�
!SѨ���E���`!l4>�-Y�I$3ot؍�M�V��^��8A5r�Y���6�u-�˒8�e�����g&�X[ش�6�J�.H���7�����Q��H��ω���H,�X2!�#o�/�H$�D,��#�9�]|�<k��{������ZM;���ɗwƧ��dko���������.U<�_�l	E�Pc����N��8	�\���gF���}cC�O
i3�����*V*?��u�L�D��^ڷYF�>��������/��`���4�T�C.��ô���oB��`���b����Ύ�C�D��߳ ����
$�ǋ/����Ds�{T��    IDAT���$�ˉ�T�L������Fn}co�����w8Jg�'0z�΍�V0<*%��Zic��OȈ����[bxj�m�Lh^��`�$�]p �66�@:�V��I��C�������P2��k�'�z21��&o0`s�� �{�8�����	Z�T��1]��0��$����.�\@�R���1v�5	3�����������'v��cr�)��V���N|z�~x��b쮯�������ϴ[��A������A��FC����Pʞ�Za����"&����ǰ�>���.	I�Ώ��D�����/~��ϟaai^�u_O/ΝFc<� 6J�hB������ߓm�F�DE��vḔ����Db���L�R���/�$.«��}�zN������Ü�����\M��9�2ycѩ�kY�w�<|���0"�{���oe�*Mˊ�NԎ��"�qи܅C�h��9e���������(�Ed���#�����
V�װ����Ў�䞘ϓͅ��$O��46�����:��ܿ���."F�ea���'Y�N�?J��32-e�R�H���C�W�.�Dk��2}���LmK'�)�T�i��EO��M�f�7��/ٷ�d�*���0�U�2!�\��H��q@Ř����AM5r��d�{r"�7�#j�����HN���z��/��g>^����JQ��a�Cـ�r�JŖ�Ѳt����MN��8ĜQՠn����
�]tMR��nd�Q3|��Ҷ�Թ@�����6�3�>��;\p "�i������q����J�,M��:Vf��iu�� t��n�	�c�43������s�5���/�� eb&�;2�0mH���s�������_��>��鹥?���=30t�Ϟ�`g/�"޼y�������4��P��
x�!YM����P�`������PW�����+�'[*�����A8�ĺ���"LX"��zs��ꄑ\��')������qZ��I�F�ds�2���.�^���W�j]}��*A*%�H�/��B��<��I���О�\�";򊚉e� Cx�?��嫸s��/(ğ����O�g<���d���<\9�0N�$/����K�|�90��l'}���%=�\�"c��N��`���Z�X�ign;�9�UK�$�󂿋�Rk���L'�y��-����v��OF�嚊`S]������hko���L�tJ��,<��]Z��o1�0��׫Ʉ,zu�̡�9�Yߊ��_Ǐ��Bk<���-�}�?��ϰ���t6��a��Op1M1��poD���b�	�!�Ig�x��_f�lNE�l� ~��m4�b8����{_���[���~3����[O[�^��\1�s�frQ):9B@���` �jYьl:��VDN�]ʓ9]�H�f1��ZS���PzS�dQ+�;ɢ�Pu�<�H�$�9oE\ ���'��E��;QbB��0.�����mHtG{�@H{lMƉ��&Ѥ����"��{��H�ڭY�ME&����2h��3��B��捫��p�GM��ن�h��B�!��8AE���M\��T�\U�f�0���>�;�p�q��fe,<�;�UUv��� \_gt܉�8��p��i�_%�����Q��h-bO|<DV�}Coh�)C򷦞�n�9�r�&��d.~���."6���JES��Ȃӽ�eY�	�f�Ntr=��'�Ֆɥ�\4��f�s{g��v҂������X�/���E����H��s��~���}�b2��Ĝ��(98Y��z?)M�UEHc�u��H�:��PH:�Ӷ��������<y�k�Ow���ɍ�=	�������ƣF�IU�k��w!�����I�����ٸI�b|k���ۺ������{��U~��v�q��[S��vsggd`hD����^ŷ�������biy^�v��O�����`T�Wt���hE;]�8%��"ȗx�U������}$�v��ڪ���u����A$M�X;����*v��t��a�I���сn6��O;:B�;�d� �DN+b=���
��E3���:2�ޓ�|n1�d�kU@��y�$�L�Lk?�u{7��*�$����IG84|W�^Eoo�Il*�����INR�Q6-a?���!�{?OjB��#� 3����,�v^������)j�g1�����W��EJ�JƊ�a^�j��B�����^ռQ���xwv����Ε�;!aj�>^�pI��L�b��F�И <5��I�&qx\H��X^]�ӗ�057��!B�$� �\(��c�����p{}��=�{�
?��ϰ��&8��j����o甔>Ih�VD!���R:�;C�@�0܁ �vw���,o�ݹ��?���=|�͗�����޾���'���@"���l��j���t C�wN�/��D��'qD#~���Z�zx�KE��q��,r&#1L"�� p��(��4�f�O�:�&���&�"��޹,�ۣv_Zb�K�2_3��PA��d�]�-_�`Zy�ވ���H��'tNv���A�{�J�eA.B�Ti��uc����#q$Hأ�܆���i3[��o��H�־n����)G%�a��f����W9����N6wQI��@rI��@�y��e3�t���͍��#�z�~Er��8*����d�ZX��R����=Q��&��&�*v���(NVt����hOˈ��sk�,�
�<�Xȍ����d�rz��[��b�/6������ЈL*m��3q�4FD��\/��Y�W���;�bf�mˊ��w�Zw}�#��Q-�a+���f�ƖgZ�W�K��W�����W~�4�Z�mkR���6a���;>���B�ͭ$����S=7i�ɻ���Jy�$3���u���5�I{���	�����$�H�A�N՚�IyO������*����D_�w�������_�{�"�W�޻�va����?�;0�ё�8��-S��������d�@t��]f\����ӣ��2���=��k0�h��Je���=8��e(B�>��XX^��N���d67�����r^��ڎ)�z��d/Hhv|⍼��!�/+�o�.e����w6aq��+f�`ѢN�<��듍"���Κ��01	X~����6D�1cX,�|���Wx��!2�._��"L�:ulS�x��9������z-܍:D�8]7����=�X<y�����$SXD���!�V6]��r��L9�m=Ȁ�$���cJxp�<��ʖ��?�U���DV3B}��++x��ӧ���b�o���ql��I�q��%�S#���ku�(��i�s����4ӇύL.���-�|�+��888T�J_�L�2������z\9�ܺ���vlo���'�{��.'��,ǃ��.iػ<,�8*y9N*�(��� �֊*c�|A
EɎ���ik�+W�����}�w�o��h����� B�^�ɹ^%ZQ�
��$�_, �#L9Q8���o^<�	���ZTH`�5���6��2FIFh|V���{��Ϣ������T��m�_x��[@/B�u��&u>WNQ)F]z}�Ɉ4�!r�I�T��x�������0�$�Uae�����E\	FL$��{h�K���ȉI�����/0:ͯ�h%Q`����i�Y���2-H�5��)�k8aE��+����xx��A
��m�sey�K*zZk� �N@�Z��hlo�~�S0w´���MT�����+(+,���S�,�c�Y��KdNqS̽m&F��y}��@6��(��3�T��!P�V�sD��O��{Xޫ�������S��UD�N��T�/d��'k�\аA�$vӤ�{c�϶��-oҹB���������K�f�%����Aq��l��mb��v�&�lO�f�����s��"��Y�0��3����!�#Y�R�ޜ�����w� �\�?~�>��t�M�:��|�S�Ǩ0Q)_Թ�)��7�����/Ow����:����.�-������hW?Ν�HW�����gF��4#:���C�č�71pj�\�L��0�ۃ�d�XTP�:�bIF�ǺQiI�ԅ../`v~k��s�?�>р��p�ŋ� �́�/(�M�i���������*[�Ei3&{G����� )!jjk1i>��J��!���irrRP5/��9���r��4������}i����@���.��?FkK��"���\9�k׮���QR�t�G�{��,�ܯ�@.��[*�;6��5	�O�E/d3���R�W�����I�Ɲ��<���c˦��4b'���KR��=���H	[�9�s���zF'.��*K�tm�*�o��cG}�ЙӒ<���R�Ģz�Q�!�q)c���������nʉ�
�\�.� O���h~p�
>�s�-M�������w�����]��gH6e���r?JȾB�a���!Ӥ���8!�p�����������@��B�x��/cva{���}v�����qFꑠV(�0���<�S�H�f��h���1^�L!G���k&�U���d����)�@��ɒ�դ�%]��T,�4J���2M4}���b��*#� �AI��4"�%�}����Gv���s9�t�k����8Y��K)N����� 1?sN�ԀsR�#:=^���$�)WTX%�c��r W��|��ˊ�dQΔ
���,��Z	�4t�!�� �xE�/�$�eCJ�OB����S8^߆'_F��Jޠ(rݣ	��Og��ނ��445jM�B����L�dF3�xp���e�2YpO�8��n�i�Y1�RM��Y�ݮ�Y;�0a%�o,�D�XXK3~PyOr7.n�=��)�||}6�艜h�[S��؆�M���ey�K��(f�t�;����4���ő�L�\:3�g@�"�5��ưw����Qq�'k[JR����Q�<�l~�D!�w8$�(��:�Ɨ�k&�[-�(�+"�,�)J�4����C$�U��[�A5#8ia�ح"L�=O�ni~��7~y�����������ͅ�S�������gό�lO?��^�|���caqFTq��I ����퇣iR;;t�-�H�c�g�tw|b���N�Z�prЧ"L����4V�����#;ƈ?���Ɔ�t�LɠKU�ִE�#�_~�<�L��.�>�$x�t&�����S�$i��?���eO����>�:uJp�4w�t�j�0��vvΉ$�d�*A����M|��^�}��j��E|��GhkiU<����=y�I���+hiiB���vujzB1u�B�\��EM�,��<@SCښ�������,�����A��lj�k�z5� �;���"j�\�܉�a:w}u��s%��"0�I�zbL�9ʱF�G�O��aic��ں;����^Y'=���ĮJN!�]䌯,����f��)Qc�/�}�v�Ƶ���t47 ���٩1|��]LMM`�###�~�&FN��Z��4�⠗:ꪢ�8����X���]|Riٜv6���i��!���1�N����
2������vt5����gN2:���0��W�V�^&-w���,nl`ugN
< �J��})[a�=���aw}/���J.1^��J.'��B �f
㵡ݤ�%/]�K��kN1��4�75!M��BH�����0��3y ���bEBɋ�ߜ���J�Ƃ1)cb�K%@���@ �hL�?�1M�0n\������F�RT����,���{HMc�"�)�pt}gm͚�K���E�jZ���*�q�7�˫[�*�Q�P֤,/wB���ɓBN�]�zE��a�	��ϩ[��@�;��R�;��3�W�&ZU4S�m[�B/��=	��m�RY�$�$ه���E���ʇ����Φ7?����'JM���E�r���4˄�m�^��%�"���X,�\iq����ks^v�:���q+4���忳�`��x~Y���mhZ\����4mM�Ĺ.㺲d�EI�#;�+�P �(I�!�-lΉ����9Fb���e�JN��ݨ�nUN�
Z�r��7�x�����Xd�P���\ׂ˃�����m����:��{t���٩?]�ٻ�yꔊ��SC��L&�n�{PNçNK�wy����L�=�����DSC��(�[�{��?�^,N[�����R��҂
����V7��t�_d&>C�i��ɛ?�����o|�/�r�v�:��$G'i47�"���u�Ԏ]�zE����.�s#geIȩ���ʊ �H4����F��1�䬍��z�F;Cބ9�}����Y�߾~��zx7o]Gkk3�v����k<|t_Vn��4�]����Ύ����S��\�X�uwu��E�
'���=]���{�.Xp�1�wir��L�~��J/�x<*��ql����ur��/j�m�=��ۇ�|ZI7�={���y�9�s�Ϣ��];U�}�Y$����H! L�#'x�(�8o iv���>��/bll\{vBњ9V�h���+������nmF1s���)|��g{�ZA.\��[wpzhX7�C< #� 
�2�!cyT)a����V�v$�b��?��ۈ�V{'�|���y9�I"��hFiҒ�!�	�� ��\jO]�>>����I��<�d��(L��-���>E{�Q�A�oRG�c�mNݹ"�Gvt�$nF���<�}4c�H�a�(�Z<�i�Rߨi5�i��k��R��.'$)R�����`�a�6l�vwT����s��i���Ʀ�cQ�77#���^��[0P=B���H',�
`mGҭ��ul����>��Ϊc�mͨ�h5�v��a�)t��"�-!D9_����%��Y
�G�jѩ��:�%����c�Y8������I��<p6>$a�J4
0�}r�Ss�Bl�����r�"\�A����n�ڃ����,C�lN�&޷$։�a���GV4eK���Yp�Z��֟��.���O�k��X�j�X�h{��n��Ւo�&��?^�,��b�x�qn֋6����������j ��0�9�>[�d���д�K�i?o��4݄�e)��e��}D ���{AE��0�~7�=�u4"ܘ�I5o�0�U�Y�����k8����F�,ǹ�p{}×�m]�k)���ޥ7����w�p4e5�*��������w2�Pr:��8���G�OJBD��x$����C���.r����=�bq4�����͐8�E3NMarl�����"q��t��=j����M�!H䃮�v�?~�P����]8�?$�����S8�~��w�81vf�����M��@�f��Ό��\I̊�T|	���?��q�)n{S�}��\�&�RWG'v�����E������G�T������cܿ�5�ǩ�(��C��8�޸��/�:8�Y���}]�x=�Z�����Q��1L�%���gR�դPkʋ�7*'�S}�r4���VV�lv�.�O��E-���>4ExzjgϏ*6���;�Mj�I/�?a)�[�3�[0:%"E�sr�b���
:���2&'�������a1�����틗��۷��Ձ�I
��*c�pr�A?�^��"L��lN?�0^0B���.'v�y���`���ۻ�Eb�m��a\F���R�S��n��$����|�ɖ,��HQ{M����#��v{]H
X�ٔ3�u�m[="�L��R�L�Xu� ,�r�ˊIkL.r��*I�d5���;�(�g�"o�9}x(*Q ��i_J4��5�|,��V9KL��kcaJ�M���̞��P�csu���ƶaI�)��!�ԠX���&��t&"I�>�%�[�&��x�EӠ�����,V����F='����&Է��8ړ� S���Q�=���&<,�$8�&e�W[��	xpx-�m�����M�7��XԸ�"Fw?���Ei�U���V�䈐�)NڗѲX���)n�,�=d3�9Mʷ�L�B�,0[֔�4f���຀�9%Nl�������)6�t�c�dg��3��f&nQi�|��u����u����c�f�t�i�E\��Y�-/i�O�.�|�����&{Jf����Œ 	�!:d��������7��f}�bA�j0hiK���4śשF��P$f��B�E��	E`    IDAT��z�Ӎ��%������&�ev����f����/8�GS�*&��6���=z}����W��_�����޻�jz��Vv������+��c����C�L��H�8���։��3�j���I��(� -@ҿ��i�S�����!rJ]S#�O!ZW'8�y���Sx��-֗�t��5��%&}��\*�����Q�����A��������[᳣�h�w��sZ_����2���084$r�h�Pç12tZ-�����s᎕PV&s"��7jli�{�RHx��A:���QZͅ�p��Miei/���k<�}��p�������L����x����XF�tGjllE4V���^�wu�3�d���t��J��f5�~���4���!��v�P�%&w�=]��Q�{I����m=�\ 4���͕+W�=���5�g38Ȝ`veE����6n޼)�<����2�wЉ�r�"�OrP��WV�PΕx-d���tN�c�ǘ�����$�66���ԓ�p��e|��G��@�� �����ݻX��Uf1 O���E>�~Jr�j�耟��N`���,]�*%gr�m���e� q���9L�L�ū�x���Ѱ
f"QC��?����}��S�R��I�(�a�#�|G���'3�4�u	$�!��S�Ā�
�a��3d��C	yr�`�G&�|*-�4%54���I{e�r�lV�d-u��X=��ܨ�_K+��Xk�H�N�����=<|KE���X3��E�ϋ�)�y�d�7�4��T��^~�,�r�Q%Y�ij�`�m,�B�E���f1ɨ��-1Q�)���f$Y�i�i�Ś�TIj")*���+]@~�'˛`A���j���?w�d%90<��x�Z$-Ky��V��=�_����,���Hy3
Z�e�N�~���D9�h9jY���U��>�R/bF�a/[���az���*��M>�	�9�\r��_��_��0��ڃZ�!k55�lh[�dO�r2s��l�zn��S�!��M��:l"�c��EA���KKI��X��r�ˆt�"̿�jQ�y|	��)cqK"��p���B���C��@}_'�}m�6D��u�"̮H,p	�)�t�}�9�{��.(�.��%�_��v�������.�����������~����[�|�SoQ��$�h�o�P�0:�;��Ҧ}�DՄ�j� r*bܗ�����E�I/��_����v�F誳�����i�ќ�$������D.}bE�uI~�������+�ya�9{���*&;��Z�%Wb���T�澗���ޞ��\��3g�h��̄������I�0IF�`mgOE��F88<������o`�o G�x��%={��S=�y���ڱ�0�ׯ����o�Q�&��Ճ��A4�4�!��P�S&���W:���t�LL����tQQfG�M����8���S�Z'���|>�s�#�v}c�8�8'G���e�/����5���iϻ�Ej���+h��0�JE6���4�n�p��hFS��_�T����7�h�K��VVְ�L��*��v��q��%|r�&�:ڐ?:���8��w�3bԓ���7��A��X ��prx���!tvw!�!�r`�����>vK���CwK'�t��G�^1������3LNO���$\��S��d�P����n�N������&���=�{�D��K��~�G+�x0�D8�x ����M�-D�J&[��/�&�?j��Z*)��
���&goG�����T�5��c�$G[Q���i��IJHmdY�	�ӈ��m&g����a  ;?��R'GZ�:����(��soG�qK{�vĜ4x8�!Ɏ�i��$���BW,�|(y��V/lmbfm�;pFC��4 �� x?S)��0�1,&
Q62��"�Zބ;WB�hz�"��0�b�]:w���!����+C[$���">^��*���[
S�x�Y�.����=���ԣ�U^󖇾�V���ӆ���ELa���\(�g:c��1�؁&aH��,Δ~�@��Bݹ��}�~��q��b���<5������Ţj+$� sW�=6'�v����of��wr*��P<y����W�Җ#I�|��ߖ@);�<���9��T���i��csXd��a7��q��`K=�mI8�Ȼ�(��ɠ�3��I��6;����"L� S�x�9h�'��$���\��~�N���ğ���j��YܗZExz�L&:[�0�s
�}��jL4���h�OtI������a
�޾�-�a\�zݽ=""���bsu�h�7vL��-��`�\�JAa�4��P�b,�_�f6�ٳ�p��9�݃C��j�(4�E��/��g�������;w�4�a������E�+p�9V&MH��?�w�"Q�nqwL[��#畒42xG��x��<|���~\�y�������������?W&%%�$kjlFo� z��u���_��ي~Ɲ--��V�<#��޼$b<�9�K8�?����v��F� sr"�����D�
���&f&d*B���ʲn�Ʀf�|���t0
������b�xPܸuK�$��<��D+j�]&�C{O�����h$a�e5��B�����$�D�������wcX���A{��yܹr����X^���$f���/�$�q��p{��5,�G���DK[������z���`�v�p"
���CE��а���r���x;�
�K�Cn�����B�[��Ox}����8ȥ���[$�E����Ǉ0X�AD��$�\��T������*)�,yz�uX2�TDJ�� ��,��"\��]�͂~��O���׃��6�g�4���Ʌ����4%�/i�F���\^j3� ��HPb��$"���9��9�7��`X&�*���O*?��:>_��f3¯���#�y�A������d?����
^�� ���*�� GЇT1��ם�G���	��Ȃ�I�rY�0q����ו�Md��/'B2�y�R�H�X�qܣ��i�B�4�4�
�
 ��*��NSV����@������h�]�(�f����|~�,₣?9�u���'�ł�_��ω�E��y�D*N���!϶�|��R��<!�!�N\D�8�(1`�\�b��>ɶ�鵠mU�x�:�=l�'|�l��Ž�=m�\!۞υ�W8���I]f/V#`� fd\$�)���4 2ɟ�ǲ]ɢg���
~��"�&� r�����Ei�U����p����B��BK,z�+^��)���˯&��luw4��"��š��K�3x��!&߾Rf>���l�BC�a�X|��$���vaso+�;x>����r,���(g�l���m�-/aiv�Ô�ԭ�l��"	���	�MM�g�P!�����)/@�.]AgW�)��ct䚞�D(CcS����g039�s��	�li�c'pd�l3�������ޑ|�$�`,��8��vgt)�p�>�u[�	=H9a�p���On���+����۷H��$��ȽK<V����ho��ޚ�!�=__��/_����7lGo��N����$�r�0==+�p{k���6���l_�>^��&�W�^����"i���FE���蒼�TA�ZV��<tnݹ�+�.K�q@�)-3��w�{d��R�HC�����UCt1{#�qDNU�[_Y���*�6�dzn` �=]��֗����o���+E�q���ݭϑ����u���h�^���h^���:��n�=nl�2���slJ6�tG/.�9��b;X�X���8&��tpW�ܮ@�9]u�*�_�n�㼞V���\�0��"��j�w���&���)3��*�f�01ϖY���0�er���q�)�6�|�I�ah���DB���v�w�����H�p�{,�o���8^��D�l�r�;I�>5AƓ����~��-�&�
����3f	n��^ēI����g�g�Ƹ�&�(Q����>���9f{G�%�\�B�
X����Ζ�z�d\�'l�)���V�|&ސ��,�H��=���
�'"���C��L�ܝ�7p���*|VX�>���=SH���t�q���U�C>��:���*xOª*-L{UKw/(�֝N�y��?�A���5�lwmj��qﴜ��Z3��"Rytk�H��1r@��eA&���ME�E��4����e3��b�=QL�%���ޛ��G��ʚ>}~�>�"�dmsӰ�-5��of���>������gaN�D")��ޚDTj�y�XZ`��V��D��~����-�cJ���>'iZ�)�I	_���j��,���r~
��"JQrn�!�"�!G�����j�������WĈ�{
!/�>�ےl�����ǫ��*����J;����+�'��tm��}>������y�{�c��k'�"|��4%�e��u錈��	�?[��*¯������C�֝���F4�,�Lc��;LOLc���]>Y�-�2��EBF/�}���}>}H,v�����c�͋��B{�jEE�;,^0�nWr���ԇ��E`ymU���G)��0����l�锜�X����'L�Y�}���n��`_?����;|��>�{q���ho�����^����gG����444�.ـ��f��Q�?H�����S�]�������ҔN؟d�����Exwka�/�.,/.!���p��(��u���L�9	��������� �g�Q6�T��������yD�as�}0o&�,�,�r�"ϔ/MB�|1�tG	��#�Q�ɀ�yEř�L�.?�?�Q������mAO[3j��V��Sc��ڕ��WؘQ�{|�����u�����|p2@� ������fu+^�^��cOyʡj��+ofᅧ�U�z1#{fe׌��w|m_]��RKԁM��9g���|߃��$�(6������y�����P�����I���٤O�R����Ţq�tf����;�}P�U��¬��x���)UIy�-y*?��>�q�ͅ�.j}w����¬*Mkr��1�T�Kj��+I�ԕ���GͿڒ�d �Q�!&$%Q|	1��LQn6<��+%7f0�#պ�IG�P��̱cf�����Y9�-���rfN�''�lfNK�ht����&�Lp:,5I$�L���=y4�)��h~s�uT0H�4�V��I�����)�5b��-�k��g��2l�\|#�we�eT�E�^�hvg][��R1��J�ݶ߅M�6fB�A��1������9e�a�a6�F��$|���u�u#_���g~ڇ���+ޙB�*W��H�j�{Z��w��C�I��o��қ�v�.>�R@�BJI���k��m��iIU$�FX�ts#8��o�]	�0O�;�J��#ސ�9��7�ȉ�d��1q��b��C��L�ތ{��rnl��M&S�י�y}$Rn.��o�\�h��x�)�L�,��܀�9e�ߋ��L���Iq�t;�]�f�0�ɡ��bn� ����dU��+���!@�m�_����ão�X��^���#a��n�w;�s&'�yjN�B����Hļ��t�#�������/?�v������u�{pPׯ]ӹ��5=�B�n�G������Sg���mO8,)����Jfȋ��nn���d���J���L�\*����=kk��7/
�b~��Ψ+�J��"���4�dHb�c��ۯ�qYi��d����F��A_ʍH�cxi��ʊ�g�zM�g�����ukgυ���O�=���V��T.���s��[o����u�����{?uRo���&Ɖ�[ѷw��G��Pk>{�F���BJB�]6o��I���W.[�EA~��;L>���ޞ౉�:����={aC�y5��{��o���#�n�0���1�{��)������n,p"���49;���A�:w�$��t�t��5x,"�Ż�Dt"���fKl�Rls:4	�2�_x,�0�@sL�ݙ�����?���VV׃$�����EK�o4;0�=��.��+8����[oj����
���z����7��9�Oͼ��涚�e�q]=}�S�$��W�je��=&B&zB*�ʇ�R��]5���}�`@��n� L�V;�z�R9 ��h%o�Q�n8y�V>���Ο8�s�z��̠���w6����g�����f���T�����:�P�h�L�% ʞ����U��Q$�)	����}��	���:���
2F
<�����u|���뛛Z�\�V�l��xL�\V
qWF�TB͚�*{�k5�Y+i��0瀢��uBG@Z���-���dS�	�	�N�"��$t��y�}�Ξ8��L��4ﳢ��WY���	�}0�5�uC�ryu)�\�F��杽}�����N��Т��?��u�A�x�ϮTpk6-���R� ����6�*�{
����l:�"�/�R,r�?yd]�/��O�]:�,nz��0�I���`�ơ�!|��~�@� ��֜�W������@��������Y��%KPu�@��)�|�����a�%ց�^� $)��}�S�:oh6��{�����4[��NBje▩��`]��"�;�Y_�}|�[^��� �>�/��h���_������0	������W$JxoBf�z�5;f=�|��>�DO�S,����"@?��4��#[8��0�:���O,�r����-�l+���?��wj�����7_~����J�/�|������D���d�{|v��q�07��{��\���tT���}�L����B�-�"Y�t�]łS�p¢�{����Q��(ڷ�l|�HE`��y-��U_�K7��������U�O>�Lc���	���hskUw�|�_~��,-p��NI�s�������N�0��y��i��PW.�O������:~�68W���w����MrA����絻��SgOy�!���+--/k�Z$Dm��Z�� ��2e����5��ę��N�j��RX�J#�vt�m.]����� ~��{�fArHY���G��4P.�
������V�4F��8!�Xx���t9$x�pez
���i��i�	�j��aw�ӣ�~�M3�hz~F�^�,h�BS�[�����>�LLʥlPQiմ�����e<�qH��嚶���j�����M�g����6�@*C�%��$�@ZV.WT� )�ҩ�o��-&U�4�Ng������JH��6���fϿ��MKw��]�y�IE�� ��p�ZǊ�(�hĆ8�C�;�t6erEx��1u���liuwWS�nn��%m�l��%"u���q���^�k��L��q�!�lZ�Bg]�|�nӅ�ʞ�`w��U˞��-0�ᕗ3�s�6���h��ճ�ލ�t�w�.�+�ы}E��sav�m3�9��Z�{)mm���/Ι���<�^�{�;��uja��C����ޒ?b�q3~	�������A|���tZ��>P_O�'B����-ܔ�O�����,������Sk�m@#鄛O���7i6h�{��X����k���;l�)�1'ja ��Ղ��C�N��a�K���!{�P�.@�{W�N���#:���=�ł���\S�� �v����V� 9g(�L�9�����5���/4����LDʧ,���A��I�8o9g�F���Wq��9,����r��?10���,Ĭ����o���73+�W�.¯��d��ɗO����1;a�|8�����w��-��{�{H,��"��!/����Qm�[�D������Ą!���W��n߾e}!�&đ-�N�@붵�J�XHG���_�4���f2���z=ة��1�P�)d8`9��Cχ�
���B����pzt��q�=���"7���Z������>x�-���M�t������ǎ2<::n��ѱ#A���>��C�,/��m&�egΎ�N�fV��Þ�Ϝ<eO����2�[�0�xK�;vn2R��2�V*&y�=�f�t�v�ӯ^��ύ=��=O8��`��?|D����ʾHu�)쎶Cʀ�G&R&tϬ](*c|���r�    IDAT2�v�y/@,� �"�
V�!��_���C�@��ޮ��_~���U��9d�2�N4�	8��Z6ץc�Nh��1E�)'(�+5�/��/Wй��z���n.k���N>׷�51r:���s�g� Ԁ6��1� g6�v�F>�7��  �t"�m�C��MFv�P�����Zq`<z�0�'��zS��y�������^U`չ��yEK����s:�_͖ʭ�Ӝ����
9̚u��֐�b�p WV�`��0�x��@����U� ��Jɤ*�J�[��M���{��i�fyc��,Z�H*�|k���LC���/2C�&�!1�F��nԵT�1�L�:E�C��Z��.�nj��+��c�f��:P� �t+�7�_��o�Й��� ��.���n�3Y�4�;���Ƚ�L���f���QЦ�ʥ]�nnx�\��P������4�@�L��	�n�~�={�/'�RsqE�<3�2���x^�l�3�׋�)��@��,���t�ۻ�d'ܕuscr �0����N�)E:�P_W�FF�}ZY^����?��u2��&N�Iޥv,S�Ʊ�Lx�3^(>��(�|p5�%f|r��#F�c��ɇ׍i��49�WV�}]���ĭ���>�㜱�h��\�yC��^-����[_j����DX���n\�[-w`���W�����I8W&SZ!�g�{�{������3�(�͝�.�{��߼ZZq�v���AS�s�t��o�ͭ/�����U2W:���:��vVμ' �Yҫ�yͭ�*�ݣ2iF-��.b3���܌>��}u�k�>��Qw�3s�
D=�T+{
GT)��I!a�'0�F�Kn�:�}���\��@β�6�r�e�s84��P�Siǰ���v+ѕv�8�f4�@/HM((ཱུMқ�����@޳���`�O?�Lc'-Q::vD��|��~���I�IDS� ��ӊ�c����q�"�,ө�'t��qO��~s�$����!�
,W�}>��g1��K�c!����W��2I�/=��ԫ�9O(K�~��ι���=j�04:Oj,�|>�aGNp�xCw�4�.�ن���,�B���a)�5+k5$�E�Ц�@c��4�-	� <cyQw���g�/��F�m<��N���)����[�����S?y»���5���6�5�7��g.���ok�حrs_�=��|�;��s!O�}rtB��V0��\�Z��E�f����������Y�6} X��E0UT�%KX�P�a��l�c���7��4�hl�OG��4:��Fmؽ��,hiv^k+�����B�a���.E)L�D�F��)�LCe��X8��K�FF��L�=7���|�39K�q�d��(ՕS���ؿ��7q�p((�)�-�4�\;l+�Ʉ���R�=�:�$�\F����ǖw���4\#���(Zj�<��ꆖ_L+\�aR��VD�FX7.\����a�p����f���:b4�ɔr�`o��l��˴W������� I'&&���֗����fi�|&l806��8��0CQ78gн�c~���f��ٗ_�;��0��M$,;Z�b�쳗/��C
v��CM�ΘD	zǤ�����=���%E�)aH�Já��$�����B<P��H��F�47���h4���Ͼ�A]"����(Fcb��t&(��.��"�:��v�`$��Ҹ2F�`�CFc
��� ݯ��������c��t������Q7)�7<7��w>�����Z)��wni����H[�l0p4E��N������m�E��� �B$a�����pbp��o_o�ON���[�r����jq�rW_�]���M�v]K�szp��[��e_(j)��c'�&����"�4 �V��=~�R�dJ��\���?йsgm�����O?��~�����b��1�ϫ��Z�QQ�������w�>~ҍ:6~�M�_���σC�8o*\?�G;{��]��L�Ň��v}G��3��=0�z����G�e���U��\�9������Kk+z��~������ѱa�n�蛻_��_�º\v��rC��*�f�7+-��G�F�-�/�?V��O�S��/�����+w��9;p�!�� ����2���L3 �
��P<���}~�Yߵ���Ke�,/;F��b`xXgO����$�`M���v' ��0���	,
*)��pL�AM��_����T��64��G��T<b[A�W���T�Z��"�Ӡ�KA1���]4�fXO���P�6�17�d��n���w._���yGC����*���=}���>$i`Y�u�	鄶'�ֿB����t,=@.ܯ�{w���#R+H����<:~�!��.���[
�+
ժ�\�HT��.?�Ѿ�ND��L2+s�\[7�]L�:i3�A"nb�QwpE��K�83(�r��!����ףQȓ٠A�U	Sh�����Q.�"<xtT��C���R��Ǝ�VW��KLX����;F2V��0;ڐtO�(慬�=EO�[��wE��F%`�c|adS{�Zx>e�!�h�*�0M�q�7.\�o����g�S@��������^���T������/P7�l������DhqzZ+�s���Z�n��>���M)İ(H@Ս>�g����$�.�_߾�$6t�>S!�K��ď��Pw�f��Z��@Buc����夝ǐ|�D�'�f�G���xn3	��i�Ȩ�<d����=�
�$+�����ps�b�Iӂ��[o�冔�t�իW^=J�(����g
�^�t28�0�$���=A�|�, �r�(n����s��d8o8�v��922������v�Q+y'��n��
Lt�!�S�5E�Y�I��mCT!u��T����ha��3	��۟^����^\�T��wWtpP��̔�|��j�J�5�5�ѱ�q��h{�D��x�hP�q��E�ƭ+%��/��/tbb\����o߹�{h{�`υ3�(���:�3EY{�����t�6��K�����������~���#Q��?뼙��Y��Z�{U�S�@���H"��5:0�j��'�
�9dӅB:��$��6:��~�;�=��7���#��\��o��/���A��U*5CVhJ+��JX���ݫT:��hH�į��ޟ|�\��ZZY�t�G����R|�0�1�o5mx�ɍJ1O@�ù(���0!�W/����?q�M?(�h����|a��|P؟|}:m��t4�l,���kS ` K�Ч���;t��т�gf� �*�vN ��jے���ϞjqiY���FG�[5+��٘�7x�@���@&R���wT�.���q�{����f��{���[_���\�h���i��kuw��%e���{�dʓ,�9�Y�_+OK����A�d뻃C�Z�	2�Y_Q�YV�ZU��PO"���]=wFC=����AC�3Z��5<
�S]:k�{_���jM���ql�TY��bq�q}�V!�1�`��I�@_�z���MaNS�����KUO��V���w��	�����]t@z�&���7z�G;5
�-F��/�o�ؕ�� ���|e���Y��]}��ȿ:EZP���7�hv�4k���c*��m��,�p��UZ��3�s���MP*0�q��@fv�H#��ɉq��2z�⹦�>�;z⤛�|h���j����PA:����546�d���W��ͷ��oy�D��=�H�d���;y���8�������B&����\���W��&0�m�@��/��@3����N�O�=��|���ڕ+N���75�B�S/����:��P�	y������~Y/^<��;ap��&M�w���J�z�)#��lh
?�p�XPO�ǲ�/��b�Y�@��=h�	���67\�9GG�G\�3��ڏ���4���m�鉰-kA�@?8_�02�{��~��J.�T>��l6������o��O�������O��/S�K�u�u���y��BMM>�>������V���ѩ	�1�1"���ۖ&�ե������\��w��|���J�ǎjd`H{;�&���\S�N�"N'�D+VWع�U�onn2����F|�Z��C��i���1l�l9P��n��8t�A��70dx3],(�M���W��7 �3'4R��;m������-/���g���ub��{���j��������b��ۭՕ5��<��cZe܈8Ds�9j�򅜻�C�	t��<�ߑ��g��d �Jӓ\����h��M�
ˬ�6,�|����Z��>Ϟ=k��}P_Ө 4���D�.Q(8;�T{�v�œ�G"<k(�L
��kGJ3@!�=	��T��)�N�\H��f��&E�.�`@]�EDLV�J��Y��ĕ!Sx���z@>g1��}��7�[�S�����������~�i,�0��^sOB4a��y���"���
bX����)��-۲5@m�f�F"�e�;�^w~nV�uEu�J%��5���0zTg�G̈́N'qM�jvzJ˳3����29�RI7��XB;�������,t+��+�J����m;���NG���Lv\�T6m�T�?������JZA�ҕW�+�D��l_��ł!n��/-�y�U=�ƀU��DL�B�C5��d�V6�DwAIHZ���jf6�خ�������K��t�tU�Z� A2���Ķ��W�J�RM������\��ǹ�?��?W��[��_qQ���X[�d��8�9|�˛[�x�Ό�k��G��f�����S�d�2~��0M?����J>wےG��щ�8yR��^=z��)lw�����=8J4 p":,硱Qb��Td�:z�F��+��krf��Z��D�DR�0Lb��2�b�W�"��J��ȄΝ:�b��ɓ��ȥ�I8��NOz���-��x����KW���W�8������ܢW��CZ^Y4�ȳ���a��������}�4{�8�O��Y��/����g~��݆��_z�� �n<w|.x���s���?��@p)¿xG/6����"S-"U#d\C��ј'��"̔�c�z>��O<�����G}�՟���۟���'?5�|Bp4lP�*E��ݯ-S����j����1�w��8!#ӑ�^� 9n�?|��3�Σ'`�֜�����g��@���bR �o�_LX�t�� .F���#J��N\�P�($�< ����`�#:KrD#�v�˚�J1br�Wi����m��|4�l!�ѩ�K��6.웸�a�S�[h=9��a7�>�G}d������2J�]ݻW��/�_3O'N��ܬ��ww����=�Y9��U��Φ��z>_י�Iv��'��v�	l�`��4���ú������>¤��HԨ:k���`.�P���0nz�W4zd���p��IH�=X�����AX�X�7r1�c�U�0��ް�?�JK���o���	�֘��V�� #ܣJUC������i�[A�@.���p%h��� �f��K�l��ҕ��FwC����bU���l��="Л�m_�ti~��wM�b?��}�$�6�h�W]�)������h�X�0��P�h{sM�k+��n+�fMx���tJ'`w�+�EZM�R���e�6w����O&����,8�N���JE�D[��khX�B���x���ǰ��#�>VSq#W�h�ˮR���j]���RŢ���O�M����jc/�6��x�_��i��0̻����U��V8��/�]T��e'8���B���xi��N ٭�݀�[iXB�0=㰅�"����╆Ch޼vUo^y݇/��>�PSK�ޟ^{�M�ym�&�χ�9g�5de(�}�:c�Х��i={���4X&���"A�7�5"#[6�����Ǖ��֣��t��}���vD�|�g�`�10��Y���0:\�,<��Y?��S'�Y���;��ޱ1
E�f�6��b�k,��l�ΌOxG���ӧ�{��w�4K0���q,��"8�� ��N��勯9:tceն�����1P��	�����=8����9�0c�j���MG��� ]�#��$�Iu[�tJg/����q� < �����y��7�������{��)��kG���7��Z�Y橨Mb(­p�;/j�+&b�a�?�I�Ts���0f��Yg
���������?{�ދg?���"|��Ew�/&�����Nn��{��:꜆���+�A�\�jrսG��rnA�%�0�29��'?�ٓ'��]� ��xD��:c�꽳�t�����t�̴�~_m�w����65?7�����(�,����m��$5td�nLRa�2��t���V����B":4�pf-�՚ai|��I��7��,=�{��޽~S?��}?��Ү���V����7�3$�4~�@x�}�(�a�M��h�C:�Zϡ'�'�cO��Z4���,Ԯ���0��&c�E�]3qqѐ���]9%��A�I����$g�5Fb�/�8��:�1�i�I�I*M��u�Rv�1#�>��f�b
e�0]�]34j{B2^���/HH��(u���Z��I��s;dM�5�U�z���CC��{FD�A(�˱��L���4����������s&
'�e����C!��{f��,.�L������Jő��݊vO�y�E�mo۾@�r�� �B>D3��H��X��D���P\#ٴٿ�J�Ȕ���̔�����z`�g2>H1�	�c݄�\��ΞV������1��m4����im--�'�D\�X�~N�x�(H(���qUk-픫Z�+yF�Ո�L�Z�߱�E�~r���ܰ���'9t|����Ąv�+/���V����T\5��T��\hf��m�nkm#�P.���R�Y���NÄ~r E��ɓ���z��5'O���Ň����'_;��gO*_,hku]�dq�]]\P}wO�O��XO�F�=�OjciIs�AXM&ig�C�w
�����517��ޖ{���ѣn�(�S�_X�N�
Î��h��u��[C�G]��d�f���D���O�SA~4��מ"܎��	$>��vX�Hʓc��i�f?z8��h�Pn6����iV&k�
(�@������'�D����Ea� x5GF��̡�ý���ԉ�Zr�S�!��10�A*@g,���}�C�eryg_){�75�J�[�����O~�S쩡�ܿ���u��j��<,��0N�<�LÒ���+�	7ˤfE�����cП��~,����Yt��ǭO޾������_� �$|����$��<����-��]D�=���'t|l�&��8���\.�����sb�Ly?��! W/���#C�c�H��~��"�(8��Չ Cg2Uy��k@�bQ�T}��LNiueŖ��6>P�����	�ᘬ�߼a�7n�q3])�/�5�0g{�$4�o �"�Ih%�th7>pK�t���!�	y��楫�˟��>�RyG��>�����4����m�]�����c�}���cZo2��f��_ڱ
2�fgB�:�+�����!K4��Qh����tT�W<���I�a�)�ceB�,n���x�;\�%��L�D9D\�H��C��'1� ��_w���V#�'S��ŕ�� ���*�D��x���GzttpD�LỨ6^�	1����p�H��!�Q�L
m'���`���F��m˯�U��g��}���ddavF[˫��ܴ�t��ם}%B����S���Zo�Ϗ���8�51� qh7��/)Skh$����ɘ�q
K{�[z9��{s�h��nC�A�c*�BZ����Ɩ�ї��{xX=����+ssZ���>�XD�����9�/Ř\�jG�H)�ɫ\kk}w_s�kj���$��ޮV�ƚ�kjC&1�HG}��\y(�UP����АR}E���c���Q,�Q,���ț�Z��-y� `[;���xͯ--����v�2�ׅ\&o���g��7o�ʅ׼�@W����Z�&�i����#C�p�5[������t���CC^?w^���䴿�n�0Sr46B����'M?��l+f    IDAT�:� �	�qi���}>�J34o[�L�l3�?�< �U+V%�|�. E���8rtL�N�u,�a�ta85&a��@��M�,\��jݙ��?��g�)�L����zxﾑ5,w+�&�i�����	s:��Y��ft��Ο=�� ,@ӿ���b.)�|����(I�|_�@�+�G����`�0���y?�{`��x��{&��u)�=�s�q��--�3�7����O�7:��PS��wKS{A�$��j+<:g8M���ݶ=�a&a�z�fK}���C��?�o��̟���E8_(����t��%%#=zxO��!E���mr�/�SO�G'Ə��7,����bR����d�v��o�ʵ�z��t���Jň�r��O�b�%S����6j&���s��VJ���鼝���\˯��*�2ᰊ�L�	2ɚ�^V*���#�����ßW!ݝ~��OjfmU�ق]���
����5m� F~)�Z= @Db�
�m��o�����G�s̓��������8����Q�����4�M�&Q�T�ʏ�LN���Rؙv���(A<���BM3!L��N(�c=�pg�Ŏ���	�μ��yL�%�F��!
<L,]�3��{HW.t��2		�7M� ���20��a��ZM�m\:�����C6�o�[j�L.�؝�������5������Ⱦt��f T,�gj
�4�8/򨠭b�j~uV/w�$�4��G��/�4����9�&iʀ����@ɠ H�؃��Mn��k� �*i �[�p�!^�}�PW*����=����Sw<�L<�f�jr�����]�˽���V;�(���Z����֞6Ke%����*���i�]]Q����\N�=E� mˤݨ2Ѳ�!�;�+�DT�Ξ��T�Q����,��& �<1n ���&�d�i4l9R#U��㾂
cG��S~xH�ޢR�E�!i���LИ`�u���^���>��zr��;{�ޠq<�pT֥�g�+�a�_�[=�|n2SW�n�wӶ���^��4�:�ݣ������'4�7��tF[K���㨗]�!e�����V#0��Ou[�ۖw���8&8�664��dLo��{x~�ݽ���5;�5ba�5���Ő:�9R�F����׫��9=x�PO�&Ռ��s��l��K��u�B��9͕�t��K�;ȞO?�� � �'�e`�?����E�Ƞ*�����uI�������4<�AZRZ�ˆ��3X�g�U�3Ӿ�![�d�i�'�7��o\�J�����ŵ�V7ֽWF?�D�dBGG�����9��p[���+��]��AC�D�E��0~�V_���� CP�x���J�Mx'o�՛�~1���O���E����������k�|A׮������N�鳇�}�/�ww�g����z7�"$�Z�@_Q=��hz��f!il�(��jys�E�ĩ�z�ݷu��9=}�Xw��ѷ���.t;'�����'�p-gJ���0���:H?A��n��X�ts��w�=���F�$����0#�٩�#7�m�t��C}���6C-0��?�f15�{kqE��˦���aBR"����^��;�o�'�`ȅ�:����TK+��f�}��06
�c.n��V@��<�6����=g"�HR@�A�8}�8Q2��S�5��4R	�Y�t`��r> lx�βS�76ִ���Z�b�"�j�zlsm��k���XT��>}$���:0�m>7����=uI�	�� ��@s��?$��&�����@G��u��Qvt&a&�ΐz(q��ަ]����� Ӊ*���R�%L�"@輾���)�n$<5lhn�V�W�����ֶZ��z�q]+U��t�7���LT�;K����3P(8�Z͚%C��R���j��׉��a��A[���6����1�A�
���=LۻZ����Ύ�p�I��u��UcoW�����z4�WTw.m;Y$%�u���"�{�9��W֋�ymV�~6�Z�����bj[�n�y/������OQ�����U��c��W��w�Q���!�i C�HV!�)j�}�n{j[ZXԃo�hciū V�Z1�ۺx��S���YkW�w�R�>������}z��w���K�\���e	U�6\p=�B�P�+�mY�� ��:�0˗���\H�[��Z�F�|8��jE5������޽{Z�[tW�����f������(W����An��������B:d���Meu��]���'a�Y�ܗ�����	N���9�-$����m[Qbt��iO��ӯ\�==�,�i�������B#d�z	����ߐ�G�,P7��>���3.-zEg�~�1�$��Р�g��>C���~�����{�S�'wV�A�p�IS�M�eP#�C�!������e"�m%���t������৯���_���ƷϞ�����kx_�|M�x�Iӯ^����mֱ��a8�wdxT'������v7�T��4zd@�B��%���/49;�H&�ͽ�ַw��;7�����B:���?|�����-�ƺ?BÝ�ޕL��'LMm
#�(
ց�Hd񾰯XЉ�����hbd��0h/��@rbǐ�e,��&����������sݞ��|��]8���@;����VU^߰-�<@��X�M Gyk�E�G|���N+��zzy9�\���ޙA���G*ż��^.��d:��ń��D��	K8���q�r@-i`��L��L��3Iy�.7bF/0�H�Ę1�m8N2��1�7�����<��9����NE2k��ίL����=]�!�P�׀�5�7�*�'��-�x8x�h(ju�=�60�ggw���c`b��N8�y:����,&�8�)��iH�"���:٣b�f��H$��������t
��Е�LM;_x�ù�^�+~-�����r����q�bW
�a�tǿ�C�Ol8��U�W^H$5V�ֱ�nP�����uF�ݴ�B_��2�D8��NC�S��fG�Yq��J���RJDv���Ry_=鄎�i��K�LRI�1�گ���(��R���v���K���/iO�@�J� �;��0�MpY_N�w�=TH+;<��谆ϞR~�O��~E�)K���~�#q�"+�M*�2@�}���z������Kj�*
�=a�Z���ɓ�~��n�������w���=���.��n���.�=}����0AX��5�!�4Ec�����F�Ϯ�D�s�6�����A���dj���1_
6��"$����w���²6V7�s��
$bf������O&u��)��x��e<HB����ZѠ s)VfX��m���t��(���W-A����W_�]����R)s'Pl�H16�N{��3=��Y^X�Nr䦰��j��y��4)W<鮮,��}�^X#OCR��f��Lkgg�(��ҒM����@w�iOL��	�2R�~�����qU�!���z����v=�	c�d�p��3,q��^G��دyw�QG*V� ��\��b�����{������z9;���k�����+&j,�����[���O���LiM���i]<s��J�`1X]�G� �|N/gf4���h6�խ-��y}�����;7�}��W���7�u箶I� �f�pe;g������)��a�z�i���4Uw.�������.��
*��}W� =�ܣ�E�oW�n���+=�}����z\�P9�4)�S0�PD�VH;K�Z����~U�(QL��@�SN��,�������S��1z��x�O*�3R,ң蠁sv�����.�-��I	�SO{�;�0��1_���f1i˻m�r��U� ����g�+���Ç�ꛯbP��Q"���@6�X9�����OCч,��	�Ə6���LR(��ց�ÇV��������B����r@9q��?�ǎ�sz��L+h2�A��혶�{�t�I�i=���E��3B>�X0�q!M,B7�z�g���2�[�����{e�J� ��Z�G`�v�a���)@�n�����k�=��ha�eu���M$4��h8������V��_+G�Âm0�L�}�'_�����7��� ���>�<���NT���%t�H��z��&��FD��i�DxP^\{u�h�Z���f��u�Q:P�	'��<e��Qs:(�Hp2�43	Ez
�S��:y��NY�IE4 ��'KA�� ��Y����T�Ӡ���\^����\ZQ�TV�gl���N���˺��u0�����a�Ǎ�-����K����M>n��u��憹��CZs|"����J�j��C" {N����c=�=������4F3ഐ�\�,	�Wl!eu���B1c+<8دg/����ֽ����ߙR�<�X3�\"Ƀ!�A���������L����O-);�qJU4�\"a����^?{�{E�v���%��3�~?��)�N�Ja�	���z��p�� [�?t�x?�e ��W/Mf���oha}��C�C��x��������?���M*�~}�͔�<	S���0�bב(y'����Ύ�hM,jAa���~w������7�����|49�/_�-^J�3���M�u�RѨf_M��_�ޝ[���*��"S�v���Ə�����ʲػ�k5�X��D+�P�Э��u'��
�����^�����oo�y������T��F�v.�C-۝!!�7�C+ܢ���%Jf�N׋;ԏ����L�0Ѡf��L!ì>�#�4�=Qjw&���Z8�h�U�Nݧ|�9�\��J� ��icnіw��Z�����w,7߸�����:ylB�v�Lfm;[53tn"y�X$�R��*��z��$�0�.LX=�ФS���J�����<_�`꫹����5�#zd���i��S����=y�<��V�{=XݵF��?��CO�	N�^��h�aV<�<l&އvUΩ���I'�D������9���q{m[���Ɓ�T.��epV*�L���y�J���igk�D
%�0��JC��֡s�E��T'S�{'���<�C�ƶj;;j�1	��2F���3�4�� yo�b����	r���B�F��j8�'`��a�A��;Jd�ޫa`���ܬ��KZ]Yv��ԋ���KD�)���r]nL0�h���*�j��K�}] 2����JU&ڰ�ܯ����Ե�W���6�U��>���+��M\�ԙ�QO��o��2J��wbL���48q�p,�	��p���9�L�}��z�Ȅ��<��bi���FZ����b:���A���.&L��˿s�'d��#��2R�4fav��I�֎�:6��WhԘ��?T	mȣ�IP��A�g��'1�z��>��aex�Hã�p�Cr"��"$&%[�[�}�y��
�
����|��~�{UPt��#��u�TBHzr]��~���yW��.��<y�-�W�T`�y��f,g�)_C�@K2ԯ]��;��*s���3zo�q�#�?'Vl^y.�����S4��uD�D�;�jfn��3��4�\_>~x$�]_���9��d�ӿ�K=6n����Ջ�m��������	�UNy��X����Tm�<Pt��8��|�wǻ���%���~���S��jv��"�����A�z�T����o�r>-�]4z��
Yt_�6"������?ob�}Nٞ>g�n���|��n\WoO��˯�Ч_|���y����:�9 �����}����UW�����57&n��g'N�ıq���P_w�{�V�����F��X�ӕ9ݛ��\e[��k�`q��fH�xFGr�$�"�uD޵;��f�C���Z�~5;��W�E����u�؄2� *�V�(ly� v��N�
ņƣi�x�bK���.4�@����8�!�i(�����ΊL����äG1���DMn-�2���e�,�;��ɓG.�x�����F�� ���&�����	w�a`$�gZ�
&+�H^���q8�k�=����7eP1�̎�(���@8y��N�>�޾>�:������t*�C6gW#�1���_���b�fm_��0���4�6C!�+���x��h�l�ݛk���E��w��
�(l5���a�w�Hu���#��^iw��L��V*A�^���i��u O�G�E��$�گ�����-��*�}�Twv|�>�����|/5�;H��=�9�����>�%%��t��[�}E���7ʪѰ���+�ʨ�k����~U���Z�<�^S��O������@��D���HF��Τ�/(=<��cc*�����'Oͼ�U�d���|P��EѡV3@Q�9�V��`�%���{��D9��o�q#(�K���/���Y����(t��Yɰ{)F_;	՚�T�bH��5Ӂ�t�<߭C:�������R�{��Y�xe�s�(�F���ȽJQ#Y�Fx�Z�Ԍt����׍��5<<hB�/~��>�����Ҁ��xD��d�Z��!����h�L��5��M���'T
}���������ٜ�3@�=�V��5	|���3C$�(�!�	�����Tr~:g M��㍆e�7I�����3�7����W�6#�������0;Z��L�������}Mn�h�YvX�����AgܘxhȺ6T��Tu��"�u¨#��;W�|d������?�ӳ�q�z4=��^�-^��v�7�޵��
59��E��O>��O M���5��9:Jk4�Nqŵ���ì_>���ʆ�K%�{=	�u�u�vw�����Ol�M$TTIPJq��$���7e?ā�_�������E�!nM��P�� ѹS'�4#3�q!�i����̔��N��ƒ�J[Z�Y�)��j��WG{�4�3�#]=�g�#˒1�jچ=[�q���e=y�B�}F��1���[.��d�0�̫���޴�9���~��	��1�@�%�AX1Ӓn���dɻR��t�}J�h�^�] F'+P�I+���֮��L��a�p��i�\W�\��¢&_��˹iw��C��@@�H,�1`�t���z�̞�u8�P�$�t���혀�;;ndV�����冫	iG�̨X((������������m�G����҈�$�1(�%�r`�A�N#r�Tfj�}f(��ZY�h�Zj��ԫZZ]��⢶W�=7wJ���~`�!RØ���k;f�Ih�ݒ�'A�j�IKw^&o6��O��$z�R�H����n�GX���0�ȧ�&���� V�z1���͠a������zyOU�����j�X��.{��L@*��%��gsj��ڨԴ�S��ڦf�6�^���;�T� ����a�0ۈ�Ů7�T����H��o�蠺)ty� �}'�f���a�Q�AA(¤��,�
�Y�O��Q���:�/�v0�h�Jӿ�l���˗=yQh~�ѯu��CM��;W� ͱ�R���M���Z��<��)�K�>�	b�y��!v����1�C*��I�"dw3�� |<Mw
�Ѭ��k344��o��k���*E���Z���wn(�Y?�懞��X`���)��E���[vic����#ݾ}[�K�P�'�ɚh��{��l������|n/tL7xݜg\Ok�C2�N�o2�WmA�qH2eE�?�g�h�l�f* 4+˫�[Zpd�e�ɔ_���ȧf^igO�d`�<~�'�/�?���U���GS��Ji�#�d���0�u�I؞"�h(�i S��Xo�?�n�d�ON��ww?��`��ϧ��.'�Y�u��^?wI��^�L��{�����x�ؖ�y���8ݪ}9>����IB)��_��Ɩ&g���������{z��Օ��S�>����\Q._��ɤ
���c��և-�����gz�౶�6��ID���hܾ�����������OjttȨ 4S�WOug��V���+��Z!=�3�'5�=�	�M*�+�����I�l�N�����ԫ}��_i�o@�_����ƕ�F����'�ի)��v��rȲ���&g��qӅ�34;�9v-(v!w�LT�ݬ��Tx�N���    IDATA� �LL�@9@��,o�&�����0vdD�x�2����E=�L���'�h.�h��ɪ�w�T��
�:<�3�.�/�ot�uFr�q�ZMX��z�pu(�
E�G�ĉj5���9�s�6;��|�S'O�l!��5PWi���������\���\r�?;.��'a���8�G��!0�I����L���ʂ� ��*�׽�B�e5��: y��09ˑ�m���2� p3���.kv���	|ł}\/���jjonk0�ёB^]��b^��r$jL��{>L�7����Қ���L�d�Z������e�j��Ǯ�;=܁�1� B�EY���������-͐�[%���"�d=�Y�`t=�R+��A!�F�}*�Q�ȰR�J!�;��	W��S�-�l�t�;gy�&]h­�G�����nᘆrE��J����Vf�nA�{M�!�S���� Q3��s�Œ�K�%Q�L�v��
j�x��b���x���l�Yi`�O�0X���L���4�k�
�¸��<�4�@�O4��+����u�Q�I:24��ǟ�^����+X5ID�\;Hj��}�.u��6/�z�τ�/_X��5�{����9�h�Z-�/ہ ME��f�05鰰� �r�}8Pat���`R��ݰw�� 	��3ל���߷'|��L���E&:��+�׏~�#;}����Gv�Zm�8�S�1�:��Z��9�
��:����8�i^���;Gs����ޏ_�ɋ����'��|jn�J<�N�MݸxU�dJS�^���;��G�R�3gu��5�)�ʁ+��%K�!�� �.����K���u��s�I���[�ľ�+����g&�����ku�ƛ6����J�@Q��
i�T�_~����w�:e���iػ�.�����u�����˺x�Lp=	����n���G�7�B�LT��M-�l�J���˺|���a,�}p�)��T\�$]�h���`ls��([.�����k={�ĻI��}O"�9��� �&5q���9��5��_���]��I ����C��[��Δ����/���A�N���'Փ*�M����>��w����ړ�[8I{�C�Ý�!,�`��v�@���6���I���M8�� ����c�IQ��z[���f[�qN�� �->�ǵ�*���O9�4_��5 ��Ҵ0�atv��)����"��R=ᡵ�������VVTZ�R8�\��p�}=�E��I� k�HX�t�$���VÂ��<�i�r��1��:9>�n<T�jkzF�f�:ᾮ�r��
=E߷���	��������l<Q����ˉF����7ٲ���ڒ��}����]t5���V4��VL��o�ii{O3�����j��}��X��\�Ƥ#!��:ܓ�	C����
c��UL=��ң���	�F >k9�M5ZĢ��������#*���4�)�Pcs[��n�.\��]���ₙ�t+[�k�À{���g}r�5l�1v�8���~�?& i�؁�>�|Ûl���ш;;=�W)�ܷ@��OA�=�&��$}ܣ�P��J�^���g�o��6�}�Q�Y��C�%$+�`|��xKo�D�>|�X��C�/��7�/���f�l�TV�\�󋉇�;��^����z1���?��N��ix�Qot��|ft|P�]H�6Nxa7�u���v��?��N�9�Z<�/_<ҋ���	GC�ƯP78/��qX�魀��{���hZ������|�?��?������W�~o��ϧ���J}��Ε���턿���9]�xQ�νf��V������(\!g�r��si�{.�o���+ᙅE��轷oz/A���+=z�@�ZC�Ν����!�F�;�h, $�{W�^���}��~��o��bc�X��-��T^'��ҋ'�������{Woݼ���.w�w+Z�Z׷/��〉���+�Z��S+���3�����K1e%e�H
�\o2�t�gisw_������}dx��ӗ/'�����^���{�dJ=�^����#�
�}�إ�gN��wnؗ�� :J<]�ǀ�����{���SW�S��#p{'�I �%:~�I����g������ǎY~`�)� ���|�>���;�0�� \���0�N^�aW�ק��>u8ɘ��Dv�L:5����h�iQ �q0�w��e��LF���5�m����\�t�.I�鹫ƒ�R�f��'<	S��b��?3>�.��i?���yJݐ$�7�k�_���
3z;�SkwiM��M�vJj��-޷AL�,�F�jӰY�̀pЎ�0��Al(�m��/��?�b������*Ѩix�W=}����@�	O94g�r��!���Z�tY���F���v��u��z���1ėL'���/tI}��O9RrqmK����]��������ӨPt$ p	�1�V��W���9���~%���W���P:eG,6�ޓBLt�� �7������^�+�B�栤1�,��i4S4$��k{qI;k��(��E������d*?�'������r��f.��)�p���EG[8��@|_@͎��yL�M|�	4��~������$G�~ќ��
�������{�H��Wb'���0�MUVeyo����tO���H-��(�A _J�A+,Az$ Wt���j��\ΐ��3=�1=m�My�U齋�p�ovK��~&Ѭ���̈��������%y0^��.������(�]�k:�^�6�٬pMG�o��^}��p�ӟ��{��H��s�;a�ؤ�>�W�k̓h�+�UB���d�5�=��W�y}�{�;����^H�eAՄ�y�m���m�Wh&'s:���6�|O��9ɟ=52"b�O������y<���N�l��!�~�׌�Au������G;a�'��G#�����7��G��"��o�����?_�ظl��n�XX���۟���Ϥ�d�(!i$��U-���ں|FE8���G<��E�����6V7�9�a||/��^�q��(��V�t��
GO���)Nvd&�v�zL;B��.��w�y���/���hf���:��?&���&k�V��ܙӸ|�<Ξ9yh��j6�`������6����p��F��BjpGG'098��?,�'ag"t���!�@�ü�>�p��m�����`d8��ح�M����`{wKf,D&�&u-�l�n ��EL'�;�΄�T|H��{zh�.#��2�0�Mt3S.�jie�#�C�'a���=~�����n�5���a�qA�$XdkU��l���<����l]A��R���D,8��7�[��bC-��剰��âc��M\�ދ[�qv�MT\�jKA��h�'Ο>� %Rp����߇א׏ё�>}R׏��m�C�6���h�O����{;�\�B�E�Z�N6c��(�fP�Ϫ�(U���al�pny��e1��ڼ$����t�ǘ�sJb�¥Ku ��,|v��p5j�Ej8��!S���DhP��Bvc�}���Q�UX�d4�)�� 	st(��Q�����~2�d*O�/5ʆ�C�dź������W��p7\���-�ִ��<pz�����D|t��4��i��X��A��j����t����O6��5Ԥ3��2�vKEX�[�K�I�5%%�]']'F�QLD�P��P��Eh����UK��:���pL���iڊMa���TJb�����Z�Y	Țr6�E��7��3Aݣ��Y�8��Y���\�ƹ&��g�o�~��'�X��<�X��/�j~����矢LRf�D:��1ם��r1�A�E����_�׿�5�?$^��ч��fS��&G�]�������43z�۹��q��Ӕ��0�g���m��Ȑ�"��	g\�h��v�@��;2��T�C�d�D��:����N�Ѐ���$[�ǎ��s���
��ob���3K��&}l�Ӥ5�U�9@���0@�z��ɪy��T 87���?{����ῼ���G���~�IG�_��W�>��˅�y|~����3r�p�4��v�*��!�5'a���Ćh?��+ais�T�-�9����
^�q�hD��O����nZ��Gt�p'Ș$�FMS����P�ȩ�;w��ϑ��Y�˫����`�fO�Ϙ9'0:<���05>n\�@�IM��Y�Jak��̿s�*��4��ܧ�#�ƥ�wrT����E1N���4`ҝQ�O�I:�����Aqo���2zhi=�NbtxLPha����5l�n�Afd4��7�3IF�
	��$I8�nFЊ�������k5�o�T:����olf�?y���d�#y��k�Hs8��Yl��hJ_Z�8�}�8�!�}���О�J��[2ٌ�=�4_/ah^C�s�j�ޒA ,N,���&Y��R$a����c��������A~dG�a���5��0	5���������&�p�!K��J,Y%�ƽ�P
�Qt�^dj�d��e���h��- �*:�����gqpQ:�l�Y��K�#��nC42���X�,�����bhp/���萚�g�������&N�L!EW�dL�t�&�ޔ��ag�n����6��8�]�5e�����y���pC_q�C_��7:��_:g�o�`~c�fe��n�N�jU�o�>�lN���GH�������$��0z?�7.մ�6p��v�u���.��IƢ���-y��L~vW�N�hǉp��ao��Ca� 1������x�Q�N.�I~o�T,&1�f�"~�I�j3HY��V;`�M��E��g[��w�3'��(���3�|T�٨Z������ه��-W7���պ >$n�Ax<7��>��ܻ-�n"Ud���aW�aaf������/⅛ωiMb�tY�y�y�m�s�\5pt��F��!�b�3�1�#�|��\�n�
m�f2�4��4$658z�mݗ���c�����F�/���G&�͆�:f�O�'rF�Ro�����5<�la���hCr98	�(m%k�:��w;��U��0�_�t��U��ht�w��W~��/����̣�������A7�<��/>������Χ�u�IL?F|!�N�"K�V(ckyE���&?°�p�Z��X�ޕ�o%�_x�h��A�K�̗�v\���ݒ������v-�*���m�mm`goO�?�0� �j4�F�&胃HD�J%1<��~�v��C���N%��F	K�]l׋�t�8�f�Gf�ݬGN*~x��PׁAo �Ǳ�1L��h��3	giiE{�p,��`Nw�jw�Qvy���<"�s��E�P��C���g����%S	�9s
��&N�4�32�F�F���<V\���3���8q�����X-��x�	��x�W�Ūi*�!i��d����[>�^�-J&�&V���2��-`S�{b��_![������)��iR���+E ��(� ��F��RI~��ϞW��?/�|A{�j�����#;~Tf�,�DH8��--acuM�����2�:�p1�+w�l<(O��#:�F�V�n!��BVp�n[�
:�2��"��:� �X�(�zC6�L�!�CxR>Җ>�]��� "
�zѴ!���1s�w�6�ٝ��uL��qlrc�	L	�⾙�����P,�tNOO!����Da#�X�%ܺ�����:Dc�TE�u��p��f����d��0f��F��Y'�ͦ���A;�J�H	Rd8�h:	G((�������)��b��Ă���N��ݢ��ՔL�S���-(�qqo	��J�����+��x�l����g���S�+\�ɻ�9Ò#�����	f�3o�˚0�+�����H�&���a!���ɜ���~�w��BAEV�'�&V��y�/�d뀠oz�����Ϫ�!�������~�[��H�T�T�W:Y�$UI��҉���щxL��*2�I�T`�t�E���N$��"*le7��C�Yύ��W2���7f5\':�K�"������Rn���b�8�J1nlN�$ ڃY�"��v�T�������lK�,�u�ib�u�I�#YT��j�SQ��|QEX)p>?<L�r a�g~2>����7���_z��;�~�����;7{n\���.\G<����y�9>����"�]��tj����~sac}US��'�'�K�e��܅��\����<%6۫/��P����EM���g�U��v1:/x���S�nnJ?\�4=v)�i�-r P�a�S1o	Ocɤ
!o�a�xL�/�>q�B�k�SG�[��Z�`�^�~���˃�q��,����gv!�q`���#�pjlG�#p�;�9�"]�U��Ѱ<���z����=���8�]م5K�]D�a�o��6%��z}D{�h4(x3��3�ޔn��Z-R�i9%� ��� �!6�lF��� ��Ϟ�ѓ9�{ʰ�I��Uo��c+�g��n�r:�*�b�q��fO	|չ[p���n4d�]I��%���o<4)�i��i�V�3nRMD�Q�;wF�H�`+�f��z1;}TL<���!>��ށ���CI=z'�ϊ)�B��,���ťÜf�H�·�$I�-��t�q�G��o�㰏��-�Ū��Q?(�����}%-3�ͮA:hɬC�-�T'ܑD�\xMN�]�i����q���C�9����L�����q8�����:v��1X�e<��;��`N�u�}ŘL$�_�����F�(h���krV��υJ؍�Ӂ|���Z�P!'D5�G��F��B��F�}�>è�<o�XX!!���z�>�ܱ��0�-d;��f�!*��e�^1�0��>��{����vZ�R����8�r��;qjt#q�29=+�vhK�c6O;{�Rn�p2��j��b��ň�;���`a���ܠLa��]�Q˱�P��p���/[н�bR*5-r*eAa�A)>(1��O��N��!_�Ŏ߃E��Q4*=���>�P�R�,�z3��~�+
Ԩ
�&�������B"���/�j,�6�Ja=J.;�&W�E��$1�)�����X�I�j� ��b5lp���
A�g"f�Z
�9���M92e�쵮�L��_W!fs�{��lp��:�70����JN.��u�1�E��涅o�����J9�Ea�Leh�p��]<���?z�o�����u���V_:E�e���x8w�~�	*�\=�qdd
��38�����9y���89{��#�R����/��r*���l���x��o���o"��`����Dr`>rd�k ��}d�������{��OLY������d^`�(^'��:��D��%D�Mq��qAx�D\>�$,[k�������-�j�9z���0N���IJ�u"�"����83y���8}���=~�ph �#i��S��������G���P�H�V1[B5[��E��i$cq�2��F��C"��'�� �9@�@��/����-�L,�FN�}N�Y�E�A3�3$�+/.����eɀ���ܠF&���,-�bnq^��'���%ԁ���$?Xkj��z`�S�&aY�Y��6Tg��r���t��[=ԫu�K5_63|������o���WW��{���`���!x�N���+����m�aae�hH�����Wp�'W���e�qtdS��$�Ɉ4Äϝ]��� 'ǐVG��������}:�Ѫ���A���J%4�A�FWa}��P꡸Jc��fQph�dҴ�+u��hA���d!�Щ�Q�gQ�g0>����(���cbd�HHicd���/�=��rdDV~�TNm![hw�Ћ��Bm/������|>�O�(�څn��6�-T�����I��������.��m&�ћ�#���8�o�^�:B&���k军�I�4QP�C��F�{W�ψ�����6�m6	2a��NѮqx0������&����"��s��)�,���'Y��bQ�Mڒ�Y^��t;Q�V�y���%��C���    IDAT8B���A���w��=0�|&hrA#"Y�����U���i8"�,΋���3Cs^�n�p��Bx��^O�c�T�/\�3���0�n�޳'p�E{t�dA��a�ّ H�Ib_��rC$2Ò(~N�v
�=���4�ύ��!
��7�˲õl{�$�%3 /@п>R�g�LY,"ۡ���/�U+	9"�Kr���ך�%"	��PZR�Z���&����nVe��p�P�Ѥ"�k�>�,�����V�Rf>�O`y*���?��o�K/�߽��S����������_�v�r�E�N,�-�������]��+�/b0�ă������R>���q�a�e
�<V.�[
�n2���ť�����/KC��a�OW��U��=z^M���sx�ͷp��Cao0���pt�M}Lmi�����ź˧"�.���>d��K/��^����ˉ�O?�A�*&�1�J'v	�I�jM�L	����;w�qqfg�u��_-���R	O>B0��kzt�f[�����\��wC1_D�PE�ƥ�1{�������瑩	��������DM��������m�Z(�xpy5#�&�ǁ������,�$�x]H�G�ռCޝ-Y���H��
�H�����JM?W�P�͇�?�:Av�F�k�eLRYQ�˽,a{³�bM� j`I�1L*��ٳ����jnܿ���9^�k$9�4J�Ν:+xm7���=�����������2Z�+����U��H[zdIf�6;[VD��`��Q$Ɔ��Pj5������M�5��	g�)͐��-1�ea��M8H&��g���M�4��l��e�-<l��8ba�E�F�\�+���D É�)̌�K^D�7�;�r�e����PC��E*b]:3�ZSA�"|���#�0Yh�JYK�R�n���V���L��wt��!�����`��e:ѢTm*62�Ix�5cO�C�Y����R�L���L�r��Ld�R��CE�W>��~US�Zy����<� G�
_��s�GqbzZ+�<pY�I����4��u%d1)I��Z.X|� Ԍ\���A��"����������3,b^����>G�o�}����R���TZ�!P�7�>�B�� 2��BzFI{�t^P1yL�3��ke�azdX��w?�����4=��L��L�|����#Q��t�0����)�*����,~
��a�[��j��]�i���oY|K�1o�Ԁ�ޚ�5��[v�*�4|�$N��IL���{���]�N�h
�*��FU��jE7DȢ�'=h�!�Z����D�z�	�p'\N�f�8�������������/��y��w�=����/��r~��#n�ח1��5J��X|!w �C�cx|������������X���
���k�Wl��|��M���;}!��K�XYZ�A�"<Es&��(���O~�;w`u}[wM�VC~���@�%Fe�t�?�9Ą�9{P��׿&��x,�"L��:���d�%t�������.�]ن<����(A��"��ҧ�fpbbR�Yute�p��=��>��'���sv����GOa}cU�q�P��(׵��$|db
�OnK�^fg�����ZV�R!��ka�ǭ^;�}(8�eHF�|� �'�E�#a����L�o�C��C:����&�s>�S�)�h�v��a�M�A��-��D��gXo4dr��8e*����DkL6$�.�he��tP��Uũ���Y��N��~y��
������O,��,����D�'�V�3���'gp��1\8uI!x|�|V�t��7�0'��HzV[p�$3��&���QO�#������a��p�) �1��J��dq��Ut�7l*��MF;�AYa�d�i�W��q�L��5j�	#��e�//�E�y���x'�M��Ԕ�XY��@(2�H >=���(^��p����E�{pz�3�nk���C�"����`=[�J��n~�#CLN�56�n<�.IN>�~N��QB����t�38�rb�AJ���h�(�r]�R�wʭr�r墊���t�4�s���q9�7�ˏ�Ӈt0
���~��$�x���;/�,�F<�O�>-2&�-~��;���^����o���؉��L&vǸ�qW�&���sx套��9��*WK
��C"� c�q��~���j�Nv���������L(���D��C�P���Rؘ)T��Ej(m�\:�5��9�`���m<�����a�rs��F�e�clM�&^+oyz|G��%W�~�	_,�"Y~ɏ^ς�vb!�u���lX�-�z6f�:\M)R�rϳ����V�K�4�K�F�4��CS2'pL�ynb���c������,���Wzm��n��4>"�Z��E�v�<�h�S�K�F�����nO��1�m4���������/�?�}���'�lm�f��"�����<��ZÓ�����wQ,�{$���vx�8��}	;�7�#{��Ns}uK%�����_j0�n>�kW���񻱼����y��c�*�nO�j�k�{�!��ck� NJX����3�t�Fc��E;I~�Q���aM�)��u��%��H�L�B�X������m�pY'@�-/��}��Ȧ��r۰���&�C��h<���}�ի�}��]��ff���wc7���8��AU<�:hT�9'��G$�C�]�ѣ�1�!�K6&�����c�,m�!Y�6��IÈnGהM�UN��g�+�WJ�R��g�ݐ�#.��Y�F�Ā�`x�W*r�bP8�Z,6��^�X	]�Q�MR�a|��Qɓ����I��n�`Bxh֚�+*:�CCx���x饗0}dϞ�?�)>��M�)�Q���ݰ_��$6N����S�C�c�;�51l���tE��i�3SQ�X$�H�O&Pj�5}�{�D7������TX�����wР޻XG�\E��z�6�,�l��h%&�sb��&0Js(�`R�c�aa�oM��.v����U�^�����0�L�a|tJ&X>16�$=���Gt����{_a$�QZ�H�j�~�n�d�E�nlby� �=�HX݁(|c��MO�5�B?U6p�,k_����|����#ᎇ:Q	2n�T�T�hMf�R�L��Ԍ9d&q�n�<���e'K�sJIb2�@6/�j���zC�9����Y\C~y]ֲ����x幛2S��̝''�@Ї��]������s�rz-�##z>ⱄ�ٚVJ���2�l�0=6�+.��}]�,��=z D���U����ڗr@`AeA���/M|F��5a�g2������2���ǥ�`��@Bzٽ�
��&�ѱ1�GF��?���U��6}N�q8H��U+�5�x�OJ�Xh�MDKPi�,ؗ�+�[�ėwX�/�6�砷��	����bO����&��ޞn�^�|�/�|]}s�Hma��$�������5�P�=�|n��xJkm��\��y��[ɕ$y$)�ׅ袲ȼv��Ǣ�����"����G�=����կ����ի��K/+�wso��ǻ��X��$��*�DN���m$��H�"<��)J���GjZ��N?�T���k�T�B>�-�����r&&'��r�1��6�߾�M�^RnP�nL�	k"q�l밤�
=L	��K"EȔ����rWC��iGf`�(�����c$u>����]3M��2�;}!w��B�%�jEjN����?@��!�=�׉��u<xp�KKJsi֛�a��(�J�6i����Ј��Jp��%�:u�C�ڟҬ#C��2s?�l(����DNTM��-9PjhP� bB�EvU�jU4Y�^l������)5s��
,N�wj�)Éx��&=nFF����wP�5e��?S!q��m�Re,}.E���պlk�~�up��,���Kbsr*|��>�{�=���4Ý�5��ȩ�zaI��A8��X*��㓈x|�ӊ�RQ-'y�K[H?_l"����W�*h4���)��ly��6��u�X4y NMO ���ˡƄ�|M�rNz�������6�|n�q+��F�b�r��i~�^?ߛ[.a,,��>ʅ'��F���022��x��3�9wѡ��x-a�|���%t�����M���h֙��~���LN��U�P�dޱ!��F�N�H2�ܣG���b��*�1��!��i)�t�FYL�e(Fk�HM��;uF�g���c�WM<�95���率'�0'�~���ȭn�wP¥�'��/^��-]+~�4� R�w��w��.���c?�����K������ur��p���e����<r�Ͼ���%9Z]^���b�i��-ޚ̬�_?�V6�,�������k/���'Oʰ���>��<F�Nn�R�#�%S�"=:&̃��X^_�>��5	�y� ��%T]=4<�"A��>�鍃�i`�Ŧ)��6�MV��SDd����灍��^eO��Y��u��l;䩘jl��Z����F��ߒ�h��Y`5H�{�������{>��m3r�`XD-}呓cdIU�Cȕ�7��Vn1�Y������+	�ٓ0�5k��$���"�����[O�������%hv��k�������G�k?�Á�#��i�8�6&%@��yc5mA�,����ev������;;s�hH��ӧs��SG�jq9;����g?���*e�ռhY^��P�bN6e��i����'3=^y����s��磏��񅂲{k����D�GQl��uPp�iy	K��ۃ�z2��B�/_���;	����pz*�G�O�K{�Y�O�bsc}�LV�4]�z�.�8ҩA�b	dPmV���� O(�Z*�Q�	F��6ִ/��$%������k�j���6x����,�^�>�"X\Y��DŢvx|"��U�"!u�$51=��/K��i��nZ�1CDPk��$�PJ�ǩ���iT�oK��!��w��#�I����񵗟W,e����'�}�[woI>DL��e�_�3��Cf)�ZE��BH��j㞶f�����H�!��fKR��nN���P��EX���{E��D\S�Z?�ޣ�n�B�R	B����\�6<b�tW$]ᤧ�	*nD$x s���+�|>�r�(ׯN�&�Db���G�G���K�p��)D�>d2�1��U�;=l/.���"�� �/�Z�䆦@�P�@�h�d��aG��K'�f���X�I����u�@���)h�Ag.�)6z��2�D��ڎ����\F0?O�:'f�98�y��&)҄��u�.�P��a��S��D�n<�
��꫸v�&���� q��^�ȅ�ݿV���ގ��3���ƍ�����'��k�j���^FE��j�B�������?���f��G�G���͎��2�,=}S���*���<��'ψ�E���d�(�9��9�%�%> �u|^����sR�Mv���2>'�cs�xݰO�At��_��AR$U2�Z_�;L�b̪�<��������Փ�َY�c�0�SQ�WV���>��w�L{4�pld��-8Z�zR���j��v��n���6�P�f_����6����$c�A�<5r|]]��(�ѦG�����B"$�z��#�����Oz�A|��|��=�����;��ɓ?�[Y��0�^�"bV"�>�������T�z�`��MR�K�� o�h�	�+����+S�ݭ�����
n\��ӌ�󸱱���%�E�85+	S�[�߽�x�{o�Rnʋ���6٣:S�B왽��vs�o��槉�`˄�K�)X�-�D��Ut�A�{���枆)!�9��X�EGk:��ɤH,��!ܾwc���E���~f~�s���(�$K�%��j-������Νq.w�d*.6&a��*���P�K=��m��n2|���h!gNd�W������H�����tP"��5��c`�����#'c^�s�[�o�"�����Qoij��A�'[�+(QQ�dPҨ>L� ڽ��N�bt+�����5�_�%ٛ��s�nݹ�[�o����:68(~ 'p��#k��~t�B�7��Vn���'�ImK�Lړ�7�!7Z<�/���m�Y��9�����!�~�G�k��D�kf��n�r�bܡ�ӕ���1Í�2N�#�ϖ�%	[�eb(���Q9����H9@�k�ׄ���Ňd:��N���s�=w
�XP�?�"��=��e��d�o���{O��ɣ����K��8�	�Cx�1��i��FR�f;١��r����k��[F"תյ/�N���-�ڨ�ܐF0{�+.��k��9�)�"LBV�֋^5U�0
�9�>^���&���bF��9�o��\9w^�==���O�8�@8 /����mq"�;�)�E�¥KJ�Qa�sM�X��ÙA$0��r�<��=��w�*��;~�,��*t[]��糉H��cqI\����Mѭ��ؽ��|P(�JU'2CC4fc|��������g�������Jș�S�4ӴC�N����=�ri�Ć�S;m#��*�e>³�M�U1�Ҧ�LSQ`�y 测���d�[�-[�dK�߹��Z?��2&��d!j�p������C�y�֤k������2��������)I,¹��٢V&2 �ҫdJ'.z�������D��?�����ߣ��G�+��ܹ3�x��=��|�;�kW���#� ��ǳg���PY����� M 1���=�-�'�/��w �+ �w ���7q��q�NL"�b{}]F�bNٰGgO�ۮ�'?z��wP�4�i����M`�u(���U}���k�S]^���I�3#�6a�$�)4Tzc[Q�{=�[e���UM�gǍq���M��k�p��YD�x����(h������ښ��z�o��������Q�ݞ��$Z�ԢLrJ�"[BI=�g�܅���}9�����Gg)���
�V�~�h�vKI���~(!6I�9w����
ʖ^2���4�����AF�U�lж��������Eo�zK^��r��L!Ȫ�u�m�O�����5��ۖ���e�b1L���[���^���c3�.����ǟ�|�&zO4�8mA�L�=����l���+��#rN�PC�^��N���'͵�v�6c� 1�%==���OބJp�B�"�6p���3���"zp�H�iv$Y"Y��ր�0�!h��a�;���o�dj�Ƅ��`@�d���E��p.#'�V��ωH,�T:��Gp��Q�M�*�����ԭ"�g�������]<|��B�z4��T���mӃp� ��L#�J!D�,	nb��2����Nm��|d�`�=�)e���kNt>��Z��&����+ݗ��9a�w�|� e�}r�J�CD���`��
�����c<>(��y��ϟG%���Ύ�3gO�`7�������V������`bjJ�F!��]$C�QڦRGr�r6zo��7�?��"�׃!�z��2>�a��R����=����^x�3�c3��۷���c�}���8���Z�v��#C"h� ��I���kk�v������������&�Y焸|Di
B,���w�-?�!l�PM��%[�e1�����ٿ��mdL�:B��������X��%��,�J��P�+=�����5��e�B��a1��wy/�M�דr�s8��������DN�M��?,钏!0���h$�����y�_��2�����.���j�\�x/����XDE,��ǽ����
�wvTN�Wm�Eng�U����d0���F���i';9<�!܁D�~�ll(Ԁ�N�x��G�]�$���M�-���|��.$9��~^EN"��a�M#�u:��&��Xt�e�T�����O�=M�2�~��F���̿Kj�ӭ)�ߋ�{�߉�.]��3�K���;?�7����sW�����������_��#���:J=�9Ш��nzY(f.^SB
"�R�k:l	�Ue`R��k	lv>o�AC>}&a�E��?L�+&���`@B:|UBٍ:�̎��	�q���8��A��BU&��#Y�-.}/    IDAT����O&�O{[�(zt��ĩ�@LR~F�G��0s����+86sã�ޥ��Ï?���O�C�.�#��F|hP������i����jE4�%8�M%1�(�!��݄G�����NLVy����BM8�� ��
�˹�����0ƇFD���{m�h���W�ڜ��#�.�Dq�W�tl`i�lx!G�V*4��X��P*��Dt��q a 9���a�ah4�x�C~���)��ۃ�O����R�er����4��iv���#�2������'=�t��3C����A��� [�ϼGx�s��Q	��l.''�B��@�F��	����A"<�D�DFY�}���B�P�t�ǽO�I�M�Ջ�𫯿��.���bw{[�Sl��q�x��p��}�2y�'i�K��PH�437�m�L{��`�����	��\�������c�Eoj>�$j��n���'@xS���G0�diui׮]Éc'��������w� D:�|�a䀔J$b?v�c*��P$���{?�YՌ��Љ��M�j�.��P,A��y��(r:s�[nO�:TLٚM��r��=9�8[��-�ѴL�PΟi�e&�@��4�o�y�M�q���/q����[d,����-�gl�����L`��0�v�RE{~������\��F/y�.�����/��������W��j��[#O?��ŝ�ߨ�{�|�"^�|�h}�~5k���@�Q5�F� �f�F-y���L�qH�7��@Ry���N\�.b�?��X_]�N���'f13{�v?���������^�\�	M� �{Ol_����� c,�,��;mOW~В����[>�PX�<�^�ߐ@�Bǝ����Y�-�4ӭ�9~/�W6���gq���������i�7��������%�ʡFQ]���mFm�S[{n�4��NS.��J#'����83���&i�O�'�\ل�����2���P��#�@�h<![��`���v���e��6�&��?~tF�u�^��斑��9�����Jt�^��mM��%����5�Ru�<�h����f���4^~�F�i$�t�
I�{��}|~��3��4J���Ht��
W!��X@�P�+����4Օ!HE$i-f��i�_�>�n-�[����q2��Z�l(s�D��3������9A���TP�9�^��ͫ`�!x�՚r�2D�D�h]H��ͥ��I8D��TR��GN��	��D�
_�}r����MM+�P��J�����W��JkM*��je���7�Df3@�id*L��'��0�dx��MԤׄ��D_�@��S݉�4������<�ˍ�V ���%���=���+L�=�j�7�*z��� &�&e�{�ӻ(�B�	�����W�(ݍ�0�������T���{o����jy����%0W���Icf�=�Aaj��R����_�=�S�"vq������ʺ��	�6��&�?��ikcS;��O�R&�����ÇD�l��?������* ����)���i�Ei����'�~��b�NC9荰�#c�pQ�F��"P�~��<����C�|</�B�I�&3���T)]ł��<�ڨ��lZI��kU�o~	��oň�g��"�����l�5-��>,�<�%���x��9��4#6iK{�>'�
�76ń6�i����lu{5ر��^rw:������{4>�o���WML�W��JE����������o3"����x��M�Hc���IbgE�=7�(�Fe������\ݮ���hOפ㸸�b �����rI�I�R�\���Y=>+x��?~��w�Q:���t���f
	�I&`�Fx�ӷ����p(�����~�,r�����{�u�ϸ�"���#����&�a�&�bOv!���C�҉s�p��%Meo���H�S82=�˗/"��`mc����xt��X���)�1&f"�sII*��йN��XU�������Ć�Ϯ�P(��#M�!1����\lǞ9�-�m:+�PdX]��6�NM<Hx���0�����L�y�$���0�HQ�Ζ��M��|��"�e3��Fk M;�IҐrEwbd�f�XA�9�ч��P�;;ړ�@G
�.xL1��!�u�hY�����ЪԐ�?"b�_ #��`�G'1�&w{O��Z��5!X.e<n�iY���t:e2B_mYR��o��.W�n0|�T�錶�-{��Ŧ�ð���HK`å�GB(�@$"=7�_l��0��>��[�X��fD�!$1��<pS�	�M��VK�ե�50�Q;?��>|b��uߐ�V��Ѭ3�DG�$)�'f��7R�`��\���x����f��6��2�XZ\��ֆ�qrTc���

Ӕ�`C�.u�� �����T��fs�l�|87{S�xr�	��w%��x�"~�[��sW�j��f2���;&�ڃ\o�߻�ŵ%�����l4��.���2M��ԑ�	L�09nG�&E���K��_���pʉ/�&��΁���O~!E�u����'ʦ`zbZ��hz�ӥ���g�� 2�r�

l<.Y���7|d'��b8�������ﭣ"81$�e�E�0��9��ueM�����Ğ&iς͉��_���f�k`���ʳ�.�bKsP����bn���}��gP��v�_&q�Lk��a�f�{����*΂�i>D¥<���զA�H�c�<����6d�kq}�lpz��'{�_�������������^5��_��+��=��z8��<[����N�y��%�v���x��`�<(�E(;��0��h\µL("�	3FX�/��K&(�a�4]X]Y���nN�SGg����g?Qns��"l�o�t�4X>�L��;h�;f/�縉P���n�FN��4+m�� �!�ɾ	�A2E>�V7'		���͟%�����{��5��z	�d���;2�?{��_���@��~��O0?�Tńא7�p�=lG 0�ǅ��&X�Z�h�$������.����x��q�%ذ�+���~�$��,eM�c�s*�p<�	8gSbv0$��u��Qv�NMk�����f$sb�U�G�5�W>�V�U�Y�eʬ�^��Y��'��i��U��iTj�3����p"�3�� ���m>Ԕ��sb-�˽��e\�N}�Z.��ujT�y�;=$#1��A�4m�@~��ϟ5����~��%�j��X�ݎ���#$�"�2��R*��T�]��[�I��p�\B�VL�c�p�-�-R� �0b'N�`i����{�k%�1�N����_N��z�~[Ey` &�V;�"h��=�5)|���4Dy���	�Q����ޛ�[�J���Ҟ��飘��Br|� ���l��\�.srJ����f3��$d��W��ww�4(Z�Kɡi��B�])�aؠ�Z�MLY{vzן8z��SXY�������׮����r����E��0,�\��v�6�->���:'Rj�y�)$;�A5�0FӘő�1�;yZ6���r'��g�����/�[���ӧ:�ǧ&q��M�LY���U�I�b�Y�rY�,��<��ZT���=9:%���(�͞���d�I�l����S�t�(��[ &ș�j��,l<ߘ.�)����~�&Pi%c�H~Q�M����V����0]���_�W�\HS�e�dG"��.���`+�\���ۺeZ�YgΗ_�a�������5�J�|1ڔ�6~�NZ�t3<���m�p�<���WO���?8~�dX~���T��^{�p�}���{�f�s��e|��s�ѕ��Ȗ��I2�?���v�E�J�N3�V[i�ܔͪ�N�
&��L1��<�6�WE��Eۑc3��9�=�{?����Ot ��E���,fv�����V��SJ���Ֆh��-S�j >���i�ϧ�$��;����K�|�h�da��eE���5q���E|x�n\���Sp}x��wv�q��5\8�X�>���R���؁��M��.5�A�<�F��su�KU�N��/�t�ѝ��'-����im_+�-"��LD��#!ԑd�dBM�7�An��h���,e
*_��<kdv�^�hb�v�KY��0eF2?/��M�-5�2��D=pO+uĭ�aDc"Ɖ�L.����ǀ7,N�!��;���a�M�� "�ZU��r6'�*�>ݧ�C�mٶ�hAd���Vޭ�Ma#g���0�Χ��n~�kT�5d��ni�m%�d���%��6�z]�sc������}+�M�OD�_O�Ә�9������؀pGL���Ť��d���Ɇ�׌ņ2�{�M��}��2�|��W*�t�Щsҗ%u��N����۔�dZUd�UTi��s/�a�M{�z����7T��Q6�&
>�
0ߟ�ljJ=��I�qRfW(���� ��)�����ਦ�����G�h׮_�o������﫡'7#2�������M=o6B�g��j�^���F"Q�o���plb�]���Db�g��B�s�V�@�{��<g�Ls���m���8v����D H�;�<�\�|���(�{kgG�8�RYlq~_��<@7���pdfF�p,�3#���d�,�l���^/ ��.�'�etfp��^�I��L�l8�]����BkPS�M�=,v$�ZE�.���ɢbg٩G�Hɛ�46Q�RkW���g��e�i��v��r�-ח׏�����ށ��H!U��r�������>f����p��Ɛ�S
G�������^�j������W*,,D?Y�����?��l��|�"^�v��U�hV�:0�'l0z���V4;H�exSБ���3RI@�>(�����	�� �҇` [k�_�G&�ő��8r|V���>��{���a�T��f����bTN�tx>��ԉ�%M��s�{�����!w�<h������jGI(�`n6,�2���VQ�7���@*�S�/��ː�~���ǫ/���gNj'�m7d0�/v�ܭkgm1�E��$���jE���Y���8S����o�~٤�&�#0M�d*�gvL�0p8���~��Șe�Mh��w;"�$<a������J����&�n�iŔ�~Ћ3b	Y�s
�V�7�8'r�Iʢ���u&�o9��0�h�2�����L%���e�IiJ"S!��C���|�	`1��)��Z�0�k���n82`)"�������^�=�,4N'�����s��"L� ~©Q�H��yOɺ�bs� �~�A tU����֨�[k��l�0栌������A�]2��sp��g�i-Of�G�2q5�bB{E,�
�ň�
#�������b��ҥ�	�=�/d��K4��`[�T,)v.�t�
���Yɣ@c!x�:���h�akmK���1`@��4��$L�ӸFԁ�����*"���w�jU8�I�����Q,Sg�G,���+��Ư|ׯ_Gv/+���,�l �����§����BlH�S/��~�&��I1��rd|/>C������{���5:�)������!ѓ1�l�I�"����
���͛*�$���x�tN*3�qP�KNU��������̴�|*2�ӳ'pi���b+���|�6��Z�`�UF������r8������"�q�нne�je�3�;�,H�#6g�Vߴ���H� ,v�ڷ�6�L�ӶI��R8�)[7�g��C�K�H�I�gz��:�t�J�����������π\!��s����!?�����c`���ŦQC���U���]G;����Gf��?�q���/��o~�"�����������³�j�X\8s/_���T
�jID��ՠiW��D�3�e�&A=o��)-��^6iv~��-ێ�O`bl;�ܾ��1{��;�����3|���%�glo ��ү��N!��)Ȧ=��|���W�� bѨ.(g��Vh6/�B���ü\v�hr��5됦�=�Z���~�����<a�);|(6�p��s��7~gf�!p�����P��Yz6��k�L�cb-9	�i��j�P(����,d�i�m�bl��[^�>����Q�N�/���[�����x3��9��=jux����)
ۇZ��l���J�n���九�0u�Y�$e&��$��V�^#��ϱ�".wO!c���<8=6��/��ˋ��m�����L,�~�ǅ�@L�/{ԩ7�8��C�S7p0�c��>N߄�d�iI4T��@42�BE�*T[A���Q������k�P�����r��f���&�Lx64W�u�ū`�=B����=(��l���=6�V*��0KN�;�N!�#�Nj�%���.' � Z����\��q�솇؎��L�twgK�;�k�H���1|Y��	�G�������uv��Li�eЮ7�jvԐ��sme�����$0Y�����~�����Q��!�dK�˨2��P��|�1z3�����eh�Fp��U��S��4���WX���1��W����\аt�V.!iꙩ��f�2��ׇ����c����nll�Ѭ	�'�f�}�̑dF�#>sZ�O�ّ�j<��[`<��~��m���"�W�F�rsh������X$�{��9l��#���3�^��RfO�D�T�]M�,.,�D����B[8԰9���8��xEd҄J��j"5)*�� �|�l�T�9�~�x�I�ڌ�f{�����8�pl��JR�Ό́��E�
��)?u�݋<��[R$�-jӹB��=��c~e���s9q<�a�o�ǜ���߼M�����Ix�tj��?���[۷��s����g�u�X���K�E�?8����>���W����4�cjt�x�5L�����f�k�=0/��I��k,�oa~~����>�d"�Ln��������BKOJ�4��1��=D��<Ŏ��,��s�,;�A���%X�9�<H� ��#�m�)Ά�y�	��c� �a�(��K�4!��l�h+ț�d3Z߱��l�I?�׾�M��~�N��@��g�RV)�]D��ecHhi��YŐR%�cdM�*��y��k�M�K[fKt8��!c�鉅���	�`����A�9��L�F�FG��	apNYސa���Y|6�=A�<L9�r�l��0w��7ޥ�֐(�2s���j����B�^I)�wa:��`p@S������xN��j��1bn ����$">c�μ�z����Ȇ1%�I ����`�N���{�8g�<*���"?��vG�~/�rۘP8:��{�C��>T��E�[��ښv~���
;`3����z���y�Ѹ��B�����zlH�����z�r�� !+��`�{��d1���E8cx0}(�c3$���N��SdT }�K%]WZ�*Ǚ�ݶ
�����D%?6]�N���a/��b㣚�y�6��2�'��p.�Q�m;�A��8Ő�J��f�r���n8�O�JGS�DD%�{;�C��F8�Ĺ+W���^åK���F�u"����_���ĳ�yd2��T8�Ӊ�hT����������b���(p��DK��׌���7��/�<�1��
B�D��N͎�ˇb	��9c�SAy���6�w�	�r�Q�A�@4�dl���� ��s�=��W�Hc�������m��n��m���(��)�	ߍ�6�ÖE%�+�	S#c8w�N=n�׽~i׉H��5�fiv�6"i�p9�	��*�.�m޷,�nQ�[k:$�����{{bd	��%)L��3���M�m����ʌߗN?�&�֢��b����]|�'?�����#|�H�{!b�v�&�(����m.4�tw������*�w����åg�M�P�;}�_��0���]�V������%9ɉ�4N�������4�n6�B�NSv�����g������=Y��=v~�{[x8��}�-l��"�#	6aY�TI�v��PY�����-�)y������u|�D�q"C��X]�����"�0�H:��Ԣ������w�q�g�]*�)�|D�Z    IDAT�����"�� ���*��ΝC<�C�R���<v2�����q�ZN U�[��	�RZ�GH�R-�˥�"��Q��)4,z��)A�S="�.0��F��+���$y͘�J#��W.�����\G�^��ؐ���G����3r]�0Y�4D��bf����A0�[[�(d��/@;�V $@ۿ�.��1@���'�}�ۿ���}AW"݅�H���r*c���VGS�������� )B�l���bKS��KWq��U$�)4�uxh�I�$���)e�?#&��'���!Vs�}h��Xg�ʒ�-��`aa+K�;��` f$"�DB1���k��=P��Y��Z���s���톟�����"g	��kS�8�
~��;2�V��C����	��9�#{��@#�?�sl����9�訊��ilHz� ��#G�T��$�Fu����7�����.�7�����}�=6'�ۂ%�q
�g��N&y;_��+6�^?Rl:�A9 I~�d^5S�rhQ����Kx��W��/��1�qbl��t�������`�'O�I���`����I��D>?�bA<e����iN�H��Zar��ȕY0(H����2�m�������P�Pc&��'+��!z�'��1:9s�������ԙ�O~�~��6�Pqt���a �C�1�E~�<?�`q"����k�0���|h���&1���I{���U4y�7o�}�##�3�Z��e�����X �XDB��Z�r��z��h��Ej�q�����ޖ߯�,p�K��n�Ír����-��;ocqk]*
N���?��Eפzy�j��<�Q���*�N�d�n��g'�O���I����ra���j���sx��ue�����G�������L(-����^���4���K��c�S`�i��2͘X�����Ul�HZp��e���t�)��w���k9u��@eWv���R��0�R��&>vXL��H�`'�cvj�jU�x�b�&�+;5veLᇢlW0)S<�i[:�h��!��8v��7'�@,"6��ֆ&an[n�x��+��y{���,;�����{S�uuWW�j7fgG�\��H?�E�W���%)	ZIDP i)��j֌�q�)����{���;��E�P�{(Twuefċ��{����k�	xqzr�O>���"�eu0����������7;W>�
v�մO{��>�ܮ�EB���-G*��$,�{1�Pk�=�b|tr$��lX�tw��}�v>���$��ch�������Ջ��.4\&	�S'W�q��e���z�!Y�D�r#�ZUH�-�lM&�K���p7���Q/V���C<���q5h4")��l���K�}�y݃
��z�ĠWzM0�"�B���&r��$�y��m��J�cYl��'c�җ�ń�
����t�=��i_L�S�h�3ٔ ���u���^�D��g�$!���v8�Z�Y}Vl^���y�b�?��<�;�:�70���lߧ���]�E���_�CNqbEӈ�bLa$��!M�eS���"%���E91�/S"�s��߅��A�z:��&I��pkGNj�vyO2J����O`��D����B*�J&g��LW��	CG�~�|�P#�&�fs��,�<ɛN&.\��o|��^���l&�]*u�L�����<�������#e�WVl�y�0.T�|��R!/��ӒA��]-a�PUs�r_���ѳ��t�g�yƝr�C��N��ռ,,�tub��f�,��m�Պ����^�u\�r�����O?|ۛ(:���hJJ��,])�9Y��܄�/*a������t�Db��}��.�
K+odJf�D��C�����"[�����"�Z\�(��L:�D�Wv����d��9�Z:�\ܲ�%�"(����&9�ю��A���1~��/�q��l��n�n��C�e�iC�iq�<#��Vq��F����&�華�I}�;��������V���d�����g��U���	���?T!��ux���!8��ˢ��"mp���bEW-�E�V�Y����XZ���i��c�:s�6?2�S�l��/~�c��o����&����\�a���@��aG�N����tx�x�ӕ�uS@l�*�4C�R�t��ִ�U�("4��en݀V��e��[�?�C��pif�{t��~�H)?�n�����w�곷�p�������Ճ�Ū�M��RU7;:c�	���pZJ��i7
o�{�sOD��x���-0�2��!� 9�p�(Ӡ�-�~uuY�?4�X���]6'd�f�y��/����������~�N��o�n�[�I��*�Q��w5������#�J�҂rK���W�\���)bEH+�t(�d����&�>���1��9P�T�?0�"|��5�
��<��W�b�l*:�����K��b�+X��u1�a�N��5A@V����Õ~���&`bf��I��]{���f���\!+��,�j��y�����:�eP¦�
b��L�P���C��	R�ԭV����T����a�=�G��j��KgT���x/�Y����3���Y50=5���HK7YSy�E�#6�G�+o򣃸���w��Ogdl�z�dJ���*�5�P/��������<nI�B��y���!��9��t�s��.L���7�����+z�D<��3�ךP����\�޼/��xس �Y����C�� �!Z6k��C��s�!�q�� ��zMӺ䃕�&7�L�Я��J���I�� "�v5�>؜-Q��)����>{���20�L1�O��o�.�wֵ"�3��E��M�����B�U�$�H���k�<}S���ǝ"q�J���f�҂i[nT�r��VmqAZ|�$!/I������NB�U�
���:�t�$8z�!���*�!�5 UJ%���w`��C#�x��[���X>�ŏ��{ۊ�%'�͔�<c�=.T9	�2���ӐS��v6:��q~l���嗒�x^a^ZP�q��:�"8:�c~�>��=�l�>��^��b
��DW�]��>�Si?#���UQ��p�H`��;G	���Mc���]Q�s	�~�.�wv�M�L�?�J>��nȶc'j%w��Vs�ɔC�Ƥqꪪ�(F�&ښѱ��=^��$@���	nuf&��J(�\�Ġ��B��r�b����~+�ϊ�E��3�K��&^�t�8��?�s�{pWō�51k4���0�[iT���|Aw"���@����i�e�RfJ�u���Ŏ�p�]����|�u���giZY]��ܜ)mmO]�<΢y|v�_,$���r�J�&�m����
x�_�5c����Ƈ��A�a���"4���A,��փY1EX�d��P��T��]c�]��~OW�����yQ�%�&g|���z��C�����ʹQ�h�8�����_Y�����xXj�.{P�L�E��h�GBٜ:�,L����Ԅ�`x�p����=+�}� �Y��m(�N&Ҵ=�
�pP�M$��c�ȃ�;�|:%])Mm!���>�P���T*�Y9�	�P#�T��*�&N�t`c澚��%�*@-~7�y�kl
t�*��`������ц�@/½�(ԫH�2��OO�H������UpX�����%ꃺ9Xy�Ke���Hʫ&I���ϭ=05�!�W��{{L�`�?6�������q��e�y�-<w�6���>��h2�ω����c��P�fDh�`�c�}xը
�.Ʀ���C�D�I�Ϝ����؂J*cM�f�#�ԨBZ֧j���s�fD�>ԝ5uDbx�=>�Ѩ�h�;���1B<��r����{����c~cU9��@@�,¼�[�M�br&�q{094�W���gdf���=�ݿ�)~iZ�� �1�yk��߱ȑ�7ꑰ/�{�(�7V�y��I�N���\��l�Vރ�Љk��C��?�+!���������&'���#��;?����Ւ,zyͨ aq'�� ��J�s�f�e B3��ь8=v�s�?��/}�E���M����������=��7�^��7�C7���c,,Ω3��e7��P� F��1�ݯ�7���H4�@�W�ff߹�����c%����p�����v��ţ�8:��Zh�<�ܔ?1s{Ɍ�B�fC'!����
�S��+[Mpb�Cl�Z�' �K50�7����"�Z��jł���&��o���m"�;d'	g����p/��"^�q� rg��ɏ�k�:�]�,+�]��y��O�qtr,� _��/��@{^_N�k+K�k�u�|��%ÊDP.s;F6���O;ѡ!��DºY9��on�@�����A�0��D"����nm�`��)��&���!V:��7�[3�]�������(#����c�#?�F]�eJ�(����ùZA�f�x[�E�R��T��ݽC$N���@�fG:[�g
���hu��IG9>6�3�|��	&��y���4]�)�ד-���m���d����I��'N����65�3���jt�^��q2%)kyiU��<\���3�Ta$Ȯ�nt186�+���M�-�<�RrWK�&#%��g7���aV��h��q��x�1ΰ�|Ap3�	���CMR����3!���&"��a��U�4��	��(��4�F*��@6?-�R��V6�8��!b�bYy�!NA���@���Ϗ�߇�ϧϗ��B���t��[��A(ځK�n��W����gdC�{�ި!�"����f3y?R
��Vj�>��L �>ֲ@lY��:���n96�\���)�$?�
�X�e�jɁS�t辒_qЯ�:�T��q��hgLI�
x(3$T�F�P4�]�GE����?���
����LƱ��~�f}E���?D.Ϝ��k�1=2�Z����M,>������0����Y�y���$o~�˨O�&���y��eoW��-�%��H^i�Ms`Ag������f?���*ZP���1B+-�d�T׭-Vn�)�C���s��ڰ�J��x+;��V�p����i��5�k���׭u���W�lښ!��Ϧ��������7:	/,,�?<���{O����t.|�������E�H&��d^E8�:����/փ��L�*^�]��;���1�WLߓ�8f�<��i����1::���S��q���0y���'89M0aC=�YZ���<���v)���p��\�r�j`k~��s0M�v���ֳ%�j�*�DAdI��"��v�MsS� ��$�LԄ��ݲ:�Gx��@Z�M�;�g�����zP�f���"~r�C�����7�.w���)��v�����%Ν7�`|dT,�{��ƃ{�4]�0s�u;첫䮜P�29	a��Bx8�H�@����+���K+kJt�u�<�;/9I6e~@����I����/��|�]<��!\ȗ����.��ٖjdB7���Aɯ�Ý}�X���y=|�!��Q�fP���7D�L>�|��@ ��W��C:_�I2�i��>�3�� ?��}���f��DZ,oN(DE舦ϝ��jKR�}v]��Z��RSדMR��'���i��)�U���K�����6�,.ca~^�H��&��ʲ`�}̩�	V�E�:����q?���0��z��?��ɩ��yB�D���n�}N
�<F�$�R+��Y�	R�n�ӂ���u�7�(,�z�%̆�ls���_�3\6��dy�I̟cw���*�,���$�%����i1��>����Y��:Y������d0A�TF"���֎v��X'.]���/��+׮�J?�2����ʎ����j��ҷv��$ʨ����ʮ%Q2��iݢhV�SX����*�o^;�S<E����h	3�U�e!K"iY�A_H;/_b~-��\"M�j�����Z���Y���Gx���t����c��V�JY� r�������iܸt	��hr��L�B�у{"c�%+߃&�f�X�6�y��[�;-�)��Vb��t�i���}֟�ĴB.x�����o�,?��݂�u?�lm�K���gA<5����R��{���I%ꥩ"�ˠ�X���̦e��W�ot4����7����)�4?p>���_ή/�W'�\�k�q��M�!R�4Vמ��?@��������^���b|x�<D�x}�rv��w"U�"�:�4�pq'T��Dq��%\�D$�"|������*]%����k�^\��/�|��������,�(ʠꕲ��i�L-���p�R#�X�!�������[q\b{� 0d��F�a!o2}k& �>�-%�>�A�D�j����� �فT��R�!W�ɩi���¥�ID�^�Sgx<��tR���$zb1�������VV�Tܹ{�M��K���B�����_���7q��+�t�b�6��-�s������[���cnvR8������GZ녥e��g?����Q��7���-o��)����ʘ�C4B[0�����熑���v���G��Q��^�+�e^E��yԭ���!�4�" 1��F�'�l�\�T%�^��w�l�I:���u�ʄXi`�)�.cA�l\�M�?l
Xp8	�,�PЁ�)E�V�`C�cRW�� r�j����`�	��'��סK%��x��A��K/alr1�^I������SF>�)�)X<�"��������مh[�D�Y.N,��JIbk�*P�$w:�[Zy��ץ���酻��)�b����YX�������	�uxt�
��7��	��G���ˆ|���L
gɴ&3}=�v�Zm�'l&`������X%�ׁ��k���,�^�0e��߸����ϔ�X��Q�G���k����ŗ_��J�>�J)��#E,�d,n�a�s���)	?O�j�m���_��eC����ҍ�VA�"�BҨ ��UD#��zU��4!V+"sr���-J��5�p�������ߍ6�4	b��*�?7������kH7*��,�Ӥ���W�͟G��t��Q<s��;0��)� 6<��g�׉��;�E�K����Z�g ��^|Q�X�B�������s���3@�|���'[S0է�+kuEf?af�ö�v�C��g �6��Fj�@�,�d*-S�#Z�d�4./j"N����p���� �8�N��H2W�^��m��,�D�(yl�{����������8�F'�?o6�~��/l���I:�y�^{�Y�'X������g��=����p�=Cw/�����=��pqW��\��t>-�탅�2���֎�W�K���B�����:>��Kn~o�=�Hl�r��U$���ؑf�����!!L��<d�6�h�ܹk<ȹ�6���(.+����C�����b���A��`e.���!ˁ*Ҁ���{��E�_`#�"|qfWƧ���O&���]�iڋ����R� �w���U$�LCj*olr�gT87�6D���}���\�|}�"N�Y���F��)���#���F	ހO_�?اf���Y���HS�E��@Hl�<�*u�?捝�礙|D�熇:��h6��t�k�
Q��2�I,�E����D��Wag�PF2�_+��]�8�C"�E��ό���pp�.������pQ�Ţ�f���1�pbldT�5�?��$�&=21����m�iH��V�������	IYgɄ�Ĥ��nW���#����/+��ׁ�.H��<��@P0�_חR�k��8�=�!�`H� �I&���s*̣TT�$��u�������ū(FNw�k��j�c&�i!7E�/�R�0������I�Wn'Jt$��%�8Bye�x##=;������%[�
|���BqK�BY^ D�ZE8�� ah�����A��#BY�&c���-5k.O 7�}w^{7o=�F�����F?m�ؑ�i X`�	`M�ʤ�� ®|ݚ�y_�Z��z")�FA�UD�شe�҆�Ns,�d��i�A��1� �RiАÐ:�^b�2��ȉ�ʮ�Ds��9E�lq\�./��
�V���G�t��d���(K����^b�U�����!ߋ#c�FO$�����_q    IDAT5-l���Ed&2��\˫����˦�$�Eg��s����l�lBY4�&�h12��牓���5"r���133#�!m`7ww���D�!��ޞ~=W,�DC��N�C:����������!V:�X,�G�r���0�3m���R�pm���&/|��|����Y�:�Qo6#N��3��|�N�-�������������8��~��ܸ�h  �!f�~�٧8��E1[Dg8�v�صŔ�JBL[[� �K]p��(5J
�fWtoa{�4�vS��^���.#$� ���5|~�k�Xu���N��54�e؋uT�cJ���������-�!�΍��<����.O܃(��N�EY1\|ht��l�4�R�J���H������0�Ȳ�!@��:w��6x;cp��a�y�6C�{��_�A��G!����{X]]�q|_�T���Ăm8�>��Ҋ�p/�E�"e��;95�T���M��
�`'��	���4�^�G�Ɋ��=YZTG<1=�����=�/.��>G"����e
H�®�2>�Fo_�&<B�
� ��i�6�hR��3�EZ�y�6v�,�������@���H=���:_M�Ţv��t���L
��9��/����
��^�`hj�9i�{��y��x?��Ʀ��<�������9r��j����_�MEX�2�O��D����)ߩ׵�$��ZN��lmnb}eUa�$D�o�x�y>�ڢr��rk�,[��}<p��5P��k�����x�8˦�*X]Ņ�	�7���w������4(�8:���U�Ǔi�gi0�R+}��{u�*%�
9�e���c"N�Dt:Pc
��h��`5����b�Ӝ���d�-�&>�&�h0�(�}�X���6rNBz��6�vp�8�J�ҥ���w~���*�e�QbD���V�A#H�jM�RVJNd&u����|o���n�R�
��R6f��W���iC;HT%a1Y�6e�:�h~�kkӤ�{QS8�Q='6ԩi���r��x���ټ�����el��qZ+�J6��n<�� �ܑ��M;�N�Μ[/czpQ�_���K�X��w��.cX��a�3�4��籷�+H��C�)uz�����iEI�ݻw���� �_l6� ��X�^�"w��5�������iT���5\Z]����ns,�,���]�U�"��,�1��U��=����ӕ<�=A��Q��3���o���~&�wx���=�P��s�g�$��D��?����w����|�E�����o����D�����x��MtG�����\�G}�����痦/�!���W�v.��mJ�*'��q�Lh��`�	���'܁.S$�I;�E������>�+X��c��������4�ӯ�.��������	�Y�l�(������eA7�F>W�������`i��=0���8I�|Y�ExdxP��V���s�d�ܨz\Ƞ�d��2�[2�k.���y�{B��2x��k��.��p�dB!	a�}���hﷇr������n>{.��Q�/~��t�CC�����O?�Cs��E�QeRY�V�/���W�cN�l$f.�`xtH�������2�g������u6s���{����ߍ��a�VIsH��rY$qp���`,u�<̂~��Cv�$9q
-��	��+��9����6�\�"�+����Y���͗��eK899E&���]�x(�!*���s�|���?�?���9P��I�H�J8�+Q���ZR
��v����"�֦����y ���p��L�L�[g����*��/��"�C�rh��r'�ɗA�&L�H$N�}�;;���Ws4�}qKR�&��[+��(~*��z0q�,M�kR4^�$D5��'g��֏��Ȉ��(0��Z��n��F{h4��|�VVf�%땺o"z��zp9�&D�J�j�+Z��H��b����n;�]HFoGlD���4Gh�5e)�\t���\G�(������=|�;ߓ���M���%Y���_�rS�Y�]#WA��6��$g4u)��~~-r�!�U�`-��9��>�����U}��+e3K�;�-$l"��г��U�\R��ۥ"̆�P-��׎���*��70�����	�+y�YfV�&D1�h���Y��D�׏������0:�AȖ�R:����alxD�z6h�bM%�����f��3����1��v�y>-����[ϩ	a�&4�F�����̿;35���5E2%b~��E죦��^sz�!T|X�����I��8��A���t��,�,ดE�V�^�j =.x&Ѳ�t�P�O7��n5-r.}�"N�_���?��F�/����~����?:L��Ь����2�����|��;H�&0�7������C�`�L!��g��p�ER"ugw_�=���ҕ:��(�]�!�xww����"��Ь�0�;���v�W1�ُ�U���ܣ���%����j�I?�����!I`�o�T�)W��y�׊0�bvĜ.Wɷ��;)���aBA?.]<������S�a�|���X��
v�i��(Y6���z�"����No�|
�~��U�}��/�^*c�{ �����d���ҫ���+�|������s|�ŗ8��;�ه�q~�.����g� �G����&��>�^��澁^5;{G��O~���]�h��Å��ۋ`$���
�wp �C������
���� |H73j�`�!���-���e���Y�f�JI;{|e?�D#�f�`�����HT�iJ���ȗ	�Q.U���Oѝ*#8�a�Li��i�֑�\	m�6\�xI��P'a���9���m�L�:&ֲ�3��Ǣ�=��ѐQIk�&Ӕ���ϸ 9��������Oh�X_���:�й�$l�����
 	��8�d��a�����X��]�����wj�y����4�or"W,�ׅ@0�����a��n���%WQ�w�t�V�OgQ�L�,'-=k�D�0(���s�2���Ҥ�.�j٘�	 ���s�uT���?,x���!�V�$��i��ۇ���{{�r����&lD�HB����Cln� ��`ll���o�o}�DR�U��_�2ￇ��x<7���M4�������^��H~���$-5y���B	��y�F�$M4=�yV��ӌ1H!����`o�z��AM�y96�~�'|�	�ͥkC(YNN�����U��1><�"���f�V�rz��Z%w%�/K\��ࢤ�RW���D\�	�ɛ�<c)����ds�s88:�/��BT�#�.�arB�|}������#����"$t�>|���M<��M5�{#o�07�#�I$����Q��z�h�͛75	�a]Y4^<�E�oB&Ldl3z��� ���'�ã#�$��'�y���WKs��
�$Ƕ���yi:�UO��:E�%�uY{Z��ɢN��C����O^���7^����?�����O�{Ȏ~���舴�qf}u	}�.��F�����F�TGaⲘ�GB����G�IF_=z���}�I����3����*��B��?���rv��Fz'�ӭC��`�>�Ņ9�����z18�#'��'Kr��Y}�YG�\C�1h4��䀻�O�����|��$ŰLd(.�}�Iѷ���K��Z_������=�{Qp;��Nb;}�,��/&G'q��%ܘ��NO�b����+�8����@���lAIA�l>o/^�D�Ī�p���;7-rw>����K����<��F�F�������Ç��Ĺi��廙��GGW���iRf�Kk��*����h׀���ޮ���
o:i�c [��w��Ed1k�#�ˋ��b&e+��	u�	֊�M'�L��eB!V�	�Xq�+9a�?�ry�O��f	g�d��`�-w_�"ҧi4�����������M�9a��}%Ř��
��4��%�N�,�ܥ��"I����ӛ�ʝ�JW1�l��%��*�,��e�@�-w�h� ������>/ҙ����.j��2�����������I�l���	��5l�X���Y$��G	�F�)�Y��?7P��`PM�`�����]��E�UF
sX-)�������bK�9:��S-�����niL�����5u+E�2��sI���N��OM���h��S>�,씼l� _,�677���C5�����˯��F�('1���PK|��G���O1��X*��z��A�#�|��\.��9�G��6}�U�iNC�K@c�x��uЏ�j;�@M�X8���.�6i��$�0��É��f^��T@eg$�5�������y=���x�*J����:�o,a1��x5�b��
a�r�h��Xӥ�PA3S �yj6\���T���+��,a{w�Rm�p��:�N���t#�I�p&+C��ǃ��NL�Mh@�B���ه����Ｄ�[�$�a/�m;��2b�ONNbu}MS/Wׯ_�u,���%<Y\Ԟ:�ˡ��:�5н�-?zF�r``;15���1��4�.�S�|��9��K�2��< �S�ߓ,6�;f���ZiN|&(�k�s�~9�3�������x�_�{�?�[[��d��ޛ�^A,F6�Ě&����;���8:�e!Ǯ�LJ���E�7�.(W(�4�ă�E<�9�A2xC��̳�u�:::ې)�`cw�C*�V�[�?�nw��K����1v7ֱ���;��W^R�e+F��S%J�:pt�B�~�N�:������P��]��K�΃��������ը�@��l,��}�;zp<�Q���Ӂ�ӎNv.;\� FFp��e\���Nwj�Qܿ������Z���.��
�

��m8��ӏ[Ͻ�חO'��q��9��>����5tww��g��a��x�l^����.�`y}��v�^*�2�Lp��%�b=����_�%�w���ڦM�CC�� �ݎho|�0|�6%߰VfW��F��X5�����]�Fb <p&`��U䪄���o�8>N�s�zWL���b����M��(��%�H�&QHM( ��!���O��gb��D�!��4��d�U�)�b�:��T���+8��f��'�S&���M�(O��]�Ѹ#�2��*�ZS,�_$ց��.J|ҩ�|�9qЖ�~�4�ozݚܡ������Ȁ'�@����Xm�*�6neu�ZXD)�C4�Gn��1�R�D,{�D5���P��P�=_��T3
&�I҄fW�g#��#B�MF��-�-�#~txc�����0�dkiY$�QO8����ĉ����k��>�F��zem��c��ҫx������;�s����T��P�O>��<@[�*�-�D+ч:\�AJX�{��ŸgC��;�iaLrb��Z�?z�D��N�y�d�i��������������Cp�vvt���4�U�X����Ң�(��t�E���&�m,a�t�F@]	d��Up�Nx�@�4���l�<�M'��ard�X���K��u�w"��4�F�PB�呔�Ŕ3�]=�ǅ�)��w��<�3�V��^�%Bv�٬��jjVB�t���ʲvݷn�¥+���"L����H�/���ɠD���5g����>�wwad|�c��"^O�����g��P���r�Ą�^7�~�U5;\���\����&v����t��?y��;�x���{���,���Y����7o�A{(�|!���E|��;�uFb��uk?L;4�8�	*�y9����K�^�ln
�>�Qw�$%x����B�V���2>��#�1@�Ql"P�!l�"w���aɣ#A|�508؇����m�wggc����n�(�,�<w�yd���Z��^+v���|��b͒yMȉo�v��,rү^����Q��'?�%�Ūχ����ύjȇ�ہb����\�p�&ϡ��5M�s����T"�f�"�/sr���>L����ū"*%�8=9D_O/z���W��\���6j�
&��1�?��'+�|��e����ܡ�d/�e�¹i\�x����i*��>x_y���pM���0�n\C�� �z�>�g�7MX��pI`k�٤�����AʝQ��E�;� ��d}r"�1
	&M�5V��U�	o���ë���qӲ5E�h�:��C"����\���-#w���~\Sg.�E��,f��}�9�k�=���a�YP4w�N�a&sJ��B;S;�ӱӊQE�V��
'Uv����{Mag��A�,�2�g���p��B��Z��B8C'���+��L����]��,|{���U)�Z��}5S���.���:�ى��>[Ѻ����BRLre,�4�������e�����\A�F�%t֘�����V���^PEZ��/�[փ�wN�-˧��\��&^˖������ө�T6L�	jwK)Z�"􀅎���7jM|���U�IEl��u��-O�F����p����ecN����,py]Y���dVz}���>P�I_bB��������\�I:�Y�>��{�`z! ����#��~����ڊX���>���� :zzQw8$�9N��Eb��=��F�D�Z=�Ã�'XI����5W |]���&j�J��p�ʘj�Í��_5~���ʢR�r�2ET�E4j��E���
ʉ��
������8�c2YYZ�Θ�K����6��KZ�M��ˆ���Pז�����kPz��Wp��E����K���c�	\ggjP3��x�J|�&I��C
3�����\�ب$�9|��.vsgH���q��r�v���Jj�tZ++a��'����TW����;��������~wnc����>��M���+��ɎNbok���'�:����kߦ�1�Kփҿ�i���e��y�X���p��!�+!_j��^��clr�j'������|�b���i�l�R���+�,ڣ!�t�?��~��)V�,b{w̚��s��K��x*���e��˚ x����^W1����ɳ3{hI7zڻ%�!!�7���z�q���PH�Ԍ��#[�!^+�YA�=�r�_��\?�g.#Bs�rk��x4��kˈ��|�1����3Wn�/֡��iK�w�b|p�|'�G*�{����T�N%_����I��h:Z7i�M��V�r:�ca��Me�X[_G�IB�C�E�����׃��Wq��-r�85��i�
5��rjp4�n��Y��V�������Q���Z�9�5�X�ym+�\H��^�;L���R��&V*��2Y�9��NS�>;L(��{�b6�)6�	���PF�m:l)�2��eȰ�Ӄ%g#y��? �D�B�D!�ю���ZrG�d'B��&�����*��DgZ+�Qe1���h��ށh{���������(���먖P�̖P���9��;���(�X��p��54���~��m�]�g�p��M"��7�ixS!��PZU�4�l��l�g���+��/��i����d6�{!�H�1V0���w�\k�࿲:4��Ԉu��Z����|@��ͦ�R���zm��;�9،�:;�̕M�{���+�bzzZ�&����n��ҫ�������gɉ�ߛ�AG{���|6+H��r�$Ս�����n�k:�>x������Δ��;�����ۜ�06����!W#��r�*FF���"���g��k��4�9��G�{�0}�d��:�	^/�Ο��W�[��x���'�{8�fQ�9Q ����s��}qmc˕��U�n��R�nL�`��O�����?~���2ur�t�L��	ȗ�����މ��1ܸxYߣ����Ɔ8+$]ݼ�ք�	9s��?8 �Q���w�,��n��)¯��._��旁-�|�
��S�c�X�pP�P�
:z���ۍ��q����w�ۏ�J
_,�a5q�c���\rz#�B��-Y��w�}�;P�L$���|ӎ����H{�������Ƌ�����������wx����[/+�d�����_�˖;���8j9qj`GM�"���`�&�<wt�Z���q2�T���u<�ҫ����>G�Q�$����w?yO��L��C��8M$�ߣA��I�=�0�x�6��vw���G��F�*�qx���Ɲ�    IDAT�qB�TGg'G��!3e�@Ns����oml>�Qa�:�.�`,� ��~���+��9���1ʮ��Ⱌ�f)�Zg�a �h�M_��.��B�Z���*�֖���TK�VL����ǹ�I�lN���!uql��#(��a{Gt~�xd�V/Tt�p2ag��Ր�5�[��yX0�.B��CJ}��v��hd9� 6@ɿq/�ۍK�����k*2�¼N#�b@�˩]�-AC�(���<��#��~�\����b�R�Ȍ�"��,4��And4�([��d�-�Ḋe!�����p~gy'*\�H�)�I�NW�	n�vv��}2<��G�4���HZ�bL���}�ji�	��P |Ń��0^IR�Sg�����5�-X]ߣP2��'�u�*��Qi�T��H	V'��׎];�u�RF�;s�S:]J[��z}�������-�����"��Z+��i���QJE���j�\Y��T���2�Xy�E�
��5kn�óS�J'-��4M��7�\+�$Y$>�>�uS�����&\���~��˥�-KUd@�#�.���RY~���"���gbb
}�ݒWr@"%�o Hƿ�8K�"����nT�c^,i:��&߀��,�,Ĝ��?�쳊�����_|�w~�s�N���yM8�	 l���/�e�o@��'~�8G��z�-�:���I[�����J�\�Bݦ���Y�^E�i������һN��������-a%���JU�h�<���̵�]��Sb6Q<?qF��H?�{���QhVt�R	�,��Hx��{�V���{��y\:w�&�dUk�׵�������sj|�2ط&a��ؠ����P@��%iA��o��n��}8�O?�D�$M�ϊ��dp�)�]E�r%br#��r������,֎qXʢ�u(���g#E�4�v�L's|p�k���S0ymv�磑����o�;k�x����ͭ-���Ó.�9	w2�Ex}o��/Q�f�m��������t!�E���a*�U7*�r��l���,��I��_�w��-LL��f�ci}?��?KȜ�L(����
��R�X��5�w��	ⷿ�-��>�<��G�J�́|����	��
z0B��C�,�1��J�����;ٖş�v)��eG����$�z:p����Ǐ�����_�E���2�Q���Vk�վ>y/^���P�j�+KX�^��;;vx�RAŀwL7a�ɉ��Y*&�˰���D�[���c$ɵT7!�d;�(��(��Iq�MP��b'k����C���*MITę
���Ego.^����u�pw�i��&��J�6��~Y��;�}����&���f��>߄TT�)��)�{>�-#�8�)衩I�]1m3�;��v��
��n,�k]Ab>w����>�BBW�L�h==�����dʩ�̼fʅ�d����D��I����ѼoZE�r	AH*�.���B�,ob�k$�J���$I���;���>��9Lb�6�����Y�rҥ�1#���!���E D���4�w4���92����"a�~�q˞�k�p���
*���駑+��l�bId-����
u�E-S
K��]�1��絑�(w�E��d:��al�Hnb�7�	'ϧP���&���6lTZ���x��� 
P�yS���B!̜?/r�řs�z*�4��s@4���KOp��#W�Osa��3��W�N�O�E*�j����ffp��U���}���"FRfÉ��ż�X8�m��ؐ��<c�Gi�¢x��-�Ǹ*��ޒg~"q&60�2����|6h�cpf
�ӓ��B����v���-�n�`�,.������p�00����&�ph
�Gp�gWF&1�b�x�P�l� �>I�\AÕ��i�[k��p�#Ԇ��nL���ʥ�z��ՠ<ian֤1g=��sA9�r�	�{͞�E��ͽ5	�\��|�U��}4��N=7Y�d��� �ˣbk��rh%��e�sSӘ���8�N/Nk3	�㠘F�mS�+"�<[�\�j���5H(��愻֤��󡎾��_����o������m,�w;��C7n���/�&8:�J`sm���'h��
Og�#\D�V%��Z?�T��d	��,8�88I�4����/��[o���f G	Kk���O�͝m��Ʊ�H�+��	9�lQ�F�nCoG���oct�O�>w�?���~�u������&�HH�D.f�R��J:�d"�wN����C�9���9tD�Tw�"f��,&]�h���	�G�l��wk/=�7�K�Ӹ}�2��b"�̮,`y��`N1o�4(�rU��`��r�|QBs���Nx��Ag�C)!n�8�&��'#�g���ܪZNI���3�HА�Q|�y:�}掄���̤�zN����f�>��O��ǩ��5� �A�7�>��ɒHj��a0J���M�<�rŜ:]�tz"�Xep�ɾeh�Ԭ��wƢ��do_����N��ds��P-�"JS
�t�b�e����r&$Y���<y(�SM�(6� ��YPfA%,�cljR��hg��V�����I?��L�78���ƏeV�i�߇E��B�lA�aʱ~]���M�s���p1M�4���;�pE�h���'b8�Z����'�GW��Uh)��i�'�|�jڿP#�^�ҍ,)�]��S����Ց�"����B��PE�-���*��t�$J����3�!0įFC��#�_NM6��j��"�Ѥ�w�L�7�^G����"��D{D�������a��L�tE+�u�YH�V96ɢ�;M�"���,Y�,������v��\�x�\��9GG�������nrlۛ[�jM����184��.�TԌ�""��ӕ�,���&"ݝ��r	�3S��'~x�#��|X;����*���4�(�k1q��
��&����;O��������+87<
�݅مGx8��rN;\��HRFR�����0D��hLŪ+ڎ�ϫ!&�`��,��H��>��Y�:�������%[�����k�z����[��ءm%]ٲē��=9B��ݶ�P N��T��012���Q̌O���!]+��Y,��T��^;*,�D�,�D�UlV
\����#�/��8�pi�����7���7^�����������ag/>B���[��#�:���2~��O�Q@_g&G&��J�e�R�"W|*�`'��EN2�<���0�����3���Zǋ/������c��$J�46�W��cvq;{�5��ZL����,�t���g��+����n>sM{گ�����u��y�ad�5lƏ��˜[	*,P�&JL0a7Dc�~��4mǵ�Wqvr���M�ڂp{]���B�P?�����������D6O{��n ��=7\�=C8?<��f.	�g�[]���&��g�%�Hr	o(B��y؊e��Uml"�{��iJ�B�yN�*wu�*�N�f"%�Ž�1v�Mr��QNb�@ZlNx� �<g��x������\MML��+��QWJS���[�'_x��CÛ\+>l��%ƀ��5�l)��2oYו��Cs�bQ$f���eu΄�85�x��X$�1:��>�(��(�F�T@�#��"ma��S/J��$C�-�N�S+I��;�S+]��X��xЪ�`���-Å��qt����@HB��!��}'��;�.�������U�{���y�g�ɔ�
<�l$���SM��sE�qjcB��g�H��x࡙�� ��F�
���&1�+��n�N:PJ�9�� �8�%!���Rמ����BANNz��[�x>;DZ(�i84��mK_dI�Z��;����ӠO��	ggBv�
�7�x`��E`�:?#�T\#�d����M�l��K���n|�\�O͆�Y
�|V�H��q8�[x�����|�wq�I�#�1}�i���g,&��ɉ	�~�7��͟�a��8=����J �͉�39>���ɀ��w�>G����Y�ؔ��YN�lθ�~��=���uc`r�Ã�B��PgL�8���-����q�⁊M�T5{ˠ��t��ز%��t��W���g/^�y{��=<~� �B$-ݥ�n��	錚V"[\�q�䢯��!����o��W$��l�����V��")�;D�TZZՠP|x���/>�T#�+ S* �0�8TpC^ =׉ �d;�ы��A�/�T���f�r���Be�I�����'%{i8����<��oBEO0_��,�gc������ML��򋏾������GcW�\��WE=��2X_[�O�CM�Թ��F{0"M/w�,�YU�y�2���T>`����N�&��+��[��f�M������>������������%B��
��+X���n;��z�V�S���*<$\>�e8H��8uf���I�ౠ����9v���rDb{WN�C<���1ɮlo���5F�\%��h�$`)ӎ�p�L�ǋ��(Bm���%<�\�v∫4= ��\~/*��/NA�� �G����S%�p''X�la3��7�=	h����rY��6�Lv�,��� �\S�Kbw&ͰfQ��r�t�{|~M �R~p��Ɵ����)�P�J=!j@�i���#MH2>�W���h���#[ȉt$G*�	�H�)���A�p	N��sZ/򰒑'Z���gy�'3rZ�5�����PnM´�k#

*�tE�0a6��XGZ�?�@���D����Dɑ�ý0{�\��B��Ⱥ��Q���J�r&!�md4>`�>:�N�GX�C�_���i�hs�I��w�$9�e8��.S؝f����or�CCp}ڹsb��)�a�C(��H�c	���IG�4!r�2IY4�!�	�9��M�-�2��Q���C���B����E�B�6�l:ihB?6Xd�Ҫ�f���9*���`��
�s�dFh��M�혮{�T�Ťx�g5	���ё�:T��v�_YYR����
����B�����h�N�X�$�`�xY@6���o�տ�A>55"�'�8�wv�����q�T����!�Ã=M���^{�u�=�wv�������ٛ��T��i'"@�6�rN�
r�Mg���m<XZP����(9(Н��2M>m:qա�o��`Á�h�z�e�r�9�'��>���Kd�C����^7.v��ZҐ�\b�����crNhq,kVr(c�o�C��!D�*勄^����阤?�K���RQ֨�o�P�E���I�i71����v�[/ML+4"]+��'sXN�㰐F��@ى�E�����]�B^�"̐_Ӯ"uz?�����"�����l���;{GcL�>s	�]]�W
�X_�/~��ꆆ�{156��?��%�?m�X��v��f2��}q���ul%?ˀ��Wo}�MLLr/����*~����h~�'�#2z�TBBN����vU��V���	�����M6Wӗ޵���e7��h����!�E�ҋ�7b�R�ѡ��	8�ҁſ˩^׺�ch'J�/�=n��Ş@v~M+� ����9ܚ����v�؈�b/q,h�Dݨt�)���v���I���N����P.@wjyA]�Ĩ�kTjbt�iy��C1{���ͼ�y��k��(T+���!'��/�������/sZ0�cS��a�\��(�����Ø:@Z�yi�����")�)U�-d%+��bϲ 2��]4���3s9�sY}��jn��E�GR�ۭC�v�,����(p�/�$"'���;i&����t��!~���c1�ӗ�:*U万*��F~��C��������>���2v�*�#����H�%C�S�af@=5�ĩ�0''Bvd�sZ׳D�D���6;JyDʷ���j[٬��Xh��ً�����i��1B�8~��`%)e��
S�h�X�c�p:�D5�MV4�j����Ô���ԗ�S�eB�[&"�RQ�*�.l�x=�w�Uh�*�������2��+�N�A�/��X_/�?�l���$�f�泷p��5D\>��o�����K^__�.uk�:I��$,iAr�=���;0�g�W��e���$9���տVc�b�I���@�_G6ql�)ա_2�N������{���W��-qr���y���s9u�D�R���\6N�W�/![N�w��Q���˛k���]��G��I�j�Ip�1ֵ"�j�9}�\��C1|�Λ���o `w����w?x�TB
�Ǆ���X�{�rC�F+c��I�ju�R�	�Ŭ@�8��0��Z��&�4����?7�P7ɠ>��PG��.8C~��h�l7�o~?rc���މ��1�h��2�,�M�R�<%�i��&�n�"x�򬠹I�8!F4�#'������ݿ�������X�����w�'��t���Q��w��1�������#*�8!�k�ȡ�ʎ�N8��$�q��Y�R���������Y��X�x����_bucgI
�=�����N�7w�,N̄�����EL��v�n���"w�ԅ�A����ÜP!�_���JG�����`H��R^��Jp��x;1�Y;}x����p*�(���OE�?szr
�F�e���iC�VA�Y64aZ��GpWG�P7�ݭ@u����M�PLg���	[�k����Q-���RL�!��\/I�K9�ث|�Ƞ��88��)��k��ØA0l>?�Y�H�\2	5�e����=&���Kh0�����N��1�|���(��L��B��B�t�x��͞���a&�*��� ?7_^{��i�Ű�!��$x��mM�,l����L�}�����"LD�60���(�f�M�&~�,J���ǌb6V��.�ptx(���^SRO[G�}��z� ��Ct��k8��W��9�a��ke]�2��/T(_?CM���՛z}<`Zd[��_��ܴ����=v�"���p�xd%��mB��P�ņ�Rd&kY��Dg�Ts9بæ4�E�%�
�U�n��_r4gSf��!�t�ǩ6d�_�|�)��H0ҦF��"�gL����ִ�Øv���ˁT�LɁ�ņ��7���~xۂ8cRR��@[D��[Ͽ�g._��\W��eC��o�W��y~�3��� HЀ�Y,�U�]]�mu�Z�R�W3���؇����y����y��5��V�j���Ѷ�-�N#u�7,=	�$@x���l���^w^F�PB�.��y�9�s3��}���y<�/4���H:�"���V �I	c�����q�؆{��������Y{3O��,����"�*���T�P �ty�/~�Kvj����RE�~��-}Of/��X�*�VB�.�&�!��׾f���%�G���{�΅d`_ /��Z��Ԝ����^9���zے��M���_����b�`���g?���'���f�rQ##�rug�KDw���nb�YW%k$&c���!R�S���:)�I87����;g��߯4j�?>.�> l}C�����������l�@g�̄&�GeD�r������=�l[��f�0�������������@�c��P+W�������o�����]z�������,�M�8q�^y�6�۫ L;��~�e@G�l��qK�ڌ�&`(��\\́�A�pmٮ�߳՝����,Wl�k_��ұ��	7l����������~^6|�;����IB�^��[��d���
���K7��||�,�O��7�xH���D��o�@��BQ�p�Z,Hf�/�j~�E1�E'u�����P��
��X�2��y��ٴ4�	C��ѸE��h-�N�U�?�sI�1Wp���ħ�Q���F1��D!6KAw>+Y��%N%
�A"s,���M�)x�n�������B�$b�/��f�õ�.�f�R1�w���atg�W��i�[&�w�#�Y岲n� 6��5$,[�6I�Pr�J٬�����gN���8:���: �P�� !�i]�)GC����k��YϘ�!yE��8AJ�D-��	�T̃9�_x�E��I���	�@�&]�x�1���S�������4�go�tR��{
����r���gIB PD��&�w	�əˮ�} ��CZ;�cT    IDAT=:iǟ~ʆ�S�=i4��oTX�xf�u���`�`�i��mQ%�VEnb@v��=�03`�DI����	�$x��V-�x��9>-�~�YEp��C%V��yNz�ՒHiV���鴒j�!����A�i����\�]B���Ϝ�N�)�����h�������]{�������4?�*���m�JEs���!̈́��_y���
�������)����v/jmR��^eёAȂ�1���O����e8P�T�ڍv��%����`�N&53�Ym�mko[�er�}������⑘ݺ��x����g���f	k�BVA_ɱ㿋Ϗ�;��Zv|�}��_����Y�@�y{o[hd�}?@���p��<����|�e��=�� �� �DϳF�*P���v��������[	����a�FF�4�����U����~�PR�0�n���S/����\z`˹]k�#Rs���Di�s�w�k�Z� 0��$�C�O������o��ԁYz��׮�����V�	¯=���X���l%bT�F��ء�R$��=��H��ا�5�\su�n���Z&gۙ�e�u{��/�׿�u;<9a�P�V�tpb~����ޮ>��j�u�;�-���R�a�SE��Yg,�����0\B ��] �����LX�]\1d�|���L���Z�����?$��F�W* 'ڙ�0q�v���u����q<���,&!�i�km�rQc4��p�p��6���Cu�Y���84� ԙ����ʖ�����T�jǻT+��kO�]p�n��o[[�7}P�j[m8��jqB	�6qH3?u�5#cXg��8t���d^[}�6�K`���NR�O�H��qhUr���9'�pM�|�UU��&0#�P}�ݷ썿��ݾ=�k�K����q����۲�S�3�Դj�h	|T�8 Q}sRWk�e�I�[��g�U�|������=[�p-i�qLh����8��O%8�wo�V�}���
4��[VAh!�(�5��W��˭3��Mݨ;7�!�I��>m�Ϝ�xO���H����1n �(����� ��6�9�܄�V([%W�8\o� �@|BSc(�/�N�y�x�&�L�E�d�f�1���)��������+U[͚T�|�B|�-i:8� ��ez��*nT��I�>������G�J&	���׷��V�n*�>���ҽ�N>ٝ�0T�h�ҷ��=������,����9�[���4c#�
��6����^@�x��	�!�P�����ٰtO��և���Z����_y�^������ݵ�>|�~��O-Ӭ��c
6X��<�"�$J�,$��d��}�˯ۗ_~Œ��fs\Vjeʹ�վU�aΝ���q����Q���^�!��Ru�����t<І/9�D��Ѩ��
Ѱ���C�f�C��u�+X�wzy�r���6�yn��v��]��8oŬ5QO� ?K7%&Zg�J��x�0A�=�J"Z��v���у��{_��[�z�/��ꥻ7wnqy����}�3���I�Z���w��~���X�#ԡ�5��ߩ�#�����pP������9[�ٷ�s�������v��!������l��ڥ��X>W��'O���D��aPk��rJ4x:\�|<�1*b� ���[��4��!3V0�?�Z��R&�"�@�"�!�K�^�+��5ᤪ��@��;���d���.�d)x����jMHZ99�1���<��D;�%�mP���%�1m�p#`��,�>�Z�������g�`'��@���ґ>���Ă�:Mu�,�N
!�-!�B�yF �=ҡ��%��)��� ��}�_���u��Z�O�#�������Z&g�lN�B�q���N^~����o~�NM�x��|�g��o�쭛���K@��i1� ��>&���*U�� �J����4�5!�^<{����x��=�/Q�IG�s��8(`b�����nY��f�ם�9sCGh�SU�9�[�<ZR���P_�>#����hWSeT��Jm�!��A;��3v�̌�	(&�/���*~��%�Y��;�Tp�a�r՚t2yiSS�8F �f��OӒl�fi��.�tmY��B���=>% ���y�={W`7Y�0�!�@��|�It?�t� ��<vLr����P0���I%��W_�ހ���t���o���as��R7C&��K�t��yu�w�L��ތcz���~I	������o
�nY(���YAPv�`A	�FH�����\b���w�֜"�nF�K2����a��TwZA���Y͜�}����+�}I'��{�����w�PnE"�@�E�&/��!uU��;-h���/~EA�`��bpA�ټ;���z���Y�磂G���+~$C��~�����fvNv��x�}t���a��GE}�3�W��!�CN]����(h4���>?�`̈́ז,�k[,$n1E�$O)f���,�5,G%\oi=$bkWꖶ�����{_���O=���}�򝛿{���	*��~�&�[�U���N������>zL�`�8�BG����0͢�}.�lj&���g[ْ�jf�����W�ԉ)��Z����~�W�J��ɗ����9sV�wUU�}�ȃl�e'�G���D�1` ���k��d�	����8�
P�Z�����72�Fk���T^�!�bӡ[T/���*B�ZT���l�0߯���Ʋ-gw,����� K�O��kB��y.*5�hc0_����r� ��@��ׄ���C(7���VsY�>�;����yU��2f�1_��?t�t�#�Ñ��{���v��.C�v��)�#�e*o*\�����Ύ��@~��Z�����cD`9c�p�����B̃���lsc�^{���׾.IA2m�7������[v��=6Z��}��5
��� $N�u�?S�,�B�	Zyl�@Kh^��#l!��c`M�ø��R�tg��1)��n�*'��9���a�`� ߑ�A�o6���������<dk�붛��^.+A	�X֟�Z_�J۱3�������a\���m�ú�  Q���ܴͭ����]�m*QNX9|��+�"W�J�PQ	�:�+��4ZjK��4sGT���I��j���J7~jzZ^�T�w��)��c U.�`K@�J�9�f bO��\��`|Be4<0h/��j�����oh`��	��G}h�_�Ю\���θ�
�D_�3u���.��D����L���C>�V>_����{֍��I�gJ�QCf4�}��E{��9�	�PI�zzm���~�e��$�x�k��_�����ܜ}p���Ϳ��zY� �<r`����E��*4A�.�|��/�f_x�e�t1y*ʚ��S�Ӌ���]�~�Em���4�?��ǿ;�w�ꄠ���y���	��n���*�GE���$��
��-v��Se�W|ڥ V��dZw8oזl��{̭'kd�g�@_��7a%���jK�w�����~�;N�����/�������z����{�h�$T��>���cᶭ,/�_~�/$[9>8dgO����N�� Q%ж�2Ug�ɡ
E��ڢ]��oK�{�_�Z�ܲ�_���gO��h�iK�쯿�=�3{�bє}����le|d�,h��`Zr��������H	Z��VH,}l ���^p��Dq��Ǩi�j�H0������\��5) �dӏ��VK�b,� ph.�n�G�l~oݶ+N�G!ւ�B���!q#��3
�-	��8R�v�-��m��m+m攽%��m�z-���'�!x�UA�K:�]&�22p����c�ܰN1z���+�
C:��w�jMGܦ X�(p��!�����E����e�`�,�p^�♇�����Oqk��9 k�\-�5�K|�s/���{�Wu}�̞��?�;�n�r o�͉�_ɘ�WT��Q��uC�\q�1]�x�O �3��̮�}O_�*Ԁ����Z�T̡04����3뢣���Ea<� #�L�Z�{�>�.-�yp��9w��^|�����[Z�;swlcc�Q���,���1IL<nc�����q;~괍O��.�Ҽ�ԇ�y�n�n)��_�/ܱ@�S�1����-�+��t )˺��DL뙟ת.Y 
��K���)�����Sglj���&l��]	��"��x ������- k�D;V��0C�޹�hf�k`j���^��gft�"�jt<"<�w�{��x�-�t���7�-�g,��BHF��U'�vx�:��D�&?qCx�
�g��r�7oж�4�wT5�#YY�q#�� N�C�~t/��0)�����TŌ��7��u��k�i=?x�h�]�h�w?��j�Z���p�NO�ׅ������\ޞ;^̿��U��V�ͥݟR�Ut�)�:1��Z�P��w���.H.$�����tgB!��0�0$e�s���J���H�G�����m�T�Ę`ׁ+�p�e;��;[e� �:_Yߜ����.�k2ޗKm~&���"����?x��?�����?w�.�����k����ʌ�Y/|^B�X��w6�G?����)?u�>0)�d�C�h��fMU��}ͺ�_\���nٕ{wlu/o�r��2e;s���9*�x�i�ˋ�W����;o�`¾�_�D������j��=A��� `����)�T���*����F�Æ�[#2!W[��c���H,���!͡�D@�G�p�.�AQ�(�� �e<���/�����1�*�2IF�W콻��a~G�y*Ḩ9h��֩(Ua�GGY�=�	Ph�j_*6*{�[\����ś!��Z$��1j��3+ּ�-d7ǎ����i	�Y3-�F�v����= $B���RD#�f��2$��f7��ZiG�ʥC�����h��y�MKPl70��,�4�->�9��LA�<m� �RMN68�0��«��9��l�O�S[]^�̉�"\Z�t ����z�"$��A��MpH�v&���q�����$��2X�z��G2�H�(��t\F�|���٨����� $TqT��x�]0sdf�AXn.���^�<������L/޸l�~𾭬�*��dCk��E1�{mt���:3c��A����b������@6��zM�LX 82�L��Zy?g�\���u\�!&p��o�(��.K},��d_	�r86����kǎ����Ӗ�첥�U�;7o�����G�-�j��3)YS�ϻYI1�T�u)�7K�HZg,eӇ������˥#����˲�%�j��w>x��z�m	�E`�i�p^ϴ��ԭK��U%Mt�|�o$c�Qr@�3na?�O�k�L���1�3�1�=�o����hع�9^?��u��A��bQ�;��׾� �z]Z^E���7
:����p(�x�ɉiH5d0�(Ul���Ɔ�l��ϒ��L"�(Vu-0å3��\���t$? ?/��$��LQ�{��R��Q�c�
ߝ��ءS���!a�q�P�U�;��_ݫz~��Wr�k=q��|�JH�Vs�_�(w�*ш�^�YN��Z�[Π(6��� �g��9���?���t����Z�o��wV)$<q��1K�:��3xg.����rs����;vg��kVn�l?W�S'g���<oSG'-�������S�w��a���_�gv��sʊ�H&�ֵ��()�B�v���5�
C�G�<QC�W-f����c�;ަC���/F�W�l��Ӈ�Y��P���wՎ����%e��
L�R��
�}o��2���~�,틯�֍K���m9����������d� ��z�(����jy[@���e�.�[}+gi�X:W�꜅���T�\> �J�-hF�\�_�:��R��kCG<�A�*��pH�Fy���D�/W�1^��4 `c�M��I� �����g�В�A�@M�۬6ĝ�uhR�\@`uS
G�9d�F�b�^�ݭm��Q)b5�sN/���S��-���<F�������JK���҂�o�8��,��	�T�PQ�� �!���N�/��K�5ь��f��h4p� �,(��Y:-��g����]��ao����,ïm\��L?��4����\��M*��T��`NM2K�o&�>&xz�^��Zqg�j���5̓Q�b���	\|O��܋�
�� U?�F���ѩi���Pe������x'��jr�Z�1� �%f�$�$5	ǜ�C�'�h3(vo��Dr'Z[^�5�b�<�|�}��E�t���c� �k2�U j;�	�u*2�t�p�b7��W���Rg�p�;^<���`$ V�O"f��"Rѫ�CACE�9X�c�v]X�>��N������BJ4.\�b�7m�弅RI'��@�/�'�)]�m��

XP���"�b$`-3\�sb�����FV����&*�{�o%��㽶�F���H��J�a�vC"3�Ξ��@e$3����_�%�$���`j�x��]�VC2�/��uG;dO�A�]��I)E�n\4$'��P�����o����}�S������O_�u�����cE%L��CV*f��ޱJ1/�сa�T�/fpN���) +E[\[��+K6��l����!E���3��s�m�Фu�h�l���?��nZ$����߶��3q�s���O��G�U�B��A�ꊮE@��D=�.-���n��Sq�}%��{�#�B$���	�~L�p�M��v�m��C���V����ԏx��#�:@Eb[)����h�';l`h����-��W?����Q��ʢF��T�U�Z(\���τ��P�̦�;�y�f���������l�����o�*C�&s ,��wJ�9���Ϯ;�x���t�ZD|V��_�c{-*e��E����4�v43`cn�+�w���Ц��"��4�X4w��6t�\S%���Ցhy9�Ӿ��d5#���m2*��WXy �ki�+�֔�(Px�y{L!�8��a�豽lƖ�V����Fl��a�3� `5e{c[*#��i����Zo��	wt�8�Oba?8�y�����ܼ*�N�A�I�h>d�F��|��C��g�ˠ��<���p@Q!>rԆ�����!��Z~�*m�:48ZN|�Y�[	0����Ѵ�^���᭪�y��BI0 $�HX	��.�A�����G���P�:$Ź
�c"�J�bI(oTԎc
�Vҕ	V�HMZo��b�� �1���ĺڮ�Һ�5�����#���-d4��V����U6�̍ <��H�moMSI 6^������j������N�i�؂�VP�u�N5 V�BbQ�x"�0+7����[G(f�GI#h�]Lr:24l=йBf��v��U�����rRI+�E�2�=I}�hm�� �A�%Hk, �k$3ҝ�>N�>~͟����'����j���<*��:��� ���qw��i�<=m��ٯ^�����"�F5IS�?9��h�����OtC��G7�N!�U�EG\End�~���I�;,�hx�����#���~���|�A���w�ڝ;<;w�*�/�����Y4�͝u{睷���W�����>�M���
�i�#Ps�2���m��
P�L�v�5�GϴR��g��W^��M�hFG������z������_�S�NYG"fW/_���yî~����T2!C2Mf�����"R�:~���?#��`<H��d�JE--GMqU"т����xԆ&'D��4�g��jcC*]T&(�����yQB-J�6Y0�����İB��Y��f/ۭ�e�o�ew�����dV!6�`��iƨ}�DDX�l ZI����V6m�����-RA�%f!��2�pmѶ�ɑ�.Aח�Tu�3���>��A��8��h<ꂸxپ�X�u���v)%I7�fp����C6�/1`~A��8*V ��e+�
BD�y��ɬ	�f��>
S,d��BX칄PmF�̓֕L�`U��SBG���?{ �.1!�����{J,wr#�GL��3�%�P�5����OM�� C+��h ;     IDATmk��T�:I���̜;`v��Iݿ��E�tᢵKUw���X"��B׋/�d�+��Ï.�����I�J�� %�aZ��*dJ%?�(q�CAqj��h	�x�y�7mh0 hJ��źC�����'s:�I`iG{*F�{ѧ�l��[��2s[�4a���D���a[U�u�2`"��(zNe��>sW��8�p�D��q0�@5>>j�������>N�������� @⿄��W���ޡ�S��e4_(���C � ̙"�=����f�������?2)1��6�6�|�z���
(1▐�	q�c�{��9�mm8t�o{ż���I� o�K�/l>ɀ��Ǩ�P�����c
�����J<%�ޘL�':nrz�2��E�f��yRlY8� �T܎��L��/;ߪ�#f�o	�0'e��ģOQ��&���
���u۪قU�Y��B�xh<B��3e]C�nVlm��֠�;�!�@8��z������߾�ῼ����w���;�󟛚>i�>��t�9H7v������L�U�(��%y���#��1��z��M�q3���
�i�i��v~�}��svxd\�,�?��mv��2�_��/�铧��3e���ù����f#Ãd c�f��0��޼�>hG=uzFAx`tX׳�����U�W����<^7�G�RQ��z�v�ښ� u��������!��!�Ws�"6#@��ݬ�����ĸ�N�X�*6��HA���e�u+��֒{���ʠQ�!��ޣ%�܄���{Ô�������7E�O[�"�x(DHZ^{��\U��&���9|���������tGqld�:���-@ә N5��u�A�����Y�'˩���;��������70�9RЩ
N������3\�b�u��vt��I����uZVf�uA�Q�kM�Li�zj��Cxr��s@2Ao�X���+�����lykUm],��=vhj�U�M.��?&U!Ѹ(Q�@�9z��AP��*	Mf�'PU�ݓ*���js@��������r���ns{K���ͻ�C�$5H����+�יp���q��5Pu3m_O��J�^iu�Ƽ�G���!kK7�b<!u%�d��H�ũ�^�#ǎ)�#@��@.�4\�P₨#�$I�t�{�����_�=#
�؀!�w�tO�{�9�'c�Vc�.�	 �%]#��¬+鳇]�@G+SUU�!�9�f�%�Z;��gNw܆�o���-�<��d��� ���G�^�YJ�2�!3W���%��`_�"�t�E$�.[�D�3p��n�s��< ��%�1!TдyI
@�W���tư��ѝ��y�>Tmd��� ț��Ȭ��Z���3e�Μ��6��=���^�k@+�B�g��oC|%;�	���"kdrf���f������#T�fn_m�����`$wP��G$�)�p-h���������G	�߻���kw����{s/� 80&���֪]�v����[����5��^�F�����J�D�bj��M�$b�,ڹ�g�;6qHY,�6o���-,>��/!p~�D�WPq�X�n��#��V�L��*ts}Ӯ~|U(Q����3�k�Jb!����ҌP���,bi$�M�C�bf��&$�R�Ж��Y�U�U3���R���2���� ����C)J6y�;}�:��,��ۃ�e{��%[���>�TЎh� �IP�H`,�Ӛ�z3���V�����`���ֲ�]�#A��O��6���1!>���Ƨs�lߵcE��ޠ:�mEg  ��;�:�?�>P��T��Ħ��ku� ��y� �n�P@�J��<㖂1|`�,`��B(�D�j�y/όM)�hȺ��֝�ZT~Y3.0d��#o�Tň��S/h�Zӵ�&��Kn��3�Bs֣A�u��{p�BH�R-'�@����Զ <���%u�c��	p�=�M9b�[�%��}G~�,�ӝI;:y��y�h�G�RIk�� L�T�� �BA.��>�deM�h�?�b8���$�R �`$h�h� L[Se�K�\A����M@��%PN����5��-'�a����{T���Z�#�%mP�ۄC�"�9GZ�x�RY�)f��έ�4#��L�ì�ψ��������s�I�X+�uI*�,��=!|9����,���_�"��djy�-�)�^�_Z�`SP{��Ʊ:�oW���<;�O{4��K�%�^k��dqu��ڃ�GJT�P}Pl��`)8���լkh~b3���"����tJ��%�cl������)ºT���3�7<ʦ�}}xY�R֓���vh�"�G�lT�	�f>cۥ�m��C�#&	�?fsx���u(ԩ��-�[c�*��lמ;��li�|�m[��0�G,��+���)y�����e8\�����������.�����w�x��q��˯J7s���U�q몭����ڪE1V��j�7J5���J�	4����'�twZ(��j����I{��Sv��őj��U&GE�����ã�Nu����ڲp�i�&ɥ��*#׋��{O�F���(n��:E	h{sS�E�-��1{�z���F))����uxH,��l�n�U��m������D<mC�c���-�hKp���S�NX�U��̪�w㒭e�-[Et� �:���2T�6Ί0zSo�w� �\FJ�GήnZym�b��%����e��h�U^귎$��D@@	�E�,@��_��v;�d߂L~�I�Р�fc�Sy���W;� Y���k����Ek�Ϛ��}�~cx�rm��ة�/9�w�PP ��ǧ����74~j?��9 ����!��ݹ5kk���R4�D̞9t�me� ����O����P!�,ִ�����<�v"��Y��G@(�t�zA���{��'�B~��`���c�Ц��ǎY%_���e��A~`{�����@�>+Z�J,������FBU����=P�/��|1z��%H"%K��q���a���ZM��P��OP�!b��Z�a�x��������K۟�Nz;�S&�w >*J*@��'�@���Ǻ�[{�h{�0�(�:	y!��Y$�I8�T�^���>3c���%�=�����Ċ�\����]�r��PԞX�?�P�Ev�B͖�@ͮEU�Z��
^�J�o�|����O�c}��3������+\��y��z:�&?ia�)D�Q���������tB�=�g(�.�"W��=Zc2]g�$K�ϛ�@x�=ɍ�yѸ�N{mo񿱍�+�j:f<O�D�"��e��e�̫����=�Z���l���Z"lt@NK��1G���\�#h�Y:�V�(�{_"%w- ��]�P#%��@"�������G�,�G,�hYo0v������s�q�����MQ�����7o�э;w�v��q��&������a��^�G�����.�d��T�C�q�ҨDA��'�
/�#a�XX3��c�v���L��h8d;�;v��%���T���3�ڡ���D���۶��vv��ꖊ��\�qf�i�܈�h����' �CiUP&�.$iȡT�2���<��c�Ѱb�j�Hܒ���4����B�(N�^~_t%�n�����E�#�i�x�b���T`�:|�N�<n��+Fk����ms�
���[��`n��7� Ԃe��x�J���59� �g�K5��ܱ�Gk�[Y�P�n�@Dҁ���P�^P���~ˉ���9$9��������
��� ���j	ˑ�Yr�\{��}��d)
����{����9����Dϙ��A�����%A�j�Ҵ�@�#���O���3�Q-P����Lg�#��C�^Xxd�}�U+��&��k�K���z�v����>���0�=�kx��%z:-�ե�6��F����94 t�u��EĂVÙ�޲��a;y��=}zFZ���v��[ZY�Ÿ�DR]!��If0����M��P��/ ''��l^��T�ܮN�P�|�2�eHO����3T�o��8M8���ѧ�ц�+���n��X'�����ĚB)��+sdڵ$�$�B���փRX_�S�j:)G�aUV�g�Qoi�0��h�c��*F�R�x؇Lx3Z�9�
���e�
Њ 瑌���%��$�����5[:�d����%]x]'Uyʒ1���;9������ɀ��%¬�_����i}^�E�c �A{7\#�Ͱ	R���Ҿ]��M��Ob\��p�Lymj���Б��P����^��0	���hDi�Z�_���}���m��;�Z�A0���Ϸ�*�Bf�./���ΚeCM+�LjZ�0��B�{���@��9�{�I�f�.;<qPIt��rA�s��g�\/�,�!�����u�7���������_�2p���߿y�M���=��M4���}p�]{pN�Ն�Qɗ-���6�,0�ghl�z�,�j�V�j9�+;1u��?mgO�(e{o����[�\��s�<m��5���y�ݻg,0	K��\������q	2���.���km�J���������e�N%�q`!���UmK��K%ThE�Jym6���}pᢕ+lR7Q��&&�r��Q�>y�����,���#���E��ߑ.n@sD���2	��tP�2�.-��c�t�2���J�(��(��-��²�<\�v�l�&iSӒ�`��$`�'��S�W/�%�{
I�y4:n��eNˬ�1�	�W"�3�y�Х�N�9�֢��}�g��V˚��y�HHk*��p�EH^�N�	�3s>�N���|h�PF��1
�5s�d-,9�`/�G܁�����bթ��[���͚�f5S��r
¹f�"])��v���9diWv��d8�5IT���//>���U��{�b��}vv�=7��sE{����W�7u���kޕH %�fɐ��c�H�iA�sBM��T��Z��N��9��=��N� ���}>����'ڦ�:�J���!ϝK�&�G�D�}�� g�٤�`�|ˀh�5���t�:E�?��`8�Y%���ѝQG5c,�Mص�ᜣ.�H�������_�3��$�S�Sk�_O52nQ-W�=9��W��*`9M���i�{��0�6p���q�.�	c��gN �[H�	���6@��]�\_E�G]����n������(����_BGN�A�]��'nf2ˁU������j�g�����~��v��X
���S2��4���х��_
��Y����vec�2���"�I��u�ydfa5D%��gj4�3�yH������f�d��4�θ��_��2ˇ]@RTo�ƞ������~�b��裾k7���{�<u|�>s���i��]�p�{�`�ʹ������R5jT�e!����<n��C�����6~��m򶰿m�F��M=nϞ��3�'��w����wmimI��8ć��v����׵�V��X� O�#���a���������u޿�XĆ��V,���,��S�W���N"4'c�`�WQ K0j�Ŭ�T�p�AKj�Z�?��67w,��[GG�8(�ܟ�>sƎ����C�-����#�[���̮\b���l[��b��8v�mٖ�K�Y�����f����/��I<�ְ���YX�V�dI�d����H{Ź� �Q���F�а-�" Qu��#��p�A_|���e�������C�)e�q���ţ��0��V�'a�6� ��ô�\($���X����T�� 'W�A��0ɕf���f�R����_��B���d�yED���s���9@Z�s�7�C&�L9gk�]!7U	3#OD�CPR"a��8dG���~Z{;���m�χ����Mi���֟�S����3OYi/k����͛7-Sv�c����CR^��Mno�x:���̛ۻ���b��#�gP׃���=�p��s�}:��
�6J�9	��h���<��Z2�z\I�2s�{ȸ�T�ݫ-��]�u����[Y�l]��<w���T�	�
鵋�U�Mt��]�|Q%���m��p�	���9o�#��Е���灳T�;c 7��j��IZ���p��4��7?�'g��x%N�O��r~.
���0�BZ�U*E�����+��{���F[����*>�&u}jg��ϓ�F"�$ʛ�!W�H÷��(���w�m�z�up�v�	��37������K���e��S9!y��$��O��*Dr��=,�ڻs7��E���V��E�˧$�|:Mā���s@{h���VJ�:(� Z��9�.�&�0 S�|��b͖�FwN�����w.>y�!����z���[w���콹_<>}�^y��6:<����ݷ˗?��G���V%���%� �*��L���i������){��e�7�hZ�V�Ƀ��矵��O������G��åG���g_x�&��F<�u��޶{W�Yng�
{-L��y�̈�%��F�Ri�UF
��#�� `�	o�Q�~�1njV�K�R�d2-�t�1M�";�`Go��$�q�=ܹs��®o����`$��]>82`��M��E&p�����5p3<�8!�F3`�
�����S��1K�X�#jŨY1زF�U�p7��7EU
�B�A�!���0sk8^0_�9yU����: WP��v��y8\��fV����_�w=@U4� D�?W�xT(o.	Z�S�~eP�T��2��#s��3��N�������_�n[WGJ��iO�S�F>�U@B�Q:\/_�Ci���b�N0��⋙�ڝ^&�&��+a	�[t�0�K�,=�o�g���"��={Ξ>}��;�V*l~i������F6�$����?���!L����A���sV��m��=�y�me���<qlJ����݌���JD@asPvB� L�M:ܾ3�4��
ר ��?��T)�mf�3U�g�$���LdU��\�}�n�O��C0CA7����� γV���G���u�l�n�{�f��R9C�����s�����~��F�N�7Tx8�nd����N�����o�k�k-�5�J�Z�D���<���ˠ�$8w6G⋫���P��s�؅�+�KWѱ)�D�u$8�ԡ��!�g����}*��C�����mb��L�s�4�h��q�s bO��#���r����9�Ɯu�}�XU��iE+(#!�}ٵ��@M�~�n�g����5��(�1>:�I��E ζ�I�YJ��k��Aq�ޙ�iW��-3+�Ú	�$*���u%Oy������*�����*�liћY/�wh�G#����[�8�0��~n��?��?18�[���w>���'_�s��^yg���7�h�޽_8q���K�0��ٶ��X���;��p�J٢5�u�9�i+r3iÍ��� ������l�J�K��>xȞ=s�NNW����mo}�����^�����؄u��6?{�n\��ޚ�r&�P��d���:�s����(+%ب<Ģ648�kwc�J�a�z,|�!�;҅���ba��NZ�Zr-NT��szx,���.�Lu���m"��ٷɉ1��C���,/�鼉�q��m7���kv��Az5�*�
�^�[]���=[�fm?д����z���NY|���}��"p��������f�V��,��!��H̊uO�O��U�>7��Is(�Tu�a跒@��=�b,��0��G=P���kR)gE�D$��p�:�D_�h6@���jC�`�[+9 �'y��C�$���2��^����ż�!�� D��: ��+����*a�d��c�l-}-Z&�Y;0��,	���m�N.eՎ��8+J2�*��瞶gff�U��=����~������d���i�b�1�=h�'��s��Ze?��~���$8��:{%/H�:��- � W�d���^>+
Z�3���hFº6Q��u}�/g�k�$U����:D#�ٙ��4)q^=�Qw��\�T^�i��Pϊ@)%:O�=�{��g��;R60<�%f��� �ǣ�WRdC_��Q>5�d    IDAT�̏�����(PS�� *Q��j���:k����d��JU�'�d\�V�ɵ�֭�������Ob�p����K<D�7�g�PҸ�'v_YM�C��3��Y��
.T�b)|r��fኣJaL����ą����{z]����z��Δ�d(�[��R�]ZZǝ �s���X��(Ja��Jֿ~���P~rO"���
�(��I��T5���P��GG���P	�w콇��ޣ9��$�	Z�V�LٍIܽ��5�J�ٻ.�f���č�~�K�|A����p�H䲻{��'��O�d��������Ư���a*�k�n�������<�Ͼl�M�����.��B[�R���Q@�EӇ��V�Z���'����H����I�,S.�
���8vTg���lys]=��^xQA�y��{w��ŏ�Ү�� & t(=�|ffΨMԨ�,��5�����ʚU�9U��1�F9����<�!��\P%Ò�+ʢBe��:�ɠ$F����f��M4jv�������^�=Y�T�
����$���C�	Q��x"e�H��͠�f����kk��jT�Z=�P_��>f}�-�B�n�+:��#	K#V��-�����a���*5d��/W��7�r�!�*<5�:�&p Ti�Zu��|�Z<#�g�a��P2������@z��T��W���_�C�[Z���8I��H�V�Rɤ<�G������ݼX�Me��N�r]O?���������W�&4+WE�E�Ń=f�e�> *�<�s�i�JѶr۫-��m=Ã���u'x履zƞ=}ƒ���sr�fneo[Hw��4pkj�{�w�N<���sq�=���LfO�o��rU�*j�Z��TR�~"GKs_�1��@� �¾`�c�]7 |�0A1!	��Swt5�D�!U��f� �bфC���z-C��ހd�;�_w'�v)�,(�R^S���{����x�AO�գ)1w�-2�란�5�����ۢDěk�cy7�t���O:�l�gwձ����ꗵ��4bB��{�Z�/�0��y�z������%��{O�# �嵫2{Ba��5$K�U�<su9h��c
�C#Ú�S	�� �9�����H>��ڊ��������}x��RE��W�KM�N�� O���xq����p�Ft����K)Tw�.��X/|�@����PؒhHh�3g�(q�B��?��r��W�K�}��t�>\��r*�p�oCx�`���;�O2�%Ѭ;� �[��Aj{��]
��HBϚ}�yR/;8�tL�ӭ�����?��o��S���ƻ=7����nޝ���S���ӟW��hgg�>|�}�׃4}��̧�s��Ӫ653P�~��	�Zz���c��LJ2���	{j�Zm���M{��mekC�g�~֎��ގ�-ܟ��.�ͫ�,�횤%i�V��9�6v8вAh)����hW��3�\�����B+�I_:O\f� (]��BQ���\A�N h�b ���4ԙ�bfǚ��%#;21j�i8}Q��ٗbk._��R^D&�m���࣡c݁Bª*�m�em�X��p�]�F2� |��6~jں��ā�l�����+u%+�xl���/����#Un���t��f[�`i�x��j��9�
��Tb��94�c�ɱ��YT��3� $���k�}���t��x�d$W����mon�"&X�)|$��pKzGV.�ܹ����a+�e�s�قj��R��8xi�1��e2Z����'pnt8�/�C�~�N�ª�@�ڢ5lf�-ۨX�;e�c#C�� Gy��9;7}�ҁ�|iWv��?���-�[�^u�M���m�o؎�N���g������ma�r��C��V3����ͮ��cQ+�JBa��p�8y`:ޏEAأ˸`��GO��=�8	*S�9�9���LIL�n_WT���ۑ{�ڝNŭ��3��:+�3�Q<�4�]Ã�=�o]��j���'Bׄ�F f��{��)���!�����sb��ͯ�� u�3��$~�g~�@h�셖*��UR�bL �G�����ԸG��R�=V��t��DA�iG�q��rk��)��B�]��D\I�ǟ���I����ú�{���������#r��􄟿��bo���}�!Q�_7�w֋�8�&[�>����"�&��eN�wE�
�gý�iPn$���T�ǎQv]��@�O=��t�ֶ��]\�k>�k٘Y&�g�Ź��I��om����\{���5��{B������:8 ��4e�w��E��1l�m�l�����O~��ڴ?���ݎ���,��_����w�G��^8��M�.������'���#}�Z�Z�unX ̆����6���uvX�����{$Op����x�1z�م�licM?���Y;sdJ&	�؍������Z�T���� ���#�Y
�]�.��щ���r�{BFSi!0�6���.Q&�x�;Z6�E�]�J�ʥ�T��X7t��.;4<h�f�zQ�IŬ'�f�,@s�]x�+U�5���HC���*�u�,L��s�*�h6�6)k�0J���6q������ʚ-=\��֮g}�L�6�֕���&�̥ ꣓=^���K������%ҡ��� a����[R#�(s�|�k	�z���AnX>5�
K�HܢB�Z���a�kC�\t8ӎ�gjl`Z���;���t�C�o:Su�Q��^����4�M�P ��ߡ���U�K����=�o8d���6��8iI͡�3{B�ӎ��X2�J���C�mfz�R�t�يW	?�^�Ij�*��=�vx�0��������m)�q�e1����I�xsH0G��{!�Nɱ
�	F��P�M��B��0����s�3QF�����,��:��� L5GNE��#���
�Q�xO B~���z�`��P� ���I^���=�tʆ�G-��%��R�bZ��Ui�6�:���?�~Dbh?�2yI�6�%}��x���$hZk���|�?�I����j�����U(,7�p�8$q�"�� mf:����r�7�}��%���	�*v�n��y��:%��h���j�{B��3T�Я��������	;=3�{���Y���{pA�$��5����<77�mxɦ�n�{���S���&|"� �}�t�]���XS�y3���P0(Eħ��R=�ֈ�l���+��ң��O�a�T1+�����FD�BJ��t3��p	.�Hi��	��Z��ך���mM*a�!���������7�{�& ������p�Rǥ���+�f��ġ��+���?6%�����������c�Ri���C���WMm_��!7�A4��H_�|S���<l/�y��;�m�o\�PA���K��'�n[ZX���Y�3wWm�l./�(d� 0>��a\�[G8bcvxhL^���J͵�%_�K���&D��s,	�1yA{L�[l����K%b�ۙ����v'�'�a�=i��LYG$h�bIp��E�X+�jV�4-_��YQ8��L�Y��V��9 �O��-�R�-ttlx������C�����Ҋ�R�7�%推;HY��R�"�]�Il�X�,ڡ@]�/@�ِ)`hN�y}1��؄NѰN�⚂�KJ�9�L�#��vh`H�yÛ-SY3�e.�f����>�:��x}��d�i�&��pT*Kz]�m��H0ƛ��q���i�Z�z�����A7�θ�X�*	�'?Hі�3��5$�Ќ8,$"R*���f��Y,��do�Ei�vt���6<u�%�f�r�V�7���}ۖv7=��Zfr����6u��}���ݜ��.Z&��(.��8�h��s���V��=e:]긂~�9O�X�Vo�}dT@B�Q@޵⅐������U�֦�cG�*�v��?|��戮v	K��D��<ɍ@@H}zjM��q���x��D��kQ*�2Wٹ�C����;��ŬԬZY.Q��dqc᨞c9_�(�/��`6ͶuF�+�ֵW�� �(J2\t���
́��C��ଙ-�$f��6�yU(�VA�V� ?Qg�V�l�;���RU&:�ks;�J�Ni^&���d������'hd/8?N���jMv�X�N�ͽ=�626*~�ݻw���?�;���VmhC����^N�ʡ�y�$����RW��*hVM�F%�#���K8uN���Z|�6�L<�>'@=T�>s�&��[�;�����y���`����tۍ���a���V#AV��^c$�p�.N�x~\�P�tAK�����m�"W[t�x�,���9�/�����/>�J�ͅ7��]Y�חo���c�=���:1� ���!�T�r��AGX/*����kOϓ���q���Qsnߒ<qtʎ����=8��o}��-m��=uf�N9��+�����>���ei��KV�4`Ɇc�sk�,�,�hJA�7��v�q�w����sb�bq�&GȠ��&s��%�i�ұ�%�aK&�֙NX_w�F�l��Sx��Ӻ!$��v6�����py�ֶ�V(֭ܠ��u(e�������v�b�`S��H�a��TLݣ#6|��9dA�0����Qk
"�\^�+�c>�D	��NX�O����PO�^��ղյ"I%�^�K����.����� �͖u��m|tԆ�-�L�#��[�j��.w"!ʛ�ohE�ګ�eV�����Ʉ~��:��Db����(8T�f���|�jǽ���:��_���u%lFG���l��L��TJZ���}��E~�a�����X��:�]&��d4��pdhКͲ�x+�jG3����몦 AH�ډCG�_|]�A�.������-z�d��M1�;�E������4 &�I��D�>�vf��v5��G��ha��C�&��> C7$��.���꺒(��ylӶ�x�Ҭ���t�e��*�>�kw~2�u�Z�B�.����c�1(�fq�Hcʨa?�6/]_x��t��D=�I�S�s�K������'��#N4�_Ry��k�kv��1�%	CG�	� Rì�.
~�$o�坑̰�R���R�z�,�k��:R^�g%��7�&s]~{ׯ��� �U�q>׍��+�߷(�u`cR)=�G�����:�����grhe��pؓ�z"eO)K���<K�s?P�8�y�?Lq*��S�{�3s���Q�V�XG$���`o��B-�֭@���C�U�~��-5����F��._7sV��)ΤT�U��ZӲ[;
´��<��Z�n�W���W��O��S���;;}0�_^�q��8�:w|��͜QX����¢� ��dz�phU�umJ
(t"���R<n\��p��1yR6�?`c]}��Z�^�l�ho�-��*� /7up�z��mmmU�� �!i8x�ea6B$��ζ���V�۳f�dHvD���n�X!W�H�	�|#�T$�P���a�P�:�XXEl�Ö�ۓ������lh���{R֝JX7��R�ʙ��wˏ�mv��-�gm;S�J� �e��b���i�ctQi�sY�Z��ښT�\�$��>y�&Μ��c�m�Z�m�-�lZ"ݭ6?`}}C%0�r-,|�u��`�,ݑ�b��c���^F�Mk��x�'��"�!P\J~@����%jU=]���'$t-���є*mQ��n\�� ,:�?��7U��RE��^��eɴ5��J��T(��H�O�ǀ~"n�FK���W�;�ܾu�fo�t�]S.D�� L#���A�$5���^1KvvY�����ɩ���P�kR�)�**p�x������ۏ~�whU��י Ը��m�]�2���o|K
t7�ܰ��xC����N�C�fT� It����؈S����nmo��'8�� LU�SF�<'q�确�qmS?����ёUр���r�l݉P(ك��
g���͡���φ�J-� �Qm�ݩJ�F�]m��`#��}��Ʉ�0t��8=zP�{����{�,�A�,G������}���	�~����y�����N�'U�R"s .��ĵ0�m��sH����\�>�u�% ��2�����*��,t{ֵo%r�N{��m�l���n�L�T�r�adz�� Dk���Gb�x�*4��t̐���S��P ���T�Q�Q'D�w�y�k��<:�<q�=�XȔ�.<��PHcA�bkU�_�΁Q�	�@��C=�����\, _v�:S2�P&���}�̚�ٰ>�q>J�� �3�hsT/T-�nE@A��]>u`�_���+��ԃ�o��0��?\�5�o�&v��:iO����&��e�t I�AKn��y���$��=���d�S�p��]IKXF���0+7*������ʒ��3g�ԑcB7c�v��{��f���vk��p����d-��M�l�Ƞ�/�m�p�o�l�[v7�f�T� G͹�T���N$,�xg�����H������h�����;M&V�%��b�j;[�_���meiݖV�l'S�|C��E��H�'��� �Ył�%+�K�8�">-$6 B���'�sl�zN�v�b��Y�ް��?`�ccV(�ʕ+v��E�9 *-e�ڈ�yŵ
�F�� L������,�U���hA?ªhZj�0��L�A4��o�]����H�2�	������]Vjv��1����gm��=�Xd���Қ��
�IH�%J�0��E%��h��~֙�ˣ5�����agW�~��~CH�����29��!��&] >�z�Ƭg%�!w��9S�HF����	;�̳6}��x�� �@4 .e�a�@�6�{������?HoW��=�b����i����+:��n���y�e�y%v�z߾����������lR�LQ�%Y�D{$�@&H`�LL#^�1xl$��1�d�$�x$Y�$RII&)���}����W�����{�9�{�;F�X@�Iv�����}�w���������ޔ��^l�p3㓈G*��RńW$bA�:quc����>Tѕ� e�T�n�!�H�`�w��$��ڈ'Ff��<�闹�����b/Ґ��xp��L���3o\���v��94U���f�
2��FW�,���v�T�E�VךAn}��ds��F6�~>5�]?�X�d�ڰ���=�S�y��<`�K����q�5F2�3�/�O�aD�A�p�Fݰ�{.���L��le���3��j&MK;E��_���rO�g�xI�2�VZe�q�ޟ��m8.���@�Ū	B1-B�f�R,��\g_'L�31�V:�晭C>��{����c��AD���0s����k'�TƟ��Slh��R7�'�Eޣa��gˤ����	�H� �(j�v�%"�.#O�>\v�f����M�"2ed'�����tNb�i��T�Ґ�Q'w[KO��'�◿���ѿ��=���?����&���Ǐ���#O mE�8(FS�M�'=����ٔ�c�pM.��.t�{���(�غ�A��mcuk������
��'���# ٨\�9ܸw�܃������"�Ш�M-��hUj(헙+_ۥ.g ��'<�i���j�������]I�b~��i��cht ����.3��-UQ�-"������`}m�{%*M��|�~�=d.F���Po����sY�?�@�Q,E$N�j!I|h7��{Q�C��G��� ������H�s�!kg{K���n��e���Y�4<P�M~`��)�Lc>�EB�dTk
0�>��@�~�L���������^w0��m$E�,����L��߸�+��C��`?n߼�ٻw��Y�6��S��F�R,�C�2e�
j��e�Å� Z�z@�%9��ĳH�ݍXqk�˫Қ�{���k�y��b6>$��6ӱ��uv��@H�a$Á�q��������Y���	�����K�&W��ƛ?5�n����/#/�'��ٓ���(��[7n��w���ܼ�Č�G��>�tNR���e~�,���+�kذ�.i����M0x(�XE�7��D��͉�$y�q~-Z	E��j$?1|����urA�By��AG?�O    IDAT "ߑ�i�u�2�S��:+���Af)D�8�0��^T?Lh"��Bj�	� �����U8� bh h>_��<��+�疚({%�Ɓ�?kM�������?WS+#�����;D���-�='iH�?�e�]��G�1��iLL���m~��N�[�lP����mxvSe������h�c�0i����j�!O�8�����`{�hV:|_�\�P��Á���BG
(�� .@ѿ�R����@�4l�)����L�Ō���sa�SG+�+�;��#;������繣���L�4J+k�O�良@�kT<�jK��DMy^��F�ʤ?�|lp���~����'a~����o.ݽ�Ͻ�@v��!1���C ;e���bl�=�v�9��Љ1���q��G�؊��:�>�ܬj^YYӎ�ږ�G����L�jo��[���2���=��]'�����ֵT�GH�BÆR�0����i�Mvr�
����c�_���B��F2D<�8w~�-LF��e��k�U.�������ͭacm������ڠD���W4��*5�<��71;Bn�XX6n�hXd(����4��Z~�R�.w ��-!B��� R�H���=��y�..b}su�������+)oHAn��v���9QУ�,�4F�l+OYI:��y����L��f܁�2pw�d��a�^�1֑d��:\"�G�04Ї�7oj�}+�L#�H�eQ�41�`^^˞�e'G��B��P��qjKR8y�0�D���U���fҢ��ċ�~Y�.�3�#���΃G�>jX��+A�%7� �����Cةo<q��hH�R�g�<	 d��h���_ZY�G_s��	Y����r7>40�3'Oዿ�E%�ܹ~��3�//Ir���˒�{g�:��s7V�F�ncB2�.]A����%X�6r[�ɭ`��4����ȃJ���97��ܽ�^��_+wj�u���I��$���'������EXM�}����@E�òF�x6ݶy�M�CCLcNOmN�*���d��`�ec��y��u�ٽ��5�u�(�b��� J�rރġ��.��t��^E�����]�_��X�Z�Z'b�/]?�V�ۓ+?S4�gfZ��"��	Pn8/�V��`&P;��.̂�9�W��~�J�7?A�W��� Q �8�T�Lm�D�fZ]�������r�[��v��q9�����C�Y8)jl���RqYdǆAg�\��F���0Fp��wO�
��1���9!#���dخg,O��K$�G���2��Ǌ���ql+׎����ғ��Gg�ړ�sG����wfG����|���έ?nt��^й�5!)��89P|/��er$�d |���|�l;�A�;��	P�ώ���z��v�zYlgR�}^�x�ƹ�#xbhJ�`�mrvlc��b�<L�j�=Xt$щA ��m�A�
%�z=�E
Zw��jT��6Ѭ�V�G�V`+"A/�ɨ�f2��i���}h�	�屳�"��{��`ua�k�D��x�M�o@E�I�{|��-ྒྷ���"4�ُ�a$+����Z������=p��F���Ȍ�`h|SSSr�!C���p��a�d!��"�o���XQ�B��e+-&�_u��Õ��$ev�$ݐ���b�o�'U�i5��ԟjU�G}�'q�����Inp�ׯ^�N�1��>���I��w?�H��� u��C	�9�b�:�!����=��M����=2eە��0'�N���ۋ�l��m$k,T��I��w�8x�z9�a"����14:"��X<i�ݲ04�0��^qO����EM�|]�ܦ�-,�p��=��d���翤�J��������
0M�GL�� ��HT��^~_��N�Q��5;L>�|o��`�-lmoŢ�^�d{2t�NDj��P#������0�yp+��2іN.���A7��	�ϱ&f{:�t�!.C6�"���2E�mg8;�����Si�	�����Ƅlug�lX���g1T�`�s���A϶?TCeQM�6��iz�
J�����!iu�B�Y���r�p*�F�>��)��f�ip��o���&��I��u�i2���^�)y=�ܱ,{���%���u�/���
�������sϛf��߫u�L�`,ou�ѫ�ps�T���~6,���v�����P6W���!FJ�}�3}�"M���XV��0z��1�xͰ��߃��D���`�����$N)י�ym�]�	Ż�*���pvu�"��;:�nȎ���o�Ӌ;����{�?x�?�������n�<��x��IE�Ad�J�Ё�����K��V~�O�	,��>Ī�EIE<~BЕnC��:;o.��:�0�9�xr�0.LƱ���͎I�	(.��m2�"������R�Lm�!�&�zA:l����Z.�v7*hsZ/�U+i�|H���H!����J�7onF�m氽����l-���W��n	�j]o m��D�2ݝ��M���H��l�k�CpG}K�Z�����\�cae;�j.�����va��D���ءx��I�>}Z�Uժ��=����J%aA��R��G�44�X����@0uxB>:F������{7N>���!$3���ʸ%|J͟􀭮}�`ѩ�ב(xp@)A4}�C;15�Gcdr\��?{������O��/d���q�K�7�� ۚ�d$�P���(��=&!��Pk(uj���&��B:����݄g�?%����1���D��f�Fq��N�,���O*"=��B�	i�i�et�����|�RU���/�����E�~�ɐ8	��?g� �b%�L2+$�e�~�PM�H��ǵ#H6#a�MMn/o=(ómP��u�l�D6wcC�R<�-�(���v�|>��g�E�Dۑ�l0f*3��,"b��)n٤,B�2�`���	5�����eT��N�&�+Ru�0�?cB���Cܙz�lr��(�@��>�f����⫟eLj4h��qM��n�q��&g½��~w�(�Iڄ0�����%p�g�e	Y�y-��M��3�ƶٕ���]�0��9��oas�X����N7-s��}��6k 51^�~gL::�y�s��%��+����U�x���̛�iұ(�r��j��(�EX׮V7)|U#��D�rK���ky��a�%Ѣ���b��Vد�\�g���aTn���&�ȭ��4���p�0�U֕@�����9���ә���^�P�9���߫��+��o\�;����Q�]���
�&�% =��O㞕I>�l�qB�c�Ǘ���s��=a���zY�H�oM~-�R1��ϩ��i���cxj�0�����O�;���������v_�Td;���n(Z��U���)�U)���mBp�z�\�
<=j\�H�CH�"�&Bpq���Y��J>���
6�����Ge�����]/��z�j7{ܽR��F�U�n�7+!f
�pX% =�KM�*$#T� 2
	[�ܨV��&鈾�L�aQ`�9ܠ�wdf�y�y|�S��aI!6ED+6�r���5,l�`s'/�������0��7���RT���r�^cw�f�B���vK�ŉ@g�Ӫ�?�Ӗ$"��Oڐ�i�R(�����	�����
#2��DvpH9�\��]���rY�N��t��>�LΈ�D��"�d,��4	?<4���l��ɝ�T+汿��'r@�6�
C4�i���������z�,v�I<�'��S�̪���E��(�!�$9���$��w�@��|��X]]Uc��/U��{_y�,-��s`f�>+^��Id�IA��tM��4ҙ�^7��~\/��;�����٬P���u��T��<i �=�x$L2��_;uN�+�*�DIX�8�U�T$�w�2�0d,����N���[f'(�#��f6EA�Ǧ=��v
��GQ�,��	fߨ0Dֳ��3�;E�;v5L��y�fp����D�U3՚�)z���}y�;Z�]��)���#�|L;�{��2?~��ִj���$�YSH���M���u��S�V,�%SP�}���5,f#)r�z��ku�xa�՜N��S���S�h�j�	��/���>� Hff��BjĆ&��"�J��_�$��M8\ȁm=�5��AEr�P�jY�] A"�����QHD�d(��m4�wwP{�
Yh|���Ӹ��*�R���p�J$뒋V�n��TLs�3bS�{V���˿?�����ك���/^d�����*¿��_|����?Y�^���j��H-w�v��3x��B��F��B���Z(JF�Vfno�2�$�p/����p��Ut�^춪��@��#����8�?���a��P�?,�q��.����_ԞR�|W�߃�E˷� S�]�H��Ь�Q/ᦜ��o��0ZyzHF��&0З����m!���.�,c��]l�_E!��n����At=,�*�6���y�z��k�z�}*�������q&��,�NW�:j58���g�9�^O ^;�U���2&�{�PgΟ����x�駑N�ǰaQ�|��m\�w��n��w~�J�.XD~��v��!��Kr��,��ӕY�z�&Bn/I���S�@*%����Y�y@����.�~?¡4Ig�2~Q��׋��	L�L!�׏z��wn����5������A4=s ��8��G�K��"��v�,^"�hgg`G�lL�Aܣ�L����ۚ��Ǝ�C^/����I�iX�<�+=���;T���$\F3��: H�kʭ!�h��;�����)���_}�UE�����/E�'���G�0�C�H���n� t�[{=�n��P��~�ŝ�c����6M�2��vw���'�������v5�ΟGr$5�ԣ����h@��X���6a���
�~YTe�(,�M����*���%�F�;|�(����;_B���n_,&�\�(������g�R͟+p"F(hc3��F����*�Ho���F��~p"��VD(�8'&�ި>���ܘ����y��fڛ����l��h�jyD>U�ӝ�9��*I��V����ò&���"\���ȵSv�iN>���b>Sl�����&�Fd�A�6N؉]vv��v^�u5�'�ƩOM�mZ�3OS�}��=���05��XL<���aË�|�h�}� ˍ�R�ʖ-�ʜ�u5��2K{�v"�i2#���?�)����X���.b�}������ϼ���+��w��^}���ҿ���pb�QCl0+�f��F��Ԯ��Ѷ)O��"���{�W+_]�����5F/H�B� �C8���Fa+<�lU�Q+�L8&�(%�6�6��LË�TV�":(ED����#4�Q���p�X[Z���"v�WѮ��*���6qa�4�"A.���VB��T��bn�|�*i�����$v�U���ѥu~��B�}A�<$y#��
�m� ����B	�e]�v����֒�41s���o0�[.Zt�#@��� ���x�3���C��P�A�F�^jT�oVq{��ݺ���%lR�ͦ��@�������@�6Ƅ��2��Tq?�N��D�
arhON�`0�A6�.т�u�.��tV���⢊-�R��ӟSNE8�E�����a�iS��1����b-�*� 'N��ɓ'q��1[�e��|X�6%�b`�v%;��<"�Uj���M�*Jn�޸��Ak��x�I*c{\���Ȥ�}�y��bdܐ�2�s��;pJ>��3h��y{���"�`_�&h��^{MF4<����2�_ZYV^�{ ��&��Zm1}yh� 3)H�����h!	,r���)e��^a_"?�KX����i�a��d�<%C���1���:�..i��vhrz���pg''�3g�	�ʿ�05�/�u�jNf)=�R����_vLb8M��<̋�z��[0���8�-�#f��j�T����l3�t�ӎ�W6;�6��zlm�%�4��-	�ѕ����P�c�bB���㖠��y�;�W5z�<*r�������122�喜M�;s�KLa�+F����Up��(�z�@�|�Z�Ab���(��pRN���LCÁj`�f�0>>�T"���aC��5b��4�Uz��YO��p"D�y�(���mxE�#/��'��D�Ȧ112�ϊ�yw,�}p%��R��}��Y	0^�H̨�
��g��)�3Z���ohE ��kt�L�Y�)�>鄽��d߿?5z��~��7>�"�g7�yjn{�_][����&�})�Ը�4�T��(&�R�#��!��8� �rY�u��:5w$���R�@u��N�L�tW;�
w�Pb�K�������m"�H��Ŕ�J[ʾx�4"^���a�����V���~+�g�b�o���_��Mm!��$��k�H��jqOW�ۏ��v�s���T��Mƕ��C"[,B8�)8�ˇͭ��_���*ַ��_��+cڸä�,�pOŹNRW�!�4�7�u=�%���G�/���sHg3��(a@��{ɮ����yܺ���WK(2��Z���T�왉��X�����g�}�C��ZM��829�c��L�@���Uln�iO�&$�I+���ܼ�cN }}A���k����a`�K- Q|�ooaqs�;ۚ�I$�!��S�e:?=9�״KwB�]�K9��)4A��hl��?y��<hTj�����&m����.�b��<h�;Ib��l2O�;PK�9'�h2�h<!��P�w���J��v��R������b{��-�o���+R�"�蕕%��X���R���܊(��(?�vr
 C��j�.r����ƹ�%�b�񇃸sKkk��+��4#0U�I�������#)O����եe�'g���z�w&�ܪ�ܢ|��h���kg���2�[=�v4!�m��%n�!�f��͘k`UN��g$��&a�jQE׎V���"�a`�c#C�{�Zk����m=�%��l�o�P(�~��jBFX�Et���UP�n�{fju��Pe?��U|�"�����2��XSS�7�a���=�ys�ʵ��ʺ���r��[ϿM�li��3+�e��
��)�p�ц��|r+�!���V���Џ<�ɩq$bчtA�JS�i\XX�@�N����i�����l�m$E����3�"l�c�$�L���>erA/��.�V9O�����O�#�'�;5�6b���xv
��lH6%�ȥ"��p��p�yk�����������V>�"�Vn����g7W���[B�
8Hp�� �ª�����*T�+��!�_ y���<4��t<"i���#�T��zQ���{�:��y�06�p����XF���@,�G����E��P����c��ټ��#e�J>���7p�㏱�������L�C�^A�YQ�s�V���k�A�=���:�C��좢��.-�zmD�)D�I�NObxlDQv�X ��j�Q]ݯb~a_����K�*�2�:1	J!����_�:w'm4���ͤ�~-�J!�?������p��L>q�l��t1�:�&
�26���za�C�.�����;$�7�}��u}o>��G��h?L��:?;v���l�0OcrhǦ�152��ۃ�7o�NA�sفxAܹKHհع�d�'2�
Ţ
G8�T\�+H]tG��v����M]g�h��8~
�ΜC&�U*���wѪ�PN�#ݚ���Y4E�ٟL������XCN�*�<�zQ� �~���IS���i���Ј��I�V
��y��]ޅy�(&�G%���P�{w�?���C�t�|������ה1��_����V�V���~K���Tkf��x����4RѤ��غ��U��ln��E��v��TV$�щq��B�(��`e	ۻy��`����Y�ү?�E&�Ԯ��L(bCc�\�[�f:��:Cf���#��>z*
��&gD�-c �Lg:�).�bro��}8��c�K,Ԇ����nBT��c6>��x�FBf�94Я	����ϲ��D�8i�*�m�ml���l�)2"\I�������"�L���~��w�^���DW    IDAT��:��ɦ����JA�Z������op0����2`a��]�ݻ��%�cG:;ua�i6���h׫��fKE�^5Iaj�ms��Ƌ@~^�#d@����(��(։��p��AĢD��|fSb�eF*2tn�K�e�axw�d���8f���@����H�Z������8N��y�6���jU��n��"^�c~t�,���ڦQ&�����u��A��jή����4�0S�H��N��C��o���|z��?��S������c�����s�������-aQ��(dp6<���J�����!��N0I�:�MQT��:R 2W{^��m<+�A9�TȜnvt ��P��e>��6�"Q�e�pr� �R��a�	O@�	��q�Z,�����.ܺ���e��X.��nJ�&*���VU�f��B���eWI��X(�DY��6|����76���1���H��S�g0�JE4�Pl尼����:f�ֱ�SB$}�F�X��#	�ŗi�nNB,c��TZ҉*���ظ�fϞ���Au�4��Β�/�Fy�n�ɍ��1O(�ˋ�57�{�KX�\�Va_1'{v��;�'7:?�LU��J�_���DS�#xbb
���-�6%�D�Z� �ߏx_��>Pq��A�MR�,hO^�|���9��#m5��}e��"��6&c���8�)Iz��6"�;�L51�tQnT,�$mq�<83���!i�	�2��4�6ޗ�`Qpl���&.6\��,*9�S1p��}ܺ{�K�2A�����I�N��#c����k�}�B%`������n���W��ʧ]������=ܽ}S��ןLځ�>�c	�����f�9��W��#�/_ӽ�v���H&q��gl�D�g�ɝ.�"l1��~0�X���B> �y�E��;�ƢF�eCξ��G46�
�<�Il�,��H�dM2��D�t��w{���i���H�j�;����1��P���"����btlP	mcc#�ǲa�}#�%�u������=}�����&�H���S�eT-ڷ��.MUn��p
y�V}����DrP��A�E��3�h��h���~�|TD�χ��}���oi�%�M��?'tF��#w(~��B�iT�V����tR�$oc����c2�)K劇�=cbl�N���I>��N�.y�s��lj|��}��8	5�� I����NVN��s��f8E�� �`@�hO9,U �Y��y�5�ȹ(��(G}hD|h}f���/����l3��ღ;)�gm":C� ��:���*R���7G���<7s�w~����?�"���}�Ե��wcu��j� R�ʈ?�Pσ(�H����D��B�o����{٩�+�-�i�p�+Lq��!|�P�w��d8�lZ�%,�P�U�s����1������ax���B�
#F��kU�lnb}cUZԥ�y�VDS�[Z�t@%	Pnt�54�x[-��,��1v��ei�����H6�h&���rz�k�,[)��k�E�Wװ���͕�\ۻ5��ĉ�pYA�a�8
:��'*v�<P���	�k���H�pT��#cc���ఁn�Y=R�-�����5�fF���KM"9�w�2n/.`a��xj�Edcb|:�ёJ�nO&M�	L�`��Q��3�7�e�;*���>�}}�f2�ԣ+�1uʄ��;��h*!/�ͽ<�67�W�(Qk�{8�%(o��ϝ����_PQ�w�&3��pg��JB��b��v�͓��y��1}�����	���I�a�Bx�a(�c�J<�k���h<�X:)B֭{w�Ə��.}�?�T_�&g���TV�G�cc����r���$�b��~ 8���k��5}��܆&��s���^�}��A��|݄��îHI^cp<.A��s�$n�!Ǧ���<0�@4�+7�cuc���:��5I��ćD�ZSnBR$ԛ��s��S΄��@�i�uL:�l_ZE�DDG���C�[�lB��1yr��$�qU;��q��m�'ኑ'9EF�О�59j���E�!_�̦��p��)���(ؠa�U)�da�*���Y��>�'�)�>��cv�I��bu��d���e!��{��!�i���%9	�a	�/T���Ko�s���ȡ����E�0EQ�R����ʕkX][S�3[daۘ�F�u��o��?�X�<�A��z]E�v��9(nRf8^��v�p�a���¹���ɣG&	}�M;X����q�nݹ�B��������$Hj��(iI�-�^[&,D�d�i�1����C019�H*���r�
�v��v��0��^t�����*�v<���xb=+~���%͝p�,+^fy3���l�����<=s����g�>�"��n�������ۻ�K��"B�(�0R�w���Ç�˯�4s�u�S&�;����ŚH$u�e�������3��-_�/�Mzt�lk�;X�m�)��l"b�����0K �P^�B�
c$�9m�q�p����Ϊ����D�X�����/Y�2���Lk�wt��.�#�����cuâ�U�d�'F085��@
��ш��"��_����߼��[w�zoŽ*X����Zh8�� Z��@"���";YG,HB\��a����db�h\���	�T�uM���v˱d�O����{N�SBO� 4�Bܟ���������9��1M(�%-���]��p���!ң�m�Cau�9���蓴�s��[]�NnSל�jfxX;iDLOO
��}�6���S�013-쥭uܜ{��JQ�|�n_�鲷!���ᩳ�����Μ�q7/_<��DЗM� kq��v��̴v��pDS'�Pܹ�ɉ_N�:s�w^��IV��"�oBKX�H�#�K2���2�~�]���{�1'�i誴w�Иd}}�F��*v���$Kq�������:��"�SngKE�����3t��aM�������~Qfl��s�ϝw�L|"/_.��nG�N<���)��oa���n��,�����2 �lr���+��b�!��f������A��î����<�,��.Jt������u�K>�,�^�J�2���H�loz;���q~|��sCr����ԉα�g���CS�T�����cƤ�e�h�B��w��>��MǺ�o˨H��ШDǎW���5E��<~߿}O�ɳ����fX�"���B;>��g�Yg�q�d���ʰΫ���.]�s��5����eַM.�w�"e�(����F�ar,߭-�����Z�RJ~��Nd��#8w�N{R+G�6=3�a�\�|W�_�$,�O;:Uar"s���0ƝFX�o��Id�z�P��������C��7*��Q���F��rЍFȏV����M�3ϰ����0�٬/�(F�(���A��Q���%J4xb�p�mu&���yz����'��~�E��������z~{}��Y���PN#��R�^��Q��)�O���f�#�!�f۸�D�������)E�t |�9��M�;@�TJ���ҶwwP����K��l8�C�I\*T�Qf�B��Ji�ۛX[3f;;�������P!���;f"{�� ��,��.H@�,D,7�3����2���$ID�	R�h�m���ͅU��/cu~QN]�T�hR������v�C�R/� �|+�����4*2 =u8F���(�?�d�W*�պ�_@�w��'���L��$|��Y�8�$�GG�����s?�t�&�s���7�����U��!�$h�-BSANC4@!���0�FK��@2����F2���cgc9�yK���"�����6����|���c�d��081���-5{��&{l�Z2{���'�h��}��}�ݾ�����HS�H�5���A�R�ufjR)@�x\���"k�˲��{�LY���*���Qs���#�<bDd�G0;7�b�އ!_(�Mؖ��ܵ��"2� V�J�#<y����lZE��k��j��~�T
���v���Π�/�*rrlpX�4#>ז��N]#?>��PP,���U,o����l���uM�/��簙߶rc��L���2�-�y`�U��),��dg��
��S���60 K���q�<tpj(��܎��[�o�̺����^�D���"�9��C�q K�ސ���ȶ]�l��WH&����҇F��q��!�<~L�`(`��eXB�/�L�;E�σHEԟ*��;'�L��D!`���H����&w�W�>6`&c�pe�51>��~�p��A�Qt�5�Ih��b��*~���2t�����X_:)B|�*>nc��0������J� ��&V93A�(k���H�p��i<u�4�=fǝ������v�,�|t	�/_�fn�V)0���儌M���-�AR����SG�50:���)����������z%�Y^�-�=T�e�I�y��/'EN0�m`"F�\�\��^�a/<�xU}�ׯ��x�g����t��[�x��7���W��t��3��/H��ƑD����B��A�X�(�`�kX�s�i��I-M02�����5�}�׃D:�=��2�P]fx��"�0䞇�����Э7050��?��B6<�YfZ�fn�ul�sb52�m�<;���F�+i})��ni���3�v��H�1�MbrjSG ;֏P:�6�ը!��wP������5�H��vd#H��	��#��B��qОNͣ�u��j�EX_^���i��Éx#��M�4���%���ɘ5ᛱ�)�;�f&5� ���.o�����i�Zx���\ƍ�Yl��s�P'�C"wBπ����;���s�O�c80<���!����SgЫհ����{wM^m8~�H0z(:aj����S��dE��ەK��hY	+��CX�S��q��I�}A,ߟǝ�ױ��(�eH�p�d\�rm���'K�B�B�M~kK���w��!���Z�y�������p PA��������{�kz����%�p+��.�������� �>uJ6H?z�u\���`����We����V�{��&�p ,�MʔM�(S�����w�:vjrh �"L����.��y��PC�H���O�}�<ʢ�-.bk;�	Z�׫�H֤l��M��SH�z�v�7��̡G��߯�Z�Y���u�8p Ǐ����^���*��dM���el����]��Mi�Qkv�a��.Nv6���)���nOt,�j��O&K�e�����IT
3LOL����x��)��@�4��ŉ�\��1�^�&�s�]S4�mӜ)+���m;ʶ�d���M�3��I`���e?K���>��<�.A�G�8��^z	��B��ƴ9�G|l
H�{��wp��Ui�%ݲ#�8%+F�LЯ�1�1���)U�k��*�}���������я����_ʆ�}'N���:�_ӻ��f������K�%A\\^7ӮMܢ��?���x�^�t�O��%��>F�1r`
�3�(3K���V����>�~��������Gy�ԩk�k��G_�&`S읾]�i��0������^I���@�����y��'^�����ח����NٞdFD�����B���n�Q,kyM��}�\L�`�}d�Z���a���]l�,�d"f�8�,�TZ{7�zyC/�����*\�&�fZS��.�{���]lnn`ys;�]9{�+�1;.u�z��K�:1�a��C�V�6�7h"N�#��ġ�����)��Qj\(nJ�����]�a��V�/csi�bCŗ+g/��ii�	�P�t�#7@�g�����uX!�#q�KG�fCE���>�H���:Vs9�5�H�rk�����V�-��x�����?�C��TL�����(����.ݾ����������n�1�=�k�Mຓ���%c~rz/<����Vq��\�q]�9O�<!V4��E�.dO��Z�_��L�r�}�F���=��Y{��;�����*�BQ�[�c�H�;qi�\^{�3�O�(� ��t��^��CڰUm �~pTf�х-N����@`zK+kx����;響
�c��\��aww.��d
�dF?��'�\�>�Μ9���ڏ_S&Q��گ�Y����;��kܹsK�u�|n�VO�=��I�7�M���i�D�ذ јE��^�����٧D*#����]��M�Xmr�--Fjv��dK:��{���:��7U�IxS�m m���i��̅g00<���erlżu��صp�V�E b�<u�tu�3���C��^��a- �v��?�����K>�ԣ��*$��o w�=�,8q��y�<N�<.� ?e����[X��λrt�^T�5ga$�ɍ���p�|*XAE�2&��Iޙ�U�m�
��5	�����?{�4^|�E���a�7�N��4�]Y�����p��e����s{,��N�V��4��e���0ҍ���|:��,�b�s╆ڋp����������3i�7��T�8�%����%�K&l����6�� ~)����v��4���M����A��(�S�(�z�w�j��Q/��w��C[Kˏ.mOiڡU���x8۞�N����$�F�����2�g
!�Y_��������~��O���O���ks��t-�3�����X��8�� b!�W�y~'gL8���k���o�H}_7�ݞq�O�I�Z�
�,��Y&��ER��!�+EMΜ\P�"��a$����T�6���I�Y�ma}'��ZQ}�V)����ͬ4!��T��)����w�b�4����5=6�c����K �E���.��,��xp��kۨ�VQ�4�������Ӽ�Xk��i�	���h�������A����Y!Xޠ�V��$��ew�����=H\`�s�~�������v�jMZe"$\�b	�{��}��$�eK�2FN�����x��U��wVӮ٤�x�d���R�Dv'�"�<_ޤ���#	�=v'������x睷��G*��?ӥ�%,//c����q�앋�|��&5�|�[���Y6\'t�x��i<��y��z��<�q{�-5b^"1��F�I��d� �p��y��e �sc�{�uݗa�������L	�2���H:b�S�''T�>���~�]�������	��^��5�Nr��!��Y��Pp�y�ǯ��+(W���_�5�������/���+�����f�#*�$f�ll�ޝ;�3&�"&� �F�y��ӡ$�T*�'O�oxP��;s�p~�{��H����
>��`� �jFU��)����m���U6=Q�������O=��{�9;��v�����za{�o������Q7�l�}l�Qm�Ԑ9E�Ϯ&;6�6d�v<lНՁ�wͿ�x3{��b��}q��<��gq���#q����m"ރ�9���{x��7���L�r]ڻ�K]�_�S���f:�7)ir\�%;Hs^g�@�q���!C}0I�/|ҵ�T ��z� Þ�f�.]�ի���sV`��R�z@֠fv������yV+����y`17�H�G(�������_�2fL#��)���&��4"^�y ���G��_T���D4�o����DR�ڸl�9Q+ͶBV�De��Gl$����|��"�hú�6�=������8Y;�f���4U�\�d�J���eݞ�Mt�k�_��*/��Н�c�����?�ċ���/�vi��n
��V�X#�,Cq�[��.�l-�EM*�hX{|��th
�k�q�X�L�Ӎ�	��;K}>�����I#5��ha_������Y�����P��v~��]�K�+WɈ):�#�gx������d�Y��.�;m$�>�%��dЗ�`x �h��&*͚L@�
�6rhr<��N�����C�7@��A��D�זg3	���X6,����Ѽ�\�� ��F�XE�RC�Q�{`����=^�
%
n���Xk�F�$#3�=D#x�#ڣ�U����j"��#=2��Ǎ���3��:^�D1��IBW�XBf�¸C'a�:<�	]�$?��V2�œ�p��qd�1��ӟ�o��,�� ��H:E;;NǱhO;"F/�ue�    IDAT��ł�Q6-�m���(HJ~^8��	<{�F���q�2�������'y��C<�Ȃ%�ǝc:���e������?����ð�q����W�u���i�R��UM$��\l$}A�mn��vB�!��&�ɖڜ9sJ��/��Y!z��_~�e��������kW>RAv�}dӞ;sV�.'ҹ�����S���3 �u�R�~�"d������"�]�uU�\[��m��W)?�TH��Ra���L� +@ԿXTnc�v�Zt7j(j�2��Y�1���g�K��EC�	��G��ljrm4��ߝō+W����BW,T�f#���;#K4!毶{����b�WӦ͐v4���2�Ф�����>�O�ۨ�Rc�OgoJ�������
�7��n�\IL4�K'5�p�~�/�pɖ�a�kՆ�_�s|�l����E�����'��ً���ŋH�b&/���N�ٻ�i(�K*ro���]�a�05�.5��bg$Uz��xhmI��f�!����mw�����5�Ĥ)�� 	�Q���ֽ�Sѽz�*���ܻ{u��L��=s��#�����C0��4_~>����<f��&ыPrw�ݪc�[G��B�<�^�~���$�@�I"��"SE�q�"�ms]:�
R����*�Vr���f���'���g_�ċ����_�:{�_��+��2}��U�3� �t#i��ϡv����܇�|E��,�BQ�:�8aq�R����[�來��:��r*��dJD+2�<�;� c�AX�3u����/a����¤$Z2��!�DL�@�W��_��hR�0��W���~/R� R����7���q�[E��J%`w���pB�^�|���N��d;5�5J�1�D�.�3�h�eI<!���^۹=llnc7_��4���fM0t�2���������a�PF�Vq���h�l-7�OB%��������Y�ehj���C������be{[��*	ETO�z�#�l�љ8�ahtx�dBv�^ʅ��M�H�<rs����^�G�/c��Jjj����Çu/l�T���.��ܻ�]���Ϝ×^z3cc�~�c��?RQ '���9�����Ζy��r�>� �����;ylon	�q܁Bf�1�hJֿL���`F����2�߼%"
<B���2���
�ff�v�RO�>��������?ԡ�?��W�*f1�o}���}�:6��up����RnE�isc�[����l��O;v�b���+��ˈ�G�:�C�2=�?���2�p,!�<��cnU K�h�R�;��\]��:�k��W��H�D�C����_�/��sl.�>pZ���UFm^���_��z�bY(�i�K��	�m�${�2;a���5�����2F)���\(A��Sm<Ĺ�x��������������gے���\�v�������.���&���cճHڡ"u[z=2��G�H�i�M|mNlnY"�Q��g/�>��!G)c�i$Z#��S�/_����ks����VD?���ai70�4�����R�)|~}�m�av�r*T4���R:533��~�+������vȊ�T)��_�w61��>���=����eO�j*�Yo�r���P����gB�hT�f8��+B��3��^Ef���*�ݠO;�1���+��G5���9&l0�_�o���� ]��Wc��B2��g(���������������/�����^����ܘ�h,���B�;�j�F[��eպz�Ʉ�u#�B2���׻Vn�O&j�>6ZG{��F�3�G����_:��j�t[x\�d,\�"Hl{+���M��՛h�(�w�M�C���4�p��|�(W��,�
�3���7��<o�v�r4�E�:-1���rB����� �ޒl���Yl�Q��!\�����M}٬�GjG3��8��R&hn#���e,-�aeu��:]�ܦ���$<D�$�`Ba�BA��qk��b�Z$4M�-�VDN���NX�_�K�4�I�?#�<�w.�"��s�D)�!��!�=�!�{�������Т���~.�����	���������4����d���:x��������"c�� 1��S���=~�l�>}�"~�K_������;��_W��d�Ӑ�E�ؓO����I@��80=-�!"�c���$��L�NΔ��n:���"L�I�|n�#�$iq'LM�۷m�˃���&
6�V)�$�ϟ�W~�<󌒯Hv�$�XG~>_��������7�3nߺ���EA�z^!5q,�;��(����Z�OS7�ϲ�#���A$���C"M�fL#C=�#^�m*�X�Q#2��Y7�p7{BB�Ѹ��|�hO�j�T�-o�dJ�N|�3�x��TL�x6f�v�0�����q������X_�B��t��	Lb��+$E�y1�l�t��k�a���b�y���@~5g���U��vf5ߋS�ںq�����4���M�,}z��^a��39;�f�3�%6l4�q�ht�0��=��t���<��y\�pAnTlM�50��q]���dO.},āω�t�$����`�]��v��4+r����ux���5��D�����"�˿��*�1�]XT{Ҙ˜�6����ˆ|����Ѓ��"���G����v�A5�d���)U�e���υB��=4E�jҦ2T!fnr��u��c��&�s���r����"�g�7r_:��lwټSQ��*#�D�>+2?�?��'.��W_s�������)J��빫��w�������^���4bfl��8�]/b]7z<���"�C��B�Y��aR���M�_�}q_�g���/q�ף-dL�^)c{u^�K�2���S]�	C5h�A?�k�=��T�j��Pj�P#�C8�ٹ�@ah�n����o��BAB$��T��(+�G�X���uX�I������aAdCDk�2RN��c��v��B�(�&���K�/��^��@��ɟMG���=X��{����`�fQx�K.�-��S:k14��A��M�W�6.Th�FV��'�^`l{�D�u��T��,�D�n^�:}h�,~&�,Q�1L�R6�1�x�3�/�������l�܈[��<D6xX2ʐ��(�?f$��h4������$���<�iP඄����l�.^�/}��'�7o����lo������&�g�"���q�����BN�t��ye��줟�H�;�fk���o�UT}g��VX����ʪ�r9�qb��I�S	k�o�L�LZ$+�9!��.`|b?|�5a^���: ���o�Ƶ+XZZ���EM��a��D�.s����i1H~4"X:����HO�̈%M�3�09���� ��E��	h�� �A�o�D���ʚ��<]��𚦀�<<8�?q����p���&�������bH�kkaׯ\Ǜ?y+����/����Ҥ�(����C[���:Eٰؑ��c��a����AF"t��܋��3�\D��4��P��xX��� �������?�ll�t�Z��y3oX�]���4"��t�<$N���� �ɏ�����xY�Y��
��V�f�=-'O�}�I8E�7ƻE`���	�X(��������B8,��|�),l|��Xғ�u�m��mG��GM��=�����cV��D�s�b\��OĬ/|�8tx��>��춈���������᭷���ڦ�e��+��s�1�К�C4�nd���7�/te�����"oi��k�����d�x�H ݐ_C� ,�����N3щDU������{�+R�zv�t�����jMx*M������#�}23�=j>�����U�+���׷���B��HĒ802��pB�t��P#��"��Y���#�Mj{��=A�H�+��&��)�@�{r#H��f�2�0� �~s�h��ww��<��"c�Z]�s8W�]��(�*��F�u��\�[d��i,��5����I�C{8ހ�
:�:z���8=��)�A�pY��Ё��E��{���"}e�����#=8��0%1��A��Qk3% {;�o�h/���"*�с��'B0�D(�p��
`���/S�s
$�O�%�(�����mQ�	I����a���ᾄ<�irk�v+�w��N�}9�:>u��^��d��s�ZWv3� 	+ݮn��XX�����nX�c}̮M7��}�5p
�*��;@����v��>�/��ұ(���x�W�|%����|~[/5�J�QJMD:WM����J�$�J䌤�'�UT[g��kX�5Ή��C~�{�s�6���4a�u�2�^����0¡�+����Դ��s��Q�ko�.&)��|�+������˿�6�]���C�}���u��C &)��(Ж����~�%��H���5�M�9�1�G��y��~-./�Gf)?c;��#��w��Q�sG�������1�JFmr��g�ן�S�N������'��$�TÿU�s��z�*~�ڏ�������cA�co�zES8�c7h�^���񽳸�>Ra;X����"O���=0=3��|�Ӹx�i5
z�9�׃����0;aa;W�E���#����#�t�i6h��=���'�p�f�Yِ��,��l�����?��tF�afP������WG_�|E+��~$�C$,��/�L^�x�H�c��GGu�:�=�p(�4D.f�����|}�x���q��A9��M��7]�<z}~p	?}�4X4rH�7�g�#i��W����PQ&JC�7&��W���;a��p��*��xH��,�<#6��=[zx�������b��<%~�����P����吐��5Pp�$���V���ֳ�3��&�����;a~��~�������t�RL2]b�o���Rio��[:4�T�V��h�RQ�O���~ƅ�7�7h�j��ڕ12�N���̯t�Q��5s$y�ۂ�t��Z���~^�(c�^U1�6��%�U�����̂d,u�^K���!�}C� و7x�MC���\���;����=���G�>��/�ofX���l�!dƆ�@���}qx|�t�'�Fy�����/�c��"�Vs���W$Y��|!�I)DRicI�����u����C�c�'�3��M���4�~&d��������JÐ��~7\A}C��#�^���͌�&ev*����Y�vp7�}g7lL h9G�)�P7�Zj'�}�U��W�L�9a�]�CȐ��Tr�w�)�vqWo��.�XA���������֏�W���(z\5ЩHNDѨ���)M��ZM�I>���"��H� �i<����e^�q����@[M^�߯u�T	[J�TLb��������{��r�����h������/����w��||�#��wp��#�y�� �!�_<8Ȭ�{�;)j�i��k����a�M��L�+��_�*�j�$[�%[�˵�C� !��'@!f:�&���6�IH�TL���Nf�$�L � �i @(������V�7ɖdm�������9���J����y�>O��Ⱥ�������=�yρ��0�@�ӻw3�x�	y��cr��%���u�Ra�	Y�}�ml3+a����x*	+J��l�a���[n�W�������
NY�a/Q��2m��E�/��U��_? +:G$D%b�>H���^q��������ܠ�hV����zt�I�w@:$��T��ǈ���9rZ"�G%��O|B����ת�R#;xB]7$�������oT�H� ׋�����%^[-3hAi�햛r]@�#s�.�^?���=��I��׾&�?q��S��f����Y�G��Alxp����p=XH
�~2z�x�+�D�V�����ˡ����cc�Tu�k����ۑf�.{T�q��d~a��H� ��A��o튅j�Z6Ќ��u��E&�8�X�;u�'/�@�8C}�#���]e�uOz�a�*�N}�-E��4m���S����l#1%�2b�����������zރ���w��p�?W����l���BI����7��0�A�o��*|d52oKaA �@%�����,�0�,<h9b�U���QV�&��&K�K�R2B��k������A]�&ҁ�Z]��Q��-)�j&�q	�@gYY*���8������\3�aH/�Pp;��$җ�J��Ȁ��^���f$�bFzK����,�R��MCb�'N:��mJe�"�s+2?� W/]�k��Ҭ�x���+N�W2�^q{�-�{��Q$ϣ<%`��1;�E�fr�|��!�� �(�2�pn��l6x8c�	�d-)����V�;WVe�Yc����j+�*�
$.���'�w-7����c)�|1��4��q!��Js���1���0�J�����+��l3�-VKB��j�?��W�%p�+��?�9q�鴄^��P�0�GI"�ӻ��S�Ƶ��O� �Z�G�J'��d�) �f�v��ՙ@ҽAx
� ��B���D�*�\����)H.\�@a�[o����Xр�V��^�:�mq`~������=Ġ;�c�<�u$��@H�~C������`%��5YV�U%m%+T����<� ����� M��`�羑���yp�L�DS@ ,W8�nv� �]��B��z����w}����d�Q�"�+bV����������/�>�k'�#n�@>@�i�-T�ZB� qW�[��G�AK��y`a�vO�oaa٨4��f���S^��C�}r�E�`���� b��sK\G���5*Ciέ�o9V{�Ng��9G��u����5�K��W,i�#8$kUV޵j����]�\��u`䀴
�Z��kw��ӧ��ѣ���Ӽ�b��Y��j�_1 mT�`u�@H����s��XW�S�U1�^�Ѫ�8>��Yב�u��	Ȗq�5ʆ`�:��D������#I���k�sި�UX@�\��Q8��mޓ�z��H��~GfV��ނd��.��6�hX��� �Rtf�(��I�R��p-H��`1���{1^h��K����nyס���|ރ���G�Փ�����Z�T��Q�(0��lQ���HוF�������q�2އ�z��e�΅!�i�;�*O96��D�'�t]�%���hT$naD������dq�m�����~$62��^���ȸ����ŗ���#�c ��R�P���A8HI&�[�"�cKy�I_1#�c2��lٹU������@pDTH++�t.^����ȕ+�R�0 S��E)a`0(�R�8�^	@���-�
w)K	�οa��lp��Joi@J��	"hCD��nK�ӖryUY��?H$�_�������ڊ\[[�J�)&�)�fr���&fI�`A���V�5pA#�	T5)R� �B@�K8��諩Q5��n=�_�?L�`�Z <vV����+�~���W� �Q�����!�Zo���dc�@��ò��6n��Y/^e`��\�PT��
�L�V�'�C�A��		{�L��%���Q��X��Ͼz�*��/}1gi�VFE� �p�0�t@�����ʃ>@q �o$�Lt��AP�X
K�w��S'T)xfx@� ��v�Y���ߒG�8!Ϝ?��D��!�!zrt����%��
��Z�E��tZ>�=�� Ÿ�y���N�~�!ʇ�*��7<�:���z�Iy�cr�cO��p�C%��Jr]w ��Q�\1�dbj���QaS"�ܐV�z�N���+5Y����I����n����%�_�0h�kՔr�Bb��������E�<T���7�4��V4m A��D+\#GB "܇x�9���5�x���'�F�(C&�Ң�Yc#���Ũ$a�'?�NWN�=�9��'� �	p4�0�@����f/#yo���3k3�CСXԹ��t.>u����{��w�)7߲_&'��D�㓉��*@}miQ~�ay��#�\���9�\��7�>㚍	W#b�@#��6��;J    IDAT���m[�ot�:觯\��ZY�R�G���)d���c�c����p�ԕV�)H^�J�B�;�CWLx�BN�e·���zWoٲ�?���7OL(�g�zNp�o���9s��*�j}�Y�?5-�vF�n�@Ŭ��!�-��a�_���V3	��s�d������t�@�E;�xP��t�ff*�X��
GQ�g����~S����D^G�x:m����yenAj`G�:��-����ӫFK�Xڀ�;�۬�������a1ef��D��q�c$�?kJ�Rl�g�c�둩�mr����"=�"C�j�&@�,/-1�._���k�2��$���4;���-`��K��+�B����t"��V�}�ѕ66�a����pm1�/�f�LNy�"�F/����ģV�J&�G����͒�Z4��U���a��l�.L���-�1�&�ꂖ~���;D��Z�?f��*}n�G^���]�9nD�1_exO6&]Δ���9s�6�)�0�T�W���_�jټiD�����׿�e��
 �% �u�ّ�C�,z�b�F��⽩Ċ}
-����A$:���~qʜ�c��6��yM�z��P�YtF�z'��!�~�w��~资����X02�*A㗿�ey�駨[��Z�����~�Ǎ�������#���}j�3ۏ�8.��x��8~6	9hÀp�D6���b/e+�s[F�@��B_�y�,����k�嵯y��-��@b��!����O3?t�C��R�L�(��l�����U��)��*���G��ZF��a(�1�[�$2��h��d�z��}$@톓��S��xݗ���s���:����*{�	`Z:e�R
��W뎤+"oJN�����2Y�+�o�.�#��p�q:$١��^�'�b0Q:��o}KN�>���|���K6�^��t�J��z��Nd����)5C$��,�2RȫF�!�F<��n;x��yQ��h�m�~��	��IH�¤�4�HcE.T$: i7��]��Мf�לB�[�t7:,�k�ryyAf�KC����z�M��?F� ��@��]#nJ)Q�"Iʂ�=���4I�~N���R�Lt���~�����jpY��z=� ��{?��S/�A�^�E_n��n:�aBפqd��Ut���xCgf��e��N3j��) Nv�	�Q���.�e�� s�$�>4��`���$����:�4R�����5�30����$�ۧ�_�&A�����識]�LU,uln_�+���%f��`H��X��Hш$'E)0�b����عU6m��/*��E'���ۻt���]�"��5�WZRE��s�W�B���Z±a��Vo�
�%���C=��]�^��o 5X\L�w�7i���v$�p���Cq�oErT�\���[5i������!	.4b�,f�<x��6N: ������%ͬh���"ц��u"TڇUU0�� 5g+�L�ʘ�R$��m�P��Ҙ�y�+erb�<����_�O��Y����r�RJ<�Ԫ�!��Q�橤��W���Pc�����7�����+�hQ�� V�$������NB��z��{� �讻H`�ܺM��巾%����~5���H�ʕYN�����D�(�,
�x���'��.T;�|��U#a}2�i�j_8�!+����*��ǽAr�ML[���9Ͼm�f�q G�'\ʳ��*����z�+�5��A��X6;��	q�B�����c��o��MY]�J��_z9�d"8�����W��:4U�c%ՓO��p��d`
�>�J �
����z@F�	����(�1�TD�O���JAx��Qt<3+(pqNX��ྥU.Зjm�p,*;$´r�ȴ��Q%�9�2�ρ�0{�X�a$�%2�wNNqL	Hu�i��T�H|z�MP��  �
j���հ4��iO��d�Zf��F�]Z*�u��"F=�DV&4�0�P�yٿou�'�mU��P�3� �!�g'��Z�L��`�ox$Z�gfe�� ���%�*w��#�7<�3kf��\X�� ���=҈|�]E��9�XP�VS�!�9��O�|�^�3$ꠝ��k�y �0Ȧ�Ȕa���7:�ǷN���7���<�����l�[�o|��������+7�=88���#��A�Ili�-QKs�X��ʖ�1.*��\����U%����۫Rx���l���Y>,:B� MaF�ݒ�+�Ҭ��,�de ��h�~W�pE��*�Wgeu~�Tr!�C�GF����
�֨KymM� ��[쩂,�4T��7��Ċ�#�&}h1�ԗ�K��0�
�U�<F�2�4T�ɉ�2�}�l�<*�����#�	���̌\xZ���i��tR�$=#����ߴ��,�U��� �knv8�>1��l�!���Eu�]�Vu�{9�z	��σ3��@,J��+�%��Q�Z�-!�Kͨ%Z���F�58x�!8R^U�q�E=�V��URdW�WXat�bW�
�#�!�恦*a����p G"Y�|A^v�]r��C�zZ.�{Z�����'�<!��$� ֚f���Ce�7������x���S��.� Z�^���9f�g0��Lb�_W�A�E?+e���*3d��'�@�:x�~�'G�|�	B�Wfg���[�����e1 'j{>�lUҀ{��@G�V�U�Ið�l����*M9��+- �o=p?�p:������g�
-�B�+d�4 ;��ț@%�D��^~?Hx`�c��Uw?Y���3�#$A]���*����Y~�ޯ�Z�.�b�K��@��&���h��X%b0i������,S���cֆ;+��*hsFݐ��ۨ}�o�.VTx�\)�ȩc�Y���g��*�S޺NV%����| �Mq��Wdye��� �MV���n�d%�^ɻ.�)��s;����,S���X��R.������f�t�l`ps���"<���8jr�.�R��t&ڎ�qc��$hs���uHP�=�l��;dzǤl�:�m�g�������������E��Ş�꥓<-�0�j�&��4>A���\����
�xH�'W�Krf������c5��MI�b��J-K�l�ܧ8�P<h�o�d�Q�'i���CA8F.�{F��r�ض_��&v�?۰�W�I�������3�/��r�^��XvN��M���\��b֦|����t��	><d@W�H�yG����U��|8F�0`̮�U������9��S��M�ٵA�puaAVg.Jcu�F����
}dh��DV��>�"T�]��Q��p����=��p�����ood��3@��D���H��H1��@_����@I2Yh��҅D�ߖz��B��J���qhI6�'��+��
E	����H*-��)7�� d�"\Qr�Lq�C�#G�� #F����#t�Ƹ�jY�^���+}�}$n�`�w3Ʃ��CC{��@+'Y"+�	z��,��
�X>�`��B�$1\��p}�7����Z�k��B��H&0*�W*��J�0�����!(`9�[o��_rHn?xu�1G{����47�BZ��N�~ ��<�s����q)A�L^-��n�(T,Ӵ�ş���H�#�Ԃ��POB%��t0��Bf.���)����³�g�!4��dH�u,s
C i�zux6�/G�p/(r�U%3��|$z��7��������9G� �+5<+-����oߺ�����N0C�9y3��y���8��}/y����Ioo��/�g���ZBU��w��%9����}]ʕ�Z��#�;n�R$Jr�v���29+&?<�q��ύ�� Ǒ Cy��b;&?�a�zT�\��� cX�u|��/Pޔ*o);zC%��>�}��EY*UeyɖI�Z��&��E^#� }}��,B�3�yշ޾u��J�����H{�QB��'OS���Y��u^d�U�W3��5��x&at/�~TR��z|�^O5ң�
�@ ���˖�����m[&������!�l�����/\�!�{g?ʔsVʉ4���y��� ���D�?�g@v`82�iX�^[fW婙���Hio��8��LX�VMF�:�փ.n�`
�%�������$�ML�A7��́-;~�m�S��o��#��K�~g��(��PF7���歲�X�f�%$RLZ١7�c�vj�"KE�Cc8?��$*�&���H�&�""{uaaN.\|F��:�80b!�ѭ�e�3đlBVY�M��< ���UY�vM�����pEǲ(h���>�ApR���M�}���E0wu� !M���<67�([���*���ltۄ 1��H$�g@�l������o͏�
��V[�����M%��͊ED�M@�j~U- h���W} *cs�}U� ���Ijs�C�*&'�a��E���A��Kg��Y ?+���`��(��T�}^�'�����bI�Gt�cG���s'���"� �WJU|OV��{ހ]!�D޿��ɫ��n��ҩ7����2;s�kOU�*��X�v�y
A��7�c~S�Nu�M�%*1 �UY��hEHM����z��i�>���� Z�
&��S������y�}��S�<M�2ƙ���P4����K6?�/�#��1*6��5d����K�Z�;"�R\�:M� Y�v����?������$�z$�$�V1��j�E&�6��90E�x�K�C6QJc`�V��*�����|�|�[��j�Α;��W�\�뜕��� 2���ϐ< ���8%֡(U�><�p�����b5���3==��A�"-�:�ˀ �����5��c����G�D�T�Fr�� ~hp6Wϑ��@B�� �vT_8CcV�@�rY�[�,��6q$(O��4�R�#؟9���}�i�2;'v.#\��sY��Q��ӦQ
�v��#�:SZ�k+��pO�҄=���2�
���ϋyٳsZv��� ��ʢ��\�W�r��S��y�?�{���_T���'D�4i��W2��+���&�(�BeU./���ks�E[���>?���r`{Մ��
n^��D�y�ga|���>� ��-����.$���vzl�z��=��� Ŭ���/]~�b��kD�̝��mhT�՚8^$v�g�x|`H��e��������ua�7*SL��Y
g�Y;}hV* .�K�Z��k�+c�7���(I�%�JY�^�>Ӑm�r�A0W!H��H�RU�	�+L�|��3�rռbu��@�"6= f�8@�{M �����2\�H>c����z]�p�MV��%��H ��!�Q�LOI;+u?��zKV������Rmu��=H"^�׋5:ל�8�X�O�s�
�U)��Sz�
�I\�A�MB�g�������Re�9n�,�|tN٢i%��Q9^�n�}#�V�.�cիTN(�NqyPZ�e��;C��u�=���c6,����eS�_u���W�R��%�P5�P'!;�ٲ�G��h\��|fz�D-5��z�i5�$1���ͬ*a���5S�
1*)� ��)H4�d����������]"�f��׎~���[�n�t�8\�[d�Hv GS�LLP����ʗ�C͜f �i<��B�ZW�xv���1��ejw1��Tp� mt� ��qn��x죣r
`�ޕf��*3���=r���r��e��1�ύf��5iV�v��<��r���Z�EV���J2��,�<܃�.j�Z���h5�0	���	+b���H��9"�	fn�	tƱej�$+�];�$��-������p�v��~����ߥ7�JL5c]��q��<aX�c�z!�s?c�~˚������nE�_w�`^� �^!�1#u�]��������+�j �'[��X�XHP�Nk&A��,`B�!X�7�K�0�	ԅ�� $���$���~���d�OMNR ���XJ��i�y���䙳�R�����Q6$�tqR^� �*�K��P1;J����[���̵y���(�ՊDYE��ș�=z1SZSBL亁+^�5�{$�)MR�1��k,�E�-�S������7���yL>i����/��4�k�z���vd��&��3�H�N(/ <=���P���0������Q�q�i���Ք�å�	| d���j�n4+k+���$�{�O�%Ԋ�5)D�L��ȶR����d�D�����t��т5~h�����/����a�&|``�r.� �4H"q�{
x��,<@�k��� � ���Q*I�W ��`P沜��D��h�M�,��!�Z	"�qM2[�jӢ`$����tS�>��i��"5_p��V�:��^U	�=;"3Tګi�H�UX�Q 	{gZ��b8:�g��wR�)�lNt�D���� t�5L�Ϡ���	FT����h�`�#CW��J���>TZ��a��3�W���ԏ>�k��LG	�lp�I�͔�(��]kaS��ٔN[ap���*�T���;�{<r��Iq�;�g8t�~aj萣ʁ!:������0�H�� ���W��Sg؛��+G�T�UUZu�TJsʃ}X(�1	�NaD.to��o�c�Ki_h,"��f�����E"�����$�vL��9bP0����*uv1���������Ėq�DI��1���;{iV}��<��q�a�=[$/u�e�������+�	�Z@��H�
P�z��c%
�@?ۆ^���~�`��t`���=-=`�C���J��?�A�ر�i,���d�,F�"؊�*�Cc����A�\��O��E5R��7�<���^�c��аLm�*w�~�l۬��|&��I��� ��~��I9s�izCc����:#�sj)�B��Ң(e)cM��y�jU<F�0I��P�jئN�K�Sn9x��ܱ�#}��l���钠��#����S2�{W.��F������PgT"K*�hE�2>���6hQ`���nJ&48c���q�ƸF���H�ғ�)�	Xx.L��S�-�#��K�x�Н��!EӁPUes��Ϧz����������|��O]����z��5��0�+�v �0��b?��3��)�,p�i�B%�DBe��A��#���XB#��K����e��c� ��O��I&e���d_���CPoJ{�*^�M�mT8��`��NJ��K���AHh�*�A0�q�!ӄ
��$$p� �̊�p*e��,X�h����� /9��V`[҅~j�-kݎTڰ��
ܨ�H  �Ǩ��5��(9�@���P��"ԕ$gr53�8�2z�Ȁ!��*e�^Pݚ"m;�L6k�&D�%X�8|�W��D\�����-���p��*T��rA�F�����fP��I����{`��D\?L0(�	�h����,��Ƿ�In޳O�MM�-���UT���8�������A��!�s�'|E�Qp�� �{�,aq-F�lZ_�o
�C;b/�q�
��
��h^mY�K�|�DhB�N@J��6Ǟ����9j�O�sc掃�k?`�sz�|��lC�.��A��`��<�WJ�1����<�d$5��쬌o�}�v+�ɪ�d�ZY�V�Nq�RO��z�ٿk���m����X!�z��K���G�z�C�Q;��b��u��Ġ��Mb��^�PGá��t�b
C�j�������{�0�z�A9x`��z{h��A� �bq����1���Y��W���k�2��Y(H6���,./&��8����d�����s�/���w� �ͩ��;�b�>:iM0$b�Ԕ��%�VSN>yV=���=��4�'�H��h(�>�_�����|�p�N�� �kù��q G3������9j3����q��r� QQ��la� �D�s�'��0F����۔0�3K�����K*�A�c�@�V7���ז�6iJB��T���>��6�"f���Q�SO{����3	ׁ��1@D:jH��;=f��L�]?�����m �y��|3����/x�tb���,uZ�V�m�y��������&��$��: 6�Y�    IDAT�x�YY[2�<+�RQ��#�=f��w�X=�}gݾYjey���2��H���+�c,�<�KS���d���bחb7�Ֆ�ِ~�AH"R,j8ZYk�ey�%�NH��+`=�������/23-��IOĨА�����%F7����+�C����Ƒ,�k��Z�5D0ZFDMS*�p;��4ɀ8�������d\E*B_�R�jS�`�nH4VaZGc@h�+�4�ܕ���@�-<�R"f�� �Tg�i��yKX�E��7�)�٦� ~@��B-A����2�P�hM���sڑ�3��"�(���W��X������&(�4�TAϊ٩Ƭ 7#ت�[�|����t`M�R�փ.�HT��е~p�B�8�*)����j���o�?c_,w�?,��a�H�	��R0!�p2���N���g�!�ĥY�+ L&���V|*��/����� r���=�)�L�;��/�X�J�%;�z򐮄���@?Ek ����/�j�)Gff��c�?!{T�eJ��z���p�`�#i �ι�n�ɋ�gfٿ�duЩ^&��ɨ���)�p��.���[��n��c1XXKvb�Ѵ)���O�W��5��M%��;U�:�l�d����H��ΕV]�ol���'�5�R�@U:��}%�z�LMMI��H4NoE̲�Y�'?��3��1(C����+[$����Y�,�S���z�^��w�����S� m\���^^ i���̴4G�I�	�HB�|v~A���0qa�Y�.IT���\�����5���F]9��-O�q$�`]cv-Z���վHQ-a��H�ya���������4��c״'��nl��b�r��nA���=�� �|}�A=�����]��E��Y��m6+#�z�!/�ER�c)�"�ZK
�3π�Č�'����X�=P�*Wm�]A�8�8cR%�ڲ�mȕ��,����: ����ϰdߦq�Y�Bۗb�+n�+YT���ݎ4;M�)T�k�TY�%`���P=0�].Lm�%ʨ��ze��F�(�=��6!#E� �V$dH�fH���Z-)C>�ِ�v��m8� Nr�W��n��+�� "�n]CE�*��F2�kx�kЂ��Db{��k�E@W���<HVOQ��P1X��[��
��nDQ±��¬�e�K� ��Y��J�沯�f�UN��*��A8(���s�>2vm��|�H�4�X^7���66T��խ�f��S(�C��}� �^��
׼~p�kf�)�]9H�#R�<(��m&Q���~�B 8A4�e���P49����i���"h�$4T>��� �d��P��(���4p#p�׍�VA,f/>g�2�Wb�q�p���3��pɰХ��[o����"���IL�/5����ȥ˳�У��7xH�VY�!1����ډ(esӃ�3�Z\CW,�5#Y�+u��Z���X��ic���r���:8�'p���{b��ܜ�:}���h��_ H�B�04���m.${ZZ���p�p_��3�Ԭ�le��Q�A� s�/���ܾUJ�>1�6��;�:�8��e9��Sr�Ҍb�#xQ�D��������� �G�ք�I`�@P��p�P�R&���N�d��I�D�z�h��L �_�Td�PK�я�gT�'��ty�(�z�d3L� �@����8��I�
X�V9��RM�8L��s|�0�b[]�0=1L�4ͮi�m˲�b�P�P�X���-�l��+q�����җ>k���s�Y��m���_���ً���r�+��(�n�a���ё)�0�R�H����? ��N��h�	[��A�؇h4��XBd3=y��h(p�Q�K��+	9��=�-��#�n�.S��b�k�Ԛ��z�L�jK�U��ZY�W���>s�F%-�7%�Q&χ���6�U��G�s:��C7�E��1p��G/k` �J���4dcQ�2��&GV�
ʷb	S)\i�,N�E\5j�7� ����_�NK��X�M��I?)�[M{LX�j3�t_n�|�A'y*5����d�����Bt��u��^_(i�4�QL���ՙ'�:��_ϼكՕ5�A'��ԇ'��8:9"&.��ŧ���V�^>��4� ��@�V�J�T)H!�H����)�͘�U-�`i��<��{���*���L/�}),�3vݍ	/�NM���[W����lثׁ��e���<���}�����������~�t��8��Ĩ���
y��ѾADH`c�lR��G���-�һ^$�6�S�TB<'�Q�0d22{eN�=v\x�QYXU�%���5A�����p*'4����p(B0��w �1���A8m��s��{Ӿ���>)��Rꅢ�����-� ]�|EI��,St#5�7�Ɂ@�S�;E7�r`R�EE(�B+Uh���+�<)Z�u��r�YxXk�~�Ͳ}\��額u$//�	��\����/1S���H&��K!b�mi囎�qAK���RZ=r�(gl��ЪS-:L���:���;��z�Kh;\ge/U+����V`�W���g�&[)��q.y�q�8w�(�3+��)Ɩ� ᇑ�E�4lӎaĞiY]C�iX׵�f,]1��'k�i�MC���D,߲�Xvm��$��ˊ�@`�v���(���r6�y�+T�x���{��W>�oO\��׺�BՈ�>��<GE0��g��c����P�/q�K�gdǩ�N��j�P �f��
��1&�s�a�Rn7d�Q�7/z1A�+n7��lQn�>)�=}bU��6Z��)�&�W���܌�\���ZEÒR��/ȫQ),b0��z�lw��~�+u��A��<t�A������ ���r���@60'2u�a��q8b�(��=	]��ޯ�\�1�&&���?���\�V��m���d;e�*e&�� �E�͝Zu���=�9:�di�x}�A�Vl�TY��5����蓫5�wZ)�}��n���!�8\? �j([}��������t��)EI���Bz<�@Nkj^ξ��G)4Mt��v�+���y����H�E���dH���[_9���$+8�lx����?µ������­©�nj^O]k]����P^:��,#a �I�וt�`h����PB���J��ID�)$�轻�� ������$��.��Ӕ7�:>�9\��0�)�X,����S�屓��X�၍�`mw�6��7��D�4�����ڱ�� ��	!	��ϲ��>1���#��y��Q	�A�_�x�V��O�תf�J� Q &!�ӧl��t�12��z���T�1���i`KH@��o�s��d`��I8+Q�32�/^�"/^��/#�B�6)���$)���iR��ϴ
f�V����-""��2)e�}�f*fad	�LڒQք1���ʪ,,��}��Wl�rs��f�q���ܕEQ�q'�����ZEu��۶a��ql���g'��EQ+q��i���FbZk�Dkb��m7L��l���ذ�ؑ$r�$��,�;#��[�l�E�o��9�_����Փ���b��[�}�0�˲�d������Ȁ�J10$$���`¡��`L #�������*�
H�!M�+�c�o�[������n�Z�m�Ɔ��3�Y�J��R�b��])���eY����ʒ�kel���<\>��H3H��8�@$T�0o����6lF?־^�� ~��A��(*���!h�\B72Q��V�?�8 �B��iy4n��C���=y`Ce�1)Vz
�S0�
�)�"5(@��Щ��s�dA��K�!+e�����C/���W�ER@OE�H�3�4�z@�I��F�L�u+=eU�)���҃)�M�i]�]��1{=+F�Q��H��t?��^i��U�f������!l��CK�aT<����@��\'f��d��	piO����(:�hZ����AO__g*�������������[��� �&�!n��AW���8��]�R�E')�*��F�AXM��C%E�`����#qѐ0�֫$�7'�7����v�<2J(:�� <?8�Z,�Z�&O]�$�N���!��� ��B�q�/�����U	�gC�M��H�H��a��eA�{�n�(�1�i���}}
�`F�n8��o�%X�6��5����G��{W�P��I�C^c
���{�pו�6��g��8��<�`�Ax��V���g�2`r�<�.]�� �2{u���c��#qg�2��0��i��i��a����0�8���$1����U�#K(
8o��bA�2��|!�X(fAh#�j�+��}py �tuy�J�CA�gF���b��6�B0���$Y��h6��k��sF!��|N(���׶o'ۏ�Q�$ΗJ�J�������\�ޘ��Y��_����r�ʅ?^���5	���:8M����ۋ$%R��t.1$�I-��2�t)�eW�� �z���}#a/�h4�fG\ϔldI^�><${G�eK�G���U�|iV.>#�W�H�w�����߯���+C��u�VVde�"�F�f�p\"�be؋-�Uo��6G�u�tpDi�R�"����6�>�]���I�O���y0�����INM���@+��S�H5J��gu�T��l�ཱ�LE�XGUw)��h(��*��ϑ=a�B!� ��=Ĵ���;z��`��4��s�K\����v��%%1�>�V)K�֫2�5A(�P���ji�z[	c`���@���}��6�%`�þU���f�J��:Q�J:`T���J�9�E�M!8��WC�@nF*(s��Y@&Ԥ0K�{�d�c]�P�H&��u/�_�(�d;g��������F��X�*'3K?3]��t�RY��{��d�!~���J��� 	��l�^ed��O&�F�!����fl&��#�,!�L��tIx�Qa$°��h�^o�mF%�N�ـ��ϊ�_ʍ��	�h��l��@x�w��KC�u�'��a>6�v�I������ |��.�U�f��9M(6G�`b��Q�xa5�(�DQDn۱I��5�j9�a��i�͐�Ү�!��XI����z�PL�6��As��$�IL��@p=aF.�?�_/����$��İ�b#�l{�rl7�� �-�q۶�cYa�~ 
SA�4-�F,Y�!Q�$θ���q\�0�n�S�8����-�o���~ ��BA"m�u��V��$a��&K++�R��g�'{��>�Y�w���5'k�f7��}��ް��Fލ��*�{��9y��W}o�m&�8��-jX�{�93�I�+�X��Q�X$b�a�AfA��� G2"�=��x ^�uo�'����A�Qd��$$}�q"c}%�=6.���2 ÂZU.?yZ:�I:-)�s���_�z�����do�Κ�\mб#¡n9$����4D����A�W��^�ГZ�)�����U��i��6��ɾp���W�U�@ "�z~�}��0��a걉
ZWE hQ�P)��T�
��J׉6�ᜒqt$D浖gCU�yE�<tc�R�* �]�k��q���x����������u���LBT*c��1�������z`O+bt��윣6�����U�5��@������6>O�����8l�����*g-?Ib�%RAW1/��0�"h�Z��*tB�� g��c�\���]�8���?�|���6֯W��~�^�1��{O�nM�K+�t�x��i^�4�%;A�P5�˪[�z*b���L�lz��q��F�����,���d���>B�[�a��H\X�I��qBy�!�Οg%\i�9��`.�H TC�!+5qH��F�>�� L(_W��b�z;�Q�3��g3�0*a|�V��G�r�7X����Sg�[��}���A�t��3s(��>4C3��0�G�_��p���Nd۱�Nl�Nb��$2�v�,��7,k�4���#�&��؎�M�8c$Q.�Ɍ���o����^$8���$�0Ƶ�=u�}����=�V.t:�hxx�Yq�0�ضm�[(7�QǶ�|���F!������g[�e��iők�nd�A`Ʈk؆���Y�k�<3�ǵ&6�~d��]�nj�6�dikc�͆R�Z�փ�J���K�~�K��Ե������)��K��'g�d-�lC܂��F�`��$� ����Xp)�#K��i�`���I�d�+YXj>VhV x�����d�����۾�>�JI�ٮ�{d2t���ui/-I�ۮ##���
��QH7���2�C�W�Rm�ă|!�T�nNJ��J��K�h4�E�}_@�Уi7<}��.�$���HhanM�:` l��!��1 �Z��9��7V\�`��W����(�� �g�)���د� �����&
!���� 6��CXgL"
 �f�	�W��@��ΐ���:L|=��}t ��}�+eUE�0o
w�
j���_'g�s�N��i���d�(��J5�#k�I�(�-����:�7�<A�W'i%�����(�^��N+̍�iʦƟ�
Z����n�@%�"�� C��	��f���*ɹل��b�>�����j��N7F r�؟	�a��a�I!�3����@T�f�P�4"��8��(�#�l��@n qB	^2�ˊ*�@�cC���N��iu[k��_�-�)I�Cɹno)_�7\�����m�9�B��p��"��~�iy��R㌫)�a���1�u306Ϋ���+����9���I�J��!Fմ�eY�r�v��RO���-c�ݻw��P�:��ksb�pty��:w�O����B߅��?p\����ÇI�8r�@{���o��w�0�;���q3�<ǈ�m���m|�w����;��B[:��}"�j�g�^=u�����<���9R{��������ã�}?}`���2�m{	�|�T.�ݐ��ީ֚�����WZ��~�#)����{�?� �����g?�������r�d��=��R��(�&C�$%�(L&:Ծ嬟r���jV/
���#�Jb���bu���{,[
`Cz��x�5�<�'�2 �G�"�5[^]�P��>Q�W�lN
��
-��{Q���Zi��(R�b�~56:-�:I�"檮H3W8=�1P� ��ԕJ
��?�aZ��h8�a92}m��5�b�	�+`�t�Uy:���Y!��3��(0�!=ͲNGuTE{��<=����l��(��t>sc KG�p�i��tvr�^��F�����u�x;�d�T�KdԪ��\��p�DqlYVdF�A�q�Fkr�?���l4�E^��>�|����o�fbFlFb�f�D��8�L3f�db�u#�2#ׅ����@5,P�݌�0�?�</�汉�o[60�$�f�.b�q�	L�B��yA7J?���:�vXO���d,ò�l�qr��i;�'DV�@(�mB+2���nl�~DÈ�$��8�-�N�c*��#�.*K#ä��FM��z�O,+,t�q��/��@M���;��~a���?�oz7�,��
�U��2�ku9yF�=vB�����ja5��*^Ek2�}> �b��W��R]KZ�i\�S'gC?��Ī��c�0
��7��a���oڽ{����#��C�� ���ry�k���O>�;����?r��ܫ_����C?q�]w�{��d	�J襧I�M1�Zp�[>�ē�;y�����/�u#��k_��ޭSC��gz������� @�	׃ ��	�yҺ~�Z�|pq~�7��г�����F��s
����l��T�?���<xd��Rjc)�O 6L(�vzVQ�")d3�u���1l���!_͢��Vߣ
���y5���`�%f�#��%��K2��+#�W���P���[�g� ���+�|���g������v�ZoH���  �79��##���@��JqE��`�"<���ɍ02�۴Z[g��9Q�}U�6m��k
s�S�B@ F�r���.]`g�$�کt3�B���@�I)�D��p�}ɺ�@�@�Ң!<��E�*0��[    IDAT�G%���b�fP�R	z�6�ㄭ'T�`�n|Eq�a���0�"?Toj�)b�h&��Ab$�e��i��m�!�`��{!P��D�a�Q�N��n5ڡv�(�"?l�nP*�z�8v� ������Z�U_nךK��[��^a�ŠrF�*iA N�Ȋ#H�Ȋ+�]�1���&�c��0I";�c��e&��QB����^'LZF�v�0��4�r�'�s��-�&#+#�B��1559rd����>N���;t�P�����5���N�t�=���h��B!/�vG._����|@.���r����7�(B��� 	���#�	�����hEQ�D������y��x��G�2��#���|�7Ƕl��]��i��}���џ� TR� �1�����Ǟx����W��#G���E�߇����s�y���7�v����ΝS����Y僘E��Nb!�an~n���ӿ��Z�ώ~��j�>ϯ׿��=�v�|�];����pH'$Eq��VE�:;��W��?�8��>��/=ϗ�]��S��O�s��"�_�v��(��T@<�i������Ԕ ֻ{I�95g�#$�*@���Y�xp�d��y3f@ajb]��1�����I�����Q;AW,TǍ�4kU�9���*�K���ĖC(�Ro	�`�C٥5/$ hܹ�t�:+��c@��R�EP�D�<}�Z�h������eUդ��C��!�_j���< ��.�a�v̶���H�0L E�����d�|>oerY�qh� :��$�M�NȁL�������f�^��~��~P1��9�����u3�i0!���U=�	P�8��0P�u:�4L��P�-�5���՜�gE�����j�ڝ���h�	
�.C�8F,}��Ac	p�3~�N̸�b��a��[��fԣ�LT��8t�؉3q��b7
�����n�f�I�ٌg��dde�l���ˋ?��Dg�	垿3U�]�ɿ�.��ٟ��ݻs���NO�R6���6����љ�yy�أ���Krm��X溕���>LV���S���V3ʭ*���$��y�:��='z��ѣ���t��wۛ6�izώ_ݿ�-����7��&��8�`\��n~nq��S'���j�72�y�[���7�r��عsr��1�'�h��--ז�Ν{�=�f�Ф��{���?ݳ}���w���3c�Fa��@� b+���w)/+յ�̮,�ڧ?�����ھ��s
��@�O�f�ȋ^�TF��X�bf�$�DAd����ߧ�=��Z$�A7Є-l�m�RG@��P�9E�A����-Lь���k�q��mw �w'��d|�_��[�]��o�9��E�2V�V��~I����JjYP�Egws���B#�c(�qǉ���0�01�@��|? ��e��u,+�ضoZv`���A��i��i����� ��@��P~�q�*��iZ��8�l�0\˵m׵|ov���r���y'���;�2-È��"\��q�~�����N�_	�Cq?0����f�~^&�8��fb�mbҾ�I;��Ј��ءaU�����������v�b>oD���^���wu�2++�\.�l�t���ğ�*0�G�>�����om�������;�`��}����Hb d�( A��h���Uy���ev~�Z�ڬ�a'I2�1��hy��w��2���=yB F������֑�����G�~[q����?�c�ԯؿ�GFȎnCq/T�&�0*�k�K�Μ�͑���s�=Ǽ�ׇ��?����}2�}r'*a�0!����n�,./-�=w�߬��4e?�&"���n�����?�yt~aU	+8��n�V��?_^l��8��d���O��7v�=�L'�9b怑�Q��q���V;q��Q^<f�B�!��"�C}�c0����%v8��J���6 t�~�L�^��t;�V��w��$�H{�|q����knݷg�h	J^����$ݶ��$�.��`@S�#Q��5�	6[��6�Ql��3������l۩5��z��Vkt;+�c4��Œ�)v-1�GI=
��$�r���q�%��Vێٶ�@R'vP�Y ҤmY��yqӶ��HP�6r�8�hĮ�&�2�1�[N����M>�@D�==�`�?~<�Ç��WV���9�;<l�{� 0а+v"���Sv��H-�����?bi��O_�����-o��=;����NnU�"L�`�ĩX���:/�=~�:wm��f�uΰ��(���p�e���Y��%A�� �<j3��v��ۭO�ڝO���/}���Ѽ�o�mjr�?���[Fǆh9	�cX"����k�dy��|�ܙ{��G��F�7��-/޻��&&6�U�{;��Q	�_[X9}��{����|��u���,�G4?>��v����[7�;��Ƹ������ ��x~�������>��>�������s%��?�=_��]�z5�K�l�� p� �jݮ��zq�����4�q"C�:ɣ+]�+���u"�ۅ�Zd8�cDQdt"�:�ԍ��;����`S�"��:ݮ�8�U(�m~��7�����@_l�f�:�	6�ﱑ	64��AU�)Wk��v����r#��ӞE�,�-'�3�X�J��n��u��h4�NOO��y����Z�����{�|�;��Ç`�����[���l��c(a�sV��R�+�Kr��مٹ�O���o&��o&���$z�H2���8��>��/�_�:7����ڝ��z��9��~�s�?G·{��G�4�s��o�t��w�oanwથ�-�9C�\Y�����|#����÷��3���ͣ{��+v���UU&��gΜ�_��/��7�g��׾632:���;'���։,f�Q��d���;^P�T>��^��#:�1�_�q���x��n�s��|�`!'�Q�%&��N[Z�Mie���jˍv�b��<��}+:�DV��v�Q��{�B:��/�v��^�7�>|�Ўɭ|��7�l��F����臲��*�N��p�����{-��-y�%�����7��4l,m[\U��9n�0����V�h����/}���Aw�7��c['����}�96>l@���GP�
C���m�W��S�N��������{�U��7���7��֩��eb|/�h�ѤNT��!��_[X;{��=Q���"fa�j��ݿ�cz��S۶0�f9��:��l�9o4[�ry����g��?���X;�,o��]{o�7[��߾i�o��Y�c\�լ�߳5��4����p��v��y'�(��逸*��|�?ˇ{�M_�ߣw�o=|h���?9�w����!�-��GC�WM��Պ<���sK��R�~��8fd��-�zu�u�2Ms�v�dQ���n��Vo�m�[�
���k>�l%�l�w޳w��it���)p�3� g�r��j����3�����9r�y������w����m�&�MLLh8Z)�9�\�#TK��s��}��s���g?��0����~���~���aǎ��Ln��e�4{��4�sɳV�E�����:��G����x��՟�OG�ހ�{�ύ~lxp��\�����u����2���z~qu�t��|�.2��bL~�~���;�z�����lzz�O޴��Ѐ䳮֧V؅�I��Ғ<��#�\�t�=���Q���ձ�C�i�K�d�m�%�2]S,t�a.x��������=��>����������ʦM�x��G�����ë\�t�<u��3�μ�ß�̷%z�S?�Ç����mٹsj�h�U&�:�ߴ��C$0�������Qs� ���[��Ν��~g���~h�ÀBM�(��C��j����gf~��G?z��>}/���A��o{�������=I�H.�*�ˍf����4^��KK��k�^�o���ڵ�Oطl�_r��(�+3)����~��c=u��wO��g�~�H|��a�S�n�'ŀ�e%Ih؆&Q\�h!̚W����s�O�T�������������`��?���Z)W�O�<��3O_��ȑ#@�n��mo{ۋ�m��Ў��{FF�HF���f�C?��R��/^������w}�c[�!'"oy�[������75�m ���ѥ�s*�j(��Z5^\\�����#/��|^x���w��; ?�S�����5�'�<�otS�d]a�+� ��f"R�T�~��ٳ������/߈[H�ҥ�~��}��i�p_��W�	�J.µZ�s�̙?�4;�������&?<�mb��Ѐ������X�-�^��h���|��ճ���|���B��O����?�}	tU�����������.����(� ��Q�Y\gZeAQ������eDQdHI'�wUw���n>�o�
���[��$�Jݷ�[�S���h�dJ�fM���h�ز�����4
�#zUu��=��~�����ۺ�F����*��.�@}D H��sZ�;�ݹ�
�=H�`¼} 	C�/ D���ۿ�z��ǖ�|c=)���~C۵m7��A����؞�":n}��f,W������~����޽{_԰Q�כ5i�
H؞�n{�`W��c��z������OҾ�}��۴i��͚6·9�x����lx�c@µ�ڷ�.M�Ѥ�l�E�"@@�}�ݗ�ݺ���k��\�9�r�����7�c�m�_~�s�#�_}�R�����޶mΙҰa����\[���u��4d\Ւ?��������+'>�~��-

�4mڴ]AA&�'�q�A�0�(���UTT�_���l�}�hڴ�ԦM 	� [�K���A�5�@�X�C�������I�m]\�z�uqW�M��b������g��{����� �ˉ�Fc��L�+�.���~���;w�[�Ҋ�� �{�w���Y6h $lK �*oЃ�c�j��w�=?���/���ٳg����U�7��A�,���=��L�5�д�G��~�Сq$_���ׯ��xF�F�=^WF4�2	�I���fF��*+�Ö,�����$\o���8E��A�O�>͚�j>��λ��(��@� .�ׁΒ�_~���]ߎ��h�R���sG�sZ��BQq��99���	)*6	��	��}����.~e�R���ѣIAA����E.((���pbp�<N8`�zEE����c/^LL ����WXX8�Q��B�ǉI�r�0�'�)��'>>ZQ=rɒ�ߒ¯.�CI�.�
��"�_����^Բy�gο�>� '�tK�2WV>�C�0ڽ��������ٳ�B
���{�Ժe˹E�����eO$a�7�ط�?�8t��y�'e[�>}�y��7��
�����ghce:�C0�
�����tE��U�~h�Ćax�=���S6(*�A'X��<�
kI�g�I&S[����_xa3)���:����P�(���~���7�|�EjX� ��L�=�ʴL������B���~��-_<Kj<䐁ojР��7l$��L#�۴=�X<��Vݺw��a�g����v<����z� ?��u�A�Ԗo�Gb��c�V��w`I9r�}�sR^^^>�k��Z Z��l�Jx�4wUW���5k�ۤ��P���Bm��#0h� �ϓ;���֠� �0L��"��P���O�c{�7#�Oy��牌�1t�u���4,l$���3��`�7�	UU�>|�r���7�ڮ1cƜ�p8V���ր����X^��j�( 	G�q=�����4i1O��G�:��pL�x]��B`�Դ�i�Ў	g$k�#�k-���X׹>�����{���<��ߕ�g=}�Y͆�qY�>����U�<�U�:;x���`d¬Y�@���w���z5� ��]q�S��*��!MM�����Ǫ��|�I"=�p�O<����$�v��EB�W�1�2���I8�В�Pxu\�F?��c�r�O>9��,I3�Ng��%�.8��S)he��&��4-�X���mq�zxP���No�"�{"���e�&����
Y�0�e����C��$*��?O~��_��N�=�����-��������'Q�D��ސaY��D55�﫪k�=����:O=�T;�g�t(Jk a<�Ĳ庱�!c�z��F*�����1�>�(1��	&�&�����!��9�9>NHԨ ,�	I�,~�ǣ�<x�`ȩ�%�z����)�����������=��e��吅IH&f��-��WhG�Ϋ��ybƌqVO���:]��9��?@u4x冩#+*OS�T��_QQ���?���]�ƤI����FQ�s��!�� P��Y��_UUWEc��dIxz�����KJ�b��-L�IM�hc"��a�'��j��̤��dס$|�H��(�ӆ��)���<�$���f-{v4�L�{�.��UVW'�ˏ.JT{t��iDԀ&O��tJ��99�K=�M�@f1����L�B��Б�Oܾ}��7�xč��1mڴV@���VQd��RHׁ�lO��v.�3TU}3�&G�5�XNxҤg��,�Pq)��'�	�C^��� �����c$Ѹ�Y��	���$\O7��6E��D`���JE�����܎�$H���ͨUUU�W�/9V~����*Q�S��ɓ����jn��J��k�p:��K��탖�`(r��f�۷�YREc�&�j�9Л�|!����4�:6�}�$g�[sP��N(��C��<y��k8�Iq:��$��v�H���</�i��4}l2�z§����)��o@`֬ٝx�� 7���R��0�'�v۞�����#K����Hx	�\�����*'?�8	�킗�8a(��"�X�CG��ݫM�5k4���g�}������N�%�,�X$|<��pR&a��E��G��!�F������t�ԙ� �yMR���%����|k�X�q��0�#�i=�iu�)�LO�P(��瞛{1ˡ��\Oh��x�	@��	 b8j�k�C��,)��ԩ�߸�I��T����P^��|rs}�HpkMFf�aָ��9�(�?9v�X"��S�6�Ei��(���b�����h�eRL��x��Ph��ѣw�ԍ���&N�xÊoȲ�Wo�|��E�ݮd�φ~L7��9�\<b�"�g��O�%h8��CJ/H��s�,:״ҫ�s=�Bu�,��`ǴL��|b��Ƭ(/5�=��#��ŝ���%�������<p���xL�@D"r��za<~�?v,����3g6��uI�Dc�M�m]�d�IX�4�5z������O?=��c_Wd�B(��3�f� 䫧�d��ìJ�ƤX̵����.��%���v��K�/@`޼e�S[�s�.�A�I�'*�)Lr�C�R(FG++_�	E��3&@��'N��Pd��^��kN��x��c��$��j�XU`�cՏ���	�fM��0ť��ۑl�$�i{�'�0��@cs"�
E�<����H�k�'On����,^�G�fH^�cO8�F�aT�>!�,�$Lj��:� E !�dɒ�dJ_��^��ٞ���0��7��XUVV�E�<���D�N���"�e_���n�p4xtY��,	�a"���<x5�{�ᇉ�ʧM�V���%�t�[���|��h�M��1 aUU�F"�q�G� 6�k��\)Iq� &�G�"dvXi�z2�����"Gӏ� E�"@��K�$��b�anv:;g�Na�<a �D\E�TT�7n\%	ǌS�u9���ͽ���0��4��h�O�4��X�����0R�����Ҟ�x���6	�H�mOX����a���I��&o�*�|{�<`{t�te�#ܲ{��z��0�G���tb�'��A�P2,XP�PxϠТE<pX���$��E��h�;G��HxԨQ�>�{B^n�}yy9<Tg�<�� �d2i�<�:8<d�?�P��������s� Q�Z	�
������Ǎ�৤��S���L�N$��T/ a��"-�pJ7ƻ��*:1���u(� B	ƚ    IDAThٲerJ7�#ɂZ��S2!�)`yC  ����5��`RC'ƍ�v+��rss�5hP �W$�s�!�>UU5�Uլ
��C}��;�?37bŞ�X�(�b6ך���2-J@v��m��ՇG���#��'>ۀA����ތ��p��ǒ�^q�3�kZ�XYޣ$Lj��:� E����lqq��,kM�9��q%Ӳ�V����A������p\�o���$�5j�R\�?�������Q�����±�q\| Z�R�p���ꚱS�L!R�=�?�1c#Y�'I��:��A�����/��5M�.O<����!��1iҤ�`��y�� �pV���RD;8��1�����S%R;DסP(/~�&�Jm{uXT]ۯ4#5t�0����%�tȀHIw�1t�tw�Ѓ ݥ��04�p��{���������[����|�LKp�C���e10�+a��Pi��KB��)C�%8T�23X�՗�ˠ<z|,bP�Ϭs��C�M��ni�?w����_�^Ex�S9�c�H���ʌ��}�&����[/��h����6s�涘��1}۸�AiC�CX AA˄�|V"o*ʰ�3�J�?�6��)}m�l���8�$�������W��Ep�݄��L�cn�E�F��ږ��S����Z�Jց��u|�ȸb_�@�	�,�����]��븩{�+��b҆�E�|�.����Ƃ��>�����2��������I�,�q3AļsE�eM�3���yő���C�c�4��I׭��t��w'�pƚ�y�fz�6�"���oJ�Ԩ眝�G��.mq�P�l<&'��ɸ��y����K��#����k|�A����M��:��|��M��{7�{x�ߣ}-��kc)�J���2���&�L�=�x�29�
%��Ւ�ѓO^K%�I8�w�;D�_a�W^X���4�a�߰��N������;S�u�&m��iP�����h�U�>H�-&^>��f$"��o���z�K ��5/�U{����[����.�s�پ&�d�!C���B�#��^'��K�d��bi�Q2�����Zd�ú-�
���X�)��v��l�uP���B|?��m!�U�x�?�y����K=� ����?S���<^��(�$g3�p����X����
�f��NL�P>�c��ri/�B��y$ԺJ&�� �Z)�H����!��2&�ӆ�Ѝ"7������"F����(�pYAYl�:ĳ|�~��5���/����,{>J�]�R�ԡu��,4W��llߛ�9r$�@�2M�a��;⾴�~��+��F�ڷ��^�T�aY"�x���'�;ϸ�������2�Xtgn�I�*o��K:|o�f��`���	��>��uA+�^p�:N��flk˩��D/�9w�'_9E�o!7�j	̭��bS�8B��ZR`R�O9�I�ޥ�i�|�Cm�g�/��2��cI�BT��E]2� �
�.����u�����	���P�
�#�3 A�����hO�TqX��ƹ`��ۭ��(�<�!+c�04M�����E�>�8:M2��TH5���p⊖9�L��={��h\<���/��o�U�Ԡ��lK�w����-����(/!�n������f���s��w��Y
3�O�hL9��z�e.��l:�bh\60N	�}����	Ș*5�RNJ8qI櫓�v��dQ��4���ɂ�EE}�jR�͊]Ɔ�ĩ�����$��������/���V"��iW�}}��ǁ@�vO� �Lo��7}��U8�=��ޟ�C�Ⱥ�Y�.�h�ŧ{Oǥ��/:v=����>/�.�2����B�k�O51��å΀����\\;�P�M~���A�-Țn�	�q��,��v�B*A��;�JCF�r/=��.�Yś� 4Э	>��f'��˂<�t���l%2����G�;³Ѳ]�8�tn������Ǳ���}zJ��θӖK��I��b�f���&���1�N#E4��C�ۺ��IBQC:k�)���b
О����e���Hq�'��Fo���%���A)�"0�X� a?Nr���,�	;wtz%�U�����_�Xr�>��|6�hKhm�6|����)�� �/h��~�+2�q�Zs�]��O�H%Ԭ�Ȕ`��!���Rd[��T����������5���d0�4�i��fK�������aK�S[�VB�������1Swd��`���[">�T�������s����
�ɒ�W��g�L�e"�^� Z��'�Q�O�uSe}%͚��p��Ȁ�N��k��&��ߞ=�.�RT��t��/��մ,�ˡ火�(Vi�UK�=Q�ɐ�ETI�gL��Ao@½Ǆ��%)))E����&W:�q�o(QZ���R�H�:�$�㶮���d+�3(pч�<T�Ǘ^�E %�`�I��P���%��4���Ms5P:ʊ���E�+�LQ'C���jW�0���a�8a�-Y�7�H�n��.�m��و=_�'/{�	S`�+���`�1���VuD�ˢu�?a %�o~�0�-�T@ԡ��+G�Q6�Q�i��5���ž쪦�X��������Aܘ��f���b^��9h��n���U��_�ig�y�����.دi�`c��}d�u�{Zj)�u�#�xoME�p��g/�]�j��X3�Z]� K؉�'_�<y��{?�J����9!����_7���s��7��V�q�����hOnj�3a2��M�G�)Vה/ȶ/ZP/,���.b�_��w�׳�h�$����&�	|1�M�L�v�W=��BJ+�J�����dG�nA���ŧס�* �4,�"�W*E��N��gGky�L���jKt ������|~���F�ܘ��O��s4��{0?�Z�(l@� 	�&��M�Z*d��w�y�R��tF�}�W�������6�����e�[������.��\u>����X�֯�yI]�aV3�z�I?F�$}�"��R5�a܆��.�ԊA��e�'�l��;e�fu*j���x*df�n�K�Y�r�I����=�)�NB9""l��(�?gS"�A��Վ��#r���d�ǂ	��4�>���T�.���T\����}�y���&�
���[r`H���]�������w��J�!2���PS��Ȭ
�m�i���NK��ǎ�클e�ڒ\���z�}�K����(xu������CpF��7�gIr�͡bPm;�N9�0�/X�)�q{x��x?�cNĿ���ݹ�Ta�����VN����}��{�/*�~��?��7�0�c.�w��|,&�� ������MzX�S>���T�<��:;� 7����rX��%�A�U������p��:;�4dA��m˔���+5�s.�����Y^�>%�aW�I`S�'Z�����3q������ӏS0�=QJ�
!2a��;�y�-�~��L��o�����9��F�l�#�'h�k�J�A�G�W�5�׺l��^QdPl�U}�聥MN�g���"ǋ_S˷?R��x5?t�\0^'���;[�<o���������朥�W�J�����Ҩ�Ϙ�x�V��5N��k ��AƳ��J��l(�)��j�8�|D>� |s,Z�)bgzs�]�&ȣ�2�}�� os��Q���ݦ�����e$R��#�r�ߡ���^��{����+��	�$`g%盝 ����8M杫���_]��6T��3�E�W,��G}��j����LGƀ�J-NE	YN�3�>oϗǳx>QT+�qn#v�V�`�/�Yc]�v�
�0���MM@'��eČ4��^*hy�M�n�М�C����|j#�?��Ë"C�G���BL�L��"w��y��ñf�<�y�%�ɶb!:		-�p�]8�u���	0/�M�V�����G���b�1�o3���܏��	z^Ї'�+�D�f�������l��i tQl[<>�_� 1x�F��~��6�<�y�9�5M馋'�%�0��a����P��¬�V�� ;�5�}���]�W�Vv�q!������9;�F��ҽu�����
�x쫿	�����<Ol.��|kT2� ª�R���m�ܣ-��]���� 
�###�!���]bY��k!�1n��H�)m��'�kʉζ�x�Et�`F��w��� 
ٵ���-�Bgk�ޚ�v_����#}�`O��~�j*_X���U{��6�2w�ޚr����M,��|��'����:��toW��!���w#S�93+d�����R7?�_���������?�o��  j`u���<<n��ex���@���u+�j��w}�C�l7�{ȝ"tp���N�y��|��qh��Xz��3~J����S�_���ӣ��gO.5�a��moæ���긑d����,9ɾ���5����FY!:�t�bGܓ���n_�05Rd��GN�Э�Q�li8�WP��G$�]1 ?��#M(���l�_[؟��=VT��zE�g���9C<z	��������w�]���.xH�:ۇ(0��H��|N"|����nS����*��El&q	X�7��?�2��\.��$.�f���]@X��{c�/xh�!�2p5�ht^��iE�5`؁%��';�B\ T�1�^�3a{
ܒT���[_��P�������~x���V�1D� �w'X�h�� jM<.�֖Zj�t���-?kX��$O�ŸtK�L���E;��v���U'J+����3"�o�}��<��h��4�bR��h��SW�<\�����Jdޘ�\aFV��չ#"��i=�oR����/�����ya����sc=��}F�?���4_1�����d
w@#���xP�k�ep{���R{��V>���g9�;�.xPw�s��E�a�)w��r�kfcK�/��d�?z���<�� ��B)!"���O�M�P@1� ���j�I���TT�y�	Ɯ����_��3�b>��~�;K�WN
USS{��3�=��H�%����4zzL�&�,�S)f���R##�WQ�J�C��B��*4%�Ƈ 3�l��X�f�o�	^>'�w�����1�Q0G���ת��eQ/�m9���sT�P�*�2��:0�嘓9$�V��;Ttv��h&���K���*�\��m���M� �*Q�ؚ��f��ϥ(�S�1�b����G�ht���3_@�]贮Φ�V�"E�P�C_�5�+��h����uS����T^^{�¨�sێ�5N�����I�ns��rĽ�N��׍��0��+c$e���S���'(���|��� m�zh?���XZ���=X�@2��B�A5?���j%�T!oN���4ʊ��yt8�ȝ���-����m��.����U������8�C�6�3�#�p��
���X�s��^P��.�ꝺ�j���&'�j�tg��K:�PH3�B��*$�,S��MQ��	O�:~�s���;��Z5���-��T�ms\��*�X�Y���7�\*���Z�o�Н���U��<�kPR��UI(]C���L�o�YM�+X%SG;�ĹUz��h��x�����^��W�$K����
qJ�Ž����YY��W�r�����ۚ�X7ښX��e$�HՄ��T`!}���L��͞���j�E}�rYF_UƄ3��x�|8ӑ>;�=C����sC�I����5�
�����W����9�ҫ��;���Xd��i�d	�b�%Sϐ���W|�+'5��enw�7\ST���F�	[��b��DW������|�`��*��u�2)L�^���Ŷ�!r�	5��XZ4ɌGW)XU�w{�Eߌ��i�hs�%�)B�D�&J��J@$�_�}Qnv̑[QW���~��͢���Ή ���ѺpmNů�6�>�oU �P��?�����|=�45=�x5`�����-{��oN�i�}�c���\�`o�h���^\�0���~��Ųۀ[dE�k0�
>�+\Ʒ`}�',C�<[�v�ؾ�[�F�K� 0n�ο �y2�T��4�"q�l=]Sq\�9dƀF���w&�!��%}9v �Ʊپ�`SZOg�1�ȡFo�x�}fzZ�QE�-#���'#��g����Y��d���~U{Av�[IU����� ���V���y���d��i�N|\���Nu������u���ȑ����s�^������a.P8!�&˗8�� T��0�ҶrL<\�w�'�:F��dtb2�q�<+�c��P���3ӱT��Zt�b��K3n\ y��vX�͑�`L��kL{c%!i��T<Fq�kwd�3��{i��[5���W�#EP,�蚞����9��`�G��U�\ d��I�ıj0��q%�[6WX����N�Bȇ�4������׼ѓ��+U��1�g������j?6��+ߘ�O��N��f�2�`��e����T�,��;,_�x4�Q7
;�		��"k~��
^xwr7��D��v��;S����.f*TXC�@�&�r��^C|,�:q��y�����S�����flL4T�L�B4���0��Hn=�.x:㊣�f1,��N^��Цh2�c:\T9�P
�qLs��IRZ�)�~:ZG�~��G������^O+�4��u2{���"�vyƺ�ݼ�H�ObK��ku�-���L��򯽥U4G������})�%�E	�G��ǆ�����Χ򪛩K��tr޻��GMįq���3;X y1#*�"��dbCxP���b* �S�
�Y�ut������F)`Zu3}#h��Nti5y�R'��u����Y���{�H��[pPf�9:��2Iއo����.U}�3�����8p�����{B��u��5H�N�bAU��js܄w뎫�ł�����+�b�Ĝ�ƞ��|(����ք�]��O���t�dEǎ;����y��Fв��6�6B�=K�Z4f�L��Ɉ�_n�x�_�y�:�[�-t\�_(��VVV:����j�3 ���))����~�ν	�F{M�e��N�KѦ�|�O��э>L�	�~G�_��ҏ�2D�Jhw��e�Ww݌���I�ظ�g��o�k���<���0'�j����i�]Y��CI?F#s��u��P����S�'�B
��ӌ8}$����C���l�8_u�Dۧ���`�kG����4���X:a�[HV5���@Y��o�&��������5`R�I(��S��`��YT����Jx�D��&�N&��o���df<`����P+Y��
�I����^y����R���		FL�.fx6����Gf���[�bo�}RS�ћ����-�<�r�(%KBz���N���h:���C�C\��I�������/�&i�!�r�_"���g~5�j�����6X�`y5�b�i~b�sm��Ӳ�Y�Q�{��M=I��2i� q�Mg����Hr־�[�&,�����Gu��Ў�X�kl���k��IN��)�岎-��!)ԍ?���AW�e��^;��zc�ײ\3.d�:* �g��&�nB�p��@>K�`�Q|���"���'F��G��XЂD������>[=��p��X5W�,5wg����R��2��i�Q/q��M<|̐��XH��=um�3�cƎ�z4�[\5�@{��ZK�;�&��$!�z"�n�,���4tu�;zj����#]F���S�rR�GX��V�e�&c΁QJ��/�_#�xu���>,g[�e�qX�V����{�n�j&��jSh N�� �f�i_�Բg@��>P1̌�I��:��,�n�L����%)MC(I�A����j��W�����٠�ok!�^W��,��b�<���n=V����-k��-�����;�c$��O
RBY����L��T���a��G��/5zb��<� i�`m�QA�~���7��]b=�k�X#�v|���������ٗOc�	Nq��~���O�J`�qL�:;���js��3��?�ď@i|��8���!��R�5��(�B���ddg+�dE[W7�Z��4�o3������'>�D���ɔ�����?���>#g���p��pӼ�͵���U���B|e�oznm!��������������&t�Ii����+\�:��[�<=���䶹x�؛7�?n�*��xOɊ���/��Xpp�	qj���p05�쾱�Ba��I�^����s�1�j�d�8�V��y�����˅ɦPtz�RHƣ�����W�g���)�BL� ����������:��Іk����I�x$��v�U;����(/���(�aN�����ղa=�Hwi�݋-���sj�Wl���Lσ���2���R ?�\���.^�*�U���v7�'��R��k"��em�Xeu�[���@��o7��,F�����>GC��������.�<��
_f�CɄ�O���8���d�J��]:�sa����0��Ȧ�	�!��
�js�e���{J�>%��6�r�al�-��O��j|���	"��+�L��Ų: j�w�2���k��4��K�yzq�kߡ*'���΋b�
P�w���~�@߯���>��(�"ԕ��K�*�vY�������[d�@M�l�q 6�6��b��C#�Hɛ�r^�~���G�?P~#H�brtL��f'����/[f<:�r����s3G)�� 
�Ú�+��=5'�`" x�RD?O�
K~�<�U4�2�wrN�r�����5�m�U���s!=||�r>x"���:|�w����x+�TZxqØ�IH�;��iqY�ײ[n(WU�hK�)ff�!jC\�sZqNWVi�g�*����~;X$�j�F�L�@��2�[&�g��{�p8��wE=;��qefݦ_����+�:�J�Y����!*���:YYM���5JG�K]ٝ~�U�I�lQ#o���rp
;�\ܪ��K���!Y��U��*-U����r�i^a�]l��ny��D��m���ʻb��+��x3哥?����n��dʇ��V~D8#���)�"�w?��c��7g�W��wR0��w�x?͢',���-X��e�hAA�Q�D���5+���N��~��k��� ���5/1P<n�I%-p�l��W�-����[hR��9VJJJ�Y\�Ï���zK��f��[f&�6ڿ5��z����������;���F0,+��f��P�f��S��	�:_`�� -�65���Hsf`s���<�eP�]�T����R1P*����J7e̖h��A�+Z��۲�F.�
N��ó�oU�}�Fv�+m��Q�~G�:ߗs��Uq��~���<���n���,̠u�� ��%�mJ�r�rK�WwU��z�5�A��e�֣J�{��c�!"y�m�,��N7T�����Zwt���9��t�Ѵ=��k �`�^RR���|/W��v?�'k}-��J�t����F;
��R�7�7ٖ�?�ḿyN��G<�%�@�耄=��������'�c|���e��YA�vwU�4�q�*)KW��M�t0�����ϣ���29ӊ��ѳ�������^���8�b�=C1�D��P��Jg�����ސ�"T�~&�ǈ�|E��X8�����2O��s�
�d] 󶱸�)p
�6��i�m/N���_I�N�>�@"�>6������	�l�p�_7CU�����X�=L����m���N�G9��D�q�Lص��,j��-�r.���o�G7�*�G����U����:����++�훏f	���O`���L9��Ѻs��s��ݕ�Z�2r��	���z���9 s�����]䁏^�a#���n�����W�+��Jؤ�������P%g� PK   �>�Xy��8�  �+     jsons/user_defined.json�Y�n�F�A}i-��K�9)R��a;�Ca{M�ʤJQq� �ޡ,�FR�
	0`Q����̙�Y~ן�q�b�\��}�)/bOƟb���~��<Y,]3t1~���͗{��=�>�0ct�z�k��㽭ㇲ���� |t����� ����[�PR� NHB6���F$G�3��)��e��rc����ཨ�e���8.|���[���>�=|OIjkA�X����r�QJ�ƚ�l^|�y�/��I�
�S��7� #5EVpa-aLJ��tm?�_JX�-������l�d�o�T�_|���|1����r{:&,#Lk��;+o��tƥ�����"�s	�*ބ�ʁ<�(y��k>k&�	ʈ�p�)-�jl\�cY����ͬ�����t�uҍNZ��������.�H/m��e`m2�᧓��׫�'.n�s�W�_�QU�cU�+�\5F<��Ee��u^�C��H�'��qfr�$d"�s����Ja�+�*���@(�S��(X�1f���J	�+J�J�$Or)�p�!B#W�V����t	�dRhM��Q���DO�(��oJg�¿	�$ʶ	��1�A<-��!Ğ��K�� �znk�Us��;Ț���G͐$�ZΔ�8�w�M���>0�r���:��Tt�$�Jaf��tk��l�׍��6��d���V|��ŭ ��n�';[6O��W=r�_��C�,�g��cT����	n�o�U�?���_X��k�;��<Y35��C->�7o0g~���'�4���M����-�?��m�j��|��e@�e�`�߽^}v[S�۹��EB5�ݲ
�>C�JeQ�����= 2-�U�$�l3��a�N�@0E1AL�"D7$QM��T`��[Gw;����烞z�?��t�ˉ���Z��P�� -0�N�JxGE��
�gϾ'�@�O�.�B����#�`�`\�`l�D)��	�5�(d����$�w`�������w)���p��h�(ɘ��L0��7��ӷg{˦��8^$J�a���N�;d��HA+��U�������:	̠��i�%E�4	��D1t�m�k���,� l��B����X+�wZ����3F#�M�RĘ�~�P2����M�̌JI���}�~T�e^��w�w�v�s!:yF�=1����pl�d�Rm����W4x
'��IssBf�b��N2	�����J y�d3�C���E��w�Tf�&:u����q�"x�=!3!�v��;9:-�z@CI�HhǓ�ﴼ�x����(Ok!w�9)�Ѵ,���U�|�8�0���޼={����� ��$މ������^�����5��X�.{	d�@b�!�;�~xՆWx�C;���_�����o��f(�囓~ѵ�M�Hp���۪�D���ש�-gJ���J�"�l0>��oK��������-7umS1�C�x>�������8%��F���C�x�mաf2��h[�&���9���qZ��� �QK;j5�t0C��hG��r�����(���؝�?�ю�,�3�~��ꬆ�~��ꬍJ��	:Dm�J �	ڒ�X�����gJ�`��SdG��Ý�/f�Q��p�-/$;j4�Ci�Ez)��ۢ����v�p�|��A�=�|��A�=��z���PK
   �>�X*M��l  ��                   cirkitFile.jsonPK
   l�X,qJ؏� �� /             �  images/278ed6c5-ad12-4b42-b098-da68003ec988.pngPK
   >�X����7  �  /             u images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   Ŧ�X�i�R�I �I /             � images/5472dc22-a170-4182-a291-403007edeea8.pngPK
   Ŧ�XF|�X� �� /             7_ images/608cf678-e816-4d17-98ae-736018483bd2.pngPK
   %�X5�3$ �$ /             �
 images/8251b1b7-c97c-4929-9682-a545aa133660.pngPK
   Ŧ�X4�:Eg L! /             B8 images/840d763d-d5af-4e15-a65d-aa66cb855cc5.pngPK
   l�X��� � /             �V images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.pngPK
   >�X�&�}[  y`  /             #� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   Ŧ�X!Փ;
s �x /             �< images/c6ed6037-c211-4162-91fa-07d26f2097ca.pngPK
   Ŧ�XʀjV{ �  /             D� images/d1dcf8a6-8c27-42be-bb16-bda153483d9a.pngPK
   Ŧ�X_��.
 �	 /             � images/f557da7c-7f17-4077-a29c-07168c914697.pngPK
   %�X��%� V� /             �� images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngPK
   �>�Xy��8�  �+               � jsons/user_defined.jsonPK      �  ��   