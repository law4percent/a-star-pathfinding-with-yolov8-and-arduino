PK   �<�X��6�g  ��     cirkitFile.json�]ݓ۶�W<ʫ���ǽ�i;��6�8�<�<7 	�jt�U���z����)RZj!���gJ��o��%�y0w�������G?Ϧ�;*��n^~r�ߒ��i<}X����Ӈ����9[���b��4����A�T�pY���De\�73�PN���=���۶Ξ�*�2n*;���2_	Y��(��U�wó��C��tBZ�I�m&L�+��&�h�WD�#3�ȴcdm�`��;�3�J�Y��,��W�!����F�4r��a-1CGq#��K�hڤ�q��pݻ���q����uW��2�Ԫ,s���`�d��mf|Q��0C��T3�Ȧc�`�H�[�9��Lx�\1����=�	U�F���QjB�z�T���T��*;�h�1C�.�����)5��ߥ0EA8�a_��Lp�2Â�((QD˂)���[G��[�d�R�LPUd��.(���ʵv���ƺ\ ۘ��|��(�2��3��3��3�~Ⱥ�T�TS*XVz;J3SR��A��}EL���k3弤N�<�"l'2���L).rm����a�!�g5
q��
�K\�v��<�TR�iB����	+LxV��0NY�u7�@ˀ�LPvesFE��vGg�2wM��`�@����N��cP��b(�8������_�Q����K��`�|b�]�"��q���Y� ������V��(L6��k�rd:���/�Y��d%h��,�wC�������+��u��!h��8�cDޕ��-r �/ r���"�0TN����|�<*f���h�!T
�����
���%/�T�OZ��}j2��Ғ9�J��ST��4P�I����AG*"	���JBE'�b�P�iP��i�K�����/M`*OY<�s��
�A�I�1���p?�D68�Y�4(fi�0�Q��a���Y�X���������s�f��S�f��C�=�4�y�hv�8/�$e*��L &�r�hr��AV	xa�x�&G��44�q|F�tG*'-84�q�dB�	x9)h~�N�	��F����y��O��b�&��O�����TN����ST��?��I���<�4rI��$TT*:	���M��D�M�^��4~i �4�i L�`��1M�b��,�N�b��,�Y�4(f'Q��TN��㩜��㩜��㩜�4��S9�8��SI��I���TN��㩜����O�\��?��I���<�]����_,��?���w���s���4q�/�Ӈټ������%��
��%��Z�����2�ی�9g��0�fdL5�E��sM^?	�:��b6ώ�1�	��\J^���Ƽ����0C#�u�jhֹԘ�u�R��d��:����{���9*�t{|Xq���5��-��F>��l��/C�T�������ûu2����!qӲ-"yx�YX�.�b �e�AJ���F���N-�5b&<���bK ���2p�@
� 2�:��5�*<���(W	��`c��r�N���~G�`	8@�aG9�J8v1s��.� 48��=��hc �e�*�Q��]l���� �q1�s��e<ݔ�n>Ϫj��?}���S���?=$�����A��, pa*�;p�j�\�.U}@��V�`\���D��TL��/����NsH���Cr�SQh�b�J���X���0��Dm���\�%��	,��v� �zԔ�Z�$��3,��j��ì��gxIj��F֦�3�Hf��ժ0���Va�ׯ¸�v@\�
������V��խ0܂�\aK	�w�M\�� �q6��A�Ä�Ka;p.��	\�����N���b؁K\�ed�հ0v�e���2lɌ˘���c��ǳ������>���wb�� �#v�rF��ߨY?1�M놱%�MilKcc[�h��ءN��أ>s��,�`��=X�<��;oY �^������ 0�{ �� #Ҋ�~�v�h�޼DI+�,����6�"��Tں�
�`�#�5��k�ȋ���1��� ��E�bu�~���D�L1��&s��Y�i!C�@8_��4WeP���Bf�d2L� d&�su�3ك��,�s�Q9����uJ�!�u�n�y�-&y�+�>4���ƜĊ9s��ΟF��&��x��H�tq��A�s�1�LcTL��u�[�"�ü!��pڇYQԏ!��C?ԏ� �{C-ԯ���o=�E|?o�r?��͡G3��_�����-zx��n��[buKޒ�[��_�⇷��:��W���-��eb�&��|�]���<V�V����y����l���7��n������ٓ�/�>�q�����xQ�$�[��Z���CMو�5��V\�����"�^+YM}ة!¶L�g^n��e�+��A�nZ,	�"��`6*n����)�ϋ�_��m��Fr(9y7\_��k��VaF���������ڹ��k�v��ε�^Ge{-v������'�Z>��Ob�n��c����5�^/y_]����lW�Z�������Z�\Y���������6�<�#>��'�F�$�a�^k�P+9
&�Y�9Y��W�*N��A������(��"��j�k@�7!7��� t4.�P�(��uX�P1#��:.�	M��b�0[�ep5�;��aKqc�[f�h� !�� 5%�2)g��2Q���2Qd@�L��?b�H�"�FL�$bvE���q�F�e���Wf�^_�	)�H@��eb,
D2;��V���9�<>M�Q���b>���L�c����%~bTŝ�e:{� \=�}�q�} :����ه��~���y�O�滹���x�t����M_*W,^�~~l��f[6�R�j�2^��aZ��>a&x��d�H����`]؞q!�ɀ�"Ӛ�,���h��L��+Yh����Fi����Fۼ;����Ӱ1���/���?��O�� Bo�����L��F3
C؏VFf(�!�Q��mR������3�_Hd%��W�T�JЊ� P6  ��q�����dT���e�#�%�̮��w����\�&oj:߀�X����2h�K^P�,9 P�ڬ��^Cf6�[\-�Ż�����ggck_�ֈULK<i>��m�rO�6��]�gU�y��i��`�3\MY��m�g�t A�� ������Hؾn67�n+�V��:xT���g��F��z��%�d&|J�j�\i d�I%Le%��'P �[5����J6�{1�Ф�SֲZQgf��e�z�v���*(l��L`���!�_������:(/咬��"��-�E�.s�r^f�� �I�+�ef��Z:|��b�g��D븅��������3JVZ@Sĺ֎B���Y;�u"D��7�r��/���	{T����TeB��x�r��, �p��� ���f���ҧ ��0�T�[� ��G��qf^���@m�f7/��!��jC~���L<���d���z!^��_ǋ�7cם7�+~{?��L���?��bj�L��v��U����v����3od�j3=J>榻y����z���\W�����������(�'�uR�a���K���տ��c�52Ɔ���!\���Е���4�Y���)�aJ�,s�ڰ3�1�1<S�rNp��`�-�0��������մ����y�Ϗ�Ţޏ�i�7M���jjG!�!���rj�ښQ���<�0�QTP]�����Z��/���7����UQk�(�I�K�2C�(�ja��p��ETT��������d������_&n1����t���J�(Čjy�>�*x���<����*���J",j]��L���~~X��.���0����C$@�����v����Hkb���������Ɓ+>�򯛺��s�X�����5��˒>��#��w�kh����x�yP��e}��b皘��GI�j�kRs��MJ������i6��->Դ>���bя��x�Mm���wo�ߺ�a�h}�F��y��`�����z��~�% ��XLX1���wYLjN,f[+�I[+u�ѵpA�)�I��T�M
\�ֵl�� Sp���Zr���Z��]f�� �JI�)8l� �WK�m�����"�9�h��m���F���w�v�[�F@��OB���(��zp��0�v��ք�=sk�h<h� ���a���=X�X:8w}��Wpٵ��V�N�|��f�ݐ-�k�u!�V�ԃ�"���?	�F�C� =�d�c=��iI69v4N-T���;6�?˙�'N���a�i�hee����7����p��p�M�w7�$��d`�(���l]eܿ��D�h�s-n���Y��g�fV}��v�ʭ`փ��LkH��h�;R뗝x�V�/�|} ��r+����O��{O=ZAAVU�A��%�R��
�������] k��xB��"h��w-�@ͮ� X.v�Qb�s�=��k�4$�l�E�iu��N ��J� �=�f�!-I��U7sr�z,���j��)'����@,u�)-��y��� j�fM �n�쌽�X�����}B�h1����%a �Z��N%�`'J�����=�� ���(�K�����A�N���(�[��w�-O����D�R �`G�&�6i=xK�m�sSOG-°�%�u�%�g43�%�j���%)r �`��&���C�o� $ρP}��Qe�5�D�>���fF��j��U��e.� ��a�0��Q&ك�d��Yu���Ùn��p��~ت}ѕ3L�E��p�{l>=xK��gm>w�c���-�A�����Ɠɏ�?����n�<��8x�?�����鋛�u����?>��?B��4�������b>~Z�~8��?PK   l�X,qJ؏� �� /   images/278ed6c5-ad12-4b42-b098-da68003ec988.png�zeSL�5��ww�ŝE���Ⲹ��ݝ����ު��3S3�a��z����1j*��HDHPPP��rRPP�|����N.�=��@�k�J@�ΐ�AAQ@�K�ky�\�<':����>�������w�«P0~�o���b���F��a9�5E�5�P���H�B�V�Z 
"D2�[��B��^:M�r]��/6߶:�Ӧ��a���X�9�lz޸0���W��L5HƴSʹ߯��l��4d���}[%�7u�[����;;KW[��1̈́��0�7��0 �LN�c����UP�ǒH'�13���1���#��Y{�Y�"[Bźq�kL��ʾ<�p��������#G��	��Ṧ�aj\��L��T�6���)e�矌v��������P�a\�4��Ԭ����ŐyA�^�pMZ.GZ�)V�:�S�J��		�t�¿E��!�Ӗ��}��}s7~!�t��(t<H�У�H&�K������e���qҭ�%&�8�R�c~ꉑQO��DE3'��t���k�{`��>�'.�
�1_,B6��<-�� ���m��1*���s*�{�YuK��^�w�B@z�R��&ed`?{�J��q��L��e��P�U��v8p����a'Af�N-��O>`��t`zi#������ap1�Ę'�pB$�,Qܜݥ ��ՠ�����K����H��������l��t2}�*����>ZM����u��=�~>�Վ��ih���!�y�tt2������дd���>�kL�E�W�X`_O��N	�w��3�V��ݧ�}/�-aDX;ڢ�{�Y.f�/�����>�
2����!���(1��H0/��D����(����yA�w��Op�׶b����(QQ��O��Ó��������
��|�5��a�a�<jUMBLp��R�1��	$~�������:\@qj_X��М�7��ɟ��PL��58��_��A/]j��R�RcG\�e{�ljS�?�H�+�[�$lz��X���i�:0����}����C�y��33�]`:sd�] )Ã૞6CTE����6I���֪�I���vr��;��P#�]�P�[���,2m[N�Ay�JL��4�!$&�b�2�HE�DŊ8�TVI�Ǽ�K�W�s%��5�gz�(��j��晎����O�A�8�/,4�ح���H�p*z%�Xa��p���]$�M7��8l�[�c���ӗjt���Q�������V��G�F����[�7�4���InM��A�;&��0�[&�ޘ&���(y�DT>�x���iN&�hTw�$M[hb��:�{�[<�F���_zf�FB*���Q���=�0���Y���.��\%7�h����#P��n��PmUҬ|��n�O>�{�5���4/J=J`��� ��f,���<H���n��*�������U�*
ć�#!y#�1�6!ӧ��R9��y�3)fH7��2�����Z|�c�����}7���t�u�`&Ԋ���p`mG�l+���O�|�,W��R<���o������lV?�ʈ.�� �犣��6=<���_��153�3=l�ѵ!�:/�[:n����@k�����zhygm9�҈Vd��O/�m��R�+�7���U��m�v*V�8�e�v��G��p�5Zr- Be�|N��,M�	re��ҝ,��s��7���C���8�(�jY��>y�Py�%;���"�u)�hq'}p��'��N!U����֐��$�Paˈ��&���?��(:�{i���2��e\( 6�>��%'�g��� ��C//��\��U+��Med�C�g1�.I�v0�n��5��'�â�F*�f�J�CqIcyKJf��C��%|�ڵ�r�w7&c�o���|y%%N��Rႆc`��f�P�g�X��~�[3�;�����"��2�>E��2���Hu Gcab0�k�UG�ӑ��2SHAQ���!:�}�Ӣ�c�}��<A�O��Naz�T�kB�:��Z�HV�j�I��9i�2;d�=*��48�:Ρ��g��ҭ~���#�^W ~'�T�������p��Я2����U�Ĳh|�q�`קJ�b|�D`b��g���'��fZt`��%���c��bȬ���n�B�!|���Ma���H���"Rc[������N�7�I���C�M�q�gY�bh.g��88�2G�w�(s�:��X���9��$�eM�.�\��)�9���03܌�2�m��9B�ƫ{X�%�vhe����u�z�3i��!f"E�L�-G��XL��RFE�����\^Z�kUy�B�w�-V�V��%[�������:~���/9����X���ұ�ef;d�w�����O����ݧ�e�s�1u�g ��
��.�
a
7���D��[E$%̬,��R��p�I�bȏ;����aP�lJ-*����h9�-E�Z�H�!*է�/����~�e��[@�"v����9.����:4d��w����5L���K�˴
���a5���Y��M~��9����f����*�Z��X�n�u8Vd��C����I�.��e��|����q{`Y
�eRJ]mW���K)����������c3�Qu�����w֟l����T��B�;���^,�m�[��`������~��"�$f���euÄ�";�Ƴ���`J��7]WU>b��Љ��>�(���qf	����\]ܪ��ԣ8x�fk�h^=�rN���B�WK�8��ɰ��.`Y	�#����������b�_����-/R��cdiS#Rd�n�Ǆtq�i�nQL���S�!0��n���^5�s�󕫙�6�{�q������S9�g���Jl�wu�|�]<IݎL�{j���[ 1��p˪ҏ��  ��3`�3�ײ���1�݊>w��Ȩ4��D{�.�|9*�
"��8$�-�j�$f�"zH�����!�,�^,Q��x����K�]%g��Ǒi�j��d���j����莁�f}�t尿�-�����_�@>���5G�x+�P�_�,u�:�Ao��
 f�!S��k
�x��$�c�Kt>1�Is�ؾ�*I3�Dhpf�8��0� t �Ķ��)LH(y42�9sbZ��<��*�u�%W��R�Km.�����f��7���\��Уc
����1��S��e �:�3�'t�VqT!�7�us�a�^^a%�3v��d<����S��Ub�G�x��{gg-,���6��!�r����������Q��a�"��6�Y���R�����J�5b�kP��k[����4�:[�&�2d&�]�h���58f�w��$�]�g�h�R�!OU)�����D����x/<��{�je߱~��3�%�gmZ��'K<�@��*��N,s_�u����F��S�K�`q�U1���?1릂��MC1u�bDj���F�	!7���߅=0{P�H5;[����r��e!�}EM�jqT�1�$WS_�,N�ǁ�B#0q���wfh<GK]_=�;s��I��m}Y%�jG@E_Zo(�R �3�2Cl�]��IN�u�;���"1�M� �C��"�Ը�W���h_�+%2�Ѿ�*��43�4�1�-�(�}D�W�-ڸ�E�rS��3����U�Q�'6.��H���; m�"=.�m_���^0z�F�������@魈5U��� �u���a�g ��[�Q4돿�DXg!*��~�� ���kL[��>0�`j"�ߙ��b�X���j�9�� j�#s��M��r#��`����n
��oUt,�b��/o|}�)*6p�c����0�G%�����?�{��>�wRK�I��)���E�K�ze2�@?��+ͅ�@��/�,�"8k-�U�SU��t��Gd��Zr��)�ޛ�臆w�(��t-��m8��[F�]��?��gGnH'1� R܇0)5�j�F�X#��bCl?��H�Z��T�nh��]��#mO�=8�����[�$>,��5)���Yb��H�z��]���*�����u8ߪ6��LV���[�r�)-�b=����Mǖ�*+�����5��,��$_�u����"��Ăa_��Dj/փ��{(�yE�ܓe���G�����ť�i.�j;P$�%��;Rx0e��Ss��d��u ���)�XF�t��K\�?���;6�2�I^}����P
J�b�J �F|�M�&��K�M0>)�����P��6����|�J�\����YC��)��]V���ÏLS�[���h�Ȭ9�Q��#M�Cӳ��~�3/�ஔ E>~�_�]0{Q�ϔ|�����ǋ �	���O�/��h���k��?���g���|ɕҜ2�w�i
N+�o7d�G�z.�2)G<�eޓ��-�L�ʳ�g
��fq
K�#&��34��O�� �$�H�2�>d��p�W�r�_�on��YlU�a��,j���)����<e�CWٰ(C]'��5�M���;;���Y���f��G0�.4	�63�	��:�bT	<Ys���BЌ�c��H��>��Pz�-j�
?�10�T����e~ȳO�>����r��]�É�-����'�oX����1W]�=~[����aZ����f}A�d�n��V�S��h1ʢ��+��lq.����>'�ʴ,(�Q���V�:{PynolNa$�f���;�352���2�	��.PPB��UζGUǪ7��$a���=ll��Q:NZ��v�zַ<&�1�'�(�v���`o[��2�b�:��v5��:��𚧰D���Ï�á��@�M����5i��d�<Q*8ci�K���p.L^��u�z�VWv>v顜��K�>=�/��!�`|jV:�E��!;� ��pAx�U�.
��9��񣄞m,��P
Y�1��xґ�x�Mz{_mOM��Q;m&[8�Nq��W��H�-m~[�y@H�i�'��!��p��O�&�P, ���A�T$'�T<ݝ~�`��&��yY�F���S�?�Q(��C�+�);��d1n�8��^.L��Y#��W;�]�V�T�V��..�Ջ��}6�VF�C�t���,������m�׉��*�q� 6D�@��7�{�ő�@���V��J�t��ƅ��� utI ���ڂZrw���)�\'N��s�#��.y:���'�3T�-�����&5�><$f)R��s�M�p[}���F��F��X붣�$���%��XtCCF�m#���5O�^�+���e�~���t��c�umYȘ�}=����sk�R�c�<�����3\�� Q79�3�~��XP%�rb�RǦ<ɐ�#"�q�PKw�x����h(1����!8�S]�˱s�ӵW�m����K�$Db�>���oy�rA<�Q�(��#�>�5B���u^���m��&f��E�4#�E�7�6��+šR�0$pLPAX"
��8&�h:�D=��-��&-!�����]�l�܌�!n��Y�ڀA����j�,m��FrQ�X�92,V�TF�x(�l�v��X���G�%a������\'J�+�>�"F}�y��
�k@�7#aJ������:@�їK��>|�%�: �\ª�	����`2`��޵T9q������vʿ���Nyq���o�����dhS�ȕ��}D�]e��@	 =2(�?k�n�eA�8�5�:��L��;!>��p�SO�[�}Y�_7��4�`��/�� 4�,�/��lMd�'>O�`������xk�����g��a���
�x�sd��5�㟕��6��[���k,k'N�16�{�X�БF�K���?2&�	����N�[�	�҆ �}��)k{r3#� eg�l�-���RH�{?2W�w�Q��ڡ-|�h����]���@grS��k���Ԇ�^7���8Lp	c$kZ���F�y�6����"���hBry�j	C0��4��+�DoG<�]7�#DBe, pcߕ,9�`k�e�\:��ΝN�� �Uv$áD�I����p�9�,���M.��s�S!��p|��R^�M�t����8��u������^��j`ð~*?��� �4F�XY��M�ǿ�b#���ic�?�P
���VlL,"�pw��6l ���U�(�L���cZC8`#�N/�,�y&b�Ջ�`��S�p8�1�qRϠ(��aAF����=}�UR�.k��i8�����W	o�E��g�|�6�$�}3|NY�ӞIST�=�����Ѭ�w�[�`�r�:I�Օ������^&ͺ�'�[�(�06Fa����������6��j@.�����v��A?��e�/{�s�}�i1�[?�W�g�v���R�EEG���QM��ң�ux�Mb,َ+�8S~6 mFy	GUS�`#=�?�8�>�9�'�)����T'����!�(L ��DHp�{�m|�����2��<
}�����i#7%� ���+J�Wv`k$3
� `�� d���S�m�ϡ~�؆"�*:��4��F@p����ɦ�	&���x��yD��O�IH(���vo]�}���5i�Z�{�v�{v�|J�[bQ��`#�Qd��r��fȶg��B�A��U.h��A-I�jki��	>���|e��rm(#�V���:!.<�����	���o�	����:��p.� ����vX
�[RE����� C��?��T���(g��߮[#9�8f�&qz�����uc����Y���	y�[7�瞟�sFqxՆi2�{J�f���0e�!">��nF�*y��E�[&)R��F�sR��D:گS������l�m�ibh1��ā��xo1L�`�PG��;ZhSh���ֈ5Ƒ�כ΁r�A�[�3Գ�s=^������������p	�3�/eX��������{���#k��,����Lo�P�),����|�AAe�J'�,��R�E���u_�ͤ��	/FjN}x`�/���]�_��%_QN�;����*�f�������N?�L������ ���W��'��|�F�f��Ws�;A<-���H���$�9��]	x�լ�=�/z.D�XRK�(\�N�ᓖ!%gP�q��b��鮣C���N�&,����"2�vCCIxh�)#����~�zU�#�}NY�X��t������R4Fd��"�	@�e�ǢD5Tm	JC�5c�p�Y���g�?BX���)���^���9�J �O�w��˛D߱n�P�3?j[����3��tϞ�B�(�N�����- ����>@7йe�lߛL���TO҅X�C4��&g&�k(��Nm�2�}�-��Vg��ʂ�<�1�RA�L�s,=C* �q��`�p���-L��k��~�WO��C���HI`�]�����$�Y�����Ƭ���W�+b���&I^��`���aKT���Ǘ�<$��YW_���8�fAҟu�w��$bo62��������Y��x����{͉6'�����'�\���s��a��J���ݔ(��_vI^Yх���4���I�hP^�&h`[��u��,QZL�r�����a�T	A(-Ee���	�W��gà�����ݞ�^��A��D�����>!z�[���e����z�Z����'�k�-����HS�/Ew��)c�= ��+[��!Q�[��H�����bmI��U�{~�ϡ��:���^�, Z�M	)���.�~`��s
$ܧ/8,��O�3�P�>%w��m�W#P�)z|.ܵ:�g��+'������Ǖ�fÑ��@M됺�����ŀ�uE��.�Mza�E�X����ҏ��Wc~3{��!&�V����՛�&��r��N�VM_�Gi.���8ޗ�J@s!S�4P[:]��O�n��R1.eܨjX��P��
y*�,$���;kn(�Á��ո�@Ʀ"�z��|�e�}���~_�JKH����
�e��-9�G�4'��U�煮z%��|W7P��""�NG��u6w�l͙O�3T���ޛq{���������*�k��wxIP���	]ՂaGR�	{���}�#���9��9:ʟv5"�'�S��%5�x�&\e'5FI4ƾ~�_/ ��G���g`�43A�C�ߪ:�|r�x������/�746��-�s%��JwbyN��H܌or����v4�ّ`�#�g6t�ҏE�W^L��]f�g�r��sh�v'�p2�;�}�w��T��c�wA*KbٵޤX�<��6�mm�WS��4e��R�i�&MD��x��R�+��	�҈���0d�6�/A�fS��f���� ��Ń�g��ܐi	X�Ÿ�m���`Ċ�ǑM�75�O֤9�A.����}��~p@f�/�����:O�E�MG��9hGB��p�����i(�]Z��b��	7����-Ɩ�6��U��8��?���|/$��bSlձ�:Q�a���E��Ö�	��G=�+�
z��#
P��H;�����]���y��e���ρ4݉��S�9᲌�i,��QJ$�y����~\N�P����$؈ ��G|��qs�������N�ȣ���o����Q�(�xYj%��\ACb�=ew=E��G�Ţ���'_[}OC�O6�kG��y�?x�KɆK�=�ܥ玎I<�B��ަ�e�lԜ�5@��D��O������������r�S�=�� �� ��KYbD����RKhMq������e4Ҙ�憮(���rMJ�<դ{tR�&�P�~gx�>̫�lS$p�Kp��	\Wa����]�U�*~\����I0**!�B��}�-��|z�����f�T��+iד����A��l�r�
{k�"��b��Z�ZP�4b��������'��#��S�v	6���A�d��_1.bz�uGp��݇���d��g�g4��I���%佰3��ɉ,8�@�.&���ed�S	�d��*�/�$�Ҧ�mJHf��0��Gq7���#u��=�9�d-J8P���K�븻4�[}��6�FԘ��gbU- {MG�V)�<�:<�����3�5&՚���"�IE����*��ߵ��B�؂J��M�fH���2��b6d�R̃]��e�!��s�B�`@��mR-�,�|ʳV+]�_�F�1�|����.݂z*'�չ�~�i�W���-#PN&dS��n����hW ~"�EŠ$w������:��"bn���ߗ��*��j666UN��Þ�:϶V�N���HXv0:�?9�����p;��d�|5�e�M4CN�)D��&�����=�A�r�U^9���#-���3�u@[p��`����ҟK�6ϧ|�q���.`+,&XV*���v�Q�|*cU�-]���C`��L�;e�ўvt�Hs�3� ��ըe-�m�� �J�ƵȒ�`}"��ĵ�U�^dzL�y]l���4�I�E����=}�p��z�+���b��r�T�rD�y؅V��ٵ4���]�G��|TY�h�V�����n�ƭу>y%!���UXl�AioP3p&9�ݪ�~�2�G�ԵV�9�ӏ�Q��N�Bs%�m&���(w�h���2&�=��j��zK͘;f&D�ߐ�>N	KR&gO
�ʋ�B�y�@y�Dۮ�����Siw��Xj��ƾy�vJ�DQ�Cu������B��u�����2qjR֥�9��?�?D�!eT]�%�L����y������9P�=*��S��s�X.����55�*�q#b#[O��~|�l�Ӣ_+���J�D�ea�e��lvn��n��R�.tR�Հ6�`�4I�f𛳧��p]Ҥ�(\Ԣ�ϣ�խ~�Ⱥ�^��nu��r�� �Ξ�h�
EӮ�k�\��ҟ��d�F�����q�Xٍ��L� O�<��������7u����cOl�_���-�8��4e��zZ�����.ggI#����
��'�bRܓ${���E��OY�ѹϐ& ��pC�076d����,���^|��A~��5l+�j�?5���h���˳���؎�b�R�蘆�8(��/�g��H��f�Dퟕ֚�Tжs~�,]���}�w�
���y>ݞ���:����������;8pDGZ��]<��
��pʬ�޸Ҽn�x���謚.l\�#n�q&�q��7{�w���n��	4y/�6��zbB�B6�;�3���DJ�3�g,�M4(<� ��S'[=iϊw�c���ѴPY,��n��&�m Hb{@���䕴JN'��H��Z��=k7�50�!�s��@<n/�3�~�D�s%��!���Mپ�#��S�+N˿�Ke��ւEM�  �5/�?��
���R%��FP���8c,����	v�!!Q]p�iRP{�|GS&�FA[#���޹r;�`���N�]h=�& �8�1�nP�2#}�)c���OYnkʚo(J���h��^����g$K���m�br�ո���e���M��M^��k�J���S=E��%@�^�oVѢ#��)�[�6����s���M��}y@p��'������-0�<�2�L)_�ԻB@�ګ��%�΢f���`tV�b��4����xj= *�k:���	Nyܓ�+~�Qo����*��H(�I�b�©�PG��tH��=�Q'dʆK>�!o����Ysʃm<!D�S[@���eֻ�����	�y����y[b�y�e�D�d����SE�6/Urt�g�SѠ�Вu��E��T��ZL���H`ɀux�[葮��Ǒ�T���$��z�4T��K"�V�<")|UppԞ�\���MI�����^�{fn'n�-���zHұ˯���%`L�Q�p�W_(����~�AlW�ԝh��{]
���J�xe�1\����Ñ#v��'��<�$��j�����?��3��ߪ/[԰�.O�"J�z E>f�)���F{6�%���y�u*��;��)�I���ImĐ"15r�1��-)!�Y���`o:��Ǥ��Ь�F��)����/��ì9^y$�)Q�'�ƨm�t��V�����.�3�>J*����K�R?�i��9Lca���vdz��3FB���-���tU�ib��6�kP̉'_E�:G�I=���$r`mZ�mR��OC>M�����<"�͢�m�	�ߛ���F���,�g�5E�$�����ߦ%�D ��Ύz����A����"�0B�������_}�z�;�"��m4BSR���J:8�2�?�d2��8�|[��yҢm�Qo�zd�W7<mP�mc-��n	�T�����E��#I�[�^!�X�Z��<#}�>��&
h���0�TYjsſ�x���\�;o3}K}Y�O���}x��
�	�:���۠�_�Z�֑]}�G�^sjm0q*!\Q_ą��/��g�c@��˻0������/j�n0XKz�������_.����t�
��_/�(�&��v�yG�<��䤦��aW.�"��.�!�8�j�D��K�R��4��RG�������Դ�t�}0�
�K�j�����hm-�[�z��#�t�Wo��փ���D5}`�@��κ2L���XA)\r���J�#� �+9a��z��N�bL�e�Fp#�!�:�QO3��l=�I����=��[Ðf�閄~�\{R��
*�J���P�\+ts�O�j==��iqh6y�����F�)�`R(�Ǎ�1��b��t��Ϯ�H��fQ����}��pp�P�f���c�2�[�{CM�5��J2�����&���(�O�-ۙ<e��g��)RO�wA'nԡy/�����ޞ�co��k��N)�Y�܅�\��s�zcjtTn��#�UL��KR�UV�ne�@�a)���C�Y�sg��`�������T��4�7Md�v���1��df��L
�L����忐�3��	��=^��j��x}�cP2*����A��͜h"�m�y$�8�q
�q�����`�w��	�T��=ȆL0胛�w���)V������i�J�9�f�r�)t�rB=X̧�m���Z$_E����2�U��,̷�����)n��h���o9ʀ�")�06�|�y���qi��?^)gG�N�^�#l|��h�����7��Q3YH���:M�<��駒�e�b�%g�#V�\(L��Ǫq�n��?jw��$�̭w��n�.�~�͝{���JX�����+PXY�������}58CYzare�z��eI|�H���
��a�8��-n�V�C$\"������-<�X�Mf�{�L�(�R�}D����/+z&���Tl��4�[����nw6d@%�;��\Ke����ie��a
�qr�t*�OVՎFp$�i�G��{r��l0��"�~��}ؒyۘ尢�G[T�WH����b��<D�y�6Y��Y�x��B�O�Y	�����qԈ�|��m-N�U�g��S��Ë��;Q7����IKi�|�!	2�qK��~�������YG1��v5�ONT����9��$�ö����l�����G���Զ�H��zvP@`ȸ-�u��h��"���Q���:L6���Ov�A�	e��P%	�6M[M��df>�|+�Y��n�������)�w?:{��6�˅��ף���?ώͧ����Aɤ��p�%��*!������kve�aվ��Öx��I,0d��)҉p�#/&��B
��]`|�L�.����i��W۩x|���~�z��Ԇaw��x�Ȣ����>��v�?����g��}��nQ(}�fl^�3�b��"�Ġ��Gwr�7�j�c����yH�E$���Y[驭"F�َ��@���_�eb,#?�Z*�Yi����Fboh)�r�W<��k�h�Ƒ�؈��$X6��<c�ה�h|�c�Ƀ��o���:�!D=Q�#�b��X�"0�@S����%�uT{�̽��BQ`�\&Q���U����]%�N�z���jQ�M��<��b�*�M�g�](/�ڹ��Hg .)itԴM��Q����(�<ơk��Ü��\ٴ��Cw��T���:g>9��?��g��/%���^��u�<�y���J��E[��-�ķ]:_���IuF.��]mIi�,�}�F�ݯ/�b3<R�{�/^�"���'��U�Г����KB�%��*#�Hh�)���V�#�+:d֗c�g�hg�#�����巸H�����|\@�5%�����o?x�pߖ@��[Hwn�h�Y����:�SA	P�{�X����E��j,ݻ�mh�we���n*����d㥊_�	�;�L9�%���u��������0B�&�n�
!��K�Y�3�T�{��>̔z9C�m�=�1�J�9��������������)��hm���05�-����p`'+~���������v�:��&բ�g�tũ�Tz0�%���,p<?�ڢ"-yڲR�c,K[�p������=4���yo�^1�c{�ƛ[�ᴴqʝ��)> �a����;a��=��p��ZB��B��<�C�u&G&05���� ��N�͞U�zȝ��@Ra�%�` Q���&т+�=��t�Q�!	��FE>�H)Q���mg媜!���q.̏��%��UWs=���+{;R��w�ԫ���v�&o>�&J�uF�s`�GF��,j2=Ƙ���ՆF��4W�	�
�V�1�D���)�Zd$��G	珃����+����y�ZN�q87���LvO����˩��l�$�=]+b��-l[ �K�K:(���MD�l�'�}��}Ps0	��1*���Սz����|����8 :ls��f�³��S�t	⁨�Ih) N�3RYS�!C�o��C�.����;×�����y�m�P��Ϝ��C�d�s�Z�LـV�a�N�!:�1�����/�'��Y�c�9eA�DπJ(����YU޶�#��7Ag�3/4��.��7�����aw�|��Y7�� J�+3�$��ܣŶ��1Ms�b��G}�tm~\��Ƽ�^3[�G"rL�dO�w�zc�����[xcO��4���ZM�ea��z���������T\�
~�#ϒ�S����}�c�U������w�������؅�����V�ʆ�����!y������xg�"����Ӿ�{x��V����i&*pN$DƓ���5fp�=�V���2%5��ؤ���w[�N޼�`�M������풚.�6��T|���t&`�O����R��eK۬+/�Y��5z$�JJI��][Ӽm�A���Ɓ���(!���P0&q"���!�1Y�����`�p3�"ʛ��KY�t����_!�,�k���G�~}�?���������Y����$?f�A��aa=���:,-"�"�|�����.I
��>��hmcc��^��_���~��O����!�h�����^�9��mw �]�+O�?��;>�X���dŶ`��>ȫc���6��Y1��b�����3(O�47�@6�U���o�),$�� ��Ŀ����e�|2d)��Jј[J����X���J�/M�����-�����G�D�����<��Z����C�b���hCK��%E(c�d)7�$�ٓ�l�NR�\��dHl�-��/d=�K+<�+�7�;Ɵ+."�e7g�O]ooB��q����AW,�Z�	�Y����H�p@�[�k�_�>3�r"�r���%~"v��c��a}%�MQ����ZM�mK����� �X#Ų2��6X�)7�����c�h��y*�u��7�_���{3q�謻�$�B�Z�]9O�oL�?_ĺ��}_v�:��[	 6�-�H���� �L�+8��d�˯��mm�1�v#t�c�vN1�h,��h"i�JVW
1%
}�;�g�Cc-�Df�\3Gߤa9�t=���qB0�� �&a�ɳ�ce�♼D��U˙m�rf�?چ>������\�S��-7�s���~�x4o��)=6�Pv�	[���N�0G-l*�<�D&����/��(ntb5�dB����,le˄�^Ka��]?�^��=��T;��q,���X7����������9���`�`V��bpD�5�`J�:Su%�s��vpO-�S�ؖ7�������$�K�L,�eP(��hjB�6�c�ĝ��v��f��T���`��w9���ܷ��=�,6:���EN{���Y�XE�=v���`���>z���~�G��������2��~�`��J�&����x�7Mꑷ�1�B��|�i���W3x���Z(A�6��.7[�a��(�*w�g��mz�mm!�.��w[���]!\�`��[Gk�t���v��\(�\��²:w���#e`��
#ʥ�}p��������5�A��S�8y}�~x=�Շ=g�:8�O&³��e1Z:�9f/R�6&�W��}��'�D0g�����N�{�6f���jc�C��&��It�=����_�r9�k�!�-�[�C[��V�e{�F��l&��AK�|�:�e�1�a.8�D̑��M!�WKo��T��_���G"��
���j�����0�D��e-��H[�{�h��A�{mkcV�~��ؠ���7��7�K_�k��&qNE��x�� ����x�L�m#�r@F*��F߼ no�өA3}-�������زej�$��
���'st����z2�t<cz
}s��9��Ҕ���js"��r��EĢ�t���T��;�y��ة�,n��*N��D��;[z��e�4�f93�D>=�'��`�*I�L��K�ʌ
���v�5H͕�+J��������O�aQq_q�7�	��1n^�J҅1����}��W�7���נ���V��Օ�<�v!�u�uiuU������^$r�H�d���ŝ�/ǋ���z��`��;��M�Ŷ�Ah��>�
��hmx�$��h�Ãnњ=]%ah�`g�_pDRI��[j�Z'��`��-��+���þ�+�5p'�KJVB�3Y+�m]���]���ʢ���HB��QZ����>�P����V��+�#��{���|w^㵳��1��F����U��S��p`����=�
�����;�a{"O`
����"�:��/��/RS�vQ�~�*���u#���0�yW����֥�pR���=�4R��� �齔�N�.��[
�:��^�$��&y�M�wy���p�*��f]v�A�n��w??L�w��T��7��rף$l�~)��$�S�3�e����=��}��m���M1��9�lL?X�w�@ eP����� �'��o+��Xs�TV���RY_l���)p03�ҳI^]�<C���I.�������3O�Gb��+w��C��~S;��F@�|I:Y�����"�ӵf۬������}��Dz���� 1@ο�;=�1`����c���T�i�˄��r`�y��Oe�ܕ��]yH��:����Y�2-+��p}���dݙ��kJ��nwZ]IV�;�
w��3ߑӚ�h���L��\4�5�:�jq��y�������cL�q��IS��O���;��10鏥e�k��X۸�R,���SI�	�cW��6�[����&�,����#�����i�!s���'�h�䐦�������P3;I+�X��R�{&��J��=R�-��-P�R�̽G����x�y�h��s\��#t|ԛ-8��Mְ#�k[��vĨޞ]!� �E����}�L���Tp��p�b�T�4`}x.�@��J��oon}�o>�S_�����õ���9���u��/F�8p�lm��s(_#hT4Cd�q���>i�L���vsʎ�˲���M´|6��ux����Qw_ߺ/��茦v����p:�Q���ˡ)81�8Y-����Ǜ�b�����^����q�\�<U)*���w�Z�«���C�L���{�5�����������}Vl���s�ŽWi�ￎ�J[v��ѵ��LlPo���:w7w���)�V�]_\b<��jʟ0��|z���3\\_����ɿ��`��E�ՕҞ��%��}I�sAt�]���g�$;Z<(B�v����u2$�����4q#� ��*b!��aW�5�J�*e��?>x���P̙�1qb2�.]Wy~u6>���L�,ӞU���,��N�|("���q�eXJp3@���il˶ly�T-� l�z��T�҈a�	ERp�)�Y�zP�1�-�b�p|�z�%̍�� �1v���^�`�ݒ	�޴�h�����d����	k������h1���)N���f����l�[�U�à.a<��W/0M�X����ÚWǃ�=���2K�]���D�t?1��PVJ�����l�KX�L�p�3��H��������&�G��]��R�5T�X�D�i4�ۃ��M�sDi�rc��PG$����0��pq�Τ����MRAg�M ����_�����z�_��M����A�rt������h�x9���p�qL��j��:p��&'�)�hbx��ܑl;|�.�̊�ƀ̀�'V�����������a�ޕ��/�p1b�/�9\&�)%�T��1��H���=��w{����x8�˃}|z�/  GȉfS���MT���/�1B?��Fc�j���yI��/�p��g�n6����ob��$����O^��WR�J@統�[����AMy]]KW��Z���kaTϏ��1���v��Z�7�=�rZ������-�7�k��{��3���c	c�fx�H;����߽�Z���/�^�r0��Ύ4R�V��67k:ЉR�V^�""5�J�z��'8��2AT�1;��ϥ���kzy�F�RYa�ͫ�	�l��{|F�[����Ķ��c�h�L�ڞ��b#O��x���s�h�ݰ*QA�	��n���S_3 ͳ
WI4Ro6%�?q�N��l�-Ƹ��5~�J����6�[4��<=�x0�>��Z^�.�F��$L���֠sN��k1osc������&�-���z���|"YҌeMܘ�|��0>�4A U	�)AcG_�_�$c���p����Q)4��1��K�_�7��H���U&�V)�0[�$�qisʁ0!�y����]1�S$��}`B
i���J�
�＾��k���@��?|��s=���U�[�Ѹ�jr���Ø�o�wK��&�6�[y���Ow4�T1j(O@,%�fI���T�Fû0-PI�������lW��,��#a]l�2Չ�/X�u}�I��	,��'9�v�xsW ��x)pqy���H:,������D�w�����XX��ݵM�t7��X�8����?>|.m�x��.���oJ�i.��� ��G�/ğD��kACt��;w�t̯Lf��ȫW塿��S|J=lp-�D�erf��&��k�wP�*�__b8H��n�%M?S�����������:�T%Tz�{�����OO�N�B�.M���S\�_���L���������T�'WG����^�₭�L��dΘ!c+w۲�Z��x�s�^�4F,����!��w���b�Up�Nג�-$\��5��d2�P�]����dcUa�`����D�	��U����Q.�	�&@<7�͂��f�NN��p<���'#aml�?*9��T�fҊ���Zn ��8�?D�^ܭ?Py"ِ��N*�%��}���5����f�c� ��:��"��o��qӋ��W�)C�A���C��l^J�լ@1#��N�W�HB��ͻ�5̮G�'3�L��.�FM����I��<�YE�y��$�x��D����5y=-H��G��U��V��[�0����Vm���_�������s��'�4ϣ�o�����.���h$]Ab%�=�s���
7Z,t*]�3��Y�i���a�L�&���� R#�2���*����6�����z���V�q�	�;}!��S�Bmw�k�{�6��Z]�@�:�d&�d����Q/� ��:��h ;�﹒�����쵷Џ&x9���t�����0m0-'�^��O?z��bd���x�է¢Th2W�qy/l_�ؕ�P��>��j��NS
����T:�0��f���0��{xc�.*:������P;��z��[��g����ở��Q�/F�x{�~j�ZA��d���K����ְ��`~�Gc/�quy)!qX���֑��o4�j˳h,����pM0��Enϣ`(X���]J�2�g7������Oi���Y{�(��2��C��$������[��ye	�8��sL��Hv�`������P�\.F��ߨ!hTE�=�>�񠏓�DZuIa8=��t�H���X����i���K8r(��cs�l��D�o3m>G�f6�~����Igvz��E$�iN��YY��<7c�Ô�zF���Ȕ��3.7a��p!�$K��2ֈ�����P���N�0:�����]ӛ-���D�	=�7�&�(�q�	�9"�!���f<���A������I�BZ�qO0p��8���Z�ƃj�{o��~����������ӿ�pˣ����/Ώcා��:
�--\�r0��B�V]2�L&�NA�����s��lG�m,�V&�b�2i(�l"#�R� 4��^[��z�s�I;��1N^��Sn��7/��:!z^U��vg����Rq�3���Z]����O�H2a(�������m�6q���/�߿���ev���|��t�:h˽L��ы����sb����1y�>�l졃��k9��o��@T����3<�:���J�X)�w�]���|l���E��5�om"��G��>� ���]����:�n���}����s�fS�}9���@vJ�l1�K]���Sn>C��ss�FH���!~����j6Ģbz󱽻l[&EgCH�tT
����N��nle�?�����˹e5��	���U �tE�tK��*yFn����sY9∿���an�4\Ut}ScJ�$��N��LF8�8�97wCI@�<�z�38�0yX8u79LYk�+����34�r
�#�,P�d��4ղ�9��}�{��\$�ȩT���I2;N2���27nӲ���(�۶Gc/I��<J���<�?�3�Ј43]�<۪u�̑�� ���@P�ʜ,
�nJ�:�o�T/�@Hd��}�><�Ǆ��f��WE����$qƤkg��To�ۿ��'�s{���vpv�+�@���dc|����B!R�ML�����v�NK:10����RGl�����#�1F�p�t��N.a)e�y*��{Ua7d^���*\��q����L��~xy��Mۛ>I��w}O�{eVem]��t�,wB���	k�`��+G8º�[������1B��_����$+l�Ax����vO����^�U���9'+����^�2뗿�9�y��OMv���L�⣮��VE��Vn�)��)~��@H�+�S�����D��vqqa��u��vQ^�W�����kO?��o���(������w�^\����ݳ�����x�l2/$k���=�i�+%��"@?9ۗ�	=5�+���׮ʜ��-۫W����+�B�w�X��jG������������ V	�oo\��Rզ�����dz]��E �OE��:F��4??�P�B��b:��G�/>������3�n��C���u>w���r$��5M}Vz6�-c�x�	��QjI[o81� ��?�4�5�뒨\��XkKN`�Kv�a���·޷ʠ%[�Z&+��A�X�8����5���M¨��H���N�AcG|�`i%��Ap@�ՠ�̶#�,����mP��2+<�A��]�𺰰k�E�4��!/��c4�*6�H�T�y(�M�͓v%[��+u�QY�� ��J�T_QO� A�(:q��`�SY��V�V�>}j��<�l����t�wϔ�|A-+&���ۍ��>�������g��O=s����������d���~s�y��^�έ;w�y�[o�,�l!c�U�[M|j�nt�
J��dxp�q���,HNL�=����
l�z�����;�h�Q��ΦC;���"nx3���3�����^��H�Z�� �1a�B�r-`� ��o���О0�8mX��B}W7�m�\Ӵ�i�̾�졝t[
nd�uTPJ5���>oEN��Hgt�軹AKZ|[�{;7�V��������$����S����ީ$dFc��_ߵ��	�e{���<)|��6��t>��?������m�<�[:��I���+7e�c��u��1e]�VmhCWn�����MJ%V���������o��Ak��Y9aX̭Æ�Oh0���iPџl��d��PI�g�OM����s6��X@�&��h�qoT�z�"��&>����eϣ��t�r�50O��1�����oF@�֏|.ZR�AO?�k�QA�e�6��j�a�8D�m�����q��A.w.(j�~��)���w��P��paZ*���2]O*C~�L��6�-3�-c�3O�V�l��������	WJV�V<H%��P�ɢ2y+�+V\�h_7N��G���g6Ȧm�����frj��s��K���An�V￻u�K?}�O��zp�gO��{���ͤ��~�y�5�[g��07"�rp��^�UEX�/�I⡹1�#����E~���,�zR������jlr�w�m���Sۿ8����ڙ�d�Q�e�6�d��B4���l�*��&������^�r��k���i�JY8���MdO���M�zi������d�u5٪��j�~���Y5U4���L����}���eN=��Q(~g��X��?�e�ESYJa�j�R��zf=��.-@  �~v�����c+��={�����P�v��u�n�[����g��}|O�[]BA%��[������,��<7l��ܘ�0�w�qq���;L��i��V^����e��ũ���nO{���ՃŌ�'�S�q
��u�e�W��(��}�����k�od��bQ\`�)+d�xӦ(Ie���Unl�ː_"�QZKG/@QD�p&�,AO\�\��(�����b�F�9�H���̡lf�M�ƿ�B��C{���y�;�$�-{�FO�נ0�Z>d��T�
;}���y y�$&z�*cCEC���U�O��&3K�'�c���X(&V������N~�nml�SU��Rъż&��*�N\\6�/H�%0>1���S���c���Sq�KW����	¾�7U��ٜ��i�,�޻S���O���۽{��O�����J�7�݋ݧ���`���[6ҍ˅��R�����.L�bp�E��4��|�Eo�((K�	MJ˳��O	lL<1�`6;m�֓��mHi�^��|b���f賱֧L�
l7�v�&��vW��F�a�~_�
)��o�����Ll��'/����v|rfk���]�ز���(g���}�����q���@�ҫ���;�Y-[�Q0�x��=y�J�}ʴZ�lw���[ۻ������R������Ǉ���?=֔�MF�d�٭���E{�쑽x�L85L{�67%�������s`�
L�����[��C����ྮ��m�V��������za�^_�\*+��׼�K���i������٣��53��2*����W2$zNP��b��4ذ�u�V�xz����R�0H[�T������,��+�R&EO�^Q>#%W�����oJ��yp�8JWB��rm4�0f��V� ai��I-�x�S��w�d�l�R��^�zMݮ~Ǭm��l	n��y1�&�%���+��D��x���!1p�%��iT>��彾�_|#܇`8MR�?9�BH�3��Ԭ:q����۩���E��	u�\��C�D3�ǃ�`2���3���S{L�m8�Y!#�n���rI'���2����M&�y|�\��nm�K_}����O?s�������W����׻��%��ſ�x�1��APɠ�&S��M�de�@pSO@^wE"�qr�`" qL9y{s��"�e���xO�W�4�dl�6���Fт���~�n�7m=Y�).��;9>8�����5[��5�F�����>}bGG'��n�\U��^��h6�����)��������Vϖ� � j���H'��Ų��sU�Z��|6�fk
�B}�Rٜ����Sp��� �+HO��۪�Y:���/۳gϴЮ_�f�[[6��=�{�^�L&+H�J�h[Ud���yt�v�B��T��jkO�����v��#a�nE�@3E{��]�{����gO������n['�����i% ��L�Z��J$>�>_�̺��:}e��|��u}���q�Z�l��ғ1U�X2��D!�jp�3.�E#9D�n�����x��Z!��4��u���V�L� �����Lf(�Cp��*��+���\A)������#��Ȭ4h	 �f%���Ւ��Tt�O����WN���1�I�t���?�}�<�kZ<n�lr޴d���2IZ%�l�ꅲ��ܱjP��������:�/ټ��};l��G/���TA��%�9�U��!1Bb��bN��Ap0l+���V�Fe�����/���w?������T����L����ō筦��ܰ���0����b�}��nH��|=�QJ$�+��o���YR��Cn$YN5U�	(�G�/���A�&����k������,�tO*m��M��@DO�
K����4}%�^2��/m���:���nn����j�DN���2���틆Đ�ښ��{�n�6�bN�o�)�r�"`ϛ++V.�,��Xo2�������)���Y>�e"ŏ��P�L�X4��kkV�0��������+Q���^�,�un�g'jēa0��	p�HRYk�έqv&���ښe�EM�����/�X[�)J%M�߿q�޻yW|�.��sj��ߴǭS�ȑ�QZ��+��+��6lw��G��hHB�Lm��ٸ7P BuT>
�Y�5��P�W8-�\
K����[i�b�M(P9�sPjP�e/Y�ܭ�
{���	�����<0��~�28d�N��;�E��RY(e�P���:���b��(���C	�ó� ��lC0|=�-0�� �~7��|T-�I��n��$�LiE��n�L��,5���i��Ya4��$a��D�P%A�i�ه�`�*JIe;����ϥ� -�y1o�H�!��Z���abn��2|�����5�Q�}t�����៽��V����%���o�x�n��~�H��Ʉr�Ӌ�V��� iKӀE�i��.�n<dw�* )-i$��go728hX�7���_��fv>�ڣƞ=9޷꧅�����C�%�Sy�-⟺&���̊\�糱�_@\��-&F}I�<}�\e�c׮�fm�J��Ok����m������?�ݏ�    IDAT��sl�J��ԯ�-h9�Z�t�"�Bl��ן�ub���E�ey�U�^]��8hm�"e������p>g�L\�n��P�7��ڵ�i�M��Хs�?�MK����tfG�"ts0mno
��9�o<{$h,2#d�y������Z>Q���oOG�}��|2�pS�1=���tz��Ï�sq.!�ב˦��_�T������Lq4������C�P�W��]��jYN�(�LȄ2>���v������ԱoHt�}��s��ÓЮ#(RƓ�!N�)^�yώ�}|]�t��J<�%KE�D��dT4��De-��A����Ofn��]�{��NY��>j1�ʜ;`�U=��)j�d���C��T��׭� "��T\o����W�x��4�T��0DR�A�)�6ۓ�u����!x=~f!o�\�0iF��B%��'?����n�
�땕��������Sn��<�����c�L�_�.n��l�}a�	^��/UA
ٌ�֪��Y����An2+�d�7�w���ɪ��������}k�nW���@ے��Ɂt���oQڅ��I8 �����.��k�_��$J�q�X�f«�5/���L�X�Z�nׯ]��lA=	&���Oͬ9٣��;x.&��tz-SP�x��%����"�U>��vl�qb/����Œ�^�ت��	�x�;Q�΅2B��{~�g���
n7�w����0I�@j=ܤ����z�H/^>a͹+׮Z���W�3���'��t3.Pɖ$���7߳��!�ԜtD���G��`�u�|$��Eo�`�h���葍�=�����T�o�խʐ�P�����lw��j�a��g~A9��)n�Zm{��Lw�~�ǰ5$�*���%,]n����)<w)X?W�|��=k������ީo��E^����gM����#�L2�%G{�w�A��Pp���7����1y�l�WXܖ��(O5H&<��
HX���.�LPP�-"�y2�`���K�!�%�0��O���O�����I% ���AS*4�TJ��3Tq��1�1��@6��DJ�T��G�*�_�Ͼ��o&���o�H39���^��^�#O�J�����V��hj'�>
4��k�d�*�5 \w��E�^A	Z	�D&���d�:�<���t(�Dq��hel���/��&�.2L@��¬#��J�
��[��&z����Sm(��L�0�EE[�'�*ɤ��=;���e�e��;t��f����)��nyU<�Z��^*g��g~�{a/ώm�����<s��U��^Y���8�lzרp4�62f�"���A��:L�,a��]�o�ݝ�V�3ov̗6�F%f��ؚÞ=|�XN�4�77������.4����Q������œ��ݱ��{j�����u2�� �K
)�h�ƅuON��՞%F#e�������BS:���-�iB�S�X�B�6g͖Tn���MA6��ٹs�j�����n���VP�V����{�ܔV"�226���0(�@�n�Q�COL_�G��9�/ q��;8�����h���@;tR{ 6�+ý-�0�~n��T3��ϋA5NKcp������ z�ʋ���	{Gz{�Sw�S��h1�E��Nl��I �i�7�~�).8�f�Q��}�eQ(j�,!Ӕ�$��)2ⅼt���[=7�U�&��zꗯ�3V�aT�~�������7Q�����o|���$��{��p�z��� j���~!��hܳ� �ɎgpLK@C���ݟ ��H�i�G�"糺Qh\1ES�����w+�R2�DF�*�Z�s�k��d�V���d,��y6kyyZ&5�d�X!���r�j����K��p��˗�PNE`�k��Bߧ���w�۔we��%�̔{h��ȕm�P%R�N�����u�a�D9����K+ꉬ�V�m˄�Y�.t�Fۿ8���c�L�j�۸��,��߲'�׽��I_��b��7k��Ǝ���=;;�
�^iqA 'S��y2����u�N�w~n�t�6V���ή� .Wl6������yOFS������<?��GGҽ;��P�P��c�[[V�ٲ����x�(�eJ�``�,)8�)HE3ᐹѻ�ِd�B��|��2��@$��`���ܔu���Hg(Cxb-BB����xZ�
As����yp#�� H�L+LV�{��Kp��P�W����i�Q^^[�v��s��Kug�G��#R��rF3A���0��{e)�B��L�:��2�e<��]!yz���~�A�T%��u�KYe��+���v�˿����(pC~�޷��Nj���������u��r�W+�� nk+��q�����2�މ^�2�FzZ�|	��TdH�x��oJQP�G-�&�0`c�'��T#nzy<���3����66���@L��~r��5<�,d��JZ>�����{�C�a8��2�$�
,Ӊ#�	n(w�n(�rȣ5��  ��@��8 ��L�k�^D��Jq����h�R�g3N�W_$���k/Ϗ�=�^�R֡�x��=�C
W��ȏ�RE��R� jپn�Q �d��d�������3k��x��a7vw�R�u}���uϛ6도�ÿ��X��ֆ%�Ee�4�_�ۣ�Wv�n[�����6��t�R��U�.��^2؊�3��d�72M2y`M\=3c={y��Xֆ�&m��8s�5��k�ܖKWk���I��-�����Ջ JR��pp��\V������G���U��n����<���Y�� �i�hm�Z�
��0����� ���o�#����w��dқ�h�(��͞ڠ�'jGUk�čj���\���_x��?}(�7?����~�e�y�aK��[n���s�,
�fD�+.4q�H��X�R�B��)� �Ç�3��^� S��&��FV7�4F+q
��2=�I��_��-���E��wx_N�Мv��Ь���4��-k@�%<|6�Rz�B���gs�;�=�$q��']�&��	)��:��)1�ZY~\_6�.V#�	ƈrj0=6�g�ڔۀ�O9_�s�2;g�%�&�Z`�Z�)�`�l澱i��E!�3wK�.�������l&S]�ܺGG��+؝k���R��Ǣ������u.Z6���͇C����2+�n�k2��'��ϟڋ�#9���5۸q�ҫU7���ܝ�����x��~$�
G����0\����^!�$�*�G�wKJ���bƶ�u�;ۢZ����2�͗�c���<^�p�XJ
<#�%��⥠� χ�����%r�t糀!T�($#*i��cȒ�x�#����k����q����=R���F@=I̠ӱa���G��dҮW�>����_��|3�ۯ���/v��_��]����B�Gdn7�C0�-fnL�(����J��dL�K��ƓџNtJ��)�D	��Z9��]�	��[Ӊ,�Z�!��I��L|�s�@�`��Ef&g��Z��6����sH  ���V5�q�m�Wx�HQ�l�z�f�f��.�fZ�L��o$YXj�R�4Α���u����5�p��YRT3Q��($�+2�.�c�ϝ��]�$��Dod�Sl�&�5�;��p/��aZ	r_���c|?�#�����=4�l�Z��ߺmwn�Tߓ���ɹｲ	�2n5����v���=�1�~m��v�,��"���<�{/�˻��vc׊����C�g�M)W�5n���j. ������æ���e�8�:�| ��O�F����9�ָ^����/��9k��q���!��Ep#��L�$*�D.i���n��Czi�����we�P2(���Qr������8T�SoK�"�����4��W�!#%�-2lwl�i�`��YM��Z���W�����O�}�Z)��{��w^t[�*�!�Eb}n�<P�� ��` �x	ntAbp��wHi;'�Y������.C�s9e�}T:��S_dA?�HTQ�i��W��O��C/#��c@^%��F't������ד]�A�Q���U�?\�g�	���� ���"��h���G$�+�I�~y����d��?�e��+����Fb3@Y�u��@�Jd�D%yVp��F�fP�:�>|a��~�k��N�}ї������ū��ڼݲ��U�»o�{o�U�ot��b'��3d*c����3�Cύ�v��;��{E��?��=x �YP�U�^q�s�bz;��=�������p8����r%��:MNAHA��Cv�9_�VA0��ŀ(���I����q�iMj����������	*�B� %�IL�إ_���:��X�k�-`	Z� �yJ�4cŢ�F���a=����ٯ�=#��C��"X=&&aD��̍�k%dn�g��9�Q]���捯�������_�˙���+�ɇ_���<�+����^��
n@/<t0_��Fp�8_�VZ����$*b�R"�SvG��G�o4�U`�M\�%��ZɾI�pSq�̐����দ/Z�����m��ZY��!��g'=3~&:Zj�� �R>�Ұ�>���1�]Dk���`B�h]'}pH���zM����QFb���UpKӌG���1��鋦�I�.�!��ӐԀ�ޤ֦�_E(�b�/��S��������(��͊������O���9�Q��]���;�{�>s�m��v�����O�uz��-س���4�����{�_\���Ͽo7߽+�>����c�F��%��l���k6+ᰞ�YƁ����:���+٥?L}�\�E�_��$<p�W�3A�c��Ob�X���=�p�}�z��kn���Y����t�	Ϫ"4�@�,�Ḟb�KҸ~����D=f^�1������E��bJ��g>'TD��M=D�<Z4��q7Ț�������� @J��;b�$Q����e�vce�[�n_���}ǟ��B������{���^b������}8��t���̓��J�H�U�ג�� ���Ybp�&�nP��\.�7dqN1��`/$��θj�^%�[�)J�59���P`�3e)S��ēe�+�����\jƬ��C�CH�lU�y)�����]�pJ�ᩅCp�e0!��P���R���F��oi����%����7| r*�ۚ�G"��r��@��B�w�l̠������"���e��n�l��{B�^�Au�`3 �V�����疄r�HM���[��}|f탖��ֿhJ߂�`L�g
n�Q"[>ew���v�;޳f�o�|���{��>>8��0�p�nZ�Z�I&�iZ,K_�ܔ	�m�33��,(
4 mRpx�@�*��R�y^�F��$��	�6�qd��� ����$s
%�4J���*�r`:�gnq»Ȭ�����%ʕ�WC����дN���!H�
K٧$�F�T�x��v�&Ke��h�-��AIK����&��	l�V�R7��<s�ƻ�׾�s_��O߷��k|�[�ѯ�L����x�m��L��<d�p�_��m�Z�M��-�iʨ��S,N�����!�r����!4d/�� ��wA"�=��d���,0n:7�gt��4�r.�u�	�`Z�Ҩ}���E��҄*�I@��CEj�9_.\JB�GS& B�M��W�en�#����1�dqp2ҬE���{�R)����c W�����%�@��Y�&��ܖ�Zn�Ә<���3��b�0n\��6<:�D�k;+5�������Z�ٵ����:j�Fß��i�!5�'�:J�6ϧ���������Q��۷�?������֚]}�m��G�D�@1\h\�&�y��X�A�<$��kǽ'���t>�L%��k�S7!v�m�U��*�82]Jϩ̓���#~ͳ/O�o�<�t[C@���|=sM2���J�޸gD�Z�u�����]�{���� =�X[�[�5Fd�.������!�ܘAƌR�W����8�dճ�S�X��LY|��l��Z���ۛ[_�����O�����[��}����Ѵ�|K���2����� }<�X.����U+=zI]�r ��8�Ԋ�B��>=��s.8�+>��&�JЃ#������#HH�؅����b��喔fy��3#"��x����M��Ұ��׬�b�.'��bZ��`�MP"0�>���K�.e�Bb^�e
� �G���H;\�C���Ү�e�%;Yn�<�&�9��X�Bh�G(L,a�����=ٜ?`�0M���wtj�W{6i6�F�n��}Ǿ��w�]?;����5�N�(l}7hq#�c�O�jEKW
���[v��M;h6��)���;�V�n���6�&m�v5�jy����o*�tA��I���I��Jls0��7������u�� �5� ��*'�����F�~j(���m�����O�/��ƀ�վ�ղ c
<"ԇ����1X^քQ!��!�\�f��&��7z�E|Ո��d*C��+�b�Z�A�x�$�!3��j-���B���T�
���z]�6/�yrf��Ȫ��frv�����/������܆��h��.��^�i]���c!�fc��V)[?�lF����m,����JY[8U"R:��:pCV��6������ƿ��}E9�M?b����22�%h(��5fz��U^��Q:�9c�L�\��3N�������Q�,F��!��{t���S�#��N�O�`�e�^3?���"�����`1�)&�l�2�� 	�u�^N�dY�Cb��)�H���3;y���ggv�Z��o߲Ͻ��U�%kv�l��Nl�ș��6)�MFC�������m^ߵ�kW,S-۫�c��o߷��{`���77l��V��!�xA��@��b�L~U��J��~�2���A�L`�`4�X�`4�π���0���9�B4�t<�y�sܴ�CSeY�S]�1�����(�,0�����U!�����4�X�4�����Fp#�f�E�a�}	ؼ�>$>�Jh���Gց��� �X�|�2x���Y��N�VRܣ}��J�$�?�ҽN���;?<�$�-��5n_kc�K�{~��bL����c��~���<������'��=s�M�Q����6�v|�\�Z�l�\F���c)�pbVG�Q�o��4(�ˆ)���nUl �������e�8�W��IF�b
�I�.!{�Âۢ���~C�;�|D@�� P��AZY��`26��K�4)�1�d}���O�FD�{҃���
��g�u<4�cpW�ʧ�-���侄���_|*K	`�ȜC�\_f8�a��Ξ�s;��b���\�woݲ��mˌ��:���k���l8����ӱ�77�Ɲ�v��Y�\��;<������gr��_�j�wo�����d�Mh������~D��&��HO�� �}�@bK"f~����ʠw�����L���<���±�&{�)��*��Z��B_VW�G��<_>�MH����߅��⿝����f���2�K�9�����2Xv>m��Ot�f��>��=��c���.g������&>1�9z����8�����p�W�{����;�������}3=��ѷ��|6�GG��_v��-���7Ce���JE�~��Cp������N'A�8��P�."�aI�A,��5}2��p_ �f� ����6�����GMl���&����"f.ң���� F�C��c�B���+B�zk���%6�>`n8=J��5Ђ�LB�t��K�j�ZBp�%8��{!�r-*��n�\��Q��3��%f�.�,�2S������Ȧ�d>mw��Ş��,?��nm���ݵw�߲�|UM}TB����8�a�e=)��Vm{{ۮݺi�ׯʆ���P���������Œmߺn[�oX?�SdD?)�����a&�9���#鵮��'�g�{�ed�� {aヰ�����M
��F�GhDI�0�Jk��t�z�/+o�h@�:	�i$�+P�Q��奷`B��:�?�1\�(Gcv.�Q�;�|��L����^c&���{�o%�0�    IDAT�����NK�{9���h������Cѹ�gg�r��{�������o�n��������{(p���Ϟـ���	n��u��I.WH�sٔm��(���(K!ד�)[�	��A�a��a�-���&%�/)�.�C-��K�-D '@ؿ!_ȱ���S� ��)�`.��ʽ�3#��ǣ>��7�`x�8���<FJG��E\�M�gL`�Ld��fR���?�l%��)f�
�K�����׵�	-���i��M���/�P0/�9.��Ѩ3hv2�~ߺ۸ѰJ6k�k����v��!-~�A�ٔ9����t�v��X}}�Vjk6��%��t�Ց�?}n'Ñ6�m��v3	����y�h p�`E���@�0��x#��ǀY�1.�4
&h�+k_�*p�5qV�^��K஫����{�漃�cOX�����cЦ
tSX)����k �F��dv���,��'�'y"L��^����ơ������A������TZ3_2��ts����)�����р�ZK���45�~���؍���wW�_�����o�~�k�}�b<���Q�Ͼ�6l���_\s$�|S�ꕊ�d�M (�5�Iצ�*24a
��%���rOA�gR������)C����?i|\\��
���@]���E�QX�(��M@�c�"��8�
��¦���E���A�}ye�d�Jz�V�-�A�����M����cQ��]Y����(=�ˁ��#JZ/eǱ$�����6�g�p�����	���+���*1g����u�ʒ��D޾~�n�^�+�V@�+�p��WKTB�=���Ɖ=y�Ҟ�|a��^�)x�\֪�;�~u�*�����1cc�C*� b����db/�R�B
o�>��a��u "���C�i�(���p�	�(V�}f�����KߌCl�8Pp�wy@ꀉ�~i4ٙL�Ճ-�R�Bo�C1��lKx���ˈk�ZY�f�,�c���"k�~ z9���	h��%^&�6
b�>:�+R\"Y}N��CA�2Y�����L��@n�^[�����?���������[�?|�1������;g�n0�D7��V[)_���
�i�0(����?�=7q�B�_g,CC� �:=�������U��ei��2��9u*������,��!����v,P Y�g�B�1@N"�1�;h���Yc��_���L��Q4�q�� �Tt��8���-�/���%a�*�z����m\_���w	ЌX<�v³
�zra
F�IT��u��:x� �*n*���e���H���kW��΍[��Yw叄����|��O�2T����e�DS�\����v���* os<vK���������+�'����c���$�"BVM��Nc���B�`Ʉ�ҍ2k��.�l��=F�o*%��{�\B��D<�*h �a)�r���_)[�a��Q�(`��P��e���
�:^z3�->�����Q�Őt�Oh������~	�!�f1N�I
�풵��!������oPia>�
�M��Z�xxgm������O_ύE�;��9w~e����dn����g��T�e���)[-�4-U㑑5zN�U�%�E+bc�o�(f��i�J���ͣ�E?�Er�CRf�Be1޴es������2�t�f�hQ9�xh�E��)�xH��<<(ʘ$���(A�D���IY
�)p27Jt�^�Q ұ.], B���o�,�`�E�/ �������^���q�
�}�����̘Ž��-�"�/��>�\��+���<8�&�Ε-�zu��[u�y��|�8�B����� $O���
n��"PY�ش��W-�|�4H��/O���A��z�[>��p��t$�F�����@.�������@b�r�e�@BPQiK=�el���d��9������D�_@�s��S�Lʮ+���P�v�-���C
�D�)E���?������C\!��+"�ju��ʩ�3�P�K�zAǋ�"���}�kI�+��̞ܒ��K���A����2әU�YqKo���nm}�o}�_�_�H������t�?�4�E�̎�7�S.xhBͧ��V�Vv(���s}��-l�� P�<��c��ʦ:C/B=2nZ֋�<�U��K�?��MҠ����4��o� ��G�
F�yd�L�u.�� �%�SS���=�X������&%HJ�M"�$�,�4��zw(���*$�45������Ri�����&z>����������eE�/���@#�$��0��f�a��D�)�W�Ҥ�#k�:��}\�mkc��;�
n�ٳ��m�t��B��	���	����{2�)Wk���mk�ۈzO7eγ*�����F�G�CF�+}�{dݐ��y��L�1F���Ñ�;=yAH�k�'FP����L/���V,S*Xf�$@1$��̤�t(-�]��׀&LK�n6���Z��p іp�\ē��Q��^Zڃ��X�Z�	�'��Ik���8���
�A|�6�7V´��oCG�Cܜ�+ /\�%U����vvp�~-&�8�ߨ�������������F��o?|x�h���G�������-�*p�/�a�$E �����Ven������
S;�T!��iq��)W����jn���.M>PXj�Ƒ:�(o�_^�sC�� ��Ù��*K������~hDx�rI
�\n>����F�q�$T W��=E�m�'P�h�r?������o�qPKe!�z`���J�B�/e�
1j���@A�1�8ڏ�M���;Rsh�Ee4�%�8��xb�k�ڳ�鹭����ΆK���1��yhzc��Ȗ��e�Ik���CM�ʵU[�޲����Ҧ))�6�٫����.p���ۚ����2����[��o�??�n�-E�v�S�YHbǁ��v���:_]�L�h�k;
�����R �\����?�.l�D�/�}Ե����b���5��o����Q�\88�r�>��W�QkE ��¡�8ߏK��װ��W��F��Rp������M��w�C �g �Of6���Xx��t�Ꙝݨ�?����տ��~�y#���ݻ�O~���ꠇo�X8#` d����WVl�Zu�����P	�-"��8ʝ����F��Z�,����zhQ�%6a_n1P�����ˆ��X� ����Ұش耬�H���}�:pbȀ��p�7�-�0����3M<#��ņ
��"Ǿ���=Ì �8Q^d`l�n����M`��?���D�����g�1���U|G��,0�ܦXz����liY����a�d.E޳����׬vu�V��,���X�i�&>,Io�Xd~�_�:я_�۰;���U77�0͂��*�q�(�QZ.ʦ��E&g�E&�x"N��G6j��}xj��@" �R��Ŋ�rY���F�<Me�ݮ7έC�/�KbN`+��Q:C��3�	YSQ������ x������Q��eq��!�8���� ��$��}R;�"��z�6&���3��5&Z�A�P�6еbO�nB�Z'\���I��?�,�m��׳���g&[�zV������_��?���LY�����i$���p��K��~�Zӑ���8�K"e��x�R��ZUcp��h�3�rnd�u�s����}7��!���[���B�%BA�C��=f���s(Y���r��l��*���k��ظ��)�B��
%�f�����Z0Xp�鿂CP��2;�0��>c��Bv'��^hRD5Y@T�K�-�L�,s<�x�%W<r�Or[�=�@M�����W�.��@�D���Ԕφ��pz<��ށ��ط�鹭��ٴ��
�6v$-2?�9���RM�X�4e�/����+���kV�r�V6�%�I9:I���\��5�C�>`D�sh�3�
�9I�2;�6[�?���E�*�]��Y�#6�J�ads6�~^%�Ս�䘎��i���Cy�V�r�Z٬�N�=�M�6Ce;����5�eb<��S�����A�
Ce��{lj�Kn�:Y��L6-�2�x��h���M�.�z�ڇ<�@	n�PՒ�[ƃ(,���{&�A��&M�#�8B�&&�1�����-i����9�����z����?y������K�������IDs5�������p�y=��܉�R��O�tc�2��SϘ�)Sa���?(���zm����Η�S� ��uOJ���QElZ�6�~e�z"�`�d�X(�;�t����R�$ʀ���XP�6�`��l
T�s���)���*>i9�LEb��P�ohH��B�F�r1��\:�JT~٥z9NK�i]
�Ll\]�8:�+��:?��:��ۿx�o�W689���u+�lXi�&��<�� ��l���,� w���"��Zmc�6�]�1�����i��Z& �#OWc;z>��32�.��	 �V׆gM�^�,��J2m�\�n�����3o�ֺ�} \�C:m��TϹ?�E�k����<:�g���G�3K�3�R�&]msݲ���������鵅��Ӷ��NS�̸�
���v	�mM�CpS��χz�J2����r���r	�F�A�.ZHA��&�|�c� �s���N�@�t�2OhX?�|Ђ��oY)���b�j���V>ڭ���/��~3=��x�����ˇ��?��рi�gn���R�EP[�,����	���N��1�ի�ORGb�Z>"�'��h�bAh��S(��R�`�� B �T����A�~ɴV�HȌ�Y.#g"1���-�Tl"p���K.�3u��c�8���>b(9�A��AC�u�Ӝ?E
���)�i����ؗQ9A��~��	�JV� �� �d�:����52 �P��4i �,*Sڵ�������d�\��e%�S6e#�N3�	�Y7qh<�0KI����+;z��f��hY��+�ו�����9=����F��
Su�D4�կ;/�ٸѴi�mU��J5{o����ڶ;W��Z����#��Ƴ�@���T8��hl����N��H������;���V

n��U��Lz�Ҕu�lH��x���I �j��
 @Č���s ؾ����d�RY�a�Y8��쇣��9T�s}3��K$9Tj����e�� t��1�p�D��PYiR�e�T �N��TZ*̳nOmx�7d�7�����������)K�ɇ�lLz�`o����s;v�5C7ߧ����s�9<7����@-Z��ďL�d�@�2D�X�.��1Ê�S�(<Xŉ���Xp��/�'����,�.U_��
��4�tr�ƭ �.�G0Ҵ��	���|J��r<�%ϕ�e�(A�`Z�97�1%���2UpY��ʢ��	JQ�
3����d�;��C'M�Y!���7�?k�/��w��.prl!(3\
n���in2��љ�2�<8����ֺzf��Fi7�v�L�Ge)rn�T���徂��ƺ[%��dI�vc��)�L��B�h|2:a���ڴѲ�i�2���Y߲/ܾk_��m�**M�Aw���1�\�q���NXG��L���v����\��t��V���+�ʖ)��3�\�,�a�x;��]���שHS�@u
�X�&��M�B�_�a6���-�G�3jé�;�"bq8�Cm��co8������Ak��3���Xդ%������2۴ӵA��Vsy��NӒ��/��̗~�ߏ~���,�ߺ��ab�K����?G�wam��S��T����JE�W\�[=9�S��A�#B���=�%hT���b����z���e<c�iX�����H�^V��Ȳ"4%Ja�}B���??����)fNy�|rm* �����$I����"#y�e`�$|�[�f?|�@�T)�˩O���BiA�jv���:�^�/���Opk�����H��<�Q���b.�kl��Ȇ�9.�b�dqjf���	�g�Ⱥd��{ʝx<��e��a��{��?�B�j����qmG� �	Ls�!3Ar6��,���utj���*��eW+���!��>��A��L�ik��hOe.�M�
�������Ƕ>I�F*g�s�=���>oo�\�N�a�'�"�c�S-����6K�,�8
�ٜ%s9ktZ�vf��_��q��:���
��5���-_)�Ӕ��S5�=�:�.(�(�
Su��z��!N��^������UAɇG(�q�k�Ԙ`�׀y��uE�b��>���UV8�n%g���Hi9y>t'��`J ��2��*8:Ɠk\H��Wf�<	轒��F>o�d�6s���j[_����!���x������G��_~�:M�.��*ͽ����W�@A���F�*��D|�Ȳ\~%�2�i]q/	$�`O��+�[�j����7?]P*N�TN�t:���?@%� '��q�������G����
�|κ��BbH�=����^*���.��b�J�L����^6'�9����ﹼ7�{7��:�����r,�EIr(%�5=v �C��(e�_j�E���BH���R�'1�u�O�}�PZ]��+��DPp�i��+�4��+&�)�}h�Mgv�w`G�r5���Z�VR�n�NY75�)P�� P���(���>��t&Չ�Y˦'��~�gW�Y���i����ݾ���}v|b���ey2i���]ͦs��RE�Чٌ{��X<����+;k^��yÚݦ�Ĭ��H;]��?��#�w�f��R�2{�#!���uf���P������epsO�~K9̄��[R �h�) �������e������89ȓ�%�%�����P���H�����I�o�ߠ�i@�KF�"=P�z�yBÄ�L֮���lm}�?���pK	n�I��mn�skL�b,7��
UP���b�!�6)���H�W�'�1c�1��x�pɿ�ZZ��%B|��8-�O�F�F�߇<�N�y��(���P!�#H�?�pX�|&�y	�T$l"��`�K��OT���>�.��y�g�k��ط�e��L��B/��X΋?�p!�8e����-�=zn���[d1뙰p�Y�K�v\8$��-�Q�Nj���3���9�Ȟ���-9[���N_�[���V�׭~m���Rh&��q���+������+k� Y��-�ZR�6�g�#��gY�:����U������5W��8���6<8��q��*��w^}˾��_�d(�c��Tr<ku���U�%�� ���7�������zސ�j�Ӳ�V�F@D�vS`"�T�l;�SPbMh��l2R�«����	�XC��$��f�^��0�CBa#��΄��(xQ�J��ɡ%aWS��6����:�AȪ2��9Ӹ�J�
�@�8H���5�ւ�:������j�w^�θ��}t"�[<K7��^Y{����/}���|x���x���'��st܂�rd�s�ep��k�m��O{Mb\)+����=�8���2`�t
���O-��?z�"q\�`�;�%�W�b�*M6���6��1��2D�J�(�%ˠR�dAfH}7�SL'ɘ�
n9>I;S�^��<
	��V��[�u�qC�q�<c��:Qf7��l0)� �� ���x�r���` � ggS�>*�i�Nl2�R\d� �$!àI���@��Rޫ$��R�A�)L�
�Ol�^��[�mmg���senP���2 �Iijbv�����S�y}}�*����n�(�i~��9���<q٪����/Isx�`l�Fӆ{��k��ݱ/�y�n�n���vzt(sh̎��u��Vk5����� �ƕ�S���	i^���hbpb��s�6Ì{D�S.m�lJ"	4�a�`|L�C����5�]*�� VI0+b�]�I9���*�a�Y*�-����?�ˈ�J;��M��1��d�>Y��<�l����S���tgؚ�̥mF�W%��Fc���$ ccVD?ήS�!ӛ���[!ܷ��xF9��&����,3�[�U(�
��������Ko�����ݻ�N�����1sk�'2~��Q�s�Y[]�y�-��1�ɍ�q �^�~�i�ȶ��E��d���    IDAT%xǲzO�� ��zX����ô���\��c�M<�CL��,�2B
���(�޴e�'CM��Wd��I+��V�:O�L2$k��7���m0���)䊖�h �@RtO�D�ol�^�� &�W:m�NV,b�H�ޥC�(H&�7�1љ���h� ���NF֙e�,S�ࡊ�=R?�}�;28�%�pe�A�]��Pr��,㩥(�)�jk  έ��e�+���4��Ҭ#{�xi��uq������Փg�B�W�l}g[�3�M@�rz���ax�b27�	��KYy4��ѩu_Y�ٳ��;�{���` �/^���
E��*2/��Z�^�r��y�����Z�߷��3�h�����:���_<?����G����+d�V)t�&���3�W����1�D%�Br�(�*��e� �^)�J��k*�
zO����rYK峡A��A%a�t�JlKkvX;kw�9Zk4�TK ;���ƛ��)��V?.���E�MK����Oң��d5!�9�١D�C�	�OC��Pb��T�6�y������ͭ/�ܛ����\k���h���g�$���t��dgSvk����rU�8� ��pWS4�2T�@�K��EI��[/27o]F�c�fC�z��^B:�z�8X����(2< L�q�,�����H�f��mVj�^�Z1���ƹ�5,X��������U�y+���X6�'�	��U�z`����0�$X���W�E��8��TFY�;H�3)L�7,\�F�N�6�m6�>�w�5H���ײX�"oN���o:�b����^�&v:D|�&��@��o��L-75����N41,l��ʕϸ�t �$�x�"�Ϭbi+'2v�乽|�D���zݶ��X�ʦ�)� %A
J}'-G"����L���y�f�A�p��Ƈ�V�������}~��T����.έ�R�r��u])�ʹ�����JyŚ����G�������ҧ��6�ӒL�8��e23+p8%R6L�6�J\Z�U�>0��T�I��g*m�l�j47�**V+���Rԟ�H�3����>���;�Ǹ�&�@�&Rf��#�h��E��Z�ױ�f�·I��(6���l�d�BQC�d�ȇ�VM>�����Hj�)�L�>�We�ʰ�=k@���
ȋl�n�k��޺��?�?-��ڿ.������ÇW�����p��+O�'��fc��Ƨ���e*�mu5dn��Ud+D��PS���� UM�X܁�A�Z.G՛����g�IQ��
u<�x�OqA�5$�p$�lz��1�!��܂?!x�:I��ɰpߞά`�8i��n��������t58`�II�� 뢔�4NuE*��RK �	��M�f!�������dp��"�^(��ZD:��\N�R# �� ���U>4�=���"���:ӑ�㛣�����K�u�r�E���>��ٱ��^�����\���əӯN�mkk��;u��3��R����#��k<��<��~�8��m�붵�c��d*K���:��IFJ]�#��;����a�f�vr��Ʈ]-�X���c�i�T��b!��<��gtk'�����8<<�o~�=/��A+K�Dq#��M'*,M�!�a�+clCx�T �=)PAd,K��y+���5uK!�V�K�J1g����V�V)��R��Z�'��"��[�=�K��!zod����Zdn����{v����E�Z����c�M�Z((�3��\xm�B����K9�W*6�g܍\$��p������x��`s�������QI����;�W���ߏ����7���ۯ?x�s��݃A�=i�������d���y�):BA(���D���U
�B)�K\3*�/�@���ר��k�ޫ�}9y�����8/w��.�
$��r���q�Jl�ғ�{�f�.*H�3��%s�C�TɲVN�l5Y���v��i9zOé{]��V�笐-H6�EE��:�FQ斤w�ʦRҠ������[��ݨ�SsU
�tk2E0�8���.U���tt�P�AV�i��:}.��%ď���=ꫴ �#���q
����M�Y�1�zt>P���s���Ȅi'F������i{w�j�V�׬G��7��9�!��:[afVIe���{�̭����k
���\����\_Ӿ�=&���6h�1�[�շ�q����Yݲ+�T(�J�C'������+��ʦt��
`�����h4v�޽�lA�
%2�R�P?�Ih�Q�F㞳HT҈�f�8GW�����w�r\-8ZD����I%Xo��Y����r�V�˥�V.�m�\�|!+s9t�J$�� 6����l�T��L�?��2�s̳[=�����`]�J��%2�w^�-W.�k�P)Y>���}1c��$?�i�ܚ6�f>#C�$�t�`zhhTL�ܮ��>{o��O����;Ϟ]9�������?m���_�X/��Q�T���b榆�z5#97qCT݇M�8�����Ş�ņ�ӯ�\x/���JQ�6� қr�4'�z"t�u�?���(y:;��f����P�w��A��6�aݞ��
��md*rU�(T����x8=���ɸ��	��Kf@#f�����E�o�S����*��	�v�c�aϱB2�ť�UW�`^6w�\QpC��+&xm�,F�ܒv
υ	+Y���Tk:��^�.�;"�9�1zR���Lσ�I�c��
a~<��{��5U�n޸*U��q�� �{n���wcZ:���v���5�Ҁ�˧um�9�x��:%�M��sj����gM+��v��j���3�.U$���u��m�� ����D��jY�?�~x�fggg�p�`U�#ę���LlZ8��Mq�
�|��)9������AL�)w:z��E�O4�LNY�?�Y9�}��N{O�TT+D�R�9�N����1���|no� �m8i_��3�&����	fꕩ�
A�
@��Y	\��
���W�V�	��r�晜��A>m�b��oy�yd0�8<9V�Cp[Ie�����w6�����27�������Y�,��uf�\J��(%�Z[�Z���$��G?aJRN���WI/%R��r/����R�P��!��`d~%-$�����@�9�>���d��h|�r�)�ԕ)��POe�Lp��,��m�PUp[�V��
�4��P��B��B:��Nw6*��� �ٍ�OK9�CZ\h�y��E#�0�0�M�~O��6Q�(�v�-�� ɩ����\AGc����c#��U&�	)n�w�-�Q�A��sa��s��۔����`�MPSF��")���������Z���a�wm�����LuY'i/-ūM�\(r8մ�a���g�o��-]�@��B�Z�0�lR)��	|M��T����<�v�捖�[�NV���&��Pxr���g ��G@��Y�^�oϞ���Ź&� �ONN���H?�P sJ�{}�ӱnD�=5�(p�="ecJ^����5���pZ��%���(q�)5RR^AV*�z�E�4aʹ���B 0�eq�6��G�Ɓd	�ѝͬ��e*7��G(� �r��5�	V�j/ŁP&���z��ڊUkkVZ�Z��f�"�(yW
�^�[;�� �I����*a���!�|%������ln����s���HY�;��_9���Ѹ��=�4�7܆4f��i:�(�M8ͧ|��IJ�IK\�e��,8v �#�	u��]["�������\��$��Z�Vx�8�2 ��)e �G0%ԟa�`&ʈ��
ɤSi+�3*S����T�6
%����V�E+1k��jڠ��b���ɺ�x�M/D�;���S��dVx7M@�Ы	�5-L��Y��O��& /(\ɤ�2a�8[�����$=<7l�8�.����R����%5��N��6$S/��un�A׎�m`%�i��2D>��k@��3ff��#M;;Ƕ��i;��Պ���kM�
n��s��GSKC����=}n�fG�m��U��^�Y)��8J��1?S(zzX�樯�ĝ����Z=��]�V�mm���D����&���� �wi!PV��C��N��N�N���T����3!��Y�wB��A84��L:'�Jyɿ�%x	b	��1<�&�Pt�R�ϓ��lb��X�nR6�-QR����2���O�h*��dB�}�h%3xg{ON4�OV;jED�<�IK��N��0��?�ڪ�VQE�X�T��j�:�������u��n|ur�-�TƊɤ]�֟��y�������	n��v<��$��ʎdf���
�`�ŀPe��j�:w�#�WC��4�4n���X�JF����B�Ʀ	�:�Z�'%W��0S�9i�Y9����\4]��jジ>Gb��BY���z@��np~�PZ-���m=[�j:oID�#AB8uz:��EeN2���H.W��i���F�֌r6��
��z!���@!(��^�0���GV@��W�^�i���ܸo�L(��NOtP�*�E��|еT�h���m޼���������Y޽�y�s�]�]�}�����&G��(��Hd	%�%(����A�3E�8XQ� E"���>>=5�y^�<D�����E�#�J�]�5���Z����s?���l���0������S.R0�)$bJp:����l
oNCq\\i{oO�z����݋������7A���z^�x�܅���:y�R��Į"���v�*�̓��
�����`}�V�H~����*��\�uF~�r�^�B���(��=�&�O�4�M��<�^_^s�[��P��7��PI>C�>�&)V��`Z:�8��d� �`s�����<�p��7�R�r��v�f�̦.�\����+[��ёZ���p�:Y��{�7tmKMaF�	�/�d
�عqbF��;��0=1*CU���A����*�*��U�J��m׵h��F͓Y�hp��a7XE��v��z�l�|����������ڊ[7����ɿ�|p�{޻��2(�mx�6��j�N�|��Y���]��z�����M��"i4�j��p�$ܴ�.9�eY#s�p��_���V2U�Ug�<^B�l�����ڬ{5}�����ZW���>�����tl\ J��+h�^�v��������C��b�?�I̅�Q��ظA*�ڧ�ډ���Id:������֖�{8����gKG�2;��Eȅ-R-$`�aC�!����t��	#�ƹ�T�����/]�V����T�ZE�J�7���+s���1f S��>(e£�/Ի���ޞS�_��+f ��S-T $��@��G�>���4M�
���j���m�c��q�ύ�ր<b�hWo^#N!��
k6����F˫�r����E�Sym��&��~��E�G�F�l�.�8���Wn��'�l��0nbĽYKՊv���l�+���$�K~��w�M.r�-8�u:�D'G�;�h=+5��D�����ۡI`�Yi>[j�h<Y�uq[�5烿�I+vN�o�A�����*`n���.eyy	����FGq��)U�ʗ�~��V�ZE����2��&��^�z:�������(2���v���_����^[q륗�j��e�p1U����0��e������Vf�pAc��ѧ�`���J|���IcĴ�zt{��W�A���En:68Q�:���v���U�蠒�2�r>�Z��� ����N{]�&#��b����%��FL�- %�wXRg�-����5rZy��PI��+Z��-�`#�H�8���8l�ӯ�$"� �=_B#�> � Q�5�E��[0�LrF��j�>@uԍF}0ٔ�].FnF�ӫ'cwc�N˧7d�|��q���aj�>�ijm��@����/��g���w���:���˃R=�͚�:(��ʭ�>�?}����p��Ζ���U��xc�g�.��U�ͻ!�d�����%�':���n ˫[=�������խf��F��8@������+`h�����y��&���á�D��w6���JV�%U!��h��3p���]��[2<����<䵔Z��Ȓ�b�k��ťJ4b���ឤpZ�J�Ɣ5���Қ���.t<1y�bF�-7.����@��:D1X"�hOVِ�ˢ�[᜛�r��<&%6��RU"�'WT�VѢZQ�U�׼���/&���OM����REq{g����O������������/]-ǿ���&�7��G
��V��v�鋂Ԧ�r�غ4�(p�Y�=����Qqta�0;ڸ$x۝� �~�A01��\^;����5��E�kt��T`�Z�� ��[��GR<��n��3b���*W�,��кQ@5�i�)�\�)"A7Ͳ!gAζ��r��~�:�~6�o{�h�c��>�К��Y<��d>t:�R�H�D����8�-y��DF�]���7B�"a�1GFQ��c3��sC���M�6�az���)�kTUh54-�u3��z1V�Q>R3��=��]�������7���k������G�a:��r�m2:����3M�5�;��s��>0��^Ӳ4�Ʊ��sc�DT�&���B�ۑ&'z\mbi��٥�X�.������L�9�6�n'>W/s80���!z챽�/���;+WJ��:2N���*��>&PQ�x^���!�N�HG/����`L8�z��z	��-}H碸��c�kF��,5c<��Mo���=d��`2�-����xj#�2˥��5��i��,�iV�J�R�r��^,�SQ��P��ЪTR���fM�jN�ӡ^n������\*���[{�?�K�k,��~��Y�������٣Q�{��۟��Z��{��߁��'#�z�&v��
c�#��Ŀ��]\�J���YT/�	s����c�LN��*�ݯ4�](i+_1�ݝ�O��bͳY- })pZ�r8�y�F���E	�M�RQ=_��75��H�r����֬2�2 n9#"xl��.DAYh<�߂��tgA�:.F�N|:`:4�4ِy���b��*!�Y�<��{�h�����I�T��
�i��E�S��l9�6��Y20n%Pr'�{nl}�]���U�}�r�nS]�z���b]��:�D��������Q��5vw��l�A�ơ��J I"�7�N)�J�����?�[�ၚ��%h�Vt�ɖ=)�v�g�ǸeHJ��lb��?����딚��zG'�2JӜ�G!�L-YJ0��&v��H?_�ͺ;�`Mŵ�8F��QrV��$ �֖_S��9U+Gbfh���	�3F�ȕ�����ɩZ`A��s�Bv�N�Q�8}�QU�VU�k\1�l��	��L:{:���lK�T��ӹƣ��l����nG�w�'S4�ge��p�Ԙ	�,�5ꏔ�t�)�0*��ރ|��r��FkK��m�;��mwpjT4�t4��]��L>mX�A�u����?��~�����ҹ�_Ϟ�],F�l��/{W92�٥G Z u�Ro���o����)"�î�ݜ�lt�.�}fcd�ZG�[�K�CmtԵ�<NQ�n�*�]���	=t`�P�꛴�rE=,V�����ZÂ�'I�[�������`���9ԟL����M��`n� �v��ra�{�j�|1�1_	��kLg5��5����bv�c`W�DN�E�|��Ä��p��V6@a�׆�M�����8�1�-["]�5�;:�@0E� ���.2.��*-��M����K>��nW71S�f�\�> |��U1����7C:1�/�ya����y��;�L��g\������# 8*���Ͽ��O�i9�������=s��)��V�E3��\踾�S2=�������L�5��ղ7�Ÿ��fk��c�{}�Y��2���<װ�2]'檺�`KUx��
����h������?�	<�K���F�������a^ʶ�XP��P���|�W)�R�XT�V�v���V]�FU��}A�$��~p�裯8|����58��-M�g�������uM��bn������ڑ��l    IDATF�"J|逧����?�tV�JE�ZSͭmU)p�;ʴ[�4*�I�t��ߜ��g+���A�����?���_�B�+n�K����`0���d��rz��#}��;z�sߣ���J���Y�R���c)]���7KqC��
��@�����3&Z��d���+A -@ҿ�+�l0��9�z�.�q��7[=����3��y����JZ�rʔ�.Bto4p��؆���-�%��M|�&!�^ �}7��=���0bXL��~���;�&H:�``ƚ�1=������I�����1�9P��xQ����r!��^GRM��_��ō��OA��KW���GV�t��hc&r�,#W���6KI��T���]�h:s�JaoK��{.h��"�����y��lC���?fm�f4u����c�<�7!�m�ӳ��c��i<�|���=a��]oiq}�Yw���3s���~�".(�������7���h�1hD<�¡���c`n	$k��֒�3c8�l:�c���q@��8�nX�Q ���e|L(����N�ZȩY.��@~Usq+�r��&t'�$�$4�����B�w�ZR\Wv�@z�Ot~���`�.�\n�!ov<���;�2�U�PpJ��1���bŤ�r��ڃ�Ju�4j�Z��r6ԗ�+����&:�j:�����o����?���������<�p�?_����{W9��n��0�ֹH����7����t���<���ӗzys��:\��>��ƺ�\�w�M1s� 9+踈��r���l�s�Jg�\����Kzow_O�����g����u=c$I�r����{*�R*0A�J�	��[MK["�|o�6E|�l����ڄ9�bЏ�Ǥ�xs�!��j�yW� �˅#��+?�ո(_�e�l,ls2����()PIԠ��c;7��d�0���K<��P�
L&�cC�焦�c�A��v��Py���I½�X�RI�3�f���k�Ƨjݬ�~ת��rD�����[�� 8{
��J�������}�˘ ����g��
���֎���e4���鋗�^�h=�X�����Z�nW�����$7���VK�rm/��z>h<��Α�gջ�j6�c�@�� V
5�����pp'Uc����c ����F���+��Vn 9&M<�1Ai�
�ze=�b�DA�{t
}��������S���kCbd0��f8��hh�m4v�c�H\��(���̏�ժ�/�1)[zOV1p����մn5���5+u���x5ыލo/�g�Z�f��>{gg������3�' &tnÿ@q{ٽ�!�eC�xӢ;����Է�xG��ﹸ_��ӓC��44��W+���nE%����\���~Ҫ�5�BB���Y-U#iF��Z��X��T�s}���wp_�Zm˟� ]�\��������hn����VgW�J%H�,�N���w�7>ӨVT�x�Mr�kE|���B �JRX�� v��J
Z2f�q%`j�r#��IW�/r��E�%9�걐M�#� tfI������<G2�&l}^Gr��_���ⷵS�F�Z��	��4vt�`q<�_@��kA:�	|����ty���;;ʳ���tzu�'G���H%���Z�r�NRK�,��l��^@ОK�TV��sg(�/����5=x�P�vǣ)#1 P�U0qOGR7W�Z0��mo���\]���X�^�]ܬ7�0i���4����ļI����ӥ4�)�G���ҹ��d�Í�<�]��|�@���c�ό�yl��l�Mc�� *,�q����J��bZ��m�h��l�����j6�v�0�bI�R�m��Dn��|�$�dþ*5Вe*����R��ܘ�xc<��q���a�����X�UJ��˪�.U)U�u.V���r$�U*��j���f���B7����}=�:�l=W��|^�Z[�?������w�����:��l�ߝ�{?KqC��O-�s���]T7Y}����;��ή/��ٱNz�v��T�I�)��	7Ϡ�I",�hml���R�����s�W�&3en��]u�����w���������N|�F]�2����֞Z�m�<4{z�e�+,���}�U6j�^,`-��bθX����@����P��Ů�R����4t|�ڇ�#vmM"}#)R���(����tݠ=Ei�S$/�~�CGyVI��8��������L�����}k2ICφ��߅�i23&�g7��m�4��(�אׄi"��*͖N.�����=���(��Ъ�����Zj �L4�i��S8��ip~���S�&#����uv�T�j��,g֨�!ڹ"ʮl"�
��V��F��W:z8j&�Nf\�j>�����D~͔%c�����ȃL
���ʊ�
EJ6��x	}���U.��NGc����{i�
�M�n*��B�d��riOh��ڊ ��1�d�3�p�I٤�A5��� �/C��>&���Ɓ�������R4��MQ�~�.�I0���s�\�wqkTk~��"��-�ku��U�ke�y�汈�.7K���P/n�5[�U�e�*�fk�˷ۻ?�'~�5Y�ڳ����/_��?�t���ōu�f23���{o�?Փ�{������ͥI���(<fF�$E�i<�,�,���t���W&dR�36SԠ�..�*N�J]w��KUGs��h��ֶ�:���f�I���?PFӝ�=x����0��`4x�U46��ɘ��(�CM�x�$87��X��z}�dDD�tHN-�~���b"��T�X߸�=���9O"k��%J�d4E�̩o���yͯ����������!�x�y�&�󛍱3
�����Ύ�!3���Bm�fП�tj����J�m���������~�}o�N��,��ɬ���5˦5�nt��z����1w�lr�R%��zcO�I��W(��lwt��C8��7�IG�cU�l��BH����5��5#p����|� �E�%�D��TL��ύbu��./(T�Kc{�l5[�J����ت'���hhY�5���e��v���-��#��%�Ю&,�ت��Ce��B�5�T���*[�<�==�6��>�1o�����
to�[��w�+��o	Gk �JDu]\>�.<�K�[�Q�ĢzE�fE�zI�RQ���b���AWG�+�5�v)nO�[/�lm��?�S?�������ۻg��_����{�;u5X�ܞ�=� ��3zo�~��z��К7nH��*lĒ�����#���ѹ��6��,6�$�--��׃[]z�F�S
��S�ϯ4q������E=h4l?��l�La���0[.k�࡚�]�M��hn�Cwn�z�ap�4?����<��nGc�s�(�l�f�E��[.��ᱬ3�R����=,-��,���'�Q/��K��k-��K�/����)�ɲ�K�W2(�-�/�c�r�m�郅_|O�	�^���sP]0Q�2�#�Ya��tg�5�N�wp��i�qoV:[N4���^���A���R�rA�4��Aci��������Z�>���0�	v��w��B��T�� ��C����^:��*���;�9 �|ecz�pӺ7Rf8Ѫ7r"=KH�[��c��[p���z��X09�w�`S(Df����8
��j5z�N;o-,�S򙅭o��� �5CNi����\N\A(l��J��`G@$�is�-�|�/e�L�B ������^�!�R=A/��*��m�뀶2o��_D_����r��u��i��u�)5�I-u��{��B��	��X���:z�����������T���WT�������=�-���l���{����F��/�Ҥ����@?��;z��c�q-�e��Pɉ�/��s��e��4^�|rY�Mڔ�u�#]���ɱ.��*u�JsZA�=9���Z������u�6�z��ox�|����*S���h�Xj<�9��+���;8[����1V8S4��#_$�����H
P�o��q#|����8.��Hw(jh)l��S�3H�d��$�.~�}���2�*�@x��MC4��8%��0Ʒ0tG����t�`s���Ł�āģm�T������p���z�@b�x�0ª(�����r���@]���e��p�l���7���R%l�zC��c]�!��J�j���*;m+$�����U(+�0y,��[�� �@�	dcwX�N(v���e�%vG��,���-��w��י�8-�
�����3�'$<���ó���l�M��茭Q$P��9%rQ��=�-����b��&���vqmA=�^r� �V�Yc}	�F13�ď.oΩ�2H�fPB��0�A �.n���A��?ds���E.�A�sN.��;7����F�m��ۺXҬ^Ԧ�T��P7���z�/{W����zt�X,�U��?�;�����|'�����������?߹Z���t��F�Fq��EØ�-��/����y�T_��D��o���a^.� �gDp)0��	a|r1����R���PSߜ���K��\��WSj�P�;��g_h~t���0��t���O���k���㲂o6�~�ӵ:v�GO�&��*�u�2��-�� >��"vW��k�"T(6�67[��?�Se���G� �
�ы�+6�����B�+>�ŝN��pS�����{IA��%��p�Z%_��X��4���W� ؊Nq��Ԧ���Es��;�1d�G���/d��P=�Qe��ϼVŬ�thٴ� ���n�={�j4�g�)M�����/��h��ənN�4���q)ת�vZ�<<�y妔�.��l�c��q��ª
67��%利fd�x"�l��d��n�ZGZb�>���G\�S2j��0U�{�剢6�Y��^S�2NL��9�
�
K�H�t�k�4��&��mf�E-�$cuT�a����1��<��'zf��b��j2��'`
��@Dk�f�MG�h����Q�!Q.���&m#όm�J����m�q���j�a�:���6,��zE�v]g�>���G�ϴ̬�f��eQ]<����[����?���!\������>�l�������;�^��&���u I7�xX������<�� @i1�_�tc��� �So\�����8|��ֈ7��*��"��k��}�w�S��z������ҷC�+��].������R��<�X�YA�]p��r���(7lFwL4�Kiwxr0����6�[Ŭl2�V
@�al���΍��{4&���������w	7�3п�)���[�h��td��DRВ�3[_-l��	�W��е���\���x�����	��L�W�S� v�z�8����|V3���;���H���Y��C5B�y�tǛ���,ŀt������۞���CYf��P�����a��J�M��o;���`w��) ы`I��r������,��S�qAM4�,�bhIW���avN+�`X
��Z�v���bWb��k��RC��t��;�9���+4)��Ì�b�U	|-�W��W��S�\��x���򵢱�D[
�G�Yg��s����"�ko��x��|��􏉺�,����C�����(L�w���^����{��r��j�������FM�zY�뙾�]����6Q��R��tPk\>�t��{�_=��o}���8=�K���xy{YDh�-�Q$Q����A	A��F�{m��Ajn[jˮ 6cn)w��>k#�7��\��1Fq���V�Qr�������ˮ*��Z`e��;���_���}O�zCk����n,L0���a,�y�_�S�qf��Y���^W��(tM����F�i�:
��{l��Q��5L�>��oouqqf﯄�pВ�l�n\锂CE � ��p���d�`�H��ݛ�?jU������H���5�iB@�k�:#:���d!�Z���sH�8�1&�ᠡ�Q�y'*uW�:�5(���uC~Cj�ʇ�R�x����*d�<���-��g�}��/���`d�o�L����c:�c �/~́��ҹ���(�rQ���᪍f.v�Ñ�˩?_;Ҙ*���7,��roh20B�lp[�h"ާ��l�������j�iJ��=��3�&�|64e�1f��p���U��U/�\�y-[J�J^�r�!1Iqs�ÂhJ�H�՜��+��#쾗�&&���X�Џ"�1��&����v�!���]�S��أ3�"���To������ֶ��\��U��I����D��W����f��� ��h]����g^[q��}Թ�.�|6��7eS;�S� �%й�����O��Goy]Nh�秇vq��e�f�4xe�(���i�CL|��HK�2a��^�%-:��լ�{~�Ï>��gϔ�,���l�v�����?�o����?O��\�:(fr��^^��Mۛ��-�����o��ڧ�j��j�;>��╅���$:3(wY���=��Ҩ��$�h��%2.�W��牄�d�LT�٫]X��%�c�����k_��l�L��_R�X��"�U�Rqq�d�rw�PI����	�hS!�*_��������T�B�4:�g�k�,'�hU�?61��l��>P���щ~�{�����ڽwO��U�M�ջp m�9`��ۮ�h�+`G����ޗ4?{YD1������2�K�!D��1q t��[t��B����8�T�9`�tp`p��]e��#�|�1,��85'��m�����3ˮ*�%*� �jֵլ�ި(_�/p�L1g:� ϳqiK.�J�cvC�^1{�/�Ď��h��e���K����N�����<��%
��8���،�tr��
�����w����SikK�vM�RA/��?<~��z�%����ɛ{��{[����2��o/��/R���d��=���b5�%ǘA��9O�����׏������-U�}q�\��L�~��]�&[2&�;�m2=-j��`,0&��-��h�L��x�������O-vN���lC�E'�{o����}_O�~[y�+���~�-h4#L()M^��泰����m7#�H���8V�E��2tT�W+�H`i5p5�0r���J���J�		fFwh�-$�h�H����#� y��Dݤ�s�-�(��	��;�o4�L�IGI}��O�����5V��1��C�e:f��A�;M�.{p�TJ7}�W/5;�V��zI�\��|>��l��אd��_n�O�˰����=}��'�<;�뢓�wZ���S�QW�^����,>y�B���4 w�t��F��FM�̘�G^0��U���X�P����6K�$�
I�E#�28�еQ��7-����1���{�	���Nӯa~*�K�)U�� ��UԮ�`(�L�U�U6�-�3E!��#5c�
#j�)'hgIU�� ��r ���MOW�������y[��p�I�M��d-�Q�#��N���ƥ۪w��8�S��ֺ^Q�����Оn���2���I:�4x�����z�����Z���{��y9��٤���^V�I�F2ov�G�J��=pq{���UЧG_跟}��IO�RZ�R�Ft\��⚢�q���5��ؕ��m`��0��+��L���g��Ï4���f�g���o4��O����ꝷ���+�e ��}�q���N
�
''p&�k%2䖲H������ُB�`J�tN�������P����^Rm�zr:�񥢰:�D#J�Kp7~?�����$I#Od`����4)`�vo�ޫ�Ɗ��������dc��P�.�D�.2����6@��b��.3���KEq@n\2JŊ��nOǗ��ϗ*tZ�=�����~��P狉����X�[,�E�;Ś��[V��}}�ɧ���t�;?=�V�����6�luڦ������G�ܵǑ�s���r�h�iB�TQ]�2�(1Ju��zc�@��#�n{Zv�>�+dI�g�Z(A(�ټf( ï�WN69X.�m�pnf����2�2��bN5�9/� �Z��1���	Da�\�v��"�RȻ$b���7��x�;�E�� �c�4��    IDAT���ʤ���Q�8�-��7�Y{����*��J5���
�ͤt��t6���s�s�F��v��>y��������^Kq�_?���[�{6�����u�bе�^T��v��o�����޹�X�lA_>���>�ɴ�~I�`�1��-�R:0&H[�����A+�� �J[��Z��N?�\�~�Cm����NVf�?���O����Otppp7�����k�w�؍AFğ��#t�nW�� �-Q��8�moo����9�3�\j��[{�������<,\La���vwQ���Q��C"q���L�����e�n�dW�.�:D'&E7K�d,�
�'e1�ş�������p���N�+�c�c�h��@�i��b����e��=�ז�l��u��l��4�ZJ�l�s��9p�B����YK�V#]Ri�sdos�V�	�7痾��q��tT�5c���I&8�B6�e�+��\m6�l���q��LNE����.~��_�V��6�ㅖ�}��W��q����L��+�G	q I�J�`��m�A�dܣ��қ��U �B�&(.�*!mib*H���R�=�a�`��Wo>�UY�@�K[���v8v��{u��f1�k���=����%�8ԓJ��%y�lKk��-ձ��a[�j�̮\P?�	ҫ�D�ӑ^�^(U��j&�{������_�����[o�O���������?��F�d�����u�i6������>j�����zzp����#}v�R˱zi�[k�	�+d�<�(�-7�v8aA�.�?��U
%��ʺ��.?}�����!]�
�������ӧ���w���Ύ�Y����\�S��|��0��	"twM$_��hŖ(��|F���vvw]�z���Ł!�n -����ΎOt����s|�e5Aj�?�1o���K˘Ƅ0O���M�L��#'�P��X���y̤�s]�]��%�*��9������<�&K�N���.���1
���)\����c$�H�ܕZ`�sB��@����d�/-�F�=����hXH�6�Q/�Ҡ ��Y�
���Kn�V�{N�1$ܥ.^���\���!��
T��;8�����gG�{6�P ���t��v!�Ȧ�&���Ik�#�9qK/7gifC�6<�Pz4U~�R��t�!.d@P��b0�D��c|�/���ɇ�5A)��İ���F7��J\���l�j��q��0�<@��ۗBO�dk��,�L�
�s2�j֨6���R0� ��zc����#�o`fe��4�Mכ�Z�_�J��f$��2����#��by�.`�sqۯ��5�~�O��|�&����*n�������NF���tp۸�Ldy�t�ff����Vs�θt3K�.�:�hQ"jYH�$P�eNH\<l)PX���Ʉ�8�|�l�q�ⰻ��ku�U�婞���6�T�^p|󇾥�}��ڿw�r�$���e2a�*U*�:H�n]0�\G�zw�$��J����5Z-尿����6���/R�٠W�>ݬt���w���}�e�7k~Mv� >R)��� �r�o�rqF#Ov
�/H��0�X�Hh IK��$y<^a��(~e��~����rH����P(��^7V:5n�5���WW, 许б��:"��񁣾���s-W����V������ 2��!k!X-q��a)�c��ճ#�|`[�ɂ�6�ፆ��T)�`��G�0�,qg�d�W����w 6[w�-�,W�LC�&���ŭ�N+7[h~�Uj4Qi�Q��r���|�4{�>���V�p�r��s�����M�d�e���'Yta��gB�K!�R^K���RU����Z��>�N$�B��8v^�{��+j�Ӗv7�	
�� �=8�.c�����iTH{�y'��Xi:H�q��-���3ثow���4)���gu<����OϏLq<`!��j��qs�����o���{�#�\��������Ϝ�z��I��A�F�!����k���dzTn��WoX��Rޱp_�����K�x�h9���^a�����^(��/{�/g���-&���^Y�k)����f�.z:�͏4>�v�ս{��#?��z��wT�C0�j��+���dK'���:i����D����/2n���]����/4
r�V
ܵ~�4��� ȧ���`()V,k�$۱\-�����YJ�v�ؒ��qNqK
O�0m�����1�C�p�
��D�����h'��i	�`R���u�J�z�`�t��F2�ɽ���U�n|t��������鉾��-�y��U��[�~v�nz���.1ĕ�����$<�Їݻ��
mi�`�x�]���h��`�Pk{��ܑ6O,�Zt�����D�yP�E��.R�o���,��]�(;�'7WeMVjJ�ye��R��e<u0\C��ȯ\G��!��c�/��Q��Uŭ�ƞ�^��]B�x8�M��Es��j��̒�F���\��D�=�p�S�R� e���ب �_�P�a5�=�ڬ��\Y�z��tPL��4���-m�닧��C=޺F�)��E���G��_��{��������_U�~���������l:�#Gݛ6��Z�goO�]��ʖ����������3���T4�J]=�/�Tw�EsF�T��<�Im՛z��V=S0?�"6ã�\��T�Ӂ�N̧XZ�i�ګ��'�]*7_��������i��?��
ޕl��Q�L;��c�#u�7�uG	��/������f�����h81�vtt��SwM�hE�Q
�q�h��s�$f����O1*͛�u�Q
�eЦ��d�H��7j1�4��(&��d�}�2�HJ�+LQ�!��D�ղ t-Iq�s�!��Y�S�/��KF�����cz{�F��9�W{��R�n��ř�o�4$��]ӺQѤ�W//�JY[���6Z�mOn���q ��#�#u��J3����m��`[�jI�|�n9��/�	K����.����;��$�����_Bx�ղ�wq�{�&uJ���`�D痎��.Z���?,4�];��Z���.�u�;q�|
)��ݚzKo,�H�r�+�p}��ȼ,
���8����Ƙ�]�
ml�m���B?r(��c']�W�\A(l�z�|;�~��fp�:�n�4oT���烣gN��aQrPi��~�k�_�K?���R��I�����N&�����z��6Z�"7�g�����M��>Ճ�m��rI\m����М7V�ncWi�:z����F[�ٚ�f�8�V�h�����r��7�:�8Sw>4�:�~��Ŗv�%�F+��D�Y�Tv�7�0�2\L0ݓNd4�G|����qyy�8�*��A>$q���#�T$?����/���ёo��p`�Ð��7s�����P]��E�4�}�������y��}G;$㆐z#13)^�jƂȯ��-�����Tc8�,�Ϲ�[��mޓ▼t��a9�+X"%��ɜlǢ��l��?�xmй��3��l(W-;�_80Y�o��\]p݃���ԺY�4���[#Qp~�R&�J
�5��o�&ҿ������z��R�e|�_?����3�Yi�w��-�48����y(n\�n_��cۖo�l���U$��g�эy����YQ�����;1��@���,���PR�y��p�otm�D_�ˍ��P6�k+�7#Ɋ��;lK��D]J3�F���\Т�o3�=�:%x-�y�H)����FC�f��+e_���2����n��{���������!�\}jA{���q���<�����tn��g�ɤ���'�?qԻݹ�������(���s��}���������b',no�tL�F��zc�l�i+6�Nf���J�����pt��Wg~��QO�vM�rE��ިoiGe��ym�Zfx�Z�
ax��!���P.�<c'c	���7�&��n�[������8k{��@���>��s�v��7���"x�S>D
_�$���"�P?���J�ם�̿�$r��y���Z�L-)��"!�N�.0�~�Z��^�x%<Bw^_�B'����Cka]���wˌp$�b`��LG����(Ij*U|�����U�������JG����O�|���w5�t<��z=��;bD��}B�����A�Y'�^���L�[wb����ڻ��S��Fl�����k� g���h6"������!e�d���irq��x��V
���p�y�4�Q��� �װ�ʓR�`W�ɒ�`�C"��#z��|�bF��Q-�	�R���B�X'2(�_E6�!��l8�2üJ���h27�c<��;�d�r�s�[\�m�{�7aDu��+.Ҏd� ܄N��2�b|1��O�RS��R��вY׹fz1욢3����n�z�����_{��_{]��Uj�G�'�?y���]L{vgl3�(a��X��/���o��5���>__�{�%Ņq�~}[Oh��QUy�gc�i��tZ���fC�TF7끎n.���ݞ��,�U.k/S֣rK����o��v��3�
Ix�O7����m$���jc|����b\D.1��V���y!W��l��p����|yd.+�V��L������,��s�8$��o�8V�k��#�ω��)�B�)v�ȅ�(���y��7��$��XD|.)��P��r�H�L刅#,@��ՉY�`�V�1/ ��+R/nڤ({\�}�ƛ���I-����M�;�@��F7ݾ��=���	�kP��:5� ��0O�B���0r%����?~f�gP2gW�==� �������Mj"��ǁ3H��| ���ƞ������M��$��y]�t�LU��TZn�r�M���8�yȾD�1��v#�AO�cg�,�vݡ4t��v��VB����N�j�?7�/є�����mW�΍�/�����2���\�R.���A�p��h6�AD<� [��̖d���k�t�`� �2!�|���x�,�eh8�Dj����-�M����Uwn���5U��
����f��}���lK��=��N�����p>����� ����4'E�|���SՋu]�ouһ�gG���$�um�*zP�����,�|2]�������w�մ������ŪH?=�>�g'����L�:'^Y�ي���_lj�X�������F'�b4��7�':��0hV����d3�jm��֬�BH4[!I7�]�<��.���&L(�S�͍&][�j5��%cb���c�e�Mtqa�x�H�m~��!q��[ut�H6m���V2�&E3����\���3죏�R�ڂ�67+�ƌ����`���7v�����Q@:�7��� 1�6��b��Ⱦ|��yҳb���(�m�6N��f6�N�yͪy�8F���"�N��β��<��
�{�K���]_^���\�r9l��U�UN�]�,��(���E�)��N���y��@M��ܵ�+ՕV-��r��8�<�-'6�t�&��{�EB�@��3���M�|�V��T)�Li�)l5��_�1���V�@_�����_���l�$�G\��fs;�4�,tqE��L��D���ս�X���9
���X\�'�1�v�>�G\����-��l����b��L��y����X��7�����/��^�~�����o�=��Mz����C���/���o�c-�!�bv�Wq��R���~G_{�m�r%wk�/O�ԟ�_+�U�T՛���ߛ��x��G:���E��.��oכz�w��֎G͓ޅ���lp�t��dkSнbCo�v�_iɆ�(�؂�
�f�\�C�����u�_\[�\��]��kkkG�;�N��������ű>��S�����^t<7=�Uz7��W�[�S���q�HK��0O,r�� �ޝ\�O�����+�J������_uTu�n��'ʳ�	DL,8���+�!���P݂]�}�Mi���(����hOH�8$}\'zX�~�4�������þ��ך,&vW�8�y�b�<E�X*�M�-KN�]Sz�-ujYT˚D����Zr�ڎ�#�	!̮S�e��tu{y��/_
S��v�v�i�o7�*�Ѕ�*�O��Q���>���+n`�
͵��OTFK����vUWJ�UZY��p���J�.Q4*eg�X^�(��ǜ�I��|0�Z���̻Q`�E[��hh�Y�V� ������Jhzc�# &sL� j��а�*厎�6�R�7ֈ�h8U�������1����]��]�#W�:3�(����K{���쨰���v88ڏ�F�;�{�\�~�q���o?}�W_d�٤~��s'��u9�?`�\!)|г���jm}��z��[*�����C^����Ʋ����zw�������(���g��q��T��FGo?zCD]��������vM�RQ����5��.�]���@;�÷D�x�A��!�BZ䋳s�|���#6� ���ڍ�	�bYy8{|�7��胏���%"`|�4r�Y��;{n>d��|�Q*Y�Sd`޳�� =E#qqg�
��U*]Q���j��d�M4�t��t�
\N��~�qp���Gx,��n������
y��Q�pǻK�􊭦�$J����X�1���`ID2�M	`�� *wXu&��I_�jQ�VY6��ZԊʴ���Z��RNW�&􍆹&�B<�
Ǽ;9Ҩp��>�P��J����+��ν]���q%��3�ǘ>;h8!~���$�r�2���rE��zo��6�=-�z�^�3嵌no���U�CJǖ;؏���-�Yb�:v!��ou�WD�0�oT��m� �U�N��B�+��W%8B��e3�t�,��6E�EN,��ڮ 䂀���0Y����p:3�D�c�0f���1�� �����xX�d}	nK����w봕uni]�˹��s��/����J�������'��_���������A����?t>���t���9Ql���v���.n�x�-����*eK:�k;?����	�x��C}}���-u6�����^�6u5����k����������L�חjn�ԩ5���t��V��z��5{( �d|����`�l!�4�1��'���8�s���%�xN�D`\!t����V�/]�e���A���y����XY���&PF�D�%
�UJ�Z��)����`����\��[�L:E�/���BĝY����E�Ɣ��m5�O��,��`n��.�}�~��>)`�N^��"���3qݏ��p9���l9�p>��#NqC2�g�K:����ۤ��]�ϵ�����(f5���s�M��{ ^!�2�d���F���,E� �L���5�DP0L6+[�$&�YT���ܝ���\�TA�lAovv�����j����Z��z@?�FǶ�.n]�����c�	 ��e	4@&M
@�.�Q��W%O��[���Z5X�'�kV�0:	э��sc:��M'K0��p��:��g焳�]pLR�(\ȥx���[�H����p^[u�_1a��Zבat4[~u4�x�ӊ~hF.nolu~�����_��7~�|2���t��!�,O�q;{���7�zG_�������gzvq��>. ��O��˺������^�\�EP���H��O:�z���B.k?���c]^_��n������V���r�\��l�X���?��R'b.���Cu��5��Tr��s!T�5mmm����ay��P�}��P���[��9j� ��EA�CoaD4X�
(�I�ȟ'r�d�c�t�p��\0�aH�2^���<����$���A$'�J	6�=[�+>�G^��M���sb�!K:R(%.��O�\��+���"ctpV��q�15���JW7��Jz��ͫ^����q����0��.t�Kk\ʪ|o[�-��Es)-K9M��(�өo���q����6r����c�O/5%dh�V�QSc���N+���}!5D5=V12X.�.�7<�������Rñ����
%e�ý�k|�� _
�-V�K������T
o%)p�_��F@�6�`Zɵ�IdVV%�N(��֮B!�+�Dp;��Yz��`�0	��ʄ���    IDAT�
*�� �r������ [��k;�ch �Y�q8j���]��`��s������	���u<�h�Ӧ "������v���~�o������?�C���;���c��c�d�$��Zڮ���O�ѷ�{_�tIW�=?;����8^�����z�H�U���^t�����M���n @�ǥ�����t�������K�u�w:�&}��Uӗ0��Ѕ$`�Y���[~�r�5Gӑ>��ͧ!Aޜ�(�bM�:͖G).���}��'����ܶ�<��[���&
]B����N�[�դ��+�|�W�T�p���QCC�b#�����|H�ӄ8;CF+�r�q��L6��o��P,-�>5)�Sr1_���D'�?�u��^=�?�荆�:Q2��F�J2r���ե.�/D6j����ٜ�>���K�u���ӓ�D�J^�ݶ�vmQ��(�[�`�l~��6mj���ar����R��KM�nMf���j���mO8�8�ߡɍ�'�'t��z6k�ک�eB�m��H���������s�\�h��c#��ϝ�F����~0�'�ӂ��c),&( ��R��® A~���FvA6e���k޹���QXO%v�l�і����Z�x�	��%M&��\
�X�!�<
(�h�E,�"M�
�q��ܸ)p���jEi�>:-[usi��Mt8�鋫sͳa��o�~��}����|}��}���ݳa��N��'��e+v/����R�����7��
�(T4�Muty�����=s\ܻ�{�{���V8|vu�_~L	7!���-���X��Σ��n��� G���H�~O����mݫuT����n2/@��[�/��V�j
�3ONO]l�)��ku�+����y�ŲG�g������q��ݱ�<`ٔ�`���������������ǘ[�B�h6#/�c���r�_&��to�L�*�E.Q�X�n/bx��J<��o"�O�E:7~@E�"#ʯ?.���X�$#h� 1�]\���¿cLj�0r@��{kD�W��6��y�����^p��F�Fٌz빋��z�T����]���jY�k�������/��ϸn�s��I�k��.���?���~�&�>Ák�l)SB�\1`��=O�W&/��!d�"��̕�TYnTZ�l��tŔ3Y�Y�I��`b�zm�A� ��R��C��lP22��K�������[!�*9
tS�WD��Y�a�~Lt���̽��	u�U*�Nm��"{��T,lA����֋��"9u�j��,RX,d�^�X[��nH�K����Jm��j�t��[[�Y%�R/�������7���ײP�����Ϝz��Q�����H�	�G� �r%}��[��w��f�j<knNf�� ����Һ]���ő>:yxs���W�BE����Zz���J���zj7\4�\P[Œ�I��5UBFmRe��������\&\:^�L4��� �;�����5�m�Tno���}���Ӌs�i�DU���8�Q2&kp3�k� ��D*��.zQC�����Q/(���O����ȷb�㒷^�st{\J�me�-M����<*
f*�"�.ql�����Yx�r�P�(TIg��P$M)!�/�H�2��� 2�,rmE��h0T�wk�����`��x��� `;�Ԩ���bb�ԺVT�7<�����=sc�D:Ǻ�=6�m�i"i�o����i|��ʅ'�t�f]�z�txp�c[�uʃ���VN�V&��K��>�5�Ψ�ߐ<E�.ט���	Zah+�B������ �l.����fГ��*�[>�
Z]�5^t/�s�������#<O(�tmx�7r��2B��є�҂z��!�ti�sH�2�I�63f���DR˱~%uu��0�T��3������֦�Pj����ʮ ��"(�M�#ݩ�{�������,n���o����w�.#d>�ϧ4�m%˯�q��~��wlM�.f�9`U:��O��z��O���W8�R3S�v���������Z�(�٤Ɵ_]Z�D�q���n���JC%��%���r*��,���|���]�����j�R�������b��be�7~�Y�5�M��4�� ���2,-^-l�(<'��wQ��t`,)ҩ�K1�>���F¸�kyU��1ۤL���p����Sch�"J�B^u�M�.��،�ѡ"Y2����1��[D�J
���a�Qn����	ō�J�|�D�%㷥N��hҽ�������B�Q������@�|F�RN��]bI��y��j���45ɧ4!u�0o�� }C�y��Xa��8ʂM�U��oo8�S��6��r!8��8�f��݌��%�fq{å����Mם":U������㑱/˪Џ"�*�Ł�ӵ0��k������rB0K��3�������C�!ۉ:��&��#��K�dJ79��	�+SF(flK�P�"��1Y������uNݴ�H�@9��Âz��Ǔ{��L������.R{��Ɨ�i��;]ה�Z����֟}���dyě���wN���E����㾉�����$ c�Q3���v8�ꍝ����E�(s���p5����>��|6��}6�ڈr�T׻����u�I����f��Ǉ��*�����ÁQ���"!;{L��!#7*�2�`e��_�\k�Bt����ԏ�ֶo��vG�j� 4��>�P���ߺ�Ar�Q��:1Z�E�{�2$rٸy�0� �z˩Z��K+Hw��ţ���0So�-�A�0M�1�X>�����Մ{����(9���p��$E�]&�tx�;z��6
<�}�T�6v涱x��ű�x�>������Z)V	�8)h�2#�ɛfA����ω"g��@�B�ωi��涧��Z^��o��_ε��C/�;�;5��5��C��I�Tİ�s�	j�`�B��l�X>�D����g�.���/{8#�΍���8��0_�����Ԁ�ҙ�ۻ�jԔY�տ�	�;�r�k+�Y��lh����"���]�j!e|P�o���1�t�f)�ؘ"�r����eJ�f���)v��ٴr��J����l�.�� /�U�a�W
p:ez�BX.���_�US��b�/ju�kU���U&倠����'֢��Uk׏�;�'�����y�;�(��>����dy��7���9�����I���ӁW�"XN�(YY��_�����4����}ߗ�׭�����d�B`P"�	J,�$2QP��(Dٔ����xc1�e<��Q"G����鞞����Z�sϾ����<ϭ2Q4�sZ��:���9���<����R�6v�p�Ne2�d��x���zԷ'�g�Q��rp��r����S�+��:6�u�wӲ�h$}��m+_�jl��Z�'Kf26;8���N����XQ��ɠveɨ�V
E���67HH�W� ����O}&0D,>9wc�����>cIg\0��5X����V$]��Ӗ:5}�_��g$D_�Zn<O����~�	��^�7YS�(�G�247��@�#k�kM?i�Sʠ�������4�H�t2���a���3u�:�%�&�TT�`��xj3t� `���M��?Pp#��D~�i{�ݩ�l{���fncۘ�SQ�mTm���,���v�v^{h�zI|dR@��lZdpd~8�S�� #�
�j����]v;�B9c�T��0'���7�:>�b:���i⓰���۷j!(�F�����n��N�b�a�F��LY
��M	�i��W�7a� �Br-b|FA�����+V��sJ����YKf����D��5�����ʍWSF&��no`����S'$���7˼��6��2�:#��\��w������v���	�J��躕˖*U-U�����nZ?�g�����c�/pn�J�+7w���������sᖲ@������y���'��C����ዩ�(�R�؇��=h��v���4�@2.�3Y
����s�.jɨH�x0�#)�Wݲ�BY6�u�\��5��HL� ��ۖ\Ω��WAd0���'GjD�����E<��	��\(X�RB�� pqv�����;Η�w���V<P��^��,nT� �q�\+?��(�F27��z�UQ�2imlAO�� ƽ�/841"�O���`�Pv==2Ѵ��#�}��V $�3��m$��� RD����P�������Y�>+��F!�:Z��-4��3*�s<P�zx��^))��6�T��۱!�$,U���n�0�nl�J��|b��Y�Y����������2��揉_,���{��21\ s�_t�wݨݷ�uK��Z�&��*Ns�9S�G�u�n2!�0�wK�e�"\F����S���D�y4TP!��P��,�g�j�0C����+�P��4��d���Y�\�ݭ�~��{!M�#���1~��i�A[9�ͅ�S¤�I�
�����0VfKk��r������|as�T�½��ʹ��J
q��%u�P8ᾎN>˕r��Vq�<6;;�l6��سN����O�3X��XE��*�Νj��=[o������|2�o��[_��v�y6��lҗz)�(z%�\�x�U�2��d�0v@��E��9�`���-m��ˁ�M6��f2g��B�m3u��A�m�d�Uc��ʶ���>}�T�fЁ|��$Q�ղ�nGVb8\s���8�{sJq�"ΆD�nc��f5��>�&��%�2��ra�����¦fJE&��e�W�����Y���Ea����<��M�����r���X��W����W�4}p���w=��E�X7�*	n���[\�(����Q=�TJ�O�V����%p/J̾4��!j�Y�n,L{�C T=�pa#�����9X�6;?�
.*㶵u`d��\�b֏��E�eW��Y>m5��v,Y)ؚM�K���T9?�dt�`���)���/��ou��;=k]^Y��R��8hax��������rt2���/�U��+�-�B�l�� Ѐ�8�� ��̉\F�M9�� �u���8��IQ��RߪU�R̫���� w�"�`&��y7��� ޥlȌ�ED�m8YX��W���l@o�S�y��B�|���E��S��e���cM�0���eMY$W�����[)��b>����ɑ�l.�����Z{�\��~h��k�[Y�7���_<���y2��0����(���|��޷�틇��-(0��>��^[k!����$8�雌h�@fDZ_Kfm+[҄i3��x2��zi�2���h��֎�y��t�٤��N[��)(k����K���l��Д�l��D���c�o������W�j�8�$���i�Ԯ����R?*��@��'/{h��J�0Y�V	����L��E�L����}m|�P��EWf��J��ZCώ�@��A2�٠���1d� ��vvd���u�p}�?����h�d\E���g�`�C�V\�]: ��=E>�2>LH '�R]�'��X	ٌzm8�u�����&��Rي[u��4-Q�Y�\��&���� �1ML靑�ჀrG�)YV2-	����}��c���.�J�H =<&��d#�z.o�v�l��۪�w���F
&�ʅ%��Y}8�2�d�3��`r8�_'�3�7N��;#�Y&���{!��d�R	(MBJTO�b�2٬Z��M���՜ �Z%��Q������<.�g���Z�L�d�D��|^	U?���K�M�g���L�U*c�J�"���b1{1��k��׶��$D�JF�Y,_�)W���9���?��G~�b�s{��.�o�w����g��J�0���x��썭}��݇���+Z��:����3á���+�C�A�X#zzSѕNS�>5za�,���#-�҈����]�AL�Z5���Ɩ�����N�eن�X*����s��i�n��=Fؖr���]����B:::������p1� Ǎ�-g.��Cp�W�[P�ı\�ޖxv�D��l<��	48>*� �?��󿔉y��Y3�A)G0`S��-<I���4�����pL�9vo�	�aHA0�Z�"����mepH��`C�kt�� oN��SU1+|��)`n �	nj�{1�cm��LA� ɿ�P���$?�L�I����A�`��弱.?=?��C��ֶ��坦���C����Q���b2��Q4�Ԑ)Z��i���Nߎ?�u�-7�@L�RE\��S�N�z�wG�g��@���w3����,M���
C/!�Zs�%�a9�ش?�!>��W:H.�1�P��֖���~2�)AN�N/N���~����g*U�o0�A<�	9{6j+a��¹q� ρe������$��*�F�������^:��*�/[�X�E*i��ʞ��v:�K�r	�`��kJW����_|�k��W��ȿ��w<P��o���'�������T8w|�� �����r��^�:�3Dwܯ���.;������`=��㫠RL�sqD��L<aL�91gk�r�F��ի5ȄX��W��Ռ����M��f�n�8�]�����{��#�
�����������L5 -:��!}Ʊr�.�߼�$��-��+$�mOm�T\�@�Y��R��O3.,ж@Q�}�]S�

V�"��zo��2���[��J��M��z�Y����L Β�Z�R�&�%m��V(C.�NC��-�:!��`%t�7�	eo�7�s̅��T�+U�d�ָdm��*u�c�r�������
��ked�|����m��*�!H)cp�����;\̧�\�OPA .IiJF�}pݵ��u�Z�'F�PB�:����52���V �S����` h�T|��]7�֯W߃w.�pf�`GP�`��tc'֜ӨB����CB��n�3�g��u�&:pŦq����0�R�������j!�"�߶���>\�/��nJJ�[����gN[��2Zne˗���[,�*��a,jgө����I�¦�V�I��Q*]=����#_����?EP��ޏ�qp��{x>�������<t������-�Ca�~�/ڗ��ai[�����>�8�S��l�p:��OE��9����~��2&�3'��\6��BĬ8YYe����,=]�j4��vlӘ,�8OOυu������ �?5�K�s�������7������5��Jx8�Ar#��4�S����&����K>�J@�>S�D������D��(�F-X�M��ƢTs����||�������W� �%.s
���)AC�[�s�ET�(F��v87]{.����?��j�)�C�H���@�!�����&�D�ގ2�xRSm���9O�����t���t��LFmH�Q���vB6i����;-;���n��&y2���V�v���ۤ֞�l�,���'�����D�07ܯЂ#`�n�/����&��t��~.�VS�a��gҨ�t��t����wa��H���b�'�h�**9=m�����
,Zb8_�Ĭ�^v�`ހy��#aT/$��/!ɻT)�����:�/M�y��T� �ޗ�p��|a�
��*�ד⇞��g:�>�&�U����ɣm�A
��筛���|l����j���&��f�r�hw�O��_�c'��3�>88�����A����c"1sR%�6k�����{���Ν{�[j����{f�/��Űm��X��q<�����gr���E�e���s�'�R�PI��Z.���ba��¶#);�嬴�۴�Q�+v����J��Ϗu��˫�kg <q�n��D
������
pdP�>z��@��K���( �.�d�E���#���3&���w4�ہ�?܄�B�Q�|^����,N^��A$��[��?��|TC�Wq٘�W�Ρ���`�%��,��q%�+eC?���/�����sLO$Ž�H��g�|6�`S	Ǽ`��#7%E�F>A�ҋ�L���^�un?o2*��M�`�zA�-Z/�*��k���;���A:UL��G�t��b����Ώ�����_=G0eж��%2�b�>��x����f`��XA����=m%�rф�2��    IDATE�lNmvӱEo x���dl�9���OU�8<Z���u�(I���zr�mlVn��̸�A�-�+��S������P
�$�$�$9+GsT+o3�;ŧ��� �J��t"�����']?����\
��-S�$��R��ժM�C;�gǆ^d>�Mdi�R�����^��?�w>���o?~o����g�ֿu>��;�;A�l�S�Z�~��/)s�+7�����=�<�O�Nm]ix@Yz��o�jVʔ�3���Ҟ��(ZS*��s���mD��-�V��mk�{ي��Ul�Z*�1�Ҕ^7���T}�H4�$]nBH��*�4m%˒�j,mo���Q�R�~�����ٙz>�F*��XF��Sݫ�B��	��T���Ŧlϋ<�s�W`���ml>�-�k�j����F��ŦN����-h{57l�^�;,���o���y���W*>kp��`�V,޾?����{:BE�&�k�K�p)�8A� Ep��у���E T��q(��e� t��*Gc	w}}7��`���xdn���Ewj�\�36�G��B5��Lk4�D$n����wI���1=��	������O]/��"������LC���6�jۨձ�hl�t�*���bq����;=����E�b� *��P`������<M���A���=5¡�^�"�����gРl�;�		�M�]L3ɮb.x��J֩���e���������t��S�x�V//dz	z���%�ί�{l��%-���k�H�i�"��m��V�����G�v�k�p1�h"j�R�ug��_��?����E��D�~�3����wwO�_x�k���i?��E��B:V?��;����+�ܕt�n_��i�l�1��;[����VJ��f6�������qd)uI��6���,;_Xy���h�^+6�n�!h�U�Ʌ\�����~	�v��IY ˍ6	'/���E�
lp^�^�=9?sY��i�66��Ғ̍2���Gh���PI E�֌�5���5��A��%S9z�BA�Gld`;&z�4���K��/8�H�pm77�Kޫ~���2Q�E�
A�N���ß�9� !��F� ��,�������+��j ��6��ե=?>���S�9�iO���ݗf���&��-��fŢ[e[2��4����Z���3T9%�mig[�4�E{Ӂܯ���B�FS���5�Ɯ�0˝b.�����HԷ�����b2i�D�
@K�Au�6���b0tަ0衑7�	����}.F�7:��{8h9:�i �JγF^������̷�`^Pr��:���M^��E(T��r�808�������^�r4���)���y���H�E���L$��H'�g����2fɴ-�s�l�f�֥�}|uj'����}K�c�U-��i4������?~�ѣ�gZ��k�b����֏�O��q��A� ���V�=�w��ڝ�΄�q��?��g�6KFlIp[����{{�d�ړ�]�;���X����H�@ NF-Kv6�[a���d�^�n۽r����Ŵ����ܮ�a�~ry���C��&�{���0�eJZ(�ɓ'��.<#!d\�J��˾`EGXt�&5i������G@�,HD�MO�($�����R�Њ fU`�p �94CC���tb�!{
��@���9G�"$�C�r���=O��2�Ϝ�/ב�n�R����֕�������S�K��\*P�%U�ִ���n'g�������]���V@ �����ỚJ�,��鲒��NEr��T���G66Mկ�]˜����X�[mwK���r*��R�$����>�}��=3�v�tI�Nm��X�������WL$�Li�L+��5���|4�,�ܫ�*WZ�r��ʩiHM�ݴt�?`4���;��s#_�^>�T�Q���ڧs�����˗�8�(��8�����
)���]>�b���p$vˢ�J�g� ����*K�ڊ[�	n
l ��E�[&Cpk�U
���Ԟ�/���$l�V�����������7��O�_L������^��I�g���b�?�M��?���}p����$Qt3�iZ����mjn6���C���-I�堭�/���$��El-�~�������}�wD�"s㴄H���g���'�Y�.�ɉ���hø^��./.��T�&b:�ܻ�,�Ӈ))�!�UФ��=(q�����u�,��a���8��'�O�/�\�98�dn�z3�P�9��T��0]�6�[��e����'8�RE��I\p �X�Δ�r���C��w�2b�q�-�tW��f�6�uht�|�O�1d��\*[6��T6�qW�kk���a���١�9�=��_2|[3)�%�։,l�v�n��Ld&���/�U��yK}0|䈕J˴$��E.�R�v��C {�I5��9.��3A(��!a4����n�.m9��u���iej��-�	�x(#��)E��+*��\i� �[�\`*ԫB	\�˃�=�{T.�u���)��WbF���k	�/[A������j�u���E�3����.��b1q[��6�HXaȞ�(����
E��R��G�'vҹ��T*�z��٭T�ܗj�����W�߫$����R���x���F�?v9r�� �S��[4m_���
w�{�����=�:���6�Om��@$jo?|ݾt�5�ǲv5h����=~�\n���Z K�2.�Yz���%�~�n��l�\�
�m�+vrt"�U�Z���	�P�����7��k��dtϦ��F�4�L��Ө�b�T�7�)B0P�a�t�� ���j�)Љ�#GX��2
@��X�e�t&^���Y�%o��k��C&#d}�+���kP�x-���J@�g(C�=�t]�_���e^@+�	��hԭ�l*P�g2z�XrpU�`��^������j����~8T`�W����r�)S~"�5N��8��>��A���u�-��h���~���d�rI������Z|�a��m[T�ց���x&�r�H�i#U�b<e�O��u��ViT�P�2��P,��8=�%�N�{�g"@���̦2�a]�dКJ���A��/�!���´9̣�9r���1׫|���ޙI��0��)*c��J�%��{���T�����\�@租��<u*JT����Ap���\
L�/��d*��F�rE��߳Q�F+VЕ*�䢆	�xn2�5o�L�"��-�y[����ՙl��a�*�w+���ˍ��_pe�~�G/���N('-N�ˍzn���M����,��倅���|�o޷��}+$2֚�}mO	��8���T�1��SpmS�%����m���P?##���g��]j�K�����$���,(�����l�F�n_�җ���ߟ�8��pF�d���u# �,0�� 6�w�
婀�c��t&��zC��l6���Y��d)d{dq,�S�p�'�1�:Yq���dN�FCY(?#[�%h=6*�!]`��kJ0Q%�Z׳����-(�p]d_Loy�)����t恚y�ˢ]��J&d�g}#���|��3��!�#s�����ե4��1U�N��/�R�ar�x߫Y�ޞ-�$"bm	������1k����ĬzeOb��k+�*�تk�Ջ%��201�#A@0qa�l�>Pq.�wٿu}m�vO0o�!���Z�:�5�}EV �)S܅lG@^����2���0�N^⧝r�b:�Wc��*�F٩Jx��������|L�e����y8qs�wK�q�(��W��-��Y�Z�c�#� 7XD�(��^����hlY!_�������u�e�6�n죓#�v�/�g�^,�6�?�}_|�7?7�J
'��_yֿ�w.���<b�nӥ��q��G_�w����nlgг�jj������JͶr%KŒ6�N���
�KSW=7�U�.qJ�Ƕ������a�nw����/�x8P��A��̛!C|���4����EHp����-������Cׯ����:a���T���L� 0B�C��1xZԊ�i��?�	�� #������P�����0�$������̕�Ng���������xq*F �k��g�,`q������=�����O�/4�Ĳ�Mv]f�g)�ᡌ�9$�5g6W ����Ж㑂e�2�)z~N而H��΍�[��i��t2 T������XF"�_�l���f�dv�m�Fή���V�I&<�	�7��Zr����S;}v$�GTw�w��`wϚ(0��N6n�H���]�7Y	�.%`Z�gݞ�kf>u
)��$H����X�
P�e@����!��� *��|�ҕ�xCޗ���d�n=M��t{��a p�i� 
���� �q7�z�O	P���Ry�[(W^S��?�eq=�;mNdCe	,+
`�J��+֛�u�Um����bf<bW�����G�Q,��j?��[o��?��/�	��x���R2�����[
n��j�ӛ�-��ڿ��M{��C;��6P<��L�}S�� D�(�.-�ƺ����w���p��4v	�1zݾM�o,1[X#�mUda5�A��Rv|tbg/N��%�������l�7����f�j�Z�n�dE,`~��M�zX��`�H�zD`����j±�N� 	�ґwٍ(�Q�o�Y_Uv��	 <�(���FH��L��R�g�T�iR;���I<������� ��-��ŋv���>$z^�qTc�R���4X�����5tzm{��ȎON�g�
���w�	C�Sؔ�;��O��p�Ab"�9��T�sܗn��h�\�'���]�[����π�D,��H"i���Ʃ�-�9[�Tm\�۠��NteK�Zә!���o���Z�=���S���| )�v����tG�m\�,�����2?1�����P� rM]7�	ĔmXJ��#�y�<��$�2����~z���R�g��@���%$�i��h~��a�������)�L�cC�Wի��R�[ghc���T�ك� 	S0�[��O�dX��9��_E1�O[<��J�V@͚�ָϬX��fi�[o>�(Z���U��~��?ߝ�_����W]�w;������u��h��#��8����)`�Z"oo޷w�n���s��ϻ��j��#L���s�����*����ق��jKFf�RXӔ����XL9;7�����)���ڧ/����BZh`���6��%����(�I�~c1�Ak��*�L��g����Aa�C��SaB�
dr~N�c�Vdqd���L�Y��|1� W�P�ך~�}���ٱl6��Wvqq�@F��)LwC���ޅCZ���C�%�c�������������Y�B=�ة�B͉[�����B�ٺn�,�g3�8��3��%LJ��Ю�/����i�aj�L9A�����(�E1m��M�9k��6��lI�Ak0n5KZv���uߞ|�}K̖V�'��������m�k6�4`�	Ԩ��z1���[⩛r���k�\u� ���٥* ����P\W�1�QɊ3X̩�Y[��7��O�����T��k}�DҐ s��#� �OBU�z)�p���u��~��.�T("�a ��l%_�2Le~���{Qma^����WX���E�/M�)��lZ�`�2�[2 ��%V���zO�{�����ݭ��<����
l���E���s���{{G��7N7����+���r�N�����}��vj�W(��K)x�i�;m@e;�@E�G���g���l�;}�F���x�"��4�a>�ۧ�?�^�	K5�>R�����h
��F���հ��ݤ��y h�C�<�7��M�Z-7�L'��s�� \բƪ�/@�|��'�O��t��zi����J�^Oٍ�>"�L/C�zk5g�Kkb������B���w�VF��s�:h\��`�b^A�V���u$3�=���K����v<re�+S>iZ�7=$l�zCφ�>�n\y��&��Yz�6�67C���n��$��p�G>'0�b�֙���Ӷn�m\I[�����+]���IZ�R��,����O-6�H:�+o�i�4Áj�ZX-$��*M������s���i�OA�'�Q�{6t����(ŏO^X�۵�V[�A����%o���Q���Y&8A~�i'{$���?����,o{r�Ӕ���� _�/�[TJ�EC�C�p�~M8\�2=@�7��]N��_�	�DNId��$�45d�S��+%ySd�In�e3ME�M���H9Q��r�����Ӈ��o|n��>�'���7N��i-Ƒ��~MT�W�~2�5�U��ܶj���F��w�|p���ρۑ�lā��47i���B��ئ;��j#g���m�8���da(7?��6��(*զ�j�SpO�v}y�`���W�@��w����`&<��6��$�VR�p�o�6�A�Jwt&��Τ-,$2T����\斛Ҷ�rN9�ѯ��Lo�pa�J ����n:A�R��g?��qQ]�ǵqݠ�]��	��#P������������gx�L���[9�&=A4�5=�'tm���N�����`��;�'�'|����87�g47���F��n]����Q�&0n�9HȢ��u�d�jں���QC(Gmf��*n�������i�,�2z���6	k �zG�[{vq|b���;z��M��jV�n�9Nv�Z��s����x�����s;����S�`���0��#�O��*�|>�6A�|��@�j��TX��|��$s�U��.�0��m������$��eb�� �K�sCG�ww=n��z���ɾ��%P�a��RknY�Z�\�b�R֬P�5#.x������Bix�����{ۿ��Kp�Z�"����E�0�Yln��ԋe'/N�D��Mk���&�N �HU�ZY7-C5U�xl[�=�n�w�j��8�%x����>��RJ�bV�m);��J��Ln��n)��;]7$���;�w�i��z����G>_G��qC�,�ƽw��N���,e)7UYf����r
`281TR:���T��L^���h\�tB�M�"�qw0��dl7��;u}D�0 H����ce	x?��w�
lP��l�20�W�Dx�J�Z�9<xR�
��5
{FII-��>�Mݤ��?��\�}����R:4���E�[f��.elQ�۠��n>a�LD��2j����7K&vP��!ex�b�Ѹ�	�_�p��={�D���L�M��=�F��npL��4���J��׷����~1��E�wH�;lG���	U1�_e��fl���6���{
�W�U�"�:���&J�Jʗ�А�w���I仩�˾�G�rkL8<���m��M��[Ω�Z@��(�u�{dx��Uv�,W�Jl��YZg1���X2��R��4���r��޸s��kp;��~�Š��/��X/2s�$�x6"�HZ5_��FIm��jt2p���>H�њ_.e��29��K'��:��hn���V���]{��e#q�A�^-���������Ǝ�:�^��� ���H�o�L��ww���������Wp��*l�\��Q���q��`�6e��䄍ʍ��Υ=�&x�{X!Ɍ{�I^��3@9B���%�O�/L��d196ߖpf��X�'Fps H����)�7�{}/���:�MS�v��9g�L�Hp㥅�t}X�4�ᙼU�׷DD��m��CL0�k�ˡc��r��	n��LF�����E�hkJ�\�ƅ�u3��6�&l�{2��En��9�Xr8�u�;��~�f��Le��VS"�~�����l��~s�޽g{{;�)fe��w5�G�5�=�	��o�3�8?��d*�	���L�X�6���o�:#w��h}��Lg�P*�p��	��{b�[�I}��n~���	~�CG^��ԃc=C��d�{��Kk<�zkd^@S���l`J�����k��Pg���^��F�/���	i�b9�M+ժNg�^�x!'E��̮&��ΈGT�����n��ފtH    IDAT�w�/���k��������l�K�7?r1$����-�;�2��|p�|�BQQ7��lF��1Bk-���iÃ���	 T#��L�72��N��T���v��%*�$�$�p�������::S�������9�{������Fc�h��Ν}�x���N���v�F�M����p�-���:� )@ֿ[���#� r��������;4e6^���*�W��ټ{�+\�=2��ύJ�< *5-T�S*���l�TxCf@�R9�r8��7�!k�9L�0 �P�0(�}�Bo�ϱ��[@D	2ڝ=�{���ɑ�rM8Z�!��;}Eޗ��mPϛ�7�����P���Dٿ9f�%[gS6��l��['�Qp��6��-��myٱ��kˎ�Zc�޹��1�_���j��>�������u{��}��/�_{Ce*�3T� H%�Ě�l��|4�����=y�L=ڭ�]p�B��Y�Q+��'k�@��f��
D�E��C}���֎zr(`�2`p��K(���~�����\r��6�&�$�z��Z��H)�� ]��e	__��%���B=�����l�T�9����0k��ڨ[�[�Jc�6���6+iC�"�YN�z4t��F��J23�-������_�k�ߖ����w<P 
�b������=��S��Zzn��n�K5~�(�2f&;�����9t����	��E*|�R��t�$)��K�����n�h���<"1�����B���{_J��'	�ٔ���ĺ�����)C ��������v7b�24��*7R�i)X���I�g�>�/{Z�<o���ܮ>�
��:Zv^M#�l�����U��E��Щರd�V,�`5qP
�L �JZ����J��L��%�IZ�/q�*v����D��<�}O�՛C�����l�f$����6}0��Π:��^����ޙ��zn����X��<
�l1o�B�ɸMRQ��6�%��=7ݏU�fg-�][n���ܻo_y���q��e��Bm1�_�{߾����Q�7��G�v˙�kggK����Y�<��S{��MN�1�ؘ�k�!~� v�h�-m>�+���mT������i�k�6���B��\�G��_(I_-[�A(�c� �8��9��;Bp+��A�E����d� �����-�|!k{�������*G�.eֱ�zk����\���s���m�H�f)E�j*;�)������y����l�̮~�Y���N�i.���6"<��bIz�jh�%FB���}5�I(W	۬��3,�g/����ʡ�Y�%{cc�Z�$m;���> ,P�����T+Ȥn�~�q��f
n'/^81ß��&l7�NAןZ��ܸq�h�z79B8�T>8&P��]:m%zB^W�M!]x��[�l�����%8�`���	?+���bїq�̅̒�H��;��
��+��笪�5w�pNTz�+ZR�����^�?l� `2gwʛ�>*8�^ϕ�6�ͦS���tؐ�����s�'�q�ahA��u���h�e)��	�eЖ@v��I�0�O�lU�ۼ��~!m�\\e)Gm|ze��WV�o�^�~��VffӉ-���{��������Af�����Y���}�W�"Ƀ��L�6���ũ==�-G�iz`2���)���fe��������)�J�%���r��N82�4x�)��tN5�m����<��ՃJٛ����P-�A���(Z5E�+u�ʊ�?�bZ�V~�AB	H�c�0� 0IR��������_��i���<֞=2XT]6k��"��t�S���Xv��E5��J?�����/����	����}�q9k�������M�~��������l�@�˼��Ce�����R�as���Ur%-��|��}��3�h���|m���v0���l+��J*k�lN����f�裏l�s�(���C�٩����t�.�&HHON�5W������P"�/�	&�VS�����v�S��E>�P���ES�l�v2ɟ�lZ���4���&���|g��h�J!�a@�����1�P�qF/��^���h��B��#��&��t�(r����K�pz�\����O�N@�����`�?��-��Qו��is��	���z@���^���Ip?xM/����L�"��Ev�6,e���(�q_b����y�R����o����W�7�`��Ȟ�؎&o\�%l\'>�ֵ�����=�۱�Z�JY<6�N-�3�<��/����ߘ�)SQ���z]��Ǐ�gO���!�%R��q�C�<�q�p8#��A�0nz?^����sCI��=��|)X�=&�"䣃�����P��l�HA��!��ޙ Œ)����U���穐���+�������ﳽ�}[m"֛��ӵ	��hD#���'�wG��Uӹ��z�'^���K_�ϧ,%�]�o���A�O\L�Yx{dn¾�ˈؤr�N&��
��c_��K$�є�i��N�n�BE'�GOۧGO]�٬-��|<��Xڪ����
V��-�`$j��]S��\�T��Ɔ"��&�FB������B�׺���Wn�7�إx�<��̚�D�=�t�������1�Д��Z������dw(��+����#�a�x�a��{�	$[>�dC�R�(U�D!�@���|!�����,Np,f�F�6�Qj�i/��f�������
A~h����o�4����b�� ��x2;�?���b#	:�i;���[hF+=66Cn�J�6�UR6��nqn���fm[��-5���d�<|dwww�I�=;��/�s	r��
���{�}c��ؒэmWk�Ň�m���8P��%WQ�LW־l�B8=�PomN�������&���J�S�?�Ğ={.�X�%ZnN�ٙ��w�6sL�s.�K��Ȱe��!�Ttc�u}6(T��\�Bp�(��}qN=�C�ee��x�Lydp���ܓ\<�@�\�㮮����s)�7v��Cۻs ^H������6��,nb�`���$j*�dj�_)���������P��w�m<��~�h�����0C�Mp�i@p��P<E��`,�[�܄�����&n��m�klY�\ї�ѧ�ؓ���j�<ܶ�ikD3�W*K��-){DQ�I���%�-� N).ݱ����iZ�7%�c�s{�e`�ʅޕ�llF�U�v�f$H\�_(H2���sYAй��v5�y��jKi�6M�P2M�n�N	�-2�.�x����AHʏS�Uʮ��wF�l���υr2�p���^�^���]en|v2�00!�i2�t��u�`��@'�L�L2Y�"���%��>� �O8�{(H ,��)�ӔoD��[ωk2�%��3�G})��f��l�V��-����e6���,mrֲ�iK���ۻk��v����֍��m���A^Y>R網�h`3��ԛ��7�v!�^]li��B5]ڰ;���k;~qbWP�`Z$c�FJ�6����
Œ�^�}a���i2ϡ
^��$�����K	���2M��k�6���p>s����E�$	yR������Q��}_Ϸ,���xB�#�1` �OP��aP��{V���MD���s¢/&��=��ߵr�a�|�:���ш��&�V�k�ݲx��J��p�T�������������<�~�h���.��T	..L����B���t�ܸ���&'��J22p��ܖ+{�٧���XAI�y��G3�I�l/]��JM=��l�J4�&ˍ=��3m66J*��s27���5n�e%W�57�A\��#�'��B1���f��U�@\�,L˕���ä)��,���1B�L(*X� ��y8���L!0���^����zd9L՟�M��R"������R9J��FS�O���s7��l��(i�,P��Qzp4��Tw�$��V���ǹ��(��ʣ���P�K��)�:O8Oԑ�i2Psb>�ޠ�̄)$��V�ز��y5k�R��ٸ�Q�H&܆�W6;���pno4w�Ѵz�`�,Qo w*�\=**��@t��|�)�Y�~�fo?�k;Ŕ�f��_ll��4?NdNsѾ�.���ʲՒ�51��[Ph)���na7ܴa3\k��M�R��v%r�j�i�%쏡}�7dX�hVLs��W�n�E���;�ظ!����0+4\[P�%�q_Q�m�x�dmrd37��5������s���߱���Je�gR��A<�h�Ƒ� !���Q��dT5��K�����ʏ~�����{<~��ҿ��?�:��x��:�M=7en!@.��ː�]34�"  σyP��V�v���Ϟڳ�c5^���sPdv�y;,��N�&���x�&����9>��Cѯ��r%m@n,���t�e�/��2��mW^zV�}H�
P���$�w�fA��jn ��gQ�p��2��� �f�\Z╞O���{w����F!{�uh�kQ%^J�/����^��`�{��gϞ��`3)S�t�I�R@ǔ����n�� ;{���㲳���#�+��N��)�D-�p�K�a��L�ɷ|X��}�46~5sӵb$�G�x.4�ɔ���d<t��`<���M���f,V-Hf|R�ج^�>����M�6>o���-�bͶ�#\ʚ��\[ji�U���ՙu�M��B$�+5{��53Q畀��bc�����Mg+�hݸ�6���\W�Z�g$cK&��4�s �%��OJ��汋� .����RM}�$I<��3��Ø�%1C56�����	G/ύ���]��`�M����������e-�A��L�R�c�m�S)!�?|���2r����ƪ��D�&���)5��¼nֈe�*տ����_������
l*��E���s^	n�r>�v#K�W����&��6\Q����$��L�U�$$:y��k�jM��gG�����`��/�������*b-,�S�^.��l����\�贪V�j������u�eW����:O��͕��nT�=I|�^���Bp��c���A8<A��&��὜v[V=��ė
��6S��� 2,Q�������y�|27�k�\Y(�|�P�D��!��_K5ڝ��{8}6��{%K�O���(�>x:��
b�L��vO��_�s��>s�PS�W�������<�j��M�Cd�oZ.�����pՙ��	[4K
n������m�����m���j�$���
Ʒ�Ym,�Z%�@�5u�����[OgVJ��~s�޺�k�����f+Kn�[El9[Y�ӷc&���M	홴շ�\p+�o��:f��P%'A��l%����\�*�sa��Dw2i��Ӈ���s�~����՚�=�^�7�a0����%;�p�]�{_����&/��	`�dUI.s�tڽ>�7�mwܷ�	
��d/��f �q��"( �� �:��V�8�S���;��?���~���ngn�x������g�G��lǖ�I�����W�JV,��t�/� ������e3���B��o��v��&-OO�t�G��ܹq�j����.�^�l) ���U�r��ط��-��jic��۷��A�/�?&��~lo۩U�������b}j�n�a��k[@	Sj�2�0�r���tJқ���N�����d�xu��:��smxk<5*&�޹'�l �cҌGj.�����(в�o�obx��h�j䀔ay=��W#�{0����ʰH��H����@��:םN�}�F4DxE��o7aVO�;f����y���ZE��E�B�����i�e��t{}-f�m�U�
n�B�换��)�h�Hb�Ӗ��;���m�T��Ib���bey�Z3[�Z��k8>;��ֹ��7�Ϭ��Pc�4�VM.-��¬��a=c��О=?���/�sc�D�2�������#Y����s���BQ�"��<C��+GA�s��K��#�r]��g��V�UU�^u:vvu�w:w�`�����@YL�����VM��	eў����.�d�X
*�4Mw�=�mHa�.�ʶ��e�{{V��l�^�u2�)A�6�T\�iw5�� ��w�X=_��˿�Ɲ�?�'��������27
ǋ�O�n���b�oG�6&���
�2�7�j���8�	�2fҋ�m%r�W(��ƾ�V*�n��I�
aB��[#��f*o;���y�j���g+{��w��h�=�L�.Ps���4���r*:�� ��LU�A�����$A@ ��e����#����bE	?Zt��-�4��|*�YaS���\�ç9�)�lj��0��)����Z�E���7� �2>::r�
802Vk4�����#��H�KYQ������:�O�Ot��QfP���M���/\��p�S�\�Ec�,�O�^�h�)��ۀL�M���R�-�����;���h���7�,Z��$�Rp[6�6)�l��Iq&��hn�k[\v,;_Y9��/�1+Y�
����d(�\\_ؠ߱�fi�墆Z;��5�Q���j���%˦�vuֲ�>zl�=ngX��	n;x���/�L��S�'vqղ�̉5�ۃp�Z�0_P�Ɵ9(����G�8'kʧsb^KT1��&�W�-;>?�˫+iJU$@<�L��tJ�,mJCz������Fɮ5ϯmwh;� �s��؉ftg�!i$�d\����F����\���!��	��ŜE�9�6ֆ+���o�u(�esӝB�y���?��ל$��v���?������Ǐ�7����D�6$ݕ*-kKF�V��:uS����H*�W��D-��Xb���&a��5{�~`{���W��=��ϏU�R>�ᖞ̭h�C�Er��Ҩ�ԝ�Dnח������*�̟��|��N�������@F�)#�
��<h����@q�B����&JvLX���!�S���]L+�ޗC���>���P2�	$��SO|NF�>����WGL�1��OJb&o�뫖vĝ@��޾�u�9���s7�έ$�2�[��!PFr�`enїB��@���i�su}a�N�#d��%7Y��?�y�>�K��Px��D��l�������-C��K;���X1g�b�f����[nUm^��*��5U��ڛ��[m�tG������J�b	+D�VHe$k��`g���|ҷ�|b�r�v�+�W���X.�=p�8�#�~m��{����p��Jp�P���H��Z*Z���&���{3;:>����t�P�j�V���ҥJ�
��	/^���'j��G�f�j0�*U+�����/�4�����Ӄç"��Y�V�;w��hj�����u�0 {3���@O��.�p���ٕz؈UdE���"��D��&FJ���{S.#B��
LXs��%�[�26���V���3LtK�Id���R�_(�~��_�׮�W`������w�a�d:�sG��?u2�ۑ��s�bC���O�%#�)����"+='	Ek���*"(��R�ި��v�b���>x�}x~dXfs�O7�[�����^�jە���i��C@��߱��ʗR��2.r�KdS�AD�A�ߵ�&���Ʊ���z������t�&bpĂ
U.VD#�A�(�X��Y𹬌����c�I�J@���s*�����
�,�M�Wf܂��/i��DK3���d���x��o8p4.J 5�;=7]����\O ��=�%�N�	[8���1��� ������Ȕ��i媾��95��ǹ�v��o;ͦu;7vyղ�n�RՒm*�Vr�Nml�(۲�7�gԓ����Vݡͮn,=Y	$^\�U"IH�V.��}Hy���۰k���ꅴ�+Y�F����Y%����]�� ��|qn���}�;�`8W�|�L���s�o�jŦ}|X�ֺ��ӣ�R��U9�C�v$��C2�V�e�/���gOl=�8�DF/~�X)�VsG�S������%kS���)����={��@�(#Av~%W��֪�鴮�Zs���*"��hj��+�n\��G!o��{�-8������\b\�|�lN��B�bI������)D��rà�7Oc    IDAT`2\�r*m[���~�����~��>���������l�g�����ٴ_�F�6��4*p0�1�晰��fF��t@�eS�7
n�M�rˈ=(7��ځm+6�L��OۇgG⬊��\[~�4������+$3�;"���'�ڋ'�uܘ!̴��٬l8!��#�:
nLC���j�����P�Y��,�xD��5@9x^�x�`%l���N�!�p���5�cASXi����A��?�=�ks2��'�%�gđ�Q�e�p^a�R�@�؟��~��� O~�);��Ӛs�)>K�*Y��[�.~�j>�x���z��4���]Mpen�LƷ���T|o�+���!�i�t⮹Z��?i�1LX3���W�ۨ��U=o7TK6b;��E�3�\jj��V~����V�l���K�+~lԷE�c���ŴU�	K�g��nU����,�<=���~l�|��Mf��"j��{
�[��m��7���}����:-Χ��5�[v�@�TQ�Xw��]�\I���gO��Eb�J�ԏ�pSokgO�	2B�2%�N�Y�,�ϋ)��k�)�~��j��ŕ���l�ͦ&��%��+WJV���aT$�8ln���J��Ҩ���_S���G�۱��3�����g1�X&c�|ֲ�ެ:vM2)��M.c�d�z빝q("�n+&�VO�w��_y����쫟SY������������Ӌٰ�pc[ђ^m�Ɗr @�U|cs���R����E,��*��Tv�Ɓm�k6�M��O?��^i�Y,-M0��-�cSp;�6d�ֹ�R �����S�裏��ʤ�Պ\�,�t4(�Z-ѵ����ց����y����ɡ�l.(*"d8wbaӆ>��&��sٖ���`(���:��H<'�){�'�t (����n�?�Q��	���N�,��
}5��)���z�ۉn&�ԇo�����
�2L5��ޠ:��D��4%�����l�u��� ���^�	�n���� �)!s�q��Ԡ!�u$a�b�����kW�R������=�`aTz���ڦW�����ږ�m'S��J�*���4|�ߵͰo���j٘��	�F�_I��N�v�u��{��O��ob�?}n�9��S;8�#��^s˘�#z���O�ً�L�K&dPs���v�ܐ(�b��Z"�JБcb�I��Y��5�4)������ى�8;� ,� �&�7~��ݽsW?�`6K�;�>�]���T!tJR2���wM�'/����ɳ#'�P�[s{K�)�r����T�6�����z���:1ThhkR����Rn�G��_/�׶(�1Q�t4�rrX�~���O����?���_����x�n��/����z>�r.��7�cqy�[��hb� pJ1hM~�����ʶ��u`;��S�����'6�,%Yǈe8��p�2�N�n�պ��̗2x����޷������M�lx�9��W�◂"�v:����(M���9J��uR�]�ߩ�乐!��
�q���n�_���d��3B�{����\�8H���B�w��ɭ
�4H��6;�<��s�+��k6�
B����8j���-9�/��!���8=7u�I�krY���Ʃx��ʌ���CBd�3sL��p�zMJ{=��\�������s��l��ڸ��a)i�r�F��M�I����6qa��ӕ�N�l����É�F��h5pP/&S[�f���Vsk$cVME��NX)mvo�dw��P����᷿kG=�ӧ�]E5Y��LÄ;w�؝�}KD#�&8\�؇�}f/.�Ĵ�^���;*IU����'o����ե=;V�n�XY��V*9t��Zò���C{qun��-u��m�w���$�@�Mj�Z��e��,M���_~��Ւ�-��Dy0m��u[]�89Uն��m͝m˕�6���؁�
�)��_��UO�AUU6W��`]��ØY��8�؋�kqpS�cq�e��[�_x����}nP�����-���?s2����rV����+���fI7�Ht)���(K,T��	�,�ִ���
n��-m��O>���?��r.��xb���b�7m��+Y�߇}*眫n�ط{�gvf�\��oLZ�-��`ʆl���W�-�$�]�J -��6�֒Z�N��ps���N�S��|��Ӣz�;htϽ��N��9��	�)�l������_���M�S���������SW�t
�t��J��xRM�3ї2!|����IT�ʴg��&CvJ=ƽ2�T��&��[$Ϻ[S&,�M
�e��A]��g��m��_���>W+t���z�ʭ$���2	n�1�<Om9u�K} ��n0Z�RQVx��g+�	8�]V�U9��ߢ�ݒ�ib1W�p���f��&��}���ׁ��k1�{�E���<y[1�N<6-�b�c�*KBg+节��`*�d�#��,�4���p0�7�Ä]� bb�V�mv�B�t��)b�.&�\ӆ=[`�X `�Q
�p�J��#��㰖��QCl�	���7����#&�� V���2��?8���s-�n�����XWq�����K�k��6B�h�������u�&�{NĤ�V�G
�hS�Bg<B��dJ����1�O���	�!���h2E�7����˵H�H�&�=}�T�y����L�M�?$���`*][�ZE�QE*����z�{�e���AOrHYr� ��JIf�pca�6.�����#LqN�""�Y��ҏ�{��Á
W��o���o��n���j�#����0r���v�
gB�����	�+�u�
��b�K�pZn`�T)�Wo���%�+;ާ� �XJ[��AF�~%��)t%�}1��^�y��(hO'���F�y�L6�]L�J�nWtkj��@(�ـ�,��U�7H��;y?ȼ�b�$+�J��#�|�6zK�ZT57����B�P�Hy,oC�W����S�s���ƪR�м���* nP��ל������H�S�2�j,JR�w��Pɧ�mu��c���x.s5_k0�}�AY�&�@�W++7��6�ع �Y#�@�5n���c.�Eɝ w@y�QSLƐ��aF|J0��`��`�h+�
3eJ1��2V�5]<t�dK�s����L2|���l��v��d�D�T�\O�j8>ك/��y��~��CX����	������=4�MDb1t:]�_���odʪ��^{�*���T�{�J�����{�Z]�RJ'3ȤHr��e���?�����Z�$-�RF��l�����a@�P�+�Vg�:��5E�i���cd�I��)`R�Ֆ��`���i:��ViTG����3�������C�߅�X���7
��v�f����/o.�[�Ꮔ����b�~���ώN?�Bᇟ��Rǚ���5�[㵛X���f|�X����|'�V����X-Ŏ��y�N�c�|0��/�F$��b�rU@�����\����9�H�"�
�T���e�F�)m������W����LV�lK9{��Q�@$�� �@�Օm�h4�u���S����ܤ��Oޝ���G��W<�m�m���������M�)	
z�`r�o'���s�2%%B���VJ�̤&
�5���ؓq��Y@S�l*B�T�v˱����� ��(�g��_�����|~7�تVµ��x�<���U�����*�1xVH���X�Tv���[�`�5�յj�W2O�Ĵh�BN��-d�*1G!#�a#�u�zB�x|�G���|�bxu���D#��~�!f���r8v���f4��t��4�>zZ���#��	��Q���~�3ؽ)�s~�Cj)
���s�ud�Iѿ{���^~�
���W�^-��Y�V�*;��H%���[��>b4�!��#�N!�߉Y&�$� q���	�3���� *�a�h�g�X��P]�M�:�R����SÒל���r�4b̧��}�yg�Ώ~��Y���F��R+c�`O��������]�����������L2�|��8��ri� S)���%�cLH�FQȤ��J�N�{?����+F[���i��^��5���m��@X��q�K5� �wŐ�X<"�`ZS+ƨ.!
nw���b��3xV;D�P�^�^�M��D[G�hvs�����{�qu��
ܹ���K|?�����f�X	�юœIq�O?~&�?��a2Q�l�O��(�rӤO6�^;�X� �[<�E���Ubn޼A,ť̾s�P�jaU5�~�ؔ���5M�ǣ��`D%@���}J�hة+��o��HkM�fi����ñ��%o&���e��eR�-�E֕���2X�Ұr�"�=���ǒ�V]̨��r�k��y��htr�%�&"SB���7Ǳ��ce͍Oh�X���a��c[j��nF6*��xD�$!sĶ4�M�����br׆9��j�\=��ra�]ȹ�f<�f&�g�<9��v��":C�������b;��5�]˦>Q*�����6�e2�h�����.�^���(@�JFł�R+ɒ����j+������]��H��nq�G9�DnV^3�.p���!S*I�%־{5J"T�=����5�\¡!)�4�yrH9_b��
[_H�'���*p��2�X.�Z����j���ܷڸ��E�ے�����6�xF��r�LV,��o��� �F|���Ԣ��������������}7����_[[�����Y�~���͞eČd��TyR=�"ORa*)_g��M���(-i��6 ����!�GO��m`�<\���5���N�р�?Ö7lK���~��r[ӑ�/��|s�[�����yY�tJ�dV�hQ.E�yn��	hf[�gBg�׫�&'��[K"��\��e��=!8Of��1fR��|�K��s/��M,�d�N|�IT����;G������S*J���y�,���:"@��_�	8*���܊@��Q�/��jH�+Fu�j�/%�8��T"�i0`V���.�v������7ź��?�7.dKJ��mԽz�-_/37{�R�^�o'S�8������0`D VG�R&���06ܪR<��'�"}� �V���C�n�D\f�ܴK�I��)�B��m��N��a��2{5��#�.���/���b.��	�V�^��'/�٫ßN�������7�x��Ũו�A2E��<J{�5�/�$xڱW�����N�^T��-��0��;�����]o%�fLW��
!�[2i����),H^/rq%u��-|��lC%�
��dDfd���B���-��CGX7͇c5��UH�~rE����R�x2T��lJ��O��t1��baLC~�-���7f¡K%��z&���~�?�`�GJ8?����-1s7p������խ����1pƚW��|�(����D=�Ó�#ԳU,��Y���wbIM��-�~�B�ݢ����O�q��?��d&�A�<��B>���E2�A�W4�r}e��6��h�+DV[G��x�����<�(��
�� L^�<�@jV9xM*�.{����R����N�m��m^���:����rPe�F�vʐ��j���V뜁(�T��-9<feŴ&���)��R��;�� �)&<NE?Q�YM��q�qDv�T�'���tP�J�ƓFod�����=@g�J�TPc�~����r�&��+�vi��d�tD�y<�E��r2	ر���V2�M)'�:�T�;V&|ɱ܆�uG=�1�tEKE@�\P�;w��c#eۨ�W�[&�B~e���d{�"j�"8�ݷ�>����g�8�B��\,�C�h���@�V�/�z�C����W����c6�H'�� S̢v����	��"|�\/l\_\�����6��1\�D��A�f��:r��T��y2�#�@C��z[O�
��1�`�9�M��\c�d8!U�蟷+��ŜpV��S�ș�a���0cw;YT��)�0P�@�euH*û�9�{�j��b!#m5�!��),c��� ����1z�\���Xl^��胂��s[���9�����\���pc�a`�E4��q������6pyU�����;�i�+��T^$[�A��������Ybg;�6�/F�K����'�PJrH:@��A�f<	X���m)y7��ڂ������s��Gn�(�b.?o������Q,d�k̔�y�2[3 ��!݅'�^�D�*=?����~陘���x�E�P[O�<�6R��`
��3w�{qz��0�<�LF���&��)�J���5]fǲ�#�C��0�dO�����T*�"��I���v�~�n�]T�c@�S��T%$��7�z�A�2a�/ �����Vg:���%���c���l_,�0�l����hw�+���&�JE$_�'��ĭ6R��7~$`��c���l�C8E*�E�T����a�FڲPv]�9�� �r�޳�ky��yl�%��h��B����N��}$�Op���H��&��}�ޛto�M���E�)�P?=���H�� G�9.�\���5:�eso.��+�Ѩ`��HZO����nuP�C�(���'�*{5�E2����Dq���pvlk]V��\��w�@�^��s�K0g)r-V��x&�R1+��b���F��w~��:�)A?E��8ܫ	����U�Xf��Y8�E$��v�{s�������X�,g���O��o��ʇiK�P,�ߺ7G�I�2�O>n�v+	�l6H�CxR��ZG�!'���ib�Y
��4�����@:Fx듊j����aÓ|H־�b�0�ꏑ���K�O���@1�Ĵ7D��^�ٮV�G���R!�Ѹ���Ɍ�I%S���dއ�{q���J�\6-	�|^�Z��J��E̽_E	��9�m��ig]5S�{�RP�֕�T���y����T�u+�8�X:��e�ɡ��\K "�M�H�'	���Ȝ����e�\��g�E����C��^[Ma>��u{���c���'P{bj��Tg�w3=!��ӝ_�̡%����㸂�nPsER4�mi*���uD�ʚ�T�h��c� ��J���'�d��%����S����7P��Hl�H���>�}k8@(���)^ʩ��� b[H�&*�%
�9�#a</��=A��BqV3�;<�:Ǣ=k|V���A�^B��?y�d�Ds3�|6�y@����GL#�����7��=?�����bQ��p��[ܼ�@����h�M���<����g���g�"Y������Zw����2g$͉���AC���T.�s�T���r�ٜ�GRw"��[ݫ�x��ӲŪ��^�|8��jE��hׯ�9��|0L��w���|8�o��ϊQ,-�|����>`�7l�`-�!���W��U�f�᳽����-��gZl�˿{g�Ӷe�����%�;*������?A�'�r���
��+s:�I� ` �v�JbF@����s/w- ��pzC$�5>)5�����E��x$WJ��ZR�I���-RVtl�dV�;�ʒ���R�9�C%�f|�P%�t�M_O���.����ݐ�7Ot�(�tVGlG5�iՂ&��6:]�?SvG�ws7�iT�(3)O�O�Ἃ�R��a��/��\��en(���`��V:Q؊�����'+=����0൪��Ǫ���7�8���i"���_Iˢ���	7JR��ǿ�=��(�y-��ও$fI*gBUH��J�m� 䌹
���3�;��^qj��siK�Ɉ��l�	��9�98�ֱ �A��	nhB@h@��"��w}���-��1<�����n��4�t�3,T��O�|\*�ϞH�B��52�����W��-���[c�!�(����?B,W�a:I`ty���T�n��d�(5Q}q���c��M���q��\�<��%3c����8|v��/>F�� �Y��޼���뷸9��b4�]�N��8�nMȾ�i	o��a:��'�
s�MJy�dJ��,X�1�jj(p����i9�j�Z���|��~Z6/P#�ۛ�g�B�UPȤ����֏)Z��`�)�-E��f.�q�93L��b:��g���7>�������wg��e&��O�R6��T�I���)~��r�$f���T��k��b��ʕD�d��d    IDATmd'�}��)'_���	���s��<N.��D���pǙB�9]V.2�tq(�ZA�. s�B"�F2�FR��i5CJ������=����i?���#Vd���$8�!X���I��M&��^X�^�YϤ6[U��/]�iN�xhy�	��7-�"��+�#M�U��\G��R0�*-q��Ԕ����Z��[i���
h� @����� �w4IX7�OޗV/����^�-�~>�D�{���y�@ͯ��'�R�=:�r��&1P�5n<~/S�y��[[���L:p���I��+��-g�+g������S�\���_lO�vS#nK}�\[���\�lR�c�o�u�3-U��'�4�S)�3��rI�T�[#ܿ���+��8�b�]"�l���c�<�`*�}�l���k���0����[��*���	JO��?l��ˊ�����kܽ�0�C���
�N������@,�W�/p���o/`��HE�==~���=d�%�r�-[4���R�0]B�6�8l�!W�0����4�j�e��n�D�M�l�V��AC��l�n��^������Q4+%�3Id�1D��������ho�n���!2GKN9�����?��&��̭eM���z�Z��@�X��^y��n�Z"���໴��$G�*�����d��a���9\�%nв��Y~����R N�{	9d3�.�s�up�/�&��C!����4C�B3!�FIDś+-+�d:#�����"���^K%`���񀹌g��<��﷜Rq������ �[G�6�����2@��&��>�f���<.=S�le{I�#������ ��s�\��R%�VR�*���T��RY*<[R�sxU��u;�]~y����F$�r�J:��&���fWm�U�P^�ⵉ�hY��a���\�PdY�T*4�y?t�LS8��l�TD	�BkVo������%��]p�E���`571oa��X�$�����ā#���ʥ���Bz�@nj�f[���ǧ�
����XT6���6��9���5��lW[�d����>�`��z��ͫ��_����4��WA�g(�!IZ/P�5����~�����c��5������Z�ı��q��
�o.�24�c$S	�Jy|t�R��d���X�)eTCtzC��3�j�Я�QC��D&�����/)V����5�*2�JbHY����Z����fs�������sD�;�J6�Œt��_��g;`
a���[�֘��^bKR"���?��������~��k�������v̈J��2;��
�h�k{xRo�ImO,�C��Ba�vЙq���q6@?`a��"WR�sI��B�֎��4��l���D�Y!��!��!?���N������:���e��u87�:�r9������իW�I�Ғ�e$�L�q��]����=�S|3�r��.X]�:ANoP	���7��*�B|���d�dK�������e�w߬�p��3Co�~U���@�����}�<OJji�c�������BF�y1"@�L��uo|j�C��[&��b��4E��G^��� n��S��|1�6�{�{;df+f@�QX�(�d�l�ı���.Ϲf�na����B��h�|�bV*�Z���i �� 1���,Q�,|R,⳽^4ȳ�]Xx��K\�>Ǹ;@�V�z<Gu����c�=9�]l�h���������)����P>�C��T>y.�3�|�&_����9��7X���'�(�h<=F��a�4�~�GZ/�0�~����|�p*�\��Ƴdke$H����g	��;=��3�3��T�TD��P,�≄8�0ǖ��w���E��H�e�ptr(��k���`>�����hЁ1�¿Y	�U%��y$S11�\�ic�Nc��εqg[�3_!(��e)��g�}��������/Ҹ_N������m��lKiR�M�j��r�l ��|��n��#��"�(�7���o]���6��lmI�a@?)JP���3��k�;�_���O�B��~�$b�
QZ�/׈�H��B7`�#z��@ҁ��2��{F(�b� ��ъ�s7:�L��>�'��g��+�g�#ٍ$*�Y�'��z�}mv�!�nE�}�c,Oz�R�{G���W Y�{�&�"/Toa��PR�s9�tZ����
����E���o>�<��&�f�}�
Lxna%w�kEp�~�l�*�']���ˆ6��HQ#xQ~R	!1�4��J"��4-���.l�ʇ�V��W����	&�9� ��v�$�h��2QlRQ���*��a�2YY��]��`�~�ppG��A��C(�>�~z�-�ȸk$�&r���i�Y>����𢹇|,k2��?��g�������d��}�?9F�� ��$�����o0�~`��p܂1?OOP}~�ҳSD2 �-�_��sv���-���]x�h*�j����2�GЅ����/�0�}���2�����WQv�T��h&��d����rAa��;�О�	n۹x�e�R��6��~l���]Z�Ϧ(�r(�S8x����#Y⹮���h0���F�6��^�};�*�22�����h1y,��4ƽ��~��s@��e)���������7>���_��^o9���9�w:�"hl�f�@� ��?�dF� �\�T�t^ldA���1�X,�8<�=S�6>�P4&�O	��p�fIٿY��ϱ����OJ�Gl鸻�"-����=�a�^��X���A��9)��eɊ��&���U�\F�Q�Ko^�n�N��

����QY��R�̼��s���R�DUV)�~\�4��JOX	��7�F�=��<l�\/�2����9u�W�ɤ�X�rK7�������R��\1����
Vfo^��<gRM5��2�K~��FҸ��$>��J�y(䗙�mbm/��,ȟ��65ĴΙs1���e�bidp�V�"X�`C`�SP.�>?����h&�tV�II#a7S�!��c�gZ�
;���0k��2Waj k۲Xx���{��p���^���粡$_��+�*��e�i<yz" Whԁpk��˗oк��AM�҅��������G� $ˇ(0�q���2��tZbC����%pp����R�� 7��
��
��G�y^-M$*�}t�t�e���qʙ����G:�F�Ԍ-DF���[*�p$��r�Ao���;<�<`<�4f�V��6�nTU�H�8�k,�y�}��a���d �]�ry4M���H�pv.Lw���v8�I8�G�\�i��kozY�g��'O��-~��ͮ=��wF��u�Eh����1�X�a#�V�� e!;?��,�+��E��Ƞ��	n{��k���Zyj���ٗON:�ă��j���5ͅ��&�HЋ}�ia���l��1���:;	N�IE�Md��E*OvΏؚ^��U~=#��r�уJ�/�Ei�;\�����H�w��+�����Hd���]2$��ύW�uU���V�7�
z�-<& �	�����Y�`x$c-��n�X0L���ȹ���T�x��XL
��.��]���2ó�
T��A��&�+_P��E���_N�v�3�i�b����'�^^�䞌��	�`Q_�#Z+`�I*2H9b@J��]���Qo��`8�&��?&mdj e/M��(�>+W�Ǉx~p��k��������h?t`-LY>�݃r�b1��^<C�B��H+!���k��X��1��)�0N����}�	n�lMp�g_`pw/\��f� �4���v��D� �氚��]?�����x�`� ��
�����d� _:#�qk��}��D����������"$^Gb�,��7��w��)���z%�R%��~�JY
��a1ui�4�w1��Ǯ����♘(�掋�vF0�y(��f��z�>�i�Eg�n����ǧ/~�7>T����3�����kcZn��W��R
��[�Yz��H�B��ɇ�8(װ�� Ð�@![T��Xy=�i/��?��?��c��?���-<\\��$7��#K �D&Z`��� ��(����ᐛ�x��]x�����l<A�w{����!ĺɫ�x�2D��ƪPY�+�%���1W��o[2%�"�H��ȹp��w�M����բz�e������"�*����6���c��9>Z�{m�n5D�W:�Z�r�S-o��Ĵr��' �ce�X]�I����{���ڊ\���CW���Z����<3~p:��m)bֆ?(�\(|��wn���*���xD�2n�"��b؆����l��k���ᷖyV�2�Z�x��.6*0D3�-B�"s	�B�;Dzn��t�i������^��L����s!J���Wr#� ��(^|�\fQea7>��]�Wv{�(���nOE�ѧ/�
Bpds�2몃��3L[=X�1�[�L�z	��Q?�G���Jc�����|�G���P؏�A���l`�~3��
��!.�0��:�\�S�T��b	�JE쎸��9+�;n���4�]M��B��A�VD�ԕ`Ғ�^�`�QU�c�E�R���[&I�6/�=�1G �`��m�E��H�#	�V*��/�|��~��ү�|�q9���|�k]c6]u�c;���(������)�1׏\0*�vP�K�JYή��R,�Ew�#�c�VE��0Of1;?�m�p��%n^��
��"�YrE���n-aNXb��8��o[b���FגD��<E�j[�����Ź����H��9`0(rn	���Cً���j�J=sS
���[Q
�y	��RVn٬���څ�'���%������,����MD�������������#��0Y���z��K�N%����RTZ���0B��Rn7��^=���i�<�MW�J��$j|���f�RM1I^�z��M�����/jZ= ���$m�&��X@�/�y���� � 1jO��"s7r�)QsKQz.��{���q���'[i�d�."I�B�7F�\����;�^T�h��2{y}�/�x)���RG��
���G��|���Z�����_}����r�H󃨟���'�P;�G�`�L��ww��'��f�i-�ݹ��WP���������nm_�a3] �#�|\G�YAn�&9`n���ઃ��;�:��ͨ?:�T�5�kud�e��q!�W���Ad`l�iG��ֳ�A�V@��6�� ��C��G�.&�.Lc��������#Ԛ{�R���M|ss���0:�-��B3Ä'��[.��;��󃵥����L��v����9�+䫑U�senf�N:�|"�t ��j���Ar�G#WƓZ�bqnE�t
���N��7b������]�;�������9����9;�raJ�Z�PF��%g%65"��m������"m�"r:�s�)�+��	���/_��ؒJ�iX"���A}�"V:2{����OҢuCrO=p{��%��`0G�{|��15x�g�xdګM��tK*6GA����Kp�-��f�䴆���)+ts���4�|6'���\���MR��>{��Iɼ?��T�ތQ܋=�^�?M*?i=]Y(��Z����r��}4���g��<*]���\�@���_�HQ���\`����FR:d,�H��D�b�R�L>nX���a�v�l�O�5Q���&��&(�.��^�8�P�e�+`>�7/_IR���h�"7�y4�ѓI����8;;ǛoΥ�g7��
�HH��O���yr���p�F�.�\��?�\>��m�\��i����ST������py���ߠ{v	��"E�U2��i���u�B$���F���g��n=-q�ϭQC�^k�*|�� �='_�^2T���3��a�zYL1i"�kt�uz��X�3l6�T��j���ͺ�/mt�3|qq��6 #A�Cw�b�[cKC�Lz].���֏��F����w}�.���b��w�ydF&6���=^$��T
Yr�躻� �	�K��-��/��. �|R��|i���e�g�(��XD�a����"��׷x���?��x�b<�R*+�Yl�7�%37j�ș���h>ň!�k�B�u�
�IKGyOR�to߾��� O�D�հ�N��NƔV��+=���j� �u��7��p	n��R^�~�Xy�*�rC+x���n�Ҷ{���
����t���'��剜M���\u5x�6�?#�Q��� �cd��L�m�!����-eӤ�y���3������d �W��[��hM��ۮ��9k��|��e8����lS@��`&������'HW��.&����E��eT��@<*j�B�"�K��8�~~�>v �׬���r�4V�,�ܲEg�Sz�e�(�R�N&x�tqvv!x��7^��!?��%�+E<9<@�T�M���K\�_	��[bΓ3��4N�����2�Ak�7�����L�+[�"�B����}|��J<_n���K��|+ˇ/^�S1�=�G頎��X��X��]�pw~c>����w���ZU��T��!��n�>�����۵�h�7+�;i�\�H)��V�]*/����t�Y!����l��CXX6�c|~v���3��;tyQe���)�]�ҙ��t���w>T@̏_��ڛ�f����9��w�g;����&D��+�����p��*��1D�FX�w�掅�c�^��>��Y�Ц�n����#3c.&�wW���#h,�DQ�&��
~J
3TE��e���v��6�L�漉@E�B2�N.��^O�!RdS�S��liEs�N=�n�z��\ϩ��&����&S��~���x��X�l9�"�B'��xz�o�G��Ĳ��*7]jAJ�j���d	�zs���ya�ǣ�C�������d�_]]���n�y\\H[I�;{Tϒ]��Tk^���}�b��)yl�מ�$AY�+�K��h���t�p�a��^�d��.�ٚ�� �M�|x$�6[���0%�+Y���"!1P`F&�5I`�̎f{�����G׋%w���Fz�"�d����h����~"�&�.t�5l<�������E��o �l�2N�MĂQ�Y�}}�G.�%��+�pZ��5�t���>N\羍���x��[�R��l��*>��9�K�ŏ���9�XE�M�>ca�A4�`��1������u��M=z�s�8
t��ŭZUr1��<;�j�����P`'����}�(�b��n`�V<t1�,o>�Ҟ2�d�z��C�
14`(�]o��.o��G�`�ݠKL��4E�Ī�+���������}�PfZ��G�s���Ͷ���}~�l#Wl1|�6��+�GH���f�8�5P�����d�qE�p�x��d��VʺgG/(���_ڞ�C�pL�I6���o�#��"��µ>B�$H6%�ML��R����@�z���-�_ɟb'��[���������`iøE�]����S�w�&�7�w�K�<[TO,/���2���)�c	�Q,*��J�@(�U��yL�_�|?ӄ�����荨v'���u���Ǎ1�!%;cx��q����H��[t}U�I�kh���%r� ƞQrU�����E ��!���K�q&H��ͷjҁ�s,O5H��h���B�VA�ԍH@��h!���IiQ-�Ffr!ʯ����@���!usvg��8�J���`���Ep�"�b���?�"�)"����x帲�6Zd����IW��-	���~��v���c���@�7�.��J�u6F.�ē�C<9=���G@8���+�˟��.�BK�PЇx"�J5��}���L�%�����뷒��J��P?j���H�8�[�^ߣ{5��Ӈe�drN�:����z��D�.�]�aJ�x���Zvȕs�4k(��+��,:W0C���+���l�F�f�lЛLq���G���[o���!� o0fW��I�����(�zX��n1����L��PAn!��W[Y�7�E���׭�ɡFo~��j�3c{��I����"j��i    IDAT�C��.?��落�]���J.��4��W�u&�OM$w429�QI��썃a��d(Qj9�x[�:r����V0&��6lIy2__\���* ���)a}
1`z'�v����⼽�y9�Z1�r��ß���#�����T\<<�q�{���[q��ykZQ��j�x�"C�u˸�[��
��=x�r���1%��gn�JЏO�߭I�%�_匒*"����}^�F���N ��G#16pL/�j�4�JvG�ӠlJ�z�m�N@jAw߀O��ù�d]:!�x
�{���Ÿ����V���,�q+�,Z@����5VKl�����Y����"=_#ҟ қ�ov�C���<��z���V�����S�L����h��j�J��
W痸8��|nʅ���X,�T4 �����x����n}���|��7h�wT�R:���n�t&��|�����'r8?������Q:�\R�*{���(��J%L��܎0��,�;a�ͥ�R���X���,,�!�NI
^�e��&<�E��C�YA�恛�¸3���p��9�� �� Q� ר#S���L���?��Co�BJ����]/ѧ��	&ާ�V%���'����?�k�w[����k;������J{e��1�:��0#a!��P2����'[��rO�PNgP�䐌%�1���s��ctfCt�	�[>����#,ɝ��zY�&{���*[=x��K��.6�)B��T�\9k��x?��d�'x�ӕA.Txo�8bT.D#R���C�*~���<����@N���i	���c*�NW3"#y���S_���=��~���"{�w�6�^,o��� ��k/ס�?�6��I�ע�V*�J�ƽ����f*�զd�z��PPU�z�(8�����W���d'yL�v�.��C�p+(R��h<�~PLͥ�<6��b�"
Z	r�y�-�9���"Ǔ4V�c����.%�	�ޔ<7~� ʆ��J�$��!�-$+G���0l��Ê2��� �p���M$�r[ K9g���-0�,�z)���<�Cs��w.ұ��"�"6�77w��@�3ڏo�tK���X�Nq��D���s_|��/oE=��
M4wk,���lK��$��}��7�mY��)9.6G�D�j	�7�\<$����+tG»#RG���U��iM#���.�,�Ɲ��\�b�/Ԛ��HT�@8�����=A��KRo�B���(��,2�V�t$�����.SX��xm��e��T@�V5����T���
Bmi���G{��u+6��*?��R�'���s%|������!�>J�63�t[���04�X`�u�����Fx�1�!`�-'���r�P@mr���W��,���6������d}o�+љ���X���J���$�ҋ���<iy����z:�H��QfM��hsͶM�,��G�UA#���F�L�ו��܏?��ӼU�*���
����y�7�0��R]9�@_6�J���R��r�G�$���ғ��+��W\n雷U���s��Z�%�6��K���7�NP�e�"���s7m\)3��J����ٯBΟD*K��{ϭi4�J����#lJc-L&Χ,g1�.�[�qf�s4J��>Xۥ�c���Qy ����.�IY
m=�(��n���Vl���%���D�-n���z�S��Z�͚/1[ذy��c���Y���[���(g3��tm�v�+%f�Fd�!-l���A��c�`O>#����h���2&�W
����6�ңN���/��縼��
;��N�l
�d�j��� !�U4�|����r��J2":�b�$4�\��`$�%+��)���` �U��@4�C.���Q��:����1��п�bxӢ�|K���\�rN��cU���������̂��=.-ٔ�S��4-ؕd�wj��?�`���?�ӽ����ѿ�w���`�b�\��%
�(�֚���3|�<B~�g��NGx�ў�0�-,vK6����fxp%W@1��=]����V{T�~غ��'ҿp�/��Α\�P��P���	B�����$\����d*<+�X��$�72�ecH�O�,�M�^��!�f��ɫ�-B�[Uއ�̿5���]ͨ�[���,M!�OA��Ymi����*�N�����k�4�����W��6]!*ٓ2�d�-U3�p߅Ψ-����K�)#��d2R�恡�N��ja"�n�Z�8lzq�^�������(�f8�Zy.��q�H�d\d��M($|HJ�2{UDEL�B߲�6grB������W$��{���3����8�[P��P�c���(7�R�Q�`�ߝ 025�i�%����]k'���Spϋ���|D}@!�@"@��mY��p7J�F�@�}M���ר����{���q��I��?E��C>�F4�GķC.����$�Qb2���%��Z��E���8O�!�I�[/-���,���>޾�@�;����k4�G8D�\@�IϷ�����2/����j�����p�pp�r� ��oV��� ��7A粅��#��͢�it̒(#wPG�Ґ�m�n���_^ݡφ+����Ƙa��b �N ��/j��O+G����*�������c����վc����p�>_!��\p{~pױ��MG�h��q1��a�IF�biJX.��7�̍$�Ù.Dd��7cf2a��z2�]��!���q�0�J*}~D1C6{�O(I'�'�툶P|�ݥ��^�Cp�F�*��Y�|:C�%TT�
A� n]	�aU9	g�6.4���	ݞ���K��T8G�I���ŅG����jꙙ�OU��7�<ꅖ�)J�ڲjw]5Ƞ��ᖶ١
���o�[U~JȮ,g��Q/�5N{o.�Tj�A�n�����c:K:Cu�P>G��:FUn;��1x�3�/�!Z��EQ�.	��pS��0&[Sl`��Q���vy��&R��ɽ�(DqIbc. �QW�)���H�v��+�zS�:#�b��Kq�`p+��C�&Y#	Fr,B~�C>d�t�وj��6�9�%]�	@BLH�"����69r�=u�cI�_������(���|4�r.���:"!:o�����3Ͱ�`$�H,�L6��fϞ�`� �b����ί0����l&�p�Oq�X#5Qi��(�E�O��f���pK�(��?i"[� B��0�O0��c�ؿ�[s�p���
G{(7+s>�|l⛋Y&̃Q��"�x�&��?�d�D�h�J�q���>�p�G_��G��?<.ƿ�sL��.����wf�!�e����)^��(�F���nǀ��
��J8F�r&w�m�T>��PF���:� �
��Ӆ�����K>�RL))����;�c76_n��EP�Ƒc] ��ҭ�a����l9�G���[�����[Hr��}�e���b:�,��ʍ38�Ex�'V4���bH�1�D�����&��Ǜ�i� ��Е�hD�W�W�XL�B&�H��O�O�����I�|����z)���ŋ���oV[�#a0U�cA�`!�����[�	p�Z�����*�*���L�V�ԾO�+8��IȖ=��7��LX�v03a�9�� ǒ��lQ	����҅�gy5҄v~��E�����by�s��kdV~$�6=�;Fpb �\���%�S,�%vk�E�G|/X%�(��Ƣ2�'A�ձiѝ�Z\�='�%�	6��"�l�V�0O$�v	���l�|�2�3�F�Q�V�:3���h�EB4F6�ko�$�����8���KF!oi�e�p�R�F�2[� Lk)�l��0gS1�t
�������5z0����0팰/�����`�b%�ړ}��J�i�:C|sy�o���i�
%��q��R��"�)�����r\�������g������њ��hi�ON�+�%)�oJ��ӏ����κ��[��,&�6p�X��r�S��
���\$����Xr��
�%R �����I�B������	LLM�P�d
�XR����2)<���3e����Km"PpH�PZ�x"�R�(�CVp�VחW*$��U8����T*=�Z�o���/��Tt�5����Z%��^(3o�]z��L,�|9�Y%qF�J��wޯ̬��I��j֤��χ��)T	Ъ�'�;,�Jl���U}�����+ T35����U�xo�;RnB�.���5n�U%��PX��^����ن�@�Z*��$sXA���h�]e��N%"5����`@^�q�Q��(5����u↗��VU�a��1k���Ap0�0�n8C�^#���G�#���|_u�^���3�����W�B�
�|�88��^?n�i�J5ys\X��HJ��,X��J���\��w�'��4`v/j�'#���a��/��;H�I�UՖr�asܵ��`����u��#!�կTjb?��d%��;r/��0���YZ�C���(9==5����B�}i?���tv6���T=��&B�,�n[#|}y���N&�X�<Ņ1ǔ��8g�!�R	������pp�[���A��?|�/NZ�ُ���9\�Ƅ��p�������>ƧG���Cb�ܟО�в��.�a���JDhA�6t��ʛ�L���r ��g2�'��o�p��7J�Cd�4�����F����ȇ�e��EbUē%�L��5��Ż��&sg)՛�&b{�J��-��8�Ʊ�ͥ��F��׃ojIil)��hLȾ���eՕ�V ����rԼIW0�M����(��C��dn�yM�1ռ�0[�o�di��/�u!�͵��&N�BD~`\����pQx�����?|�q������"�z2Cs<T	Y��Qd '�*��M.U���~�g (j�M8�u8 ;��e$�Xg�21�ѐ�~(�ߐ�A`#ǎ6��M�^lE�RV(|��0jr��y[����
�p��p*�#7�;�k�.��R����������W��cZ�(Bz�$�)|�CQ �	Z;�K���=#�*��w��Œ�g��NrL��p1��/@��` �-�O$�W*�89x���}�3pG��q"�>�L��U�T����Y�$:���v���@��HD#8*W���JE��	�'*��DxrQ��mq�@�V���>�NŰ�l�����Z�d�g��e��i<���3���A�dz��)����{����_�+�n?��_���?��O~�kσ&)bK��l���~��_z�1��w��,�7p�w?��a���d��c��oŶ�W�VXa1�T|�BQq998T2�t󵃇��\_�3c�4�"�o��v��[p����"� j�^�Enœ�-O�v�����[��Ծk^(p ��pͽ=%�Z�A�VʞXz�2V�"�@<�L{����WF$�����H��#�G�ǜޒ����kʉn���y�*:N�_�Pe9�<n����4J->�;F���zn������7)�@^?.�m���xK��%�D�:��|}e���zt�;/]+���!PJJ�t,բ�@�y"S�W?lZ�B@*
_:)��n.7R[Q���2Z���2��{/e�'"��t
�jyA�z���'���!v^KJk{n�y&ň�7��)i�d�C��9b�*A�VM�ֽ�m)����b�ʙ�!r&�z�u��o8�X;��!׿�ʬ��K����[à����U?[�P���C>�@�P�d7����%���Rnv����b�ʛz��Z��L6���Do������c#&//)�������rFc��������X|��2���P��$u~�\�WW8���&����T�(��b�m	g��'R�f6��������?��_m8p3�?����e��DW
���ǈ>.>=x�g�}�e
�����ږ�Y6�qF��-��v2K�+��C�B=_D����͞l_���g��н�{���9�M`!c ,�I0�%��U*aP1`��H�|�*�hI���ߐ�\�*v� !0h B���S�k�����<��u�(�ݪV�ӽz�Z���>�3|���r�V���+�ҳ'�g_�+�l�e>���YM59�_�-3���%��j�h+�1�E#n�Ή�Dvފ�GR���0S'Ǒh��d�Q��{=;���ݞ�	Ȯ�ce����l�.���Hp�T�2x`�$�}�Q����>�JSZ��Ƕ^�4A����Ȗ`bH�~�A�^J=�)�;�LDx��������:R�BY�k,$'�������#X��^?u�0|_�$qz�pu�	��'�49�}����&p�f�F�
��ՂmZ�V�4��9�?g�,���[er���l4��GiϤ�r�����m����kv~m��=e�� r&ȓ㯠�6Ityp󬖬�6���7A�!����r�g��!�甩*�I%e,�ט�d�y"d���տD�gy��$�=?�lN%,j�U�u3�`�	�kKVY*H~��R`wOϤ�v|r�~��'����G���H��]����F��v�_AoͲ��]�\�M�+_U(]�Ȯ�sa���|���������_|�^���M�`��/����.s��kz��ig�V߾�����ݯ���|�\Q�����A����������_��|�[�^a��0�gx�t�],�Ó����qz_'G�T���Yϣ�g��������:�؛m;�5��n�Ȧ�pf�vi�=b_y�Ծ��M�g���
��6��p��<]�FfHՀ(�6�8vXm(E�?��)IeY�+�`}m�x�%�� ��SJ���6���\���s��t�X1-n��߼/`L0�4�;�gQL�M7��MY�~�L};Xt+�t�b��':�g1�L�3�=��2hq��X�:{����E�U�@���e�K����᳐�2�7=%(�-�aQ�PP�����it����1�h�4g�O�|�rG�e�6aW�GX�%�J�v�H�׫��`"d��!}��z9��3���@@�˂�)�������C�,���ϖ�R��P�-4u�"s �y��"�NALmZ-@u��]�!��ָ�ޮp�B�WJY�h���&P)){p�Yl�sm���
��%�Np#z�*�0�X�ժ���#�nP"��W���2#�E��������w�ٽ���˯��J����z�W6��Z,؝���?9��/�W��4����������
��|f�J�<�g���e��=������ˏ��hj�R�����m���6�� ���rR������������~����w6U;��?�?~�ӯ<��>���������~v���
�[9���恝"X�:�Y"��ە�լlSdƻ�
n�r�p@���;w�}h�"�%g[��lh��7��o�n�n��Y�ڶ�zŬ�g�:��:%2
p3[�F�9�Xu��rȝ:��s_�,jz>0"p�Eo� ��)����4�ِ��B�da�G-D|���.�T��h�z�X|4w���m��	�׬Tv�/�O}�}����q��`¿�.A< ?��˥Ґ��υP@��.1WL�����1
	)#�v&~���T7=� ׁ��&�y��PV{9���Z��[�m2z�AḘWE0�n�@X��mV��9��x�Z�U,[���[6kѫ6�@�f���2O�Pɲ׸�1�%0�����`f���*������4�=	4D֚����%�1� ����ue��I��ћ��A������"��d�ku�\p[��f0M"��^ؼ�TW��p��r53�i�'��H�KԀ�++���ʻ���=)��g��+���1�iU�vv|h/�kwv��՞���-�x2�
Jۨ^+{������4l4���K�wo����Vz�[;Ϛ�1��
2�W+��y����W�'��o�}������}��g��'�z��t:�_�ɭФZkCs2�y�+�hY�T��jU��a�f���՛V�m�Y��td(��)K��V�jj�n���jf��~����2t���s��糩d���(���	*�7��|Q�zSXI"�e��[sx�+�������L. Y��֨kAv�mH�vL/�e
MƲ��5�o    IDAT���b+��w\@2iĕ�M���Pa�L����i�+1�S�#L�@PT	u���2��<<S�ů9��U��V����E8�ň(U���<�o�c���z��jKQՂ0�?UU�Hv��q1S{�5��S���$��Y1#�A��a�vݲ���u���`���w�>�|��������@�UP"�.-?���U�� 1@οp�֜o���Z}�Q@pÉ+�ge?IYJ��kf���s�2��)'�&2�WR�O�zMd��)^�8��H���gU�5Vz���]JR��I�N�7���e�����&1l@Y�R��tf�G�eZ�Ygg/�a�#ț�߲'o=�0v�f9��f�;F�#�YԛnOkh9��ِ�iW�$ ���}{rym_||n�����ݷ~�j���9�۬��A�ʹ�Wkv���O��u?����k/$��� ��~s���g�aa�]KrF�g�*/�
֮�dCj�o��Ұ�����:
re�,gK�Rqn��`����A�F��avcϧ�^��|ԓ��t��"[�����N?Y�f4a>n�˞-nzV]g�
/�X���$�]�-�˞���$�=�!'e�6��� �K��u�i.=�p�w3E��N��E �$Pe��0#�Cm�����&�2iJf0�����&D��T>�k���x��x.��E�
�-L�SpSB����<�Q�iJ*W��D"yn,��K�	$�7e��F���5b��IN �7�����%����e4�rP����f����3���$�� ������H��qzNXH*H������s_d���h�:� �O�<�[c��e�t-�\��h��6AS���[��;�,���b�I)ׄ�AvD��-�-��J�x>��AV�0�� #���R�z))KD)�d�P6�D{��r�3?(@���N\o�,0��e=�X�V��߳�s�^_ʲ��z�Q��Î��tdN`���r��l�L� �4� ���hF}{|umO��ʶ=�X��ݔ+v�ڰg3��
YgVfP����}/��S?�-���/$�}����w<���l�O��G�Qfesj}j~p?�2Yq��M���,6
6�l��ם�l����!4	̠jk�	+���a_x��6�쭕l]/� ��c=x90r�#�]������s2��pj6��<%�1h(-6�"�.P>Y$�lg����'���M���J����	zIz�7��7��SI7;_�'���F�@�X�2��P����4��pŒO�.O&�&�:�M�/��|�@6A*I�4�}qɄW)�^�B��!GP��e�aŘkK�J�<��28�W��\��?��eI$��B ��ÌI�{<��mS+�K�OV)YV�T/�"�3�xvy�F������$^��6Ye7�m��M��P=p[�j��� �<3v�6*}V>��P	(���1��^!`�W���"�9������
n��@ځ�5��UlP�!���~�y��bM%�J��$݄�f� ׬��O��MX<����&Q�֠)�>!�Z-+࿱1��phJ̈�b�ע�1�=;9N��O{�aCkѪV󙛤���咵��>l�$�}��z�����Nl�nY�Z���/f6�.e3P�V��K��'������B���?�;�<��?�x2�^27���/0��B���G���T�{��W;)7�~�Hd�{�����ɽ�tR~����ϟ�Oۣ��6˛M�����,e�<��-Qf���*�L�Bf[��N��l�٦7�,����^O��X����CS�Pp�1㜪lBmr2�B��Zj�j���9��A�þ�+	K�g�p�,Nr;L��d�`�=�SyYp�����d��$ˁY��E�OS�r���{RGj��|rr�m��!!��M��&d�*ˋ�C�D�������)�.�-SY��$C��CK/�78%K���u��٨)�����ЊY�8�d�䁌�N�s�C�ߓ8%���/JS6������tO��4�4���[��S�Y�` 4a2���N�
|�iɜ	)��	���]NP�bH��������C���|%�$Y6��ua�]"��]�m�T;��a,��+�"���{KK�Âl,�*�nj@����U�L+)'�q��	n��|�?�^ P񾩐����:|׎TP(�i�PF�,�}���j��Ȥ�r��J��~��P�����زղa�*�����F[��ՊN�|����{O�}�>��|!���{/?�~�Ѩ���&�"g�]�TY�Y˅J��Z˚ټ���)V�^�H�V����q�>停�\�������wcO�.�rط��u7s�첦rx�h���
��XiAn's3��pj��H_W�&s��vX�[�\�M�Df��Jn����)t}s��7���FL@��V�l�F\�}�L��$���'vy~!�$�J4���X��i>���Q����>�/�́e\�Sq�9����	V�5L���21��E�㭷�;���W���b|'��M=�0�!$h���qdeLH'��������{ٖ	�MI�~�Zh�1�#�9=�
�=��5[�A�m�Q�>(z_<�x2��CV<g��g���J���A��\F�>�l
ZGL��m�곥��Q�f��1�A��P��pߒ�J*�S0�C��f�.���`�qJ����p)��a{�����f|j��puQx� S�7���@�R,p�W:�k��u�.��iLkc���9���l��B��X�&�KK)-A���Vз�/�u�
�\�{��f6���m��H�vrl�Vӆ�]��.��39<`BK��A�����O������'_z�����<ߔz*K]b�a�S�lF��޴�ZK"�w��vvرv�nEAW6�L�j���FDsіJ���tm��®�=�+��ci�A���:�l�b�T�?8x:]ֶ���a�J�$3�Y��58���Jی5�)C�g��`���0ǒR�I�``W8>q3 ��\4�ZՍG��L^WO�����FZX|%�#`@ ��Ni¡ �'��U���W����j���BI����*~���2"8���	�b
n��QI��@�qEl��� *�O�8z�<���m>���`�W��=7�Q�%w��me�ʢ_�d9UIFVN�Z�R<F!�˴�a�ʧ���P�`ks蹑Š���n����6�:%Y�e����^��W�b���֔��.lֽ�,�n���,���WK���\��䥩:�׌���Fr��I*.n_��`��g0�?�C��l��U��P#֍k8L%e����"б_�D�c�r0�ˮ�LRB��n��|�V���z��5�E[�8o�fS�U�ADh�-;�9���Ōk�c�<��n2��h��l���'w,-�Q�a�b׶�K�xPJy��������w���������S�N������7G��!��8塰� �R88�W��޶W�Ni�kP�e����ƞ��)�ܾ�t��hl�r۵��g�ך��ٿ����z��f7�f�����싌aD|5'sێf¾�ӄd?�m=�)�1�x�TVj�T���9�Aq��.�������|��g�S�������c C�1~�=3,�"@�' 1���e���J�x	E���$�DO�� Ϥ��lH�է�$$iS�>,^��ꇬ��3�_�l��X�4߄l(Q�Ȕ���{Ų���te��[��Rω,ǃ�U��]��l\7��evc��J�pC	dp�]��dU24ze`�d�ykɇ�Q)�y.{��{����P9݇@@�P�r���W}��{��Ҧ�.�֎�)�v[z_ҡK�\8"���8���Q�W��2���L�M4M��+e%��,�q5�h�$(�2�X�d���2f��y���c�� �T�6�H0$-eT��U<@������6���J���V�{0���r�k����'�:��y���Q}�O;V<A���fժ�K���\CC%=��Œ=h��{�|�_~����B�����y��b��ǣ�?}2����������X���/�{�bg��Y=[���p5�6���ƞ]^�h�P$�W������iw� d&o�LQ��{����o�/�h����(�'�.W�����o:�[~��p��g��e���� �`dN0E$3�ò����R�{wO��载������
��"�ʗ,���gV��H����MJӔ���~\K�wa���譄!��C@����0M0��.�A %��P o���l��q��v}z64~i)�a
Jl�Tn�@?u�i�"���@R�k�ۀ(�*�½M�,@eqN���V��-s~H�r[���V=hI3���7rV(x����4HWtf�rS���l�\.v%;kS�2&��rFIO�P��6k���V��6{ra��r(�T���.kY}���Mp�������pA�ԇ�G���Fpc-��@�a�a�:
(��yt�H
Y�[kI A����m��!l�38�D@,L���)�	�7��Te��R&gU�	h&�l �'��\J�0�P��B�HW-m:[xϊC��|FIڱl�c�r����u3[�Y�m�Y(h��v\*3-��o<���?�����i��?��ﻘ�?�l2�o����f�lHN~�XVv�l�?z��^}�ݫb�\d8o���.7�����<��,�u/C�BA�߳vG��{���V��mh3{�����7�ϟؓQ�VHҨc8�DzY�D�����[��b<Sp��%����r�]�1�����N����d|~q.<������,d�l�A�Pr���EmA���Ⲅ��t*��h8���ظ$I	�����q<��y"�9dÃY��l2^r���n�&�Y��o���u�=7��"XVk.��Є�:xy�c�������.�E�"ey*y58qXF��jX�I[���g���ռ�U��R�I�(�ls�`�,${4��K�?'V���o�b1�H��A�S�Ԓ?w`ǐ3��lyze˧����[a4�,jд8� �yo����^����L��,�{��;N�B
��4��=�t=(��Y:�n� ���(�&�TL��>�L�a�h�(�y��*.y�]��5/%�k��p �e��{d��TEFp�@������,��Q@E��-�����:0��!��}�S�.���r�Jg'V�sh�֡�E��s�͚����f3kWJ)�}��9��n��O~��v�����w>��y�L۸f4�;��}ӻ��}�;�mM�FΔ� �2����4�(/2��K�D��N�)g�oul�����%IJ��}�/��>�0����n B�ܸ������ʲӹTK�,��J���`l���֓��A� .n+���]{��6�г�=�̞>w�NN(��SH�n�U�X��#�H�E�\�jՊ<-�3-9�\���A��IC=�OF}.̆ͩ�$��]C9h\5�E���5}ϛ�^��HY� ق���Bا������	�n_p6��x�	����JQ2���ĢP��r��@����v9Uq@5+�oW�ЬY�Q�|������щ�{����^���-�E!RpUba�"���A�&���q^)�"���e�2[Y�7�����ז뢼�@j"?a���bV�{�3Q��$,`��L��ny��|������J`o#����n�����D�<;�w�֠���V��5�ibˁ��.S�B��P�r�pX�>Sp��9�/�BٮW:��֯3��e��q��oj���(�����4�V��ϡ�I��'�tڱ���mZ�]pf36ڬl*6�)�ݩT���/�9=��_~Q��'>��o�X���t��4�G��G�I7�a�y�{��n�A�j���y�U�H�����}�F
�h>�Ѳ��NG~�Yٓޕ�ś�ٗ�>�E)������4o���㚅e��3;�� �|�K��Ж ��c�/7ҒC��.���|Y(�a_e�6�\������$���P��LMN�%�@��y�C<�d˙���)?rqN�?���E3<Q��8�y	&(,����D.�E�^�R�`�����O'=�o���Z��eA&����I���dQ��>�`1�KS:J//���-�����V
��AJ�W�C^LO������u�<��+��R����K@�&8ty��o�p�����hSS�51]Z�?���\�z`���r��-�#]0���ڑ�Bqe�e�.�	�ה,��[����+�6^m2#���Y��C���(~�!��Ǘ�=�� �������U�6�}x�䔃3�x$�B�\��5��=�a��=@`9XU��L�� �P�F7)�2�է�YkTv�<����3�6���t(�b ��;GV8=��Aݺ����E�r��b&x���T*�?}������^������y�����F�o{:�~�:���H�hm�B��uT�er����t\�Dx�i,��L��邫��ɩٟ]����(W��)Sn��7����.��1)�4%��t�����@��#��ʿB��/49ː���*_��3�+�ֳ;�5U�Z(!Q%L=�68,b<�Ԛ�4�n�Vʬy:�E)��xU��vvr��f���'�)������#�PVӛ�L�T�6�C3��=�p�����A���� 
�JBʎi��}�ﲧ2��A��o
�)�iқܹ�sF��� �8i�p��u��?��^�b�f�zE^ ]��b�)hL�j�VC��jط�f�̏a�6eЉ�?j��P���i���Ƨ����le4�z�L8���e��p�'3ѝ2L	a�T�jCp��S"��4Y%h%7�s�S�+z�\�_sW )��5O�7�D�?�Y�OV���ٜzW�C|_�����L�5�at��]�������{�	.$]0^�>j�$P�Q�U"S��9����RTk�����]/�z~� �0r��X<�\��þ��`>Є��ݸ{�2'��v�5��ۗ��t�R/�肃-����'��һ_\p�,}<���[��w�φ�-!����9ɀ���2ApFo�:���۵��>9�++�=���d���*����n�C.��S��,p��A���s`JGC�)�76"SUz|���[enL��rZG�8Nz�D�� V'/�E��,"o0{&�ʹ����0���t���S$YDI��U<��d�2
΃�P��j'H�Պ�dH��qu}m��P�v6�8��W@4ܘg?���'H�i���G���ep�b:���.��Ѿ�+��(Nx2 �٭�[�T��oT�C��-�GPQ֕ \�":t�IK��$��yɯg]f�=I3r�'�# �U+p_��	ԚS��q������պ�]���o,;[�l?�g�� T���ز�L�C#�1�&��L(	9d
V����'��A�J��J��F=+�[�V��&RG���U��i�3� �C��Be)Mz
L�ju��YC�#丨,�N�%�5��ʶ�|UkZ��i�o���kѴ �ǔ�kG�e��foO甤܃�NBޑM;n[�������+Q��r,Z�wmsضa�d�٭��)�
�n��V+;��n������;�AA��g��]ϧݏ=���r1�������� �Ni��k�)�qSeT葐��)�n@�	h��`b�x%��.h�j϶<yixUpw��VCRr6p�a���Z��JTEd|1�	�� O&��z�����od��5`�j�:7�[����E��%,t�¿� ��t8[�X'-N� _z�u{��F��tI��;ׅS�������K�e�'��[���ɮk=��ؔ����iAv�̔�N����O6ǁ �c��x��I�ۨٲT���'�v	nd<�ʠ�a�G� (�V�J��L|^��d�"h8�"� uM��oC�	�L��x�S+��VǶo���U��ֵ�pd�4&�o7^�俇C)z��Q~R=�.�;|��s�R5䡦������W.��r�.�n:��m��	��0��0zy�R_!���Q�G�T?1P�&d�����ϙP��IA.\�����*�>�u?�����.��� �}>pc�@
L����TQ�RKpȫ��>j��Uu�V�ϖ�u�y�A�+�m%8�c-���    IDAT9�P�EU��Z��o}�{~�����/���}��UA>��?��lx�k�'��X�K��h�	�HtG���Z�!U�fʫ��p�'q���'�FΔ	��+L9�;nFK��`�$*��L�0K,��KSS�A`�'zv<n-���G�̠��Q��x��[��|��#�4D� Qd��r��a�'��	�v�}���>��CKʾ���I�s�xd���0h:Nm�ç��!��][�����rf�a���������8� ���t�}(��L����M� �(��:�����2U�v�6�e���N�ș�9eppG���XC�lf3Wu�v�,e��N�8��逅�E~���df��\���Y�?5{vm�'W����u����j���9	2v{}�ªA���^�ׁ�J��ɘ�C�����^Sp�EBy�5�	>[t(˘jb��b�hU��d|mq�&`� ��7���24�iQ|$��^�5|_�4���`��ɔ\���5�no Uq��t1uc�|F�����I�j����7��F��o�֪[����gwmV�X���.��bAgL�%�/�۽z�����?��o���>[���Ǔ���t>���K�L`SZ+xDޚͺ�	FZԑ�q��u�#=ήoq:�ݩ�W��D�������F�D(���se����f������
I`[m,�i�a�B���F�S7_�@^<T�~CYf��@�{�P`蚂?���" 9��O��֞�tlfe�X#��)�� sS�@s>pdpOS��sC�J��,�tm�X�)��i�% �3< �'J�ǧ��/�If��Pe}dRaD�����e��QR����8�J�l[a%7`�J��Fp�^�,W�!�	.F�*�(�45��W����﹬�B��Nd.\zo|��5�؁嬹4���m���J����f�L���2 �T�cz���]���DL�ᏂZx(HΝVC�i�!=ו%��с�5�,0�,+uMN�{AK6*��&;��L�KL�$�͠����Rs���r@y���M&6�u%ѕ/�fCY��qZ��;��`�;���6�d�O_g�b�d�j�7�?���j�f�㎕O�m\/�M1g�b��ł�;����y딪v�V��oy���>��/�[Jp��v�׷��{<�֮Q�o';x)�����"���N�����{��*������:0Vo*��p�4k
 ��f�VP�@�6��8x.�$���J�A�,Sl��8�����c��$���`� ��[dqh�!r	*�	,C�B���I=<�߱Forʴ�m%t�l�h]����5HT�B9�f�5�IX�[;Q�wI�:�d?ѣ4	���~�����70�`*��)`�,Q}���%)S\��fw����|���T�ʁ�$�s2;��(O�ذ��a������&��Ԑ���k���݈XO��,_���A�Z�U��RC��te�u�ʨH_�l��S[=���x)�VQ� �ȡ����Ź��xn�v�B:wP"Ѥ<gUDYMeodzW�מ����aM@��Y�}����P������rق�!(��X)#��	"	��`!��D=�f5�O��F9�Y�O�����Y(،���B*6Iu91'��TW���7A
7/�>�-z�Z���!���� �[��\{�@,&�׵6�ۑ��ۨ��n)g�]��|���u���T�{���K��������_��k.K��g�����_?����W�%�~�6�R)ѿ֨���.w�NS]4˫��7E7��b�7�M)��A�$� ��t��f6M�4��� ��!�(�sna�y,*&���b��Rٛ2�$z	�e��D�{��d�r�2�r�5e8=&�_}�`K��$((r�-iwR:����}��l$�s:���nXA��T�c��X~|��u�y��d�R2�� �f�[dF);������arB͊�xd�)�&�R�Cz:|�/|�eq`s�I!2IO��d^di�)X�h��W��dn�BI�N�9���$�eL�$X���������G)J�C�۪K�	�x�WSW)VA�t8���k�=~n��UfK�Ŕ���q�$Eӳ�l��!Ȇ�c��?G�Yo���b����K����=�kUeas��9�,�2�`M�ʲ��A��<T�p:v�(������|>�����5�����Y{�y�ӳ�v�����|��-7�����򔭣��o�w��a��I��Вj`>Ѿe�vƍ)p�c����VL���8n���sh�j�nJ9�*K�$/T6+a�h�j��~���g����w��T�}�{�������t�?<�����f�s �� C@��͚�o�`&�n�f�@qSPV�,�Ͱ�����USY8IEU�i.$pVϊԗI����LLN�NR���!��:�2<��&3����K�J����MI�z���L3����Dť��VP�W�oT�ϒVZ:b��sc_ߜ|����;ft��#�I���}�*���C���ی�;�؃*٢����)[4nxDSi�T�mr���ӽFX�b�b�ZEޣ��Yރ�a�Y'�+�ِ��
;Z�.�#�5�l�ԡ�ir��@)͡��%h&��k��-2+�t5]�,�Mm����o>�����f�������Δa����p�ۥ�9��&�zV�v[���hj�;���>USf��2�����<j4-M���3�XY�ٖ���b�0%3��41����d���H����\#A^�rY��U���'�\�+h e�Q-���H{+����nH4ׁCvO�]k耤t���+0��[�c�V�n
[�5�f��MV�D/#��=,��n��_wp�?�����}��ל�!yt5��[��?uK7�O��#��f�9emU�O��B��>���#J1*)h4y��6`@ܒ�n��:���R��Ŵ.�N)�� ��B���[�-�c�i�HNZMYJ�%)�R��i����Ց�1�`��WXo�U/�,Mk`"�� #'�2��O7%9ǧ�K�¥�@BpK=�0�I�C��������m�����~�JI��H�5�8]�]	�3=�Z�'� �`�	K٪lm��(��y��A��I(�5JR���d��(�������.�9ǆ��؉��qMt3�w�6d�� k�UKwp+�������.�]���������l%[<�@��K\m���3�b6J�nr;�֤L�	���ŵ]Fpc�9����6 �������ߗ�'t7�V�U�y�ɍL��P�b���f<s3���i�Q���م�rDɱ-Q�T��C�nq:��)��޷ZP� ��2^Al?��Q�?M�E6��Bpk�Y�����]f6vU�غU�\�m����|WJvP,��J���ux�G�;~�/$��
r�������������\��n�u��4y+��~WF�A|�-���ƣ��m�x����%ewn�+D��$����dn��=�	9�k����(>������Ta��H���PŰË2R�0?�DpI�$z�7��@�{� �ZM�����=�=8���U�F�P�^�.��S�()�Fp��J�y���|h�S���q8�饪��y��	'���E���,����W��}6��,��"���u�S�H٭>0`E]kMz�2�S����̆	��U�����ěۜ���`l��6ytn����[��*���M (��!�>�HP��E���f�)r�����vuu#@-A��m��D}�l����U���6�����u�����yX�$Z ������"6��]�����OBy��K��Bw*$���oHzp�����k��1L�^0��=3n�^P
�:���=,h�}��R�3� ��>u 	�:G2���l;�t��<��s��J��f�h����+_x�������#�B���?�;�\M��x6��Q��*�.�<���Fߍ@G�W��~\�` ��~�/Ђ��c��k��=�T�i���Y)(��E��y���"68ϊX��CXY9c�[��$;����)S� ��8h[ҏ#R�*�jLy)�AP ��7���2H���(�r��~�+%w:_���~�,Ӯ�}{�&:P��{x<��Y���h2�9��2/��"�>"��
�������ZYPG�&D>�:���y g�A�N4�4\P�z_쀘.'��^oTP�¢�Ǒ�q��PÉ�6I�o���_�z��噦�FEr�Zp\X�X�&�D:|���ͬ!� �Yn���� �&9�>���Ö7=Ӄ�՟��7�TO�̍5Jo	{T%�]���6k�ֳ�69]O�a�MC>���zJG*pa��ԗ2����&�^���"I�'����V�CZty)~L��dʋ�Ng��TI��2H
��|Ҝ=GVe�f�J��ЋeO����Z�[��V����O��?��?|!��7�蓯^.G��d6�гI�0خ���1Spc��(4j~������)��/�uR7����}D#[ӹ(SS��O��JRY���f�����TH��Y��2��ŘP� #s!B�ps�2Maԇ�N)���|MY	�@L&3?ф*G�	���C�[6`�g�YJ*��=��a�ז�a��R�K�O�^����bA�Tq��d��:F&����~L=�]g�1��!A�FŌ ��2�33����;A�� ��E�À���,�������#�9��T�ZVF_4Q����0=�t�9�D��3�9�l�{4�oBߊ@(tW][^�X�7�RY���f+M� YR�d�R�1L0@��� !dY��0��/Gֆ\��NE�q�V�st`g�
��2�~rue_��7ڌ��6c�͖�v���r
��tYM����/���)��`B~ QN
��{�P�5AAX c��$��$Tv����dj�� �Ei�B�J)\��\��N�*0���F�!����2�Z�i�c+�nE��d3�I9oVo؆uDPg|#%ރB���/|�������O�������y>��������M���v��v׈��sS�F���F��E,�.�O�TE�7YƢ%�J����#{��$����GV���ۂX*E��f;�c9!�h��@"�[=26�W�T(a�h@R��+)(]���#�#���[r2��~�6"'(=�oߥ
u�[�샒(�����ݺ�K	e����(?T�ǄU}��ߧ�dpd���̢Dܿ����Æ����Wv���S�^�����0�PY�/�*�H�M�3!�P5���(�e���c*�.������RI��f�/�h�re�����[,���]��&�\�M�Ǡ�i��I%�d��M�f�oԶ�b�����{����F��=A6��=�;�rv�Z���Y��?�/}�5ѯ�N����X���0���D�~����v���0�Iz�
n���<~�s��.9��aZ�ĳ��W�K+���mO���Tʼ(��ѭh�|�f˕�'�>#L��5�T(9 �a��S��9�r�m�B�η+{4�·��$.6�r���m���������������/(���;/��xk2�go�n
}[�3*������`b�'[և	�H�Mj�
�$`�������FѰVɦ�/������G�,J٢�|�<%�ƴ��.d\xR���$����b��f�E��t'&�����2��]��2�l�|��F�#�K��)�_%Ys2���I�.�I��{�/ é���wz�[�����c��11r��FL���馂�������DD�W6Ϥd�W�x�&ʰ5.ML��0���/�$"�ANIr��o�L��{Pp(i�����Y���n���#HH2Z�aȚ�/xWe&nV��!`ʤ��/�[�[A�3�* z��= R����֜��k�{G�Z�9�w�q(l����?@��A�f�����ݽu�̾��2��p�ҷP��f�:-��ւzV)�2������n�)\Q�k?�8"��(cCz�����B�[��j�%�,��%�(\��g�;d8���(S\O����봿B�l��C;�{�N�ݷ�ѱ�k%{�Y�듮=�Om �)e�TypnY��ڟ���/��/~�#�y!��7?��W/'�_s���G��
B���F��i��m���-��-PO���
�HpK����M��ϣ!@��e��UG���2'�ӗS?��D��F��5���A5MR#�dv�M��/JMACd|���J�W�@��썬M=92�(i	r S#��� DR�5ٜ	���Xh��-�T���� �kHs��0dW^����]������,����CD���|r ) �9]��	�ͼ20��GqJ� Á#�϶���இV�ы��J�!ƗT�Bz�CA�E�x����Y�K��;�E�R�"������y<&���w<e6����g�K[�a]�,?^h�����c�F����Ȼ17%Y.��M��D����H1ꓬ2*���K��T���JI�~���|��Y��ʲ��K���[�Α���+������Y�À�f �%-Wk�n�}��NFI�J�ddx,ā���5��^4�j���ߥ߆����6{9[ =���X4TK�.�	6�����<x`�<��ɱ�j{���k���5Xo��1�&�=���f�Ŋ�|x����=������(������\}��Q�p�����X�h��ܜc��d��$��P �:�}
^��C�;5�=�Q�e<�J7�@2�T�@�D�6B�2EY�r4�r��ϸ��&�p��x��@����9�K�J�CG�%�a�"
X0#8����)K���^�$�c ��-���o^	��I�S~-SIO���cD�, �0�`0 +z���@G�p���C��J#�� ��i
�d|��N �0Pa3���7ǐ!��hU�V�����+dw�H�)m�H�u<!'�8����3��1�j?��N�M��ӂ6ٙ>qE�O,�ۦ?ѿ������𪨖���g���'�� �2�q�J(Uܣ#��0[*�lΎ�-	MP>wC��zn�L3IR������=;99RFz~~n������BrLR�az�l��񉵡P!Ǿ\��͍]���@y�~@`�]!�����tj���2'g�`&c$��&S�<	s��Ғ���|C2�m�>�8�SD���������U�[?����=���|1�������̟��y~/����;:�y�×~�>���b2��|���r�ko�	nE��P�-�_�빵�Z�l�p��Cq� �9���j����0^���}�C��
/�Iu�#�/�X����k�e�����k
~����T:���Q��Bdd�Ѳ�n+N���uRG�z��/ԁ;�o2�ݮ�`HMk�?���x�,/�g�l�����P捃"��z��������h��,:�t=3cahV``ӳ�чK��ޏ��� a�R0�O�*&�L�f�$w/[��M��9AL$���-xB �֭3�I��>>�7���&���P9���Α~��Mwd���2��m���W�0���0��d��A��^�R���k�rCf	E��&���֮Vի&�R�[�m��"u�/K���7Z= e��<��T�5CFȄ�Ѵ��S;>�h�cC�׵>�}�� 3 [V~�AQ���:P�08�S�� ��K����0����@'NԲ�.X]V[-�޵��^����ttd�r�ΗS{6ؓi���S�Y�/1�JinknG�W��c(��]�g�Jp{<(�!)�@}p;���:������� ���OY�hF[/+�@b����Y���W;<��z/�T�$��())v�M�(�vt-ֆ�A�P�e��C${ �zn!���i�
J�C[�O�@��aL��EI.��ن��������a ���P2�=0=��x�~=,���tbs�Ѣ̕�2�8��=s�Sߚ��kk=�F����WG��~M�\�ط�c���'�4f��I���R�4Q�F�d#�\�x��D����$��'������u����dJ��c	dӅ���zL��F    IDAT`��X��Gp��H���v�"��#��%����3L��}TE☂��|%g�� �U�T�y�-�awF֚5�mȈU2^\\�u���[�	�Ea�igwN�谣�u}��i�1�WK���eEY�+x%z�PV�������Ԟ��O&�Tk���	bȃ�/�wP�P���V@Y�ӱ�{vrv��Z��%y�����'#�'������"��l�Ke{�� (@׿���ҏ������ЯnϦ�_{4���'�a�i�~p�H�hO�/N_�K�� ���9�4ߔ�ikR�*�p�����V�~�H�
P,8�)�fz&�)�����ɣ��[ʺ$%_Bc�&���4��t,`($pU#�C�D^F�[ew/�\��7g��Sf��	�ɵՎt[�r�P���	��58y���i4ޓJ��25��4��+�����W�ha>��y�r�{D� 4zdcSV�̇{	�S�̃�Rbh�)�y����F5���xj�\32���P���{��g�er8�������~��0&3[�V��l����g���򓥰oL�ד�O���` �����y��=JxϤ��32I�S�� h8Ƚ��a�}��AL���\�~�s4� ���vm4xƕͨ����֮���c�F[H�n�,�119 Yg��]���v�R��ܸL9$��z�r(�)���$6��g�ϭ{�����֦�-��(X1q%�-��}ܱ��3;<�gͣ��Z-[Vkvc+��4��q��g#�o�(f�����T����?����?������ŉ�U�|�����ӯ<���ڛ��|:킛����M�enj߉,�[�#p<ʔ����"8!<e"��&�66=����rP�A�C��0��0�����XNդ�F CxP;)�(��։���8 ��큉�@�bDPk{�RpS��$}�G�$<�18��y�TVx�IŃ�ۙ�Y^M����;�Ԫ�s+=�2c^b�qL��*=�iR�+r�pLa�Wi#C����۾nb���)� X�w'�ZSɤ ��
�Y$�܄#�End(�ЬN���O�-�Q�B����M��h��F�� Kì{Fp�زӅe�#�3��?��'(K'��ď�1:����g�$>��A��
�a	e������4�`X@EvG��|>SV'�Q8��|:�
$`���P3�ʑ9�j>Z.hJ�bϊ�5���:=�ć��\Q�!�&��Õ��J�����xBD��z�S�V�c���
n��#�.�?ۥ������.�c2tTb��&�����o���=ǧ?��/

����W��|��l����R?�������#�E�����M�N�36`��>�[��4T�*�_n"��䖠���CT·2&��g	t��}�?n�
dQ��yY�Z`^��SH��E�zr��v�+b����Q�zv%��r�0�^�M�ސ,߹�{�)�M}�o/K�/M;I뺹��~�*	*��	����0��*Ch3�⑲��#?��ߋ����E)K�A�2D`$�E�q?��	����9�ESW�M*R)�=6��|#���$o)
7&�5��l"��E��k7�]Y��,��Ta|��������K�L"�M�-I]�m��7��]��E�'s$z�L{�
I�h�,�g�M ΋��&CM@9�aE�_����-�ܰ�9"�x�B��:��Rÿ^��#en2��d4,�����L��4%��;/��[��x:��S��^V*I��,y5����ٰz�m͓;��@�-�h��reW˙=���gOg#�ZOm�y��V�d��
� _x���g~��|�S��R�*���������W�^�����DY:W:�t��6Cß7��m��ir���n���WHMYN�q;��\
!a����L}2��ঞI�����������5�T�:K�\������xRe)p3�M0���4�&*UC$9�{m�BQ�(c��~���(f��>Ѓ[� �i�l�BK.���UC<`2�c!��/��1�K'bg6���e�⇫�Ͱa["%�G !�}�64v��� �ei��S�[�Ȓn
,]N��mTv)�>֔7��^�7Я�À�H�m�d�SJB&��bX(
���l��ۺ7�md+&��KaS%�G�]&����;��rt;5#�
�p��bރ��2ޔ ,��T���w;_JVH~FVG��S�)O��5�{���J��mIc �P�0� ��늲�x�~[��SI�k�)�A�pv��2i-��������JJ�b�=��I�ri�RQ�4�[�^��ё�[��c�:W��Od��|6�g+(�2k)*ӗ<���\Cf�/�:�������-���?���G�ޯ�9���n�Trߡ��Z��o��s��T���dr�ҍM��۔q����$�T��x�!������O�F*�U#�$�K)�s�"�ȧi*Mէ�X�LAP��!k$��7\�nI_>�]*y�9F�*�H0p>Jl��I��5����_wR�H�k7,��,��$e:�R>�{Ġ 靥�F	��~�82��� �F I�V��A[�r���m4_��qܙ��1Ō�Ab�(���E�JYI�� �8�H�>��.�n^�*�	�6�r��	^��r�M粞]�܂���=�(N�#1��^�M? !#���P��ɻ��[�"��3<
���$,a�o������g�s����'h����\��	�����q���U2n��EP���t�@����|I�O@�</��ڰ׷^��&dn�dvx2@�*x'0Ը��Ppc��\ �s{�7�d�Z��p�sh���Vm���|=]��rf�2����n0��.l�Y��>�V��Pp{���ً��O��������Ëi�W���i�$���.��-����~��d#���E�F�%zE���x
B��+c��I�׳�T��hJ���>�,Nv%/��JM��T~
��7 $i��gQj
C}9���kK,4Up]즭~���0z��JT,�8S
V��{������2��}�� ��$LT��s6a6��C�U�[�T�z�l㛞��S�G��.W���n�l�v���34�.][��㣦�NHx7�^�X<�yL��<�����D"�@�wԳ��y^pt�� 4�߻\+�����%]_5�j��f2���M�{ܠb�`�8S9+!UI�ϝ[��5�������:��A;��{��`bZ�ս�>�����]扽 X�C�V�9)�9�A� ��^���+�1!B���K�Ddٸn�6��1Vv�z_G�ݖ/A.ABFӱ]����C98q[uk7�R!�$St��U�:ֹ���R��|i��=�m���8����j9��z�!��A�b��m��l���j�������*	��G_sY������'�����#OF��(�QpK
	�CYJ=��m�~�pQdr\Ь ��2�
:���ښ{����B�!M�H���*NW?eCH
���Tj� ����� R�Ie[Z�*-�L".�^�
�������~�{``�y<��4L�,�׬׸���=&�v���-25zx�tB��a%!D���	�nO���֮�*�1Ӧ�vm�S9�?�Xg�R�}�_g�æ��|ص�vc��̃[���ߢWSM���~�a�B@3�����PB�Hel�x*�^��d�B�J��Lsyk���;�����۔�|�������f݁�)K	�;�3�ZH$q�90�͞�{2�Z�{��i(� K�j��%a��͢��o����	'���1 \'��q��]�>��IՖ�C�*h	A�>���l��.���J�[m�z��Q��m6��{ջ�Nk�>�2�Z�ڈ#(AS�g�j�'�89�e6cד����v9�,���������d�V�u05�%;���A���W����o���-%�=�����COǽ��p�,�* ᝋ&�<AL����t���I=��փ[��i2�_~�[
h�i}Z��d75��n�zg�kx��㱪]#�2��6�oʦR�K�\|��2�·a��!)�iZ�T5d�yF�5t�����օ���	�*{/c��!��qz��j쥶^g�X
��{���+O��f}j��D�Ѳ:ÄMƮ��ۼ��އR�!:Wf־�N^y`�;
n��º˩M9gd�R�^kL	`�oJ}Np�5�K�䧑�"�r�ا�! D�t�_��y��x&�ۚ5e�p�ؘ)�Mz}[Ƕ��6����3M%��Wy�������:��;0v��NÜ���=Ā��$q �2ة�h �t5N(�F_U�И��R�gq���MS�f�a��*����/	v�2%�@���4�n���Y����[?�P�O��Ԇە�Xd���U�Vi5�ztl�F�F�݌�v3�Xo>��0���va��ږ��!J�J�sk4>�j��'~����EAA~畧��y<����7���
� A�W�R�IF�%���5Q&Ɖ��%��d��H2i�:\B*/��8%L�܉9N,�K����dS�nR�
�"��E�}7p�Ϣ,�d �-�P��`3 �+��s���+�������G�9{�/e\)�'K�JV<��*�e���҈甅�� "��;�}�M额v��o��g�?���94�[*y ���[u{����W^�gî]���[�T�
�/�M ���A[&&�׀�DpSi��};h`-�̞ W
^��J6�f���Fl�029�xpb�Pɸ�q���?c-�j8� �@���i%n$܀
Iՙ���w��4tJ�-	$4@�2�uJ��V�ϱs���������[j�x���&��9!�L#r�=��z�L�*>� Cb�t�]0$�>
�({��hZ� �r�9
�2-��P�m�R����B)�@��eq-+l���K&o���&�� ��m��H�����A��5kf���f?�r��c?�-��b���],��x���g�~�G�b�����E��[Men,<���wҼw����7��>��UHنP�܈��5G0�}����[E�ԫ�j�%
h�^�R�,������/9ky�J%�"
<
���hW>�Po�	2r8E�I�
�L��TS0ڕ�އ�r*���)�y�+�y�%���;������[���7ްg1��sx�)�l0����+��N-�DJ=��`JCY �bƬZ�w~���޻�aO7j_��6��������x�fn�Ep�7e�E5���6�26̰Ke�
�NBG��B�^5�+.{76��-�'��\
J�e9��4��RwA�rz�W��>`��'��%]E�)����^�G! *�	��W���.kۓ�O�i��A�U4�ZG/O�<����C�8Ӵ<��1��@M7���$�b��j��X�_��&[Ԥ  �V�\���
ʋ�Mfc�OFn.����R��f�"�u���l7-S-)����[�ٲ�vm��º��)y�Qi���ɱ�ZVYe,?��n��?�?�bd��s��M������^��F�6�IB?�b�l���m�u<T�D(��L=͗$P�{�H/� f�����'=��
H=*Np�jᵰ���V]�2=1I�$��$.=N��H�|����`,8�b3����1L^�M��Ty������{�l�[#CM���x���Lտ�y�pPye"�'/���M��˯��[�
@�t%���2���㛾A������|:����F���fD�������RM�[�Ӝ��}Dm�(�)�����r	rx���@�G
n���U��	n$4������uW��Փ1-�v�j+`�~��6���2���uS�T�����u� �ϝ��&g3t���o|�F��t�%�cQ6�1H
x�Jo�n�w��t�%P<�������:�L��VRx�
���G��,G�^�[�y���v�pk��E8ܔ*^�f�,[�Y��A�օ�]ͦv��ëR�����bbS���l�٪��ɩ���M>�R��џ��|12���O��b���Ǔ��=��sdnhrQ�y	��P������_n�
N�(�^��(m��)��B��WIF���?�Ʉ��Ʀ� #Y��)hi��4e'���̉�WC�O;&t+7�������	iiJ?��r&�Nl1�)�'l^*w�4MִyR�&6�A��,�^[�:z�hP��ƓPg�����*�,�N�@�ψ�GOlxy))ut�(3��	۫X������y徕Z��'v���w2�nm�����)�ݲn^:9)^m9׉s}0�j*{A�U��k੟9�{P(�X��G��l�H̡F/�=���#??=:RpcZz���M.���2	���t.��t�PYN�A �RP���^�hX!��H��g
X�.���!֩�����!�W!G'��[���q�	C�8�7���c	mϯ�'���7�2��jN�"�����}�̍���nWU��2�f�d%�0����u��W��T?2���Zm�u:�b��ZhŴ}�3���Rk>n�,͢4�\��+G�~���C�����k�����|��t��'��w?���fQJ���Ά�	�̋�
��tv<������x܅�<�qs勉�J(�J�(���֌O735g�i��#�����N��\V��)=�N]� ބs��>̇(G�4���ޔ��v�-��{z�{��
h{f2B;)�F����6̓�t�-��u�:F���ʦ�GP�4N��\kT% �V29�?�����+�zͥ{Tq*�[�����mTm�^؟�����k�2��,m�����
�n��B��� �!�����$t�j`k� �1��0�~L�)M��&In�݀����-@���{��g�#��Ս=���/�%)�:!�-�S]��~F�^��Ñ�сA�W�R%;�r��?HJ���#�r1�N�BE��iT&�jd5	иX�>�a�=��&�̮�ۋV�����/��$��d�!�~�%���x�ڣy24�����T�f�-/��YP�`����ʝ+�,�l����F��e��C�������*U,7_Y�P����?�/�����B
�������?����'�^��Ȱ��&3~���hօ��p7J�@n#G��{�FE5����J#�D�ִt��������H.g�$�)~귥SQ��]��L�x��H�(���$���,e]���T@��̌~�9��o���B4�JB�I�b�����X}�R@S�>a�$}[(m��t�o3֩7��PFӣT�m>�$ �����N_�ow��P��'7�v1�[�PpKe邀_D�l���J٢��/�*��-|+e���u�t����pu~)��K=*�5\-1��erOƕ�
'���	e�SE�
[>��{��*C��]�~zn�~���� ��kB�c�xC�.�ے	w�Qq�b�>�#c��k���g���4ݩ�DT���^����N#5?�<$�K=�[N��7�zB�Zv�*����)�K��$1.Ր��H�s��%��ALv��Nk��h(�"?_��"��Hнb��m�%�2@e` �&r�y7eF֪�/��F��yt���m�/m��ci���=7�X�ҭ\չ'��,���Z��D�暆m�-3ˤl@0d�h�$�)���_�P�,j��@n��ӱr�7�l<�9���ޡ��htw�[�}�s~�������dnn���6�
n%U#;N��kn7�c��n�:��4a�i�I�YeF�Rѯ�����Og��1���]���ݛ��؟sS��i�-��|����ćQ>Ǫ��� 7��~7�aXN��#��5��nJrn�z���� ��B��Z���������є=X½;�%�i�rfTB�[^+K�d4�l$.?i���,������TI�N<�`]h��B����nW��߷׃x<�,,��/��47�Es�G�]3`������A� ��4�q>�܄�9�l��J�F��.��ں/�6'3*d��T0";�f��z��~�0��<Up����1�s�'����4*�A�kXf�\{��w�e+���g"sr�t����@õm����S    IDATu����V����m�m����e���T�N7תpC�=!�2��Zo���;@5�����j#�n5J�� �1�Zi{�mX)Nb�bVghc&8Fբ`&��i�%��1Ml��-��o~��?��W�uZ�w�(�գF�[��?b�8�V��UARt2���HQ#���� Es�ce��T�����a��θ��Z���<	����љ�z�ne��Ȍ�43�k�������I^��6����9�@�fN�W�hvp�b��.ke�.���쳘7�g>C�, f���j���zMLxJ�JZ�g85���Ws8B&�Р��E1R^7{[d&�nդYI��	9]�9$8����+�I���s3���E.�����L����vg(��z�]���G��Ե���Ԕ&���A�g� ��
Z����z6�&xk��i�
l=�L<��t�xi���p��2���r53
����a����ʬ7�Z��px�P0f��c�o�7Nފ�E��0��i�8�G��p�q�Ѥs,el��O5}��'�5�zy� cpS/Ӫ�8��37�bq�=4��Ng*��H���2�)C��@�<31�\��L��H }�Ӏ9�C/�Rae���$��N4�Qoݔ�DD��1��-��������)K�����I������_;��(����nx��r�ǒQIR3�	E�udt��Nd�qb���B�s����LG�pm#u2s���M73P0��27��?8��vJ�R?n�/��it�<��1�uC��Qj�@�m�K�H�#n4-`��X�������}�U�}��1nO�S^I����y�⣸e91f�i���JT�!���"X�_���"V�E�>�8�	[Ĺ�<(��
pa޿s�������#琐�����!��Y���JHf�T�}�����c.ԣsRo�9�f����0�*�:�*2v�qpq�멒��aƐj�Ny��E��Y�yҒjG��nO�/�39B=d����j���j#�#l�g�V�ku�ԑ��u�b �
N�uuk\� ��֕m�;��R��nܣu����pT&Ƚ��q������8��֟1���ﱛ�OVNZ�V�NL:�.!�N�_�C;�N�#ax�a���+��C>c!�cAD���|�:)r܇H����xj����/�~��'_�|����d`����
���76N[��W�����W!ZR�"�,��h�V�	K��`D����6�S��5��tL�f.�y=�)�ص;*���ocf�9�\p��vp�Y~i
g�����8��ր����;�6�T��I7jbq��3a"H96�t���eb��v�W�ݬ�8'Γ��J�1y�5��4M�� !S�hW,������7n����������#<�|�ݣ�h�W�7�b5����G��_� ������ZkkkX[[��Ң|+y�1��
���q���{x���`G�Nꖦ�:����Y-~^�(HVq�H�R���������ݦ��b��&��NmVYvG�g�"|�֧��{H�xI��$�떂�֑J�M�Z���)�*�YN o����Q�����LVu���\TAXe� �]�v�I58J�Ś��������u�;�3)��_�e��DB��b���rf��t�v@b~��z�{n��x�Ԍ�I�J�����6��D0�ԋ#F1I�>]0�^)9�7?��
��|<ux{>�������Y����ܨ
r9l��;�˟>�\�ʜ�t�w�~�=�x2� ���x'0���<Ỷa��Lps���ƛ��fu�;���(�ܿ��މ����dCU�-	��o��Z��0!��\�����++͂�\AG��=,7%����SX��D�fhܮ���4�k��Y�!FE�<>�^���ept�2]1,,o�#�����)�b}qo߽�w�z���x��9��|�
I�T1��f6��O���2=�R��ǏQ<����{ｇ����x�ݞ�I��B-~�/�0z���Ϸ_`�`_�^���;X��G&�4�4�?%U�>\H�����x�_<�a���g���:� <"K��h��B�5"��z�J��l�A_|Kfx� H�cp�|��X�8��D��ϑ~7ܴ�&��F��7�gs�����.��+
�D����}��X.���3њ�u"s�#lt�j�3��n�3�-�M]��  ��c� �>s����G��Ǩ.�#��epQXa$TE*�4��^������� �������_�5��|���
~���_>���E��;;�˟�/_F����o��l�n�-K��$�܈OkS�M�܌|x���N������J?ʞ�����{��b�����p<�p@Z��+�6�p<��)�p@��P3��/nqO0+�I�bv��	����Y�B���B�u(�j��&(aԩJ��a������}���xR�����8�)�Ǐ�`#n-��ޭ;x��q|z�gۛx��)l�[�={c���_�q,��y��dST��/��|�3���;�S�(��M#�8��f�AK�"������M�pgm�x
�~O���ZU��G�p�S9#g���o���Ml_��U����mb�M�9����N�ҩ6�`�VwL����E�R�0�P*���3�9�ǤP�[:h�����!
6j\�\�7�P�����!��E{x�{y�[�;tݞp��5c��mš6�N.C�ai�������1���M�h�5$��K�p�h�X�x����a<PU��<�W��hL��oBw$��d`��߯ඐJܚ[����Ƃ�e���+W��[�'0��q�@�K2����8�u9����L�z���R�����5ї�p��)8ܜ��d �|�I��}����zeN`���ǲ�*����	B�9&�O�|,9���.��6v
.����{������dO���F=�Qʴ����dx��3S��qoeC����}'g*K?|�
.�A_pn�?��쬂���eB���߿���e���c��j��$m���cX�XW3�(��/�X7W���g���>�W�jT%��EE��������#�ℾ��K��X.L��8��F`ꖙXSR�-ܜ�%���rU�p���s�-���\�䂝*@w�'@'\)�Ke��*]9)�)u]W���i�:�I��+�'׹�Z�0��L?�|����a�j�H����j�wz�U�Z�3�DB��	*�I����<���n�}z���y�~PIJN��x�H��ȧ�{w�W~�s���җ�����dp�wY�/{�Y������ՊQfn�J��&���z��2	Er����6����d�7#k��=%ո1>Z�3� >�˵o���JVW�1����LНTZ�Nr��K;��`��q�zǎFi�D�5&�4�@�^�Q��7*n�����!̯7�48����pM��ND�WV��e��:L���1D�}����<L��d�#�<D�v7�����?��;�e�ɋgx��ʭ���Bͯ\"�Ͼ���!Ev�n
=���C~q�^GW���Gb��D��$�-@�w~~���4�J�8���n��k�����|��JU�?�ហc��̴6�����x���sM�4���@�3$l�sY�]�ڑ֌c��?�vk�<C@D��"�t=�QN}&������̙m��(Z�e�Xf�d�!��0�#l�Sp�0�q�c2s3��P�Ȋ{c̠�Ƹ)Ks�U�^&HP��"�5CA�� ���h������"�1�1s�&"
l�0͂�s��54��ό� ahR��&�45�����[�����7"V��<����v���+�?w\/��s�[ĸ��e)�8375�%Zi
�,epsP��{g�e�Q�M(��Mq�9��uٞ+��z�=���O�j*Wl�T�`�\L����YR1����S�Yj
]㒤	Ԅ�_�-L�פ�Ƅ��Ny�����{t}�!{��F��@��@��)-�S:�X�H��a��$���t�������{�n�F�\��-<|������2)ٯM'����|w����;O6EUʤ2��R��x��<�{�3�MM��#�Z���Q�N��W�9�YY�[�uty��}��Q��|�сc_L� :3�}�]^]��N�?k�֏�Zݚ�Y%NK�l��M��^��?�5�nX��8�˪M�z�NHV2���Zq��n蠃O��3 ��>\W�Z���� ���a��C֖�nR�CB�њ�[����5��6	$v|m~�Nr� jl|�԰�{�k���j��g�F�n8�Q�`� |Q���(�N~)��o��m$���L�R��I�L�<�9��w����ʷ?%Q��O}ߙ�����g����S��/��x��6�}��e�#3-MF��2s�Ӽh�~���Czl4����O�1���� ��>����ZX�g'�rڴ�e]���(��tSI-..���t6��IMv}>=*S(��_%�I��b �	븟*-��ev�_� �G��I����Mt�Z��	UWȩ�O{,n�����:ˀ�ЋHX�����zoݾ/������}��/���p�/~�sX�]B|��������8Vnn�6���1���w�[�T�bC�(��&)�;=��ǝ�e��~wo���;���7>����#�	?ⴇ84��aƾ���`=Nݺ���el�JC�;)�0��6087+H�������E���PMb]#�>�3���m�L?�\�;�Q��2�٫>��3���긥"$���yMŠ�N3#�L���pu�[n� �@�Vq�-{r߫�V����|�:�|񈙐��R�Q���3ȱ
�СO���	?�+>�I� ��1��������_����?�����N��V/��Q��,%މ=-e7C�C�s#z��.����cIS�p��q��eT�ҁ`πs|��0�ܒa6hjey4��0���k��+'�=A�湮�n�[<����i�;�ܩ�Ǝo�j��,l�.�~��N��&&���A�n��b�*(
�F�c�Ĺr�~��?a��<˭>Dh��)����w��ݷ5���%���!*��zf��yF�Ke����n�-#?ζ�,���omH���������~�,Q�a����Az<v�Hz|�5��;�k��qC��R·�>R`<��P��u7談�Jr����ٍ���!'+B���8\pp[��_��8�1�1�&�sS��k �n�mH�G]4�/\�Ck��cu����f�)��*��ǵh�����Dn�3[B�C���FL6iA�6�������>��jv]����g[B��ʘ�@J�y�(d��(Ti��%X�5Ì-H/}���cCp��xM1L�z�#����?��T����7�o|�F�3��F���
��i���	�fn��)h�[4Z�72��$H�G&�qK�gA��_��iw��X,݄^1^�*�O/J��;Ь߀'Ǵ�	�N>"�]&����0=6'�uN�������zꝍ{w��'7'5d� �|��k�o{z�KlW�ڛ��WNm��;9(�W{B;�~9n$�z"�j/ ����@o��W��ͻx��=e���{���C\U+z�N� �7|�s?�;�� ��n��J073�b���ǻ��'��@�?��nN��@��Al�E����n-���;�tOO�W��㏰[��9}-��e�ݽ���}Yǻ��t�_N�N"�}��Ϝx��������/co룠[{?��a����S�0���={���������Wz�t-�k�P�l��w���;�,�ϭ;D�D�'���d�$ߏ�^(�.�
��&-6�9H�+���p��q�3�G�xI���U���ƞ���"NI)�"O"O@т�Ef���^7J�����������}�������?��oF����e�z�_���17)��N5.Fϻ�m2��M�Ր5�Dp�<�\��iN��ȕe)Og�+�?)/�J��ӑ׉h�)���nd.�R鯙r��Mu����9-;W�^8����ZD���M��M9|M�r�	P�bǋq2X
�b6���i��f63��m'xƳ���f�݁����Kx��=�w�-����5�4�& 75�Յ%����iqA�_�
�C'����Z��է���E'�R%$K�>�@�> :!�	`cfN���zWW|rq��~�-��QAM9k��F���\����tDs�?bݐiVc�ܺbc�G�+Q����n�,�(ee��I�e�u-Mam6g��Tu=S�'U~�qA9�@����3��{ߥȤ���p7��q�T����w%��UI��E4���K��\�z�r@F_p���'��F�V�26VK��sC.v��[�hP � �(�W��CU>3��H33s���a���P)��j(���ͦ���P�@�1�n�W����?�fzn���/�j���W+��n칑8Ͻ�2$7-�g�J�Eo�S�&)h�(Hȿ�3��-}}cN=wB�Ū�5�D�*@����-���;�{�������^�u"'p2Ⱦ�3���il낙�&���g{fщ����TA��&����X�3nnwO�\	��(�X3�����GA&�nN��7L�F����9?{���s�'c1�^����Ul��!��[o�x{_ާ�H��s8.�xo��c��E���xk��Ã�:o��@g��lwV7�#ｏ�׏��s|����A�M��1��6�0�Q�ϡ2,qp�$�"�<�0�O��cX��F�x���>'s$���)�v9\��t�MY����$C�*9���4�7NE�I������,kf����(�U�qkV�P�Sv�����=c��p�M0��$�F�@�a�f�d��>F4Ͷ�ٔ��Ma������5��-C4���i�J����� ��h$�����ssy���#9;�B����S\������{nӱ8fB1���On�-��nG���:bp�4b���X]����~�lJ�+�N`��Gi����B��I��r��mrń	�x�e����fr3�a+�ZP�d�t]��z{�AcYb����<���r�ؼ���(�s�����^�k&[m57g�<A���k�5�)w��O-�;$oc�����1�q��c�
���`7<�|�ffpoq�Wo �)�<99���)
�W2 �X]��ħs
�J[O^h���`~q�Z[G���qٮ��1{.�����;��~���I�Z^�۷�J���p��~�8�:G�7�K�x(�I�����'�KaܸI5�&��cZ&�Ym8����v0�p������$O5�	iy��60볒G�I��~�>2ofp���`Ь1r�L��&��,��|�`0��J�O�F��+�0�k���4W<7F��df(�bK����������!��BQj�L�K�U�A��DA˨��\�d�ك%v��Š�xT��*�J!'�����4��s�B��Vq|q�B�
д�o�+D'�z}��&��F"�7f�~�����f���ou�[���V��&sk3h8bf_x��2����j�I1�1	we��V��
�.۲�W�W67w�|��pCgv��;W�!�+=u�-��5v��F�M~m���I�c���^��iw�6��x���WH�&�2�M:I`�(M�&"��2�f���7r�g2>�@T���{���븯�:��!8Ԓ�	<�G������i������:n�.	)>�uP8�@�P� �K#5=�z����c�)s#u���t�}�����+E�;M�������7ـϏ�����lV��T4���=�/��qY���ƐŰ���X.o2��{ؿ:;���A��iA�su=-��fC�� �0�i�kYe��l�'�G��2v<�t��v��>�%����L:��כ
�Z[�X��7�
�Lp4��y�T�&�D�q<��~IIџD��jU�a�FPu$�^�fx����B�P�4������A
���N6�v�:�鷒�����	�(��2Li/�����}�)�cQ$�2
n�a�|>1�4\�EQ�Pl�Q�Ք�y���5i}	��F�>Y�������_�� ���C    IDAT3���k�}ܬ��a���<h�M^�q�����L�4�9�R:x"�D�77�O&-�QnE��Z��Q���c]��Ԕ@�\6�-vG:Z��G�s  �^'2�n{\��)�z�񹀬A����`�=&���A� V*���� _��:��o|����O��׽C3�5����Y��*Q5淧����I�A���V0{�����|XHM���*�-�b}*��/$��V�(���\U '@ؿ�8)������+��yun�oݑ����gg*Cj��2�H(�T6��D>���w��j�$Ú����4�M����˃]�.�
�#qu�����xxt��'���>9�jt��!
Z`��n��*��&���Y�ç�2t� y�m�4I��+�d-�@RJVR���aP�:O��@�Z3��}��A��I��} ط"^���v�/�v��C��Х��5{k�i�-U?���#iOg6͝w)3~C{4��0�(�XLXS��&�v���<
v�m!�M�Y�@eXNWa0+eB�
����Wl��s�lZ����
�^K�{����@b��� �pȠ+x�x<R��Ɠ𴚈�<H�}O6rs���A�o���{����I�����V-VBb�.���xB�'�	c�F��G�^.s���ƾ�QV}%�	"d�a�`e�,m����]{z��E��˻�45�дb�R�$1Ϳ�.��^W����'�g��8�n=x���5�:F�S},�aޏ	B��.ss�����=Yc_.(@��E�J�r,�h� ���{]� m�u�j�"v��@`��̣7@��G�F>����<n�,cij�@X�pNL�^��:v��u�����ܴ$��,� �g�h�u�{�Ⱦ�w$EkЕ�Ь��>��~��YI*�L}Q��E��5%�X���QA�<�C��ώ��2����{�b�0#a�Mz�e(H��i��sV�k2�1X(����LY�͹�q�YZ�����VHb"u���t=���A�f<|}^'36�@$S)��9��t�����ۢ�5秒�`��tW�����V�4m	�>2׍���S�x&� �l�Qi6����۩���v`B��I�v�G�P�Ϩ~�5j���xM�$�6V��Fi�c���~?*�=j/K`<�I:~�W)#��#<�3��K�?>���<��}c�S��G��Ϟ���p�(��B�nD�3��$\��
e_�,��%Vi<�����[��5�dMnx:ܸ�Ͷ��Q�7�S�|Be��d�#k��}��LL�'��5P�	21z�`�����P�9�O^�	`��.G�c����*�p�Df6���D�q-'�ᦹcr���n�eO�qiQ��~��T����	��1Ka=����e,M�"�K �e���1��p\:G�Q�k:���S�|fV�hʌ+� `�����q^����)��x�M��oci����M+8R]���'f7�h�͢T@�mb��@��LJ�}L(��}�����<̴8�� x���s6s\Tez�K̒�b�Ɣ)��1�0p���5`��o�PTY��I�o�|�x@�rYL�rʠZ�"���,��=-��8����w�g��h ���0y��@*&ʐ���~��$ܧSD�It=�j5�DqX�5�QN��+����b�I93��=e���^�.Հ^̮-#���N�+�=�l�����k���j�A��?�� ��D��]^�ۍ���o���O���9nU~�Y���r���D�O�M�H
���(3�Lc�a���讧|�%�&�� ���ds��WP��&�6~Iz0�2���=��0H�|���izn��cl�-�^n�S��^~�ei
�f�`�f� 	�k��8+t��l��ۡk���W%�a!/NY�&�\Vfb{���Y�z��\f(����X��{#�KH����X+�y���S�yG�::��y���װ����`��46��6�����bi���(1l Z�uZ�=>T��r$N/3���y�^]W�cp�]���0�tL"�~�h�v�}v��fU�4��pj�gJL�k+���H�?35�H`�ӤT"�VA���;}5�ō��V��IƳlで��(k�P-��G��
��K��m�'�5(�MT>�������B^���h��F���y�� 1�9�AUr��F��	��V�I�� |>�Mz�R���X񩴔��
�J��LV�@�e��ϒ�!�J(���J��K����Џ3�e��� ���ߺ�A<����YG#@�=F�#����փl��A���?D��'��V�7~짾�i�����W4e>�V��q��S��Z�:����fn,K��'
��2���[��prv00�`1C��u�*p�D��2��@X��)_��Υ�B�����>N���	�e|��Th�NK_�a:��0������a�(���+G�Ӗ	�n��3�V.�)Of��9i%~#�6�9+86��taqV��&��q�jy�*���������Y8`x�93R�Ng�W���q�
�g'��z�q�ډE�7�L<����SY�'s���$w�����E��m�~\���m�Z��Pm���:6�KRP�4Z��F��?
�����Lj:�x��������>hcD�&��R���R�WC�H��T�r>��-:��V�q]�P3�` � �V[4ŋK��>D�Ĵ{�6!�^�/-bvauz|Vk�wZ
h,I;���=Y��<�x�)64��02D��+Z�>��Y~)9���p��)�8a.T�(7�h���Þ���tp+�Ʉ�������R�A��K��}�u�W���XC?D���UG��\��l;��>JN�)9E��H�8��w�V��o|�o|�����76�;�t�*�M���+9翬�F�?sp���ۈ�h�U������K�I�K=W.NH���Aӓ��±n��*s�b�H����Š��=x˱�i�p:pn2'a�rL��D+-r\�'�3������i��	"��ǌ�I�Og3=M�$XіX6�Pvh�o��\p��kN����G�?��4
���(+���S��5NT� ��K�!fN<��a꣎>G��6oo(Hɔ?�\ ��hFx�T$&:A�R�N�FU~
ln�o(|�Ǉ��9,�,�Ԍ��d@�}��E���RW�
��"I;ԠK�5�IN�{���_�-)s�ka�C��EU2����s�be�l��J�C����̏��Zs�:(]�scP7 b��L�Tk��>�Von 3=#ɦ�rI=���;�:0T9�#�zG���Ϙ�){a!b�:}�Z]�9��A�á�Y��( :��G<�A�U�e��,�i!4<T��)k� ��T��-�`ʁI�QW ���Q�vK�Vև6DC�Z_Blao�n�~J�E�F����2�öu�t�u�<^�ƒ�'��]Z�������o�C���a��;'���7�!܈��jZj�R�]ύ��&A�?%A�R 5����6��i�+KUJ���8�B�{X�N'���oM�ݤ�/����<88�Y�/r�J>ı��U9e*��d�b'�����U�5�j�#�����L�L60	j���H\���D��L����ף���K*��S�P��h�hP�I5{"t#��s��4��t��<��P� ՙ��|D�K

Z`�|�f�z��R���z�"8A��G��o�M�@�;D��7��`��@��f��/`�)*J�!!�e0��3��̬�Uo������EG�����̨
͍䋅%�Ĭ�O̕���zo<HXQ��̭�U�ff�
E�Kbv�~+�;M\'3zM ۝18؁z���C�%i0�����>Z�:zVb���N�������C���p��]$�S�FϊW�4��Y��Mã �\+��3� �üʊ��"<����ǵ"ж�аX��ZM,��`qm�T��8��Є�I
�1�q�� �u���I�"���+e��Ѹ�(����:���S��ـ/��Q���zU���(�	�۸��l4�iQ�r�Q�����8qn�����K��O��������W�ڍ�9�~�U����&dc� �><�!�Ѱ� !�v�����f�Lp3���y&?�����5ev�E6]'���]�Po�N
���A��U���J�Iܗ뵩e'C�\�~�����J=*f��p�%����73^+���^	��Zed꙰�jpM�T:MbߔLy�CN#� b}���2�
��bO����sc��n�^��r^�R��_�v�'���2��ZW�a���U�ZS�D���0V~}*?�Bh��RXDC:h�1��d�d|a�=��tkm]�7b��վ`�k���R�h���){Un�����d�����ƴ&�S��Fft���&`���ҟ���� 3�vW��dV��� ��0�/>SN7[�A��J�9
W�D����#N��IJ[!:'o�ה�/���kwqvx��I����/bznV��F��b��R�X��M���g��053�Z��Ó#�]�K�D#
�<X�!���hf60+���A��}na���F8S\n6Qn�������;92��O)�`$�h��r��z` g��k4�3����LJא]Y@�lNqV����`!D�y/[&��Z��ø�n!��[>�x�����n�MMK��?_=i���^��3g�z�:���Li:5�H�"�hZ��7�(�3>c@��Q�����k7'�勨gd!#*�/�Y�P�v��pN��������L���j����U�	�4�<�qg5�xmA>~/��!���2���yiKE� `��Bׁ�c���'@�m��yu"���{�aL����h�Hf5-�'�
n,f	.�1K`i:9q�5��a��f�YIQm��q�D�{��C�%����W�,�LH`�h�FHIw�xߧnTkaPmb��Y�pP<d6�U.���P�F�/2`�U��t	a���PD�TB�A�ߑP���0��oev�6��+SE837ra	?h��֚*�U���uד�de~����Q�XN������|�c@�^Ҕ�_��1أ"d���vWA[��� �W�����K%�)A�Q���N��$
�`��v��y�El�l	[�v��y�8(��6@���Ť�)R4��/�aiy�pDX�v���n�J��$i��Y��D��y��F�H�:~��M�����-1=�A�U���Z�^[����
�����v�fM���
*L���'_����_짿�Fpn����6/���Z��:�Pmx�����7���@�,5���z�T��(I��%K0v��J

F�I�=
6|������bIe%�i^A�}7[ۻߩ��"��ԝ��f��~�F�ሰV�f5<�I�G�o�!OpL�=�ٟ�)�t<�B��R�d�=��ya:!���d�N	�d_I�`N+�#Ľ�;t�5m��A,D�Ȅcڄ�v[�D�\��%�E�9&f��Rce��P'݅j��'����_qe*���8�d:A���F\��^-��>�g��ƕ��"A�� ���*u�
5��@��>�Ʉ�/3���2�10g�i@(�w���L��I��;�����e)�f8�6yI�Jf�H�R���O���Pe���E���ʥm�{��i��\{��gX,<0�BR�����V/���N���҉�🎷I,b~v�xR���4�9��-�!��Vp�=:ĳ��qrr����w>�{���R����prvf�`�Rq&��RvF���U�BQ;/�H"��!cf6�p4j�����Z$���wt���S��_��k�+��G�{҃t:�u���^#�-�fM?�Q�}>\v�8kTQv� ���^�W����{��QoՕ����x����^�����ҟ�����7�j��W+��g�F�7C�7����37����c3k���&	c<A�,���R��K{��q�:�2]��'�%qR��=�O&EK$v�n|]7�f����;����d�L�}���B���f0B6�d��r���bъt%�̓KR/v�TK�cc9J��7��/ ��eճK��Ć>�gg�������8�1�`[��G�V��	�S=q/�'��$����}$��ɅH-NzF���2@.�����L%�-���*k�V�]�.T�Z���a�8<8x 4��|�|V��s%��fy���tg߈�-ɾ��/FJ���FA� !Dɧ�i������Jin��Y��V*�f�pB߻��֒�#t�/~�����P���iTV0�gnl8�e�זW�x�T^ǳi,n�"H�m6�j�����8�;T%q�������k%���'�Q,����'1��­�5Ap�g8;>�����f��v:-���J�r�MO.��C4"����	����,���}���i#�8�r"���jn�]U;>?*��k��m1H�k�:�	��?Kx�p���"�E�fܦ"q,�[�.l��\|�O�Hp���uk�U�'{��O�w��On,K�\P�����KQ�ޘ��� ��˙�L�_�u��,m��}�zYc �E��48�	1.�4�fe�d�%9c�W��I�x�,Y/�`oKg$֢�8'f]1�PX���cl54]�|h�me��K����<Hx���$0�F�Ї�;(��[������l*c�cv`P-WT���[]^A�RA��J��e�0hz���R<~Y�����,�777ǁ���$	�͎2��D�w0���g�XE3q5�#��f�3�R��Z����R��f
;e>7�t!��jקdp`a�\������	�q� ��c�/�)�a��fIJ��
yM<9�`�Ȁ&�N�FK�s�2Y��l�R.��f�Y-��,��
a�a��sv٤�v7�b�zt�~�o666��BQ�X*)!���4�#O�������H;���Օ%H�51���a�:0�sy�^^Í�e�����C�_Z�R��Npxx�B�d�뤊��"��fg��qtq���:z��|�3���D�N��1�)��=�A�խA_�m�(�@�?��Z�3�\�շ$sH�h�^`$��Xb����/ߝ���7�~��|��I��O���������E�ABD�W37�o���h졠E'�RfOײޮ\ �rK5��p
'}<9���Z�.q85�5n�� }+nl���!#nk�f�t�X��DvʨbaX���b�6���5H����'�����et0Ppc�D�Q�^�,��2y��Lx���$��૶�����_h�8Oc&��;y��~� .N�T�R�a>���,�A���I� ��A��M������)���=B�X��Xi"�9Qe	�Ǵ��"a�A-k�'3)��?�� R��]�������.RA�0Γ�'�ZV�ө��=�9D�D��2�T���xR�t�x�%��D�#�ӄ!Х��<!ӫcvʉ"/�X�. Ą���2:��BH&
�̪*����Ѱ%�����Ѐ��1��@���}S�n��*��°�ѠL���d��i#�������
dL���{�垠1wn����wx�s2,���6��t�7��qsqE��U�GG���	jR<���O����Z�� Cy)f����	�g�ܶpp~�J�n�0 �0��Td#g�I�g���Lb�#���a#�A���(t�����[m�����m!���`q�oN���7�~�����߫��A��Kg�&j$�����5-�,K�0]p�_��f(@���.��B��B����enn����� x�@������{D,	5�4��q��2c���z�
^���	��FΓRN�d��g�H-4ꍯk�Lɟcpk��-Q���Y� >�^gf���x�/��)ֱ��Mc#r�$B�l��=���
ES����707�k�3�)������Q}��m�.-#��ŋ�e0i7Zf�Kd;3%�l����nJ-ҀWA2�M���\f�h7�c_:6��T�p���bp\�tBA��p���2�5_W�'~ U�����1f�����tA��5Qf�&������RY*a)l�YI��j۩��>,7Y)DX��U:��4鶞�ϫg@� ��,��e1.xk�
 �I �ˍe���L6+��栋J�#8�?]\    IDAT�uv�=�..�΍���#��n&r����'�:?�j~��n���MԊeGVO�KHOO��|w{{;q/��@<���*nݺ��TN�Z���+�Ѽ�j1� �����]��	h���BaN�M����1��-π�eND�*|�_��a�-��t����_�l>�'?y�'������f(��G_��[���Z���:�
2	Ѵ���!��\�,=�s�tmH�.Q���ˆ��4:k�>�zhV�����j|\�m:*�S���?�(�1kb���.�f�٩��������/b�T=3�����G�����0�d����&(N����G�㗱1_���S��L.���]�51����&p�~����{��j��#� 6�#����l����w�A�ZF�X�I(.��'��i9Ƞ������%������X����!./��
���Japc|�dH^������Trl�"�NW����������:
�XN���r%D���jt��P�x�*��;�5P��'ׇ�T�=Q�S���S��3� �k�Bg�~O��v#�h����*W������}���g*i*�y/n��zuNA(�t0sҘa��v&�d�G /A���[����Ю�%����ܨ�"�:�!D^�x�g/_`��Kd�)ܻuW�[-��wx �"����l��ᶆ"U�n��ծӿ��]Le�qzu���[����RSܠ���o+�6���0ݬ�(
jKSfol]�j��)`��x���IP�fߕk�U���Q�����7~����~#��w?��=��~�Y���VU�.�Zk4��[���5�B�ېY�27�����h�A�4�x�иx�&������a��^U0���LZr����)�pL�M�$r.�'����4��3"��Cm�������Y�))��d�Y}-�
���wTF���$I:����m������[}������)W�v��T�eq$�\��9��T^����+�p�r��d�>�G>D�4U1�9-��e42��'��he��+%a��Y8QA���q�rC��E�n��L	�P�,�}��`E���1Cb�Y��%��L��Ϧ�2`b�L�,tz�d����)�k[=82&B:d���癹0��a�|F�����w��ra�F���:z6��Ig]�O�X�4�031"�	˰*4V�03r^ܸ^3@�`���{�@˴.�5r\{}ӷ0����<\f��ԻF��LO!�N*�eB�a�;�o���[zН��k#�L
��R������,/�w�A�P��с��ydg��d���ob�`� 3�A�]�f��t�J/v��h�J��_�e�T��(�`�e3��5dd̹��U�h�~AtH�d2������f�{dY�![8�fp��XI���ϯ��ʭ�?�o־���gn��џ��A��������^��ϫ�-�x<"�!}K��&ʒ1R�F��\���4�(l�au�"����E�cw�i��e��/���s�X�D�DF��ܰ'BH�m֫���h���/�ꝳc\6�c�_%S�!�b1�CQ��꠵nU�$y�*ݫ��E��$�0��F&y�3���i�MZM�\��	U��*��з�L���������bs��SD�]��>d=A��^�Dc�G�0���2�ഋ����墲n&�f��'�8?Q�Li�R]�2r#Ca�':�W�UA6rӳ
����Nt~psI�KɎA�+���F;�Q������E�O�"�l��V��%!�<I�CR�l0D��l�N��o <�,y-��`[N��C�f� ��(��2vV��,ǉY8{���d]k22��))>JP�(k�i����9�1 XZ"j��WwtbQ���"�I����4��p��
y��[/^j��ֽ������s4�U��y5�yؼ|�\A�Y�;wpuYTpc�9��n��{xy�-X��#�=ݽq�������p�϶7�`�.�9Z�����p�B!M#P���z�^�1/a�B�����a���%�!&�@H�2�}�=�;I�bp[Me���/��{w��՗�>o��?Ȳ��}�?8jU��A���I��7���9�?`6Q�3�*��n2��BU��u�[R;$i� �ĵ�<Vg������[�{�j�vcʘ��Y�/,am:�$��������g��en�wl�2-.��8,_J�����NS��,f���ĕ�q�P(���T�e��r�t���,6V�8���3{�̍���P���e����#���A��B�7B7���A�$�~]��@���U�;�(��:��),�s���t�V�kq�czfƸE���SR���4��h��p��p�M���OrN�պ�)3�S��}x|�����ɥ){��-AJم���Od�[e��t���T6� �L�V�j�Dc1�P��3KJ�38*�S����K��Z��9�ｴ�8�����Gz�̇x-~�YjuX�SX,Uǔ�7��G�p4n%�M��J�b~�S`�����3���r�ԣ��[(�I.K�t:#��x:�x:�tn
Ssfj�������������T|gg�'�t3kO%����}��E���cgO�yy��O�_����Er��|xw6n�ޝ;X�/���O67�p�9*�����,Mc��p���ZC���}g�36����o��:�|����,�^�ʐ���!I��`+���[󫿱����?���G#o��o���v�4�o1��H�����A�1e�GT���(Q9����9�̴����T��1�t8.���Y�Es�Z�(W��U^����6�Z4=,�,cei��<�l��\����յ�0vb��9)�5KFh�hW��.%}Vf�qgy	OXM�z�1r*E���JQ��p���U�Z���DoH�[7N��qj���G���|OvwT7<��}��'H7K�� �.TP><Ai���2RC?ֲ�X�ɣ[k�Z,�m=��2��Nÿ9L`�"�RK4����/��h��!�?2��F�`�Z=ee-j����"H�jt�8�8S_�A�7ș�ƽ�X*'�Ò��6Í4���:Ii��l���1K�7��6��Ph��`����:���+7��.�9G�#6+���X�� R�9�yܓdi�>�������3�k�Ϥ"�@	�Gf������ngw�����W^S�K�p#�+	��$AL�L+��#QcP�W������2�S����������n�n��=��g�����uMI�����v������f����e���}��G�O�|kSW}OЇ֣����oɥ�8�Gϟk��F��X�G���z'��>�2b�x���9�`� ���>��eMP�=b �PL��j�V�n�@��V�S[��-�Z&��o�8��|�+��3��:l����f�6�[� O��#�G�fl���@����n.�9��w$�I�->0*�X�Ss�9���X	_��)������Ԭ��ܽ8�q�R&��b	��u.���T�`�~W��J�.�)�e�%S�8Qd��Q���閥�!e�j]��u8���q�Gg'r[b3xmi��n!Ok��F?a,�|A�l��@rzH<>f�����W8�A�
�aK^�0�Uou0h�Ы6�*��<�BXXN尔�	�OC2��Uh��?��a��4L 05F6��T6��}4ZM�_�Y4��p嫒���N_�'77��TV=�b��G
j�n6���߲�� b��X���mw%'j��\���W������,6n�aeuUϋ�\�^����Qk�li��1�87�7ql�F˔�v�"�˨0[%F�V�4��[:N�:V�ˍF%���JP/%ٌ��h<n��DH]�(�&\�X���+�Zt�Ji.)���]�*��P�n,�%	��/��`���N���X1���[
p�jC�ܣGt}�9h�wO��4F���CGJ�K��/b��?�g��um�Ff���w���ￏ��<O����<��B�;D�<r����k训�g��e��R�a��bY�zx�Y��� J%'h�3�ZE-
��p�F8�r*��~n�W>�c�~��kj�_R�~_��?���/�|Ԯ��a��~ܨ�J��tB��ƍ�q*�׸��ۮ{n��$ �uz(C��У(}{f7f�o����������Pel����ÀW��a����1	NѬf4o��ڈ��^\v�����<��ae~��y���Y��3Ǟ%a�je����\d���*޹s�pZ��˳s���{���� ,`s
�y"�P�5�u|��<y��l"�+��>��A�͎�*��
��%�����G�D�\R�ׯ�T�R��6��`$j�N�l;n����1����:�G�%9O]N�Zm�V�h+@0���_XY���N���K|��_���!�..M�F�l ��̆���ш-�������,O�Y�|�V�� r�)т�gsȲA�l��r�d��|�Ͷz���)�����
,�����5^�����~�~��T�S�5h�B���cpY<���,��Leǥ=��H$��C��`5�%�ym#)�*c�s׽�*�e��`�L�	���*�Vn���{�[Z�����x��}�.n޼�v���O���ÏT���r��m,/-
��u����L�RrD�K���������|�g[/��ʨ�<��m���{��̊~���3<|��nN��#�O%��$��t���*�� ��U���?��\4}O�j�X���j�,@�o8gn���˷g��G>���xp���oF��ÿuܮ�O��ʲn]&���A(�ϣ��3�$>�4�%�h
.�����Eէ!�Ӂ0nM/��5,Ħ��N��+;%�(U�&�P�CU/��t/O4�Z��Cgp|k�&��zh�FU����#��%��TLX��ǭ�%�L�a:�@MK'g�U�f����^D��i�g'(7*����훷�'P�V������mԚ5t�u6�#73�U;b���h:8/��k}_� �~��$B�?[�1I��*蝗���E�ᶊ]/�
$V*�����3�,��L3~�A�}"҆�a "��5�t�bE ����y�I����C`���c��&NO�����i��F��x�l�������bN!�M3� iN~dRi7�g�D�3@��)ezD�
�zidKK5\��&�)@��$����sxD;d`�r�U�aW\a���?<�s���(�A�ו�eMp����fP��'�L-;ԨU�KEN�k(�*:|ܴ���σ�33?����P��cR�jY�Xtcko[;;�f7n���Ҳ��'O����b[�0[]Y�ﾧ
D��
WEj*��T~��p�Ock[�:��81���o����*ҹi�����K<�z�b��QdП�h	7*gK*��#�^��/nZ�`�?�Z�z7���>�̠���Aª��� ���{3�_�b?��?p��>y?��S�{��r���e)��x�3@Nfn(0{}�nD�k����n 9�0��.0��3�7q?���7o�/����CI��(#����TN�x.�j����>�~�`��vDg!�<��ݛw���DQhV��s��;2�e���3'��VpoyK�",G���.qzp$n����Y��%:�^�Y�
�����rab$�������e�4?;���2�ݺ��?&������#|{�)J���I�A[�����x���"�CfBqD^�k-1 �8��8��t�(g���s���(-8�Ō%{<�7D�M��)gݳ̎��~���N!��Q��?�����ى~6����C�[ q��e2
;[�ꅱw&hIؔ��d2�H�\�@ȉ�2F�
T�Z�}Q��mԚ��	&��0�8n&����ycX6�5y]�/)��az�V@��U���Y�q�E-�ʸ���,�\���Mg�L��A�I�A��NO�p||*m3B}\pS�]�PP@ޙ��֘��"�-'��ܔ�1�0�q�Tg0�w?�}�����2�4޽���X�/�*K�YU�5,,-j�P�qtz�ÓCe�*��]���&��^O��6_����D��B�6Uf覿fX<���
ǙE���=s=!V�u���lw��]���:I�P(��Hb��t�W�����?p��n7u����a��뇭��9�S���4�z	��N7�ٝn��S�^y̩n��}M9�B�@�-m�ś��E�V�����
��NO!�������a�">���^�\j�T�`p��E����5m��c�hT����I��˛Ͼ�o/o`!����������)JW� |0,KhEG��;D�]���|�<ɂ!���"���Q�3 ��|O�X�Y�o�������񭧏���gh�<�|��B�k<?)���ux�-�O/�s�zCȅ�h����*�6Nn�����s��
n"\��^��X6��r��=��A��Y��ݞ2�Ľ#&X=8;���啚��dZ%ԣ�ի��
�"N��!n��Rpѫ�J)C:�?����	jT�E՛��I8�,Nس�@��8LS
�ev,f�;Q�W��p~q���=���#��F]��U�`0Ѝ�2�O�I4����E Ȯ�o6;b�Dc���>��Rc�p���9H(���"����卥����eHd��F6��$�EӼ��.���Ln
�d\��dz����@���u����|��x����~PIemi��,���q�4-�����0�P(DRw
��ܦ���J�g���K�<����).���J!p��ב�5�2X��T$6j}����g791���S����pY.j���"�b1��wy���3��>-�=�P���V�W���[�Mb[����l@JQ�ˌ���>J�����N{
nܰ9O��8�]����u����3#�X��s�jd�S^�W2��">�}���J��hv�zB��{X�- ��QŃ�x���0��u���[�e��_��]��=���7		P�B�<yr�����N[{� �!?F����B���c�	��rg6��j.�l0�n�+��l>�Ã-���!�M��]MLG�6��6ZG�vF��V�*	
�F9�1MhQd)A��w&�[��6��N���f�$�v�K&����H��9!M�����'O���l���$��o�pq�ʠ���R�(;N��L�dg���7�F>)�&�9����E�;??+ƄhS$�ǣ��*��x)Wj�����F>�d��\&�2�Ns�@�k�x�A��Qϵ��L,��3��"?р���H�6�@��ܜNr՘g�t��bo� /�w����j@�lL�:EB���M �	>�Á*�x���W1����&`������<�9��SU=3������FC����(�&���9� x��o�\���Ac�(4��X�t��}]�wC����U�H���Mw�9�|{�{���5:L����=L�x��}&W�T�VXGp _��>���n�K���4Z�&�1Ǚ�p�X�<�:����&��A}R
��C��㑠ũ&Gm�kF�34�D$\��M!MN�'�E�L�C���$�P�R�B%3M����G6������:����Q�����7��P�Q�5�� f�_k��n���ɞ���Ȉ�/B�0��CT�-Z�.�SF����12X�Vj�e$6����P��Ϥ�����Ѯ�Iv�al/������?���L���\�M��y��ݷ�;��r@}��Y��2LO���5�Y�����z���@b��d5�ӧ=��Q��*��F}�h�n�������9��7��/���z��i��ͣ}�Y�w�����ՈI�<uNƌ�>+�*=��F��g(�D���+Ȃ��D�L�����nP��t��#�>��i��\+E|��+4^�b>��sP3�"Ræ}h���}����:��t� n&qp`P>��&��t�;���3��v���0��H����)B8�+%���#���2�2YN+!	׵ڻw?�Q� �~�"Ŏ��\2	�Xs����}�BVD���*5[    IDATkc>4���Y�W%@<_���ؤ��Q*8b�q2#�kU5i��ôs�n�羟1�k� ߇��57+j52Ӗh����n���j�\�0s�Wʤ��p\:43C��E�3��H>���O�� �禦9*�����0U L�X���)VFA�j�ʨ'B*j�٠3L�ut�z�> �5:N9����,��r*Kâ�n1�=_an��(�.0yd褦,VO^�u��4	�) �M�6�JM�2��M )@ֿk��{����w,��&�����������1Mp�Ps�3w�
n�\�:�K��6�e��|�NZC�C�h`�\��]4�9_g�,1�����"ݹk;�\����#�q?��b2�T��~��޻wQbR��u�A�<���WG(-��+Y�m�Z�����ٱ$J(���5��/�����i�n��\s�-ކ�=�ؓi@�R�shog����=ph?�U��e4�Pü]@����6��m�ퟦ�/Ӡ�ap��4�0&�z	6�����ۜ��>s�xHY �ͥ��0�Շ�h�'��`�#0(�����q
���!����t�R��cWq]
����8
�-1���I����Ɔ,f5�gԩ���PL]�0�2�WE�N7"�c��H�J�	��ap�օ��㱈#�����O�^�1�x|���[�L ,��_N�k��
HK���S����]���29:FyMI,�#Ti��?�x�h��V�T�����o��яi���Ȩ\)�~�fh!/nX� #�<j&�T]�SA׭0T�|�ȥ�v��t�G��N7D���e��O����V���P-���/������:D=��'���#9��f�P�|��!5|W�Q���!:��p��$��	Pdx��QB<�>�!��x�*��Y�� e+%���m�=3E]��@��r	⛩�����j�X�;G�n�uoeε�v������R��R̍rMF��Y=S&�3Y�7ϯ�{����6��YO�����Ct��8�e*�}�v:B�f<-NFѨ���KDS��k�vڽ0AK^�4�K�!k�=}��<L�l�{=��N�g�.�tD��6^���Q�o�=l��,W��Њ�x�@&�&'��yڽk�4kRR)�Ӈh��]dKb�'Y�JӺ�=o�3h@�Q۵iOk��ط�~�/�[K	xJr/�Mb�1X�-vȝ���H��jq��iw��jP��A�87/�A�H�oL���W2�DӬ��MG+�#���S��i do��i��s�驙Yz�����[BS����yUoƔ�r�	��(����gDIHYy���uEg��ivKרR,R}h�Ny�S��ςP�U!�	'��� ޛo���m�4�����q����
��\H ;�#��n�|��ypp�����%"�LF��b^��{ĳ�j��N�Ӟ�4��!}F�fY��I�R43��͛n�6�޷��	���H��
+����g5�V�D�\��|9�Qi�FC�$�Mv�:�l���ѸBe`�
đ�0�Q=1�����*˂/��Pkz�Z3�\ !�`}��Y:����)����N�ڡ+�*��]���(q_�8�N�l�jV������~�O���u�E(d�K��T];J�e���8�rZ�{��Rɴ�p���u�o>�5��o���;�_{��T���GfKpCA��H ��.z\sc�]���� 7:����%1stR�N���P�DQ����8����Q�����U��A���ݳ{;텠��f�ktZ@ACam�Fiͤ�N��߷��ڽ��@���0�
n���T��@����ؿ�CpIx(���ӵ#�4`e)��h��;H3,v.��;s��!z���B��F��Neh]e����T�r������H���N��}��jH%$W�@�����wIk;$/t�����d�Iv�<7��� ��H�*R�,��ӣ�7:��ST*8�e��Y{���) �jHǸv�`xtlڹk}��ߠ��I�s�\E�/7��EWL̓2�L���@p&�H�Y!����G�����
�Wj46:B�|�3���1%D�h޸�#c>m�A���۸�����0�B���{!����g���I��R��#c�����V�sdT�� �%H��Q����=�y<É��<�#M��M�v����=����`\6������z 7p !�M�'Dި�q���-Y�<��_C�j�����D4e�0*��h]p,���cV�x$����Esk��in���x~�]Ԡ��V��G�L��u�J���4ow9���_�NA;OL`� �a�BtA�I�J��c����NߦV����le��7�%�V���Si���$�
 735�yl��6���uU��=|���o�k�i�w���%�� pK�A_P`i�����WƬk��<n�wbv̲C2�t�� �J��CZg&hǞ�l9��58�Gj�t̚�T��C2�Z����t�|%m���v`��m�`���N����Mw�~��|KD�Y5R�q�N��l��|�Z��A\�C��K Eְ��{��:�G�w�û�f�2�ُ����<��G���]�T�i]m��~�S�l��T:�o���Ow�}��j �M���e�g:]2I!��x�ҽ�F�,Y=���#ݕ�熨u��-7QP]6�2A���ߠ�F�e�T-��7F/z��\.������Iب
����������o'#��6�I�߉.`&�f0M��$�yx��Ħ� }���)"PU�4Ժt�֏���7m�Ӟ�L���[�>j�A>ꑚɼ���	��7���57��#U��a"�I�0 �r3]��z]�IR%�;�H���Cj��<������kuKS%Őhh�F/zыh�T����7(����	��3�s�o��Iߺ��,
[>怩B��P,r��v���,��Y��e5-gRm|���A
,������") ���K�!�I
D���b�z�}��!Z�s�h�	C��
��T����>ni�M�-���<"E��{����1��&oZT/V(�,�.�I�}�J
e$MW��N�Qiw&M����Hq��M5��󜒕�����<����J�ƣ��od���;�^}���L9]����8�- ���b����<B���聡9��>a���PUO�q�c�ax��i�K���fh��},��s!+��Fc�q��y�	ԋ��C�Y�ܴ��7��-�3�=�F�2o��v�>���޳�Z��ĉ5`���Ik7R-?@�%~ϟ�|��؁J�����`�D'mD��F�@����9z`v?��qH�kr?M7�˅�4T�њ�(���x*XY��:К��w�O��y��jDM8Juݞ�:����9�̻�Y�`�7�$�ѥ�v�{�G�-��fJQX�r\�A���
��u�b��4G����追��L? �3wB؍�.�؈^��w�K?����w��9 7�s�����?��:>�)`eL0$�������)Hq8_A�8�>���锓7���<J�sD����������R����_o�7NQ=_lT�J�o���i`@����,,pD�>&��z!$H�b:�i�5��SȂ�&pR*���������k�l���C��t�u*���顇w�?�����?�Nj�"ҵ2��@m����	�6�s!��5�@5Z��406B�a�\���d�� �a����	��ޏ85̪�\2��]��{���ER�K,DZ��9{���j�����Z�f�.-�g8�{�D�j�P���ʔ�B��d�����*�b����u�=n��c�f�Z��K34�Z�i �� �)[��G�ߺy�~�K�"�_����h���;<�7�^}����v�Ԋ�A	�;��WQD&��t�O:p�8\&ʲ_ �A}3dpK�e쫜b:��uT6KLd� ���ãN������ ��&_�z�Tc�v����Yjy=
Qc����n��t�U��M�K?;�������������	c���Lj��3}�~��!�1�h]Ȍ��Cr��z�(ȴ4=˭t�Đb��ʩ$���Ȇ8*�P&S4j�!��? �'������������#ؚlJ�Tߣ�Tre&&��L���A̍���̶�+�'FX#&K���1w��n�hE&*f�E����q�C�9���^��#��WU��l��Oo�����λ�D�TL ����B��@���]9VU�U:t��\Pw�b�NN�DO}�����=���g0W� z�-X��)\�@��ٽ����tם����p�����(����R�>L�n�f&��F�0aehQ.a���H�L��-&/�$���n����@��� n��n +���V����I��m���=�)��x���e3)2S+��Y��u�{�t����^���v���-��mp�8��<�]\�%ϣ�g�d=�Y���
J��E��
�U��K�I�OS��S��"����hb?!څ�������'�5T�iH����¤�4�p�	D�%&Mc�蠕%��y�&�[��/Q�H��%�����y���֝x�jeN��7�i��@��.7Srf���Ɓ�O�����R�����9���;�_�K����ۣf(�5(H� ����0H�0��c��sG�AF��B_f��X�c��Q�,��v�3��P�n9���ô�>N�#�^���K�ԁx�&S�0h<[�gs����V�ҽ��{�!_GA�����6L)�d�~���LН;���H� n9ՠcFƹX�֜���&�`��C�P� eB60iqd0@���w��ٿ�v�N�X�g�ԗn���PwbpT*8�s�L��Y��}VQEj
�&�#��hc��0n�,d��&"
Q� ��.�@�Hk֌�0���-�Mt�c�T_@�%�v�����~��[��;�l"��a���AǴ\�{B-#�f>�� ǆ!�Rׇ5b� �q��|������>����g�1��!��0���$�tm��ޟ��������g1�%CZHc�\y���[b��m�b
B�E4	R%�o�^c�f��8�ei̗��tڰae>�#�yC5�tڷ�0}�71����Q,t�uCf�#�P��i��"f��?�¹Q�ӦSN"���9�G�v�";���"��v���h`�g%��:f������Q��*RnD��_��{�B��m>�R1��@	��	�ʞ"d�?N���@�%�h��$��;d؞0Ǵ��A�A��&{�n~��8RtL�vL����Ys^浨�3����02�������
n߼��ڤ�|�a�u�Ag)3���HG����LE�;��*�(b�D�
�,�����F�CO��bк�0mĠ{�� �@Dvp?�:�����5.z�����o�ɥY�3u�&�s�ň�*��"�36��D��
K���� ���^�2�P5�۱cki���d��%j�H��Lc�)ep���n�����BjH�t�#4��!_^F��ڃG��Y�����~�C|x�Jȵ�XP� F��d�\*b�lAvΑF�B�Bԓ �6u���v�!%��	 �(�1�����{%E��.��6��b����gK6PpB�;F��*�f�����n��N���i��K�Cw��Wcb+����\C*�n�br�����f3���&���g���O=�T7�b�`��� z�^���{�cp��{������@y�i�ДCʎ������H�
D�A]a�� nL��5f�i�������t��J���_���	N$��ݮK{��Y���O�o�x>�n0ꄹ�f�M���<2�6�ll��FZ.M�����=�ɴ;�&hڵ����i)H���%�@�T��hDm�܌H���,�g�muY̆�QJ�PoX��)�<�x����+��}C�>4�b{ ��K���M��Z�T�;�r�Oa�C��P�@�#�hfa����y�O;��|���=xx?���n ��Y2��Ɓڇ7��� �V����?�N{��L:�8K�Y�OM����%�Y��e�[�t���Wn�������!��]��� �T���.���+�η� �m@A�V(р��Ej�m�\r;�k](Yae�5�4R��)T0#�on�xM!�D-`|`��=�Z�]�p�ˑH���!5>ۚ���Y�D�#�YH� n�� ���@��j Ԩ@M����}3�t�n��"[��.�
Ea$���Pk躔꺔u%*y2O]��BP
i�Yj���nw)t�Q5А�k�@�7ņ�u���!�]�g����I'�D�}*F�p��D"7(	7�:t��ӏo�	Gn�M�um�l�<���7b_t����"�c�����ՁE�7ӯY;��; 8P-pp ��B����y������~��A��2��2��,EL� أ���B���6����&���,�k��<0����7m�@�/fs�b���&�2d�����l�i��}��3��owP��e�u��&���Y�	\ZX��!|��Ad�(�Mц㏥��7Qa�B�'�}{vQ[����6��-�
��ұt=�-��(l��=3K��%&��K�G�	%�z=�SHͧ��t`q��:K���":�T���� &8��2P�.&4}�.�[���K�&}L5����B�G{g'��C��\��
^�� �l��.;�>��s�y�э��s[���Mx��K)NK���c�|��U�^ظ �ƪ�Ѝ����O ���A}
�R�Ų��L\�p�Q��h)���<����ɨ�<�w�����`~��?����u��(��q��S���Q��44�p�`X���xXd��l� ��3R��� �w�����f92D٣��@��4�!��R/�VG>��o��Sץ�R9P�iT�2�u�<V�8;CKaV��h�a(����
���֩>:B'�p�� 7 >Z��3"#�[�ѥ���n��/`pxu8L	�,8Ʀ/���BVp�X���Y��a��I�)Fd�J<L뻧?�����e��N�ǯ!�B���1����{��{�B:��5��ryD�B\���Gl�8��.�#T��|36���#bܐ)ܞ��r��2�bBDQ)_(q�%�v�K{�`*��X�k�Rv ��5�g(ɸ}1I�g&Y ��f��CU����˾�ir4��h"�>5�_	� � t�U
c�z8�nh4`f�iIo&F�Rb�*��:5}�&�t�9Oסn�������!s��V��F��`��7ZTʄ
)���#;4�PN���LA=�N��b_ Bl���n��Y��1����}��㞹pT#7�[#t�����-�@Y��,��!jtZ��� ܠ��mj�M�x%ܭ�
N�t}��eN��a�C! �p8p��z����s(��˱�87�h��x-��F��!��A��XX߳�� BS��� `�4s���f_F����E8u�^ȡCw�Ue9byā<� �h�X%� �����P[�M��{ ֐��t�f�N��8-�J:�%C [ߧ��#J���\�g�Bv�
�C�cp::���0��z]�P��T�;r
j����'m>�N;�4�j�: ����P[�;.A���l��<H;w���N�ↀ.����Y�ud BZ
��蒁�x����Q
����kC}5�Ye�ŧ=�T^4�M%�5�t�5ZB\����O{�d
�y+"]E=�K���2��q〹��P�eB2Go�� lEZ�(�t�f�Titd�6n\O���,>��B��w&���"@�>45ó��?�SCn�(�Ӝ-究�N�B�3���4�S=�H@�@�mϡ\���v�QTΜ� Q@Mf3��&aj�ό��� .�TF�%<�>e���R��uN�Ģ��:�B�MS�%��uy�J���Q�������l�"|1r�)v�*i�k/��$�=��L�Yy.�5i�Ӥ�~�&K��k3h�z��*�T瘁�-    IDAT�e��F��죝�~g׽�))x���>_gΚ�Cf<$�B��q�\sCH�]�`�ŏݯX�g�<�-�4� ���h7���c�j.��1/a(L��>>���=�k'�#�Pv�4AKM>�q��P#�XH3�Q�`�YN+�0� �� j�A�{,s�$'Jr<X���Z.��gH���bP�3¹I�������,*���gL��eU]�
�i{�a �!�6`S��Е����;�,�<����C��Ӟ�57�Ȱh �HT$����M��A{��c�H�Dj[3�n(}�&- lvtK��	�a�=.�Ǿ��h�N �=D�+��bq�Ӟ���i DF�B�/PIX3m�I���f��� �	0�ẒauD%��@/���x���),_
S_���O8�Hs�Y��iú�t챛��ͧp=���B� ��z @��&�]l��C,��id�̘T�Qi�ʶy>�)��P��cW+~�Yǆ���@V8m�x�Q��2���x�N`aJ����!�����j���T��S�J 8�?�4��Б�d�� ��t湳�K��CO/�Q6�P@����HU�4�!f����8�1	�ua�2e��d ǡ
pC��bY�c+Տ��n�g�^{��Q�� n�r��)�s��ά5��'���l��LN��p�C�/Ո�5�� ��T��a��1��/u���k8�-4X9��Ɩz\�)#Ȫ�N r�9��Kȅ��*�D�xf�G�s�8̻	����`|��"�� 7x� <�w�QI��zL�#�l`'��;��[�a�8eqB��G�,y��"2]�'��e<�Զ�nXn��t`o����d�V���p��gITf�}�`�s�Π��u�x��\תժ|=7�7����YM�	h��]t��$G���P�:HM@��f3񸓈� ��QKֈk��`;�J9�A�:�"Q������È� 955��0@�czs^c��ӄR-T/pLVEtp�C4ߏ:��H!Rg�7��q}�|���{�T4"ʤ,ڸa-m>���o�ʵ։�I���en�;�el҅f�f����G�HGQo+��4�v�R�"ua5��9�Taڃq3�fPD=tna���ɺ��*�v�{u�x�-��/Uϭ��l�	�C#�7s@��g�� 6<����0�l��L�:p��ؘ߯\�c��������Q���ԡ,�E�{qG[��@�m4��q�� C�f���Tkל4��?����G�nڱc��u�7e�/�ߚMO�۴�h��-���]���"���/C'��s��G6#>ҩ�����8��nӭDK�0�1x䏅Y?
`�� �NT���9�GB��hN�d
��X5��x|"
z�ٱl2GDp$��tx@E��JL��8r�k�2����Ʀ���k*2w� ���⺂��m��'�-��̎C���1��v��R\�B�
\�xnpyo�l:`���BF;�^<����#dhP�W��@���Ƙ~>�G��V�e_̙����T[Ã�X���<�L䅒")p��� ۅ<� �lڢ�r���s<��a����p:&_�s�(BL�7Hs;�ЕkC��H_���Q�%��J��f�N���<���N�r�(���O}������uk�M��ӟ�4nv`�B�3�s493�ׁ� ��^���SP@�EG��~��7m��H�f;�j�35dp�*x�06��Q�Ğ��TLgp]�;n�v���^���o��Ĵ��U��r�%@��A �2�5�O��E\�+�xE�G�[x��Y����"1�Ƣ��"%<:���t���g_=x^�W(cV)�0�/����������;X�򜵧�?����={����i����s���65d�l�"(2�����B��P��OP��c�DQT�oN qj(BMB�����ح:�$ 7N�b�%���a\����Er;x8��b<^?���}�[��:YP3V9��Dظ���Y!A��8>{ "V�����Ih�' �(d�yZ����=Y���"=��IЏ��s�%�Pk�1�V�L/�10���e��bg�\&��`��$�?x�7<:���8�'Q�\�n�0EFW ��� �����D��"��{�-.1�e�Vc�P��D!]8�c������9��k]�[3N�t ��<��rA�R��m5439A�SS<Q�v�{`��� �<�Gj�2�o�c��%�q�_� �q���p����#:[�^�U�'Ky�W�&B�nn~�S[�'ܱPD���"^��S��� mZ��N9�dN�!8��C���71=�T�{>-.5hjn�"��ajdp|�;�F1G��y��4X�;҅�'���"��]��?p0�
���$�'b�@�7Vs��Lf&D�/�~Q����މf��T���4���i."5�����m��`�9@���,�؜A?w��`�/*�CȺ��QW��m��c��p���q�J5�8�_���j�C����=G�n;tȚ�[���[�:�]��;Ԕ"�+#� ;"���Bk_�s�ƹ?O) �("B$1T
q� ��4�� �H��Ŕ����Nd���
I$_�C�w��ش���1�N4�+$�|bAv���	7`��� �DnlylN�Ҹ`��p<����\��&���X'B�L-CD,(��DB,����]�Ĝ$��p�r2�A��A��*e(�
�=���/�3����p���-ƉPA}�3<<�\-� "`lN��Y�������`*m;�㇛�;�����=,��TjB�(6F]
�w��gY��Mi��ť����&��ժ�f|����B��\\`J���
�pԤ �v@n�>i��3��2>KJ��ƀ� ��}���u~x=���`�44=$���T$*�s\�<����(ds�̪��MNqF��#m��M��D��u*�۠&�.eY_p��DM���#�D$S��E�tT���A?c��gq
q�sS�k�EqQ����k�?F���9h��W�|��k����y�x��������/D�#|"D��S�Ĉg'ؿ
��(��I&<�m��c�-�
��fH��ttl��O�W��}�1�~���[E���<pڢ�~|�m�2k�L��	P`�)�p]�ܵ�eX��wS:Ǯ� 7�)2�����!��A@c���9z,e�������f��ՎS���>��n$�k���w�Vx]���R�Iׇk`<c	�A1^U��ч���P��E�"�mL�E�'),ݠgj"��7�"���/{r����p�nذ��[h�(VN39jC�����l�ݣ
�\|���''�^��Z���L�a�����P�ذaG2��D�'�=t_�@���&�;��<�.jX�~�M�C�Nw����k#�2,4�,�� �X�N1�M ������:^��������yK�6���q�8�N���Kܵ�D��� �i�uUj5�>D�f�Z��8<��<��6����nx�K�<�`Zf�*�,���N"��.�_D��<�9pQ�74�[�4�����J�0`q16kj\�b[H�P���G�q�'���5��V�=�Zs����b�`@o�C#x��=��uR�8N�q���+�&��>�. �1�c�X�O,���dn(+ r�h1Z��C�q)oXT�Dn�i`�{������=���
nx��>������/����7ޖ���<+���I	�c7�.�z�C�|	�I�F2��O��`�'7"�~�N�4�BI�{p���8��	�~�4�8Q�@��������"P��4�'\_�
�j�8%����D���}�7�W�%��1���
`r$�C���k��ro��遀��HOḍ	�"�p	�b���p��IA�4��b���/�l6�/6�T�/"|�|Z�
���� ��@ �$����:��?���Iw�^E��ވ��K8t�B� ���NO��lb�*��Bm�J��!�� �8��\"��p�y1��{�iG��ڊ�D���dCV)(�
�v������닚`�(㢾7<�C�9iצb>+D֭��o���pQ��Z�
�t�uP
L�%��ݥ�ӧE��B��h�z�k ����GN�NA������p�J,p��l�g�|�1�QT\�fH����q�O
 ܒ��-�z9����T�5"�ľ��_�}�_�����P���܄����/p ��[�E�Yi�T��h���[_}�s�;������w�m�n[
^�J�M�s�p_��@J�MFq�n�_�8g-v�!^'>��kq1��3Q�K�;�����Pb�:���V��Ϩ�ŴN'�v�x"����e.p"c�t4�]�A�H���& I�T 4���'#���|o,\cb*�a?�d��P���S��	����<$�	�h�A��La9���1�,�Q�	��e����"���Lg��9����j��ֈr<P�$:� 7�����;@�'"�N���� ����b�x�  �DP1��'\���e�T6\��	�t)�A�#�� �"Jvuo6(0�������+<Hq��}�T�/�j��X�d�c�Ls�!8lF�쐢�]���+:�I���xx�x׌��� ��L�9}�$6��3��#��I�:9~@��?|����*�l�4��p���'�~�!�/�p��t�J��<�b6"R�^�:O\*���s�T1I�EY(���T��e���q�F<�&�f�^jl���%�0,c�� =n,h��� �"��
	�df��X�eM���sO��_,��E���'C������F�ɉ�J���L)�M�49p���(
dO�d�k���\���:3�������'�"�Ʃ��/DDH��ua��	�g�C�x�;F�T���:
��h����",Ce D�
��1�V"��8����p�Psc���Դ��r���"��S1�#���$B����Q:-��ŏ��n�LF�6�=�����q2�x
�1�w	�)���:A�(HW�fÐ�cכ�Cˬ@��
φ�}=�8�u��?:sX�TZ��I����8�C�  $n�Ğ�\���_��T�">�$�~=��B���UT��,�YN*P��dP�t	l��������rBl���m�ݎ#MD�
���L.���-�����O����)��9u�;1��J��̢����)��ध-R�ƣ&�)���9@(G ��@I6�(�hi���X\�{B�;x#!�Fq�Q�ǒ)�ԅ^߿�6�g�`��
תqء��&xo�떨Y�,2"���T$O4�pL��a��)'����B�
���AH��f�"�������"�=�B"2"����˖�?Z̼��N{h��/|�����`9���Z?
(�0�}?/�a.p�|$�i/
�F{A ��$EA�Da$G�/KR$K�SR�(R� g���9�� �P�$	߇?s�U�|A��i�dhj�HRER�G6��ˋ9��T,䇠�O	D@��x3��;�`�sp���"%����h�3O��8G�$�`����T�ൄ$�@u&�2eEaQE�'?��c�ҡ!���kp��#�? ��
u�H�E$�c�x#���P,��"3���i0�� �UЁG(</�]��u
v����czL�K	�H*��4;8��PK�'?���8���w y�C=B7���yʁ��4�d������������>`L�Ad��XByW8I�>��/�$҄2p�<�.��������?l1'��������8D
��p�2�x]��5E���+���t2�2PC�$<�tX��9!��������`,��2��gB��H�~$eD=�)�l�@8JԘm r�#�MAWRU5����n�^�L�Z>2H��� ,�=��LF��oH�qo���,��>��mV�q�q���P33_����y�3�-+�=�ŷn�*�^�b��hh��$��"��L���&���E�H��a�	R� �DA�+
ô$�iI�@�Rjbb'ᓪ � ��Z��l�J�˪�i�,Ɂ�ㆶcG��I�(]�W�0L���k��*2��X�v�ʒ�a�^��پ�9�"��/T�TUU4MSE#��"�{��E��ya�ы$EQYR�>�5���Q\;�Dx��Q<	 1@��*�H$�
8 �e��� P�#��-��'�Ma�#���K�*+V� �]��1�;���Fj��d|J��g'D`�+%�-[�!�°���aů/Zύ�qQ�����ʍS�ޜv#�øX\�\��"D|��������K�g�Ѥ>�"Ɇ\7�g  ���iq�5�����n� =ˣ�1�e�H��AR��""A�@�U��N���+<d��D��f=\�7t2�I<� X �b�����جQ<�A�ф� 7$�� ���E�ɑ����&uj�a�s�1�@�Ah� Fm�zqGTdC<��*&�']ͤ.�1c\��,�%ymű�� i�!����&�$*��D*�Ϟ<����B:�����s��_q�gK)����k륗��Y(��qT��M���1M)e�R�Pt$�5�g�Ty�43���K�2�.�a^�I��yn��8�5�0���V���iYiE�R$QJ�|h��8c ��繮���۲=�`.�KYSCWU�#�D�P�$Y5�P��-*E�燡�wG."+J�2�,�rR$E~�y��@�I��6� ����BY�d�)�*I�UՔd�B���6�} ��|)�TI2�0�d$I�R�1�*��RT��d��0���	�0�Y�x�t ;�)*\��0�S�	��x,�@�;�{NS�(�"�M>�،�����@EUU�PQ��
��%�8�BE����l
��`�p�8PTt�А $�\.�Ʀ��%5YE1��i:#��+���ZR��DH�ٸ�'�A|^�Bt�Q.�J	�I��pim�@��@@
	k�D(<�PB� �YP��\�/E�$#:�����S�eهXJ���<
��/�M�5Ufw�XNJ4�b~�#X&�c<����v�̃�	�\LĄk�WR�͇��?������x���Q<���X&��Ч��S���bN* ����*���:�/i�#�JG�hB��[3��5��s�-�����)�<���[A���i�J$o���������Tk���l6�u�����`�֭���޺U޾}�477�k�޴IZ����[,Fٝ;�J���+��<�N�Y]��\Z����Ț��2��'|�^��# �V��[o��:�NG��j���JYӔ�fS���׺����c۲$���)a *��@1$U�K�T�iHU�Y�j���5Y�I�d�ZQ�-]�j����x� G���B�)���>�?h���_Q��(�p�D�,)��*����v׵HK��AЉ°��j�Ȫ&ˑ�(z��]�=;��U����EM��"���u]��1b��b���I3H���	���呩��T�4ͮe�|YUd�U"��+��מBX˃&I�w4SVQ�G܈1,�A�z1WY�T5�d9�%92YSU�ʦSפИbQN���0���בj� �Џ�i����p:�?�%]�eK�e]��n�4DUJ��(�C)d=H�PLMC-F�A�*r�y�|X��(�.�(wSE��"�6b�d= `��J��ʎ&���+%�BsV�#�eI 0�._�0��y~WY�BY�U��� 9N�%�_\׉� 䄵�T$>P�w$I�Y��J�iJ;��yYR)��S��]�����O8A��>�ד�ka~���\`lQ`�)ЍP1�B+R��D�`6c=�2�?*��O��)���ԥ�<n���*��n���q�g;$�W	�92�@CU�%3#�u}!*�ё�H������iQ��$�<�?\�>�È�mSN�{���ZF��Q�a8���SӖyF�2��tMIa��16��%sƒ4���N�!G������z��<�w=�\�,�Bѳ�hZ)��HuM�U��5UAN�    IDAT�E�zv�v"
]D�<�'��H�A"�Җ��M�:�R.?U��N1��1�A�J0�����'K�Lϵ����7�m��%��@�����W�(G�=!��_ �����<���z$Ij�Ry,�&�n�_�X��)!��E�I�K(.D�P:�ˆ�R5v�&9� p#�q]_6�H�(A�E�7�@�+E��*��+��7�:���6~WY�4C�̔��iEU-E�o�a �{�"��<�(J����f����<וy�+]��~]PK�l�~�P��</x-z�_S��7�!� �t��SR�SJj
�0FwHI	�����1�1J���}������s���u��G,j���,��0�s*�xu|gS�ת�V���;nM�^,s�5�m�b�����|�,�c]��hD8R-�8����Y���n��Nd�f闽ve( �v�HU���.[ �[S�Sa��[o>��;��x�}�G\��a8p4iʀǾx�s�"�q��$�s���h�y�\R�O��AI1h�њp�n�_2p���Av��[Wb�f��~�o��M?��V|�ʅ��>�j�Y�hӽp�1�Ǥ�11��f���C^�Y��@��s�\K徼G/�F�o9A��۱� jT܌�TpkDxlĠ<����V4i�if�`�ns|=�J��A~�x�ߦy���p�S8SM�qշ�Zxr�յ˖QFƜb�@g�;S�E���̬���&0p���[���x��Ϥ��z2�����m���Ŕ���LL��`�~����������m��{��|p��ЅZ޽��
Z������0�T�X!���~f%g���p/����,K��ܒ�s��uW�Y����$@D�����M�\���xeOV�Ȏ��~xX��;6r7��C J1-�j\�����h�G��l!�O�����uF�^�����_�������a��5*��.�H�LOW�����3=Ehx{�EL���M���(n��8sIQx��p���W۫pm2m��-��H�Σ�K�L�WbD�A���J��r��t�O� 0�~X��p������j�� ���ŏ�,�L���y!�vw�oH[)��_���~B��J��&bgͫ]�uMzQ��5�t�[�(��|K�jY��"�\v�Ԉ��:�N�:�Ԫ&!#���}5��K�E�v�ư܈o*���9�1p�o����7�J��ppm:i�;�%�-M��l�荹6�/if*�{�F�P��	jqZ@y#�η���p��_1���oNo���8�}��Օa$}}�I�d�e�����㶟����6��a�Bݝ���e*�my��m�.�hf�<�G]���c�l�Mݨ�K��M��x�a�.�������N�|��L���]	L�1�t55���p5�r�A^��/�F(}�~����9�� �zp��=��G,��T��cy�}~�}��0�پIz=�&�)CI ̸�Ύ�ZhBG]�@D6�KPҨ`@��$nx(t���C}��E~����;t�2�u�Q+���#O�ё�l�ێ��؁�ۛ��|Ӄ��n�d��E��Ǳ�k��
u}��V���_bK)��~�Ch/6�U;��{���]�j:���a�p��1�!^	[��`������M䑾��FS�Q�Z��R��G���j���+��`i������`z*�̥���>/��rd�����J���k�4:�S��^�����C<ih=���U��S�;�X�o��-�����~Բ�������әM��r�&T����b��=ot�����[�3��˥:]Qhݨ�W���IMMM�d*�
.��n��3*%���!,�K[�疇��������T>�Y]��^�З���=���/Bs8�fE�NR�a�'��-�J��L(�^�D�J?ޝ�;d����A	����oS7}������Q��u��?v��7p�'�7�HN������BE��k :DMZo?�������O�oDз�T��"�+�!ӃN瘫������:�=�H{g����������a5���$�-@�7�^K�� �Q�G��n�:��R��`E��N#L��B�İ/%൐2�t}=��fn�6?���{}�"{�N���k��"����ֺ�Ia�[�U��NU6��&K����2�Hy��AS���}U��
�"9��Ma
��rKo^�]O�����m���i�e��%�m &����A<À��o�N�D�n��-����6�
�&����£F&�)	����O�A�
�Pn��w|/=�N���ϑ�E���{��{ա������'���3����2��sgђ�=B�ϛ�ϽQ�����S��~���}��I�B*�I?>�a��Z��a�Y����'�U`��)]*�J&���V�J�(	�E�]bbnn����gV�ˊ@�U�M�1�U0W�O	�V��/���~C<Wҽ���.��J���^�����Ó�.'1gR�q�U��%K����.��߀˿��Kϕvg6N���T׹��Sja���D�fs6�\�e]`�����
M�h���k��#i��^����}��vv�R4Q�$ҟbz���f��,��~��)���K�*��Zn���m�>+ra�]ȯ�K,���s�hYB�Ȉ%L��WbB^�-�j�GN���駦�����/���7���F\�+�P�p���j.����[�1�����{~e��Hأm���Aa43��ك��^F^.�.z %�[u�)���5UJa�W`t:}ʹ�E���[0Y�OCK�A��G�&���R��\�Q�<�=���Kxș����'��Tm�X��؄ �F����Шa4,p�,8�{YF�^/u��T�����tmQc�&lF�8�������b>ʪ���^�ҺQz���n��s���!�{]�UE�e�1�^�9f�Y��R�Ix��6.@��56t_K>��Z��jX<Y*�ϩ�5)E�*����ϐ�w�9<#�e�푇�����x����:�s��N���Ҩ�蟷:�x%Ug�>��Gǔ�ߣ��Y�?���"i]p0=�ј�erM�L��tyD�V,p�4�pP_�y�K�$8Z����7���-�� �pT�P��t�?7{�,]��(�`��(���F�Z����ڀU ҈�"#��i#""��isl��<G�+��^���l�8T]�,^���=ޡuh�pE�90�[I�Y�:�]9M�/7�m+�!�s��=N�<�~��j��v����Y����iYM���D4ӿ��7�C�*|�}8FM�}�ڒ�8ٶz���R�S59d(#5�9T0�ye|j�p�����r�$	(]��>���}c��$M2�� �xR�r!c����-�����}@����;|x��}�s	�lŏ{	l`�w�ͼj�C��s.�*M!����`<�K�W%�o��6/W�MPe��>�LN2>�6���e#6�N޽v�����@.�gc��A
�3AdMU?E�k�-���jXB�rXK�\Z�U��S�n�dt�>ޮ79��I���Y�EN����Uڅ��5��7n�r-�W��B뗡�N�'1�R�NR���/�(V�/�;PO��=��^*�tT\�)�4�׽��V�������$��uz�^E��遽e��u��N���;^ۤ�]�^��w�>\h�ԉ� �D���ʰi�`�-�fx���š�h�����_/ÿ2�UT��*��pClXW�(�4����γ��i[u���AN>�WR���������oi��|I�mR�^�F�}4ǣ)FP�[?4�&�zOm=B���������̆O�rH���T��ж����:��?/�뇻�G	�0��(��y�VA,d�/]��IW��5�Vm�t�ͤ�r#%2�r�٣|~�l^�˘�J'Â'y�6��� wh�D�͛@�ϟ���=��US���6Ԩ��GC�[�����ڼf|C"8���}f���ޠيװ���Ӡs鎣9�ޓ�}'g5�SJ��e��6S�QR\�����$=���L�j�]�K��Bij��å������ګ�!�6���B�������fɹeKt7��:���Z�
MN�b�͓|$\��҈i���|�2��h<?ڰ�����o+4W��-C��Դ�#�1�滉�͹�C�D4�.�����T��~��_c ���>��nl$ x>ؠ�8@8�(q��s=�GӾ�����5si����|$��lYn;��3]���}ގ-�<·H��t�Rq� ��"�Ns�;	7;�'6e9ˇ��`5{�Js�VQ�n�:�c3OU���p�z�Rjr*��;�)
��J*�r�?�� ZQQč,s���v��6`݂�Q��9���.���_����r���;>d��t����*瑺V)(���>!�<w
��k]������|��)O��<���:���O��wL�.��f*�DE����^2U�'1TP�Pxa�[�����ɧ鸈�^|4�n�9��5��?�^=D�8.��j���Jem�5�n���dA��އˍ�����? �{9@�x��	/�oj���ϖ0Y��>5�^y���<u��p��Z�sU��0��U����冃}es>�jx	/6�������/��=�I�Q�V�<]��:
���!~���m�\�����fj�b�\��ي�s�����|^(����!�"���K�k����K8�5{����z�1
��!�ɠ`��3� �;�q>�̉S�8�d���L`��i������k֟�&��m/x�<�¥���i:����44��b��n�fK2�4��c�7NbM� �S���	�h�ʍ;t�Ē���B+����n�W
����h�S�r�kXf��a蟀h(�kN7�U�y�^���'ߒ&�m�]d�O�0P��������gu~��uP�zfH�O���{��`>�Ɏc�`���=��if�u_��*�	$�d�7t�Σ�9-���h-�h',�N�QZ*yc/�3�lqO�x�	bTX$%��s@V���j7��Ƥ��1*��6D���:KO��ϫH��HX���d>�i���J�r:���T����Zlƚ�M<[%�瘾�t�Ӎt�S�j��!fI��wY����d:4���رi�E�A���T9�L>����9�f	6y��W� ��2z�I<�Z�3E��ɢ�0�<����Q;�PClTNoL�5j�l�o˕9̣�5�j=�~�� .���4� �c>��<h���b���乄<H�Iw#��������|��MD�ݵ�Q9���7���?YذB��P�{D��6=Z�8�a�C��Ѕ�ӧͤ�r�y��
�)q�� &B�ܫ�7�+�tX ��j�3�j*����/������'��u(|AT�g��n�)��Uz�<�|m7��f�v6��~�1�nnQ
<� #���M[���C�����D �:�.'��k�c~ƛ?��==p����i[��A�RF�7�v���j$�fO�NR!%À�e�_��[�DD�����4�R�u܄5N��ځ=)���̔�&3��b��|6��#�y���{w&ȶ7'���s: ����M�V#��������u��âV�Ť��:8���YԚЄ�����!��"��o��qTS7�@��?ة���B\�	Y�c�,�Uyقk��ZV5�S���gm��=��i�bY���n�ng�C��T.fsߝ�������	�>�n���>��\��b��)�"h�q�{�w�ׁ4#�,d��%�
�	L���������B�6��b����
e��JYÖ�%��k�7T/�����(����*.@6z�@Gk��#v�U4�����n"r��%j���u���״���tP�pxu �KE2�[����z�'�j+��Du
a�j��??��q���oxz��e�u���H6��Q�wk3��Q�$ySVR!�����*�&x���:JEQ�~co��x �
zA7*L�\�x]RX��t-�լ�yGF�������5O�𓣡#	�ƾ�S<*D�tp�Q�	��|�;�91��b��ixBx�]VGڝ7d<�9�J�J����D��T���k��ۡ�n��%��I*z��#h"�R�SV]z�E�xu5�m|�@�2YL���	�,�7Iv#kĩ�ޭ ݔ�9�`K2�"��'X��'	�$ �����leV)R��J~	 ��_q��_\�9�F�)���7�
�xd�r,��&&n�ɫ�+d�U�Ѧ"k�eғ��x��<���;�����5��
�UN�Wc:D���g�#����I�R�Y����ɑVMZ��Ú����)L��}�&;4|{���|r��f�YW��������g������k��\����LLI�����¬����,�U��I~����+c"06��XF��,���ǹ�r�}�
"9���^��ۈP���V2&�P�y9;�R��ة�̚�9?ȳW'���g/���_��P�<���� i�1@��U�T��ONq�7��_%a�z�ϳE)RF�j�:B�lE`��j+�jځ}k�3�����,��ł�9�$N�q�|4j�Mۄj�c��\q=�.1f>�p6��Z��_�} U�b��
+���uMv�Z�4��w0daM^0W�}@J�1 @�lw[�-]�[��k������_ب�K�a��m9�[������56����*-�bFw4v���@5x��O�7+���jl�'����7Ȣt]���c��kQa:5�4 ��xE��P:����������N\�̚B� ����{^
�x�+�&
 p��b��-T��+�i|K
�&Si�԰
bsL����1�pmw/]��1y��u#�����IN{�*�R����H�%]V���8�0�^�Д��Ua�c�1����&Ŷ�>ϗ8�E�|��2��d��:�� ���Uf��J����=�4��k�� ���Y}�E��tMk^�C�uL����x|���
��Z�>zS����mI$F�@~�`MQn�?AS�2�vؕ%���IZ�e����R)^&�?l5"E[$۾�v����ɿ�J�]B�2�z5�hl��aԕ� �	�l���	/�	y�(p��@�޼a9ҿ9D^��M��$�z��
V{w�Ϛ�2�����	M!�En��,x!���H����`�=��1�������M#��bŅ�Q���b���/yY^�!diA�2c_jQ�'�6��R:������RA6�T�/#�9�:�a^���B�RO[u��>6�SP����T\����l\>�@ w��\�������p���?��yFoZJd�"W���25�؞M>���8����546�Ae�����%Q'k�}�]�+��n&%����2�W�Տ�XO����j�-Я���i}"E���H�J��U<�֣���<�m�g�D�R�����W��j�Kȃhu��~��������u54�w.���/nhHY�, 3���Kڂ��bGX(ňH�D�E��%�9y�5'-[����a���xw���T�	��|]ڊЙ�dE�;U\[��(�.�]��?���Uf3�{����a˨�W�Z��ja�ɊJ$o�\�C3�D�I_��'>��!���o�zA\#���?cN�Õ�����u�,.�%�X��l��r�r+)�V�JT��ґ��<#�<��b�������b��߷i��ӯd�I��M�����~��-xAP�����mK�@�h1b���W��L}@����v3����̵ږ��&�?���鑶ӂDEO,)�+�V�ßQ����sx��7�W��ْ~��T�N�~��v��;݋ޫf�+xAyg�:�+���C�H_����\ˍ,��!���ka��V�į'����O�b0�Q*��V�%|y��]K�R>��=���۽E~���6Z�w���0__���&z8C?yC�o�v*����x��������U�N�L�U���+���&2&'�����|�&�<av	��_{��Ƌ��PNN����@*�j︭D�j*␪L�-�`��&�8{{{���W����������R��4���\H&\�(�D>�Uu/O��Ė+DM�������pDX�!
����M=��!�I=�jA'^ճ�>:.~�9^��{�1�-4�^.K�m�'��cb���0Q9w�Q|o�X�76]G(K�L��e~d�10�B����f�9�b�!:Jv[pq� F��!��B7<�d�����X(�b��'��b�(�rF)�
4��)��㣉�7j%2�J�S�\�߿yH�B^�L��kM�RsY����o�gUW�ҫ�2���߸#�,d˼)3���(c�@\���F�!^��˴�=N"�}��`� ͗��T�����0L}Օ������៾�ޚ�_��3����e56i��A�=�Ns���v�mo�f��{��<����ĉQ9�i������@2cޚ�)�@�ZU����\5 h�t�sݬ�6�cӻ_�T���d�+]��F�R��<E���[^4Ӄ�8aڮ�Q�;;���,cbU)���@+�EҼ�x�9��>��ۿ9��g��ZW�N�ռ���!���O����$�!�3:�M��:lT(�Pw�F�>�~��ο���ݫTъ���`��+d<�ĵ5���w����l˸AQ|z����^il�ջ>t���I�]:^+f�/��)΄D�Wi+����wj=��(W7�,ͻ[Ӓ8Ʃ	kfW~�y]�/�Us�o��{�%���>�Ԥ�L�]RjШ⊢����6"�@ �
�<���2t�c;��s�˻VlP$�RS����=���NP.���J'wfm��oAԋ��0޷��?6f�Eϵ���@�i[��{ݲ���ɭSNI���N����\1��q]��(����}�
1�|k�'0�d���&�X	��}7��,kٮ~�2w�L/����f��?�cߘ������`�c��9���2�N�ϊ/X��^�I��l�)G�����%��`��f��׍��1�u�S% D}4���қ}�Bq�E��9�<*�PB���v������>����-4�1Z���p��-rQt���Q, ����O�O����ؿ�͑�/pO��$Q|3ߚOi �+Pݡ����s�*���?W{��\�ț%����ǊO��RF�rF7�z���n۪We��YY�խ�\)��������}��cva u��bOSo�Uoo3�H�=�V�x	E��$������&�jf���13����{����,��VO���L��T,�LWk��r���*wy!JW��YF�b��;�ؚ�������+ז�Y���ɏs����~ŭe�s��OU��z�w�����֯-a]�*t�M����˺HA;'��Π���̃�M��/6K=c�}��;c�5�|||89�cX-vnUU4x�������S�ڤ&�ٌ��Uƙ�W��&\�b�:�£4��V���I�Q#�o}N,�%��jA�ߐД�'���,b7�N�h*+2V	��쐵TN:�֬ˈ��"LH����]�|��eNig)3��}�S,۠�����P,.n�J�!�b5%��XB�a]����*�'ņM�jAZY�����3��_A�j,ろ������1�1����MG�"�C�ȷ��B��c��!a��x��ٌi�_n�U�O544�CYG���9+o���U�;��]�^(��K�@���t�1�u�3��~�4F�X\l�5un����׮ȼ��+"<]j"�gf29wц�H�t	���Mu�"���,���\5<��H��݃!�+Md �0<�{N�l�4��m�t���[,]@���uE�C����Hu_��Q���Ï*w�F��R9����W��ƞ������wKS�?�^t4Yչ>��.��5��9�.��z�
����K�p�"� S����4����2��1��Xt�"y$O]����#�c�K�>}�e0@{Z�-��gJ������Nfu�Qʅ�����]/��\9<��m�ǉCc�*T֬'��i���2O!&�?q�)&��z�f��8)`Э�9t�b�_wF�:d���d�<�!�6�� �=p�j,�e!R��v�&�l���l���1�w��3Wo��k	+\�U��(�	p���s*�7?~�;7����`�� D��������@��n��Pb�{�<����f�3����5�/�u��7�ty'�U���G��-ł�D�<��<�QC�B>dU��E:`2�%ޠ2=;���yȞn} �=;�P�Z�>��@x�Q�[w��t��,�J
���@�=_|�׺����kl����7Ղ9�D�֧WT(��UTYa�ŜM8�R�����]�����G��57�'�n�M�V��򨉪*-j2(� BNM$8'I�C��hK6�(G�BǤ;�lޘ�"��t"��ւ��T�aUL�D峈��;�~Ef�<��}:�+L#9��������%��2�G��hЎf�Gw1s;}�i�p��2�/+��z�(����]g|�� U'_�"�v� '����������B���1�����ƃiz�	0\����,k���w�&�;҅�e����n��(iA�~ʫLM��E�pw�
uJJ����a��y�</�)���E�6� ������ۦ�$䪁��ȟY�򍭎;��l���	�Fw���M���e��3￥*��}(�L/�������1��������O\�k&&��c�QPoѶ	�4V�W{�Z�8W�{N����̎���CH&� �|_O���v{�L�����c��:�w���	�D;��Ֆ�36Ζ��Q�N��l.���%�7������ۈ��3��8�����-m�çO�r�j�bl"A&�%��J�M��<IK�'�7P��D�KCp���@��t	�$)Q3'ׁs��e��͕��*��:(M�l&�7�"Ν�06u�խj�_�A:,-*"�����6����/���Τ��w���������%��+�
�\�Y�$nc�����ޗ~~tB�P2)�R��TY�����N��Ĝ�3�Ɋ"j�K��d�v83��u����b�F����dzc��M~���7U�\�'s}��]��4,�3&tA^"Ť�=E�_Fo�����d��>�r%�wS��p�l�.ʷ�T�h����!;go3_��Pnǲ�D�X'Y]�Ş�'26Z-<�FD��{�x@������)�<m���Q�V4�9)]3r�wŪNw?n���w�ǊhÙMh�jg����/��Ou��B�������E[[i#���E���^�q`=~����-�;��rbiI��[�K�Wy�a\��CZ�BZj��k����y�����'����U�j�0����#L���=��E�eD� ��r���4���݈�d��`�B]�E��s����M��������!�d"N==�Bm�4g��Բi� �Q�]wc�����a;���U�9g��6A�s�R?|o��q'��g*6t����� ���x�^p�ҿts-�����n���q�b�B����~5	j�{;A�3�^q\�R�������ҏ��e����;�z7��m"���
��Uwu1�M�m�����??5ܽ�s	����� �^���%"{\T�k������K:N��kN����^ɿ;}7�g�t�
��NWlh����
����]�}��2��N���}��n$�[���z�����{jd��F�e���O�ӟo����l��� ��SO�^� <_�$�e�W����)���&���h�ɹ�oN*]s��,�e�uMθ-UG��@k[JZ�!��r�a�K���?���%� ;o�\�@�0-M?77��^���I��CDoƄ?�}d��|�x:F1�����sPf�m�v�L�W�ȓ��D#J�>����8���D���q*�ʂ���p*+��c�J�r|���1��>���W9�8L?�H�؞����^�St��M�~��
�u&9s�I$�y�G��X�	n%W�� ��N��Ɔ�?m��̌$ =��&]Z}:����o���4�@	^u�����+H�WG�ظ,e����!KB��FR��㑑Fb����0��U+� S���{ޭ��$�>9��t��G����|����63�s�$`��	Q8e���ػF}�k��aw(��F�YB�����ҿ�|��[������&�/T�vg%�S��
\�Lv?���^��:0��t�q�7.�Jf #];���-6¯(��ǯ���V}-�|^8��!���cP�E[�!l"��0�3��MLDp~N:&:�q���+\ ��r����c���텅��C4��
kZ]^��k�>�����Դ�V{�u!�aR��q�E����!��=!j�M���ے��Z����<�W;��b(�
33�I<�i�m�݅O�n�d����.�C��+�BV7*��/����F;y]ԊVR]�A]�d/?�_/8{ѝ����~W���(B%��~D{A��6@C���dN}��!���C�f�m*��Q�k�C���o	ݯE�A��r�\��}�VC�@�<�D����]E"hI�(	pR�kh�C6E<�2#?���ܐ�x0�_���
ڻ��jf<�	��ڊ��N�u�P$�l+JQN�Js�c4��� ��0�ǶzBH����x99��}���i	��#_��w_Rb<?�+���_���i�pr�:;�D?��:C �5/o�:�%΃���<�H!��x͆O���as���C�9�O�N���^JÖ5���vN �3|ꀜQ���l�p���:qr�w�BO�b���kf�Z��Z ���(�: ��X�.��ZIHw���y���"#W|�e�B^w@ɓ�yk�t��DK�T�Ik#6��z����s�W���OL�*��)I�z^7�>�~p_f����t=���LV���A?W~�gV#堎��Vkw(����mq����Io�8>��_nx�r�3�Eh��.
�ښ[m&l�}F��r���^���u/�������ƛ���GM6$GBJ,Cc,ώ�Bg�tţQ��FuZ`{N�-��unKQ)���M��+�������|Ce�����J9�)Z�Ş��L	���vc#���m��ɥ�LO�]|O�b�2У���D�ʒ���%#B5"b�+���Nݛ������Ҫ��+�$]l��5[�¡�Tٖ��,rxm�������3j�/�/	F�b�b*1�@�J�]F]��D��]N��doT���@��T(��ǔt��{�O���m���)��U����ݒ e���N����$��9I��`vh#�b7��0�QU����ڽ�A]<Iw%]�0f�; ��(h�W�~
�PK   �<�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   ��X�}�R��  ��  /   images/3fe24426-b06c-40dd-b590-a579c31a1c4f.png 2@Ϳ�PNG

   IHDR   j     ���   	pHYs  �  ��+  �EIDATx��W�eW�&���>��Ȍ�d&��E�XlV��R;@#��G��yI���� A�z-��R������e�2��dz����������7�LF��&�C#�c��k�oyW����\:q����=���z95i�O�u����cuk���W��0��C�/����С����}��P�J�k4Q��ğEe�CEG=#Gy�6V�V�JY��}e��^�G�	���ۖeգ(Rqg��~*W���[U���&�0�2��܈\�ҋ��9���J��DW5��9�r&��%��
�m��r���\����o��>zN("N@� ��ժ*W�#ʲ�[_��ވ���7�#n���,Ie�^6�~3	E��@���Hg��͍�g��U�k�qU(|���GGG{"�{N(Z�6�e�11�ń�_�z��F3���P.�mҭ�����sB��6* �d6q����F��~���WgG��8l[e�hq/��Rj�~2���*�� [쯨g���b��$��[*➙=')���y���N�sY����GV!
��`��^�K�	5<����*�&,t����Q���#*0a��@������J�Fd�N/��KƊ�UV=GE�D�,��m�ێ��W�3@(�[�~���> ��(��#j�E���}�&����Qǈ�.��0d����<?(�g���`��+����6�c��ս<�Ra6�[oG��u�aֱ�A�!�6O�%iL�(�}�3���@��T�['[%�U�N�ٴ�|�Q��D�(!��tT�}�	��dۮ�d�f��\����Ê�<|��{�ҝ����g�P���l�Z�F��L��`]��9#>�8����!�,
NY8?���X�z&�+���[�u�����|��F�(+�BR�>/qٻN�z�^bC��-�˛y�Dv�o�Q@�S��w���=]s8D��(��/�A���f�B9v+"m`�Yq�D����L������
��������<���8
�q�bR������Լ Kp
U*Wrv��������P&�[y=�+�|�����"�ϱ��eY�U�7��ؽ�FC岅�-���vIEq� 	���>41����~zN�(*����cǞgٽ��0���8�!���J��!m�W��sB��;�{�j�]�1Ic9�(r�{}_�y<2r�L.�`���m�a������<�V!��ka�|B�=�R��Qພ��N��j�^o�ӟB�Qi),m�!��睻ʍIۈ���Gz�I�س��g�Pd�g�C6�~52Y����ɸ-"���|�s�W���Z���Y �[�|�HJ<����y�@��8A⮘3@�X(�=��W��L��Kz���7��y�XЬ=G&C�3Z��s]�6:Z�&Gx�O��3��^B~ٸ瞉����6�0T�zwE&Dг�z�؏r�яL$�`�NOEq����O=p8D2tы�����L(~��k��o�PV�����B,�c�X�@N���n4�(�1)ێ����3A���z�/�.�7�P��Y�٨�D�b{�8�%��Ǿ�;�Y) GY��E�I%߃���yͬ4`G�\�Ŷ����T��k��5��N/��
�z��h�G�;�>��ޥe�(�D�8�8���w�{n�6��j6��z�ӆ������ކぽ��$�L�<����sB�Q�_�V�|���PZw~����s�ް]��d�,�8PD�S�c�	E +G��A(��X(\�i�X=
P	_���i�=i[ ǳ@(�F -�hA2{}G*
rae\2�� ��4{��"�qm��drP���=ݹ8��AB�G :qD_Ocd='m�����TD���!E~�Ѩ��z�y����:��l�A�]ő���yt7����z����>�D� �7�Pa3"=`���Ђ���=99�*2��C�V�����zN(�se��n?��O;���FG��]�>�k��g�o6G������h����fz.��\&��[���~����l�"n�*+bn
� �m�焲ju+
ђ.b��c�egz����"�{Ȕm6����>��ݗ'NY�qˎ�����sBَ[�f�&�C`�B��tf۲�<�]8h��z�l;*����&
�ȸ�� {~Oq�|p^bz���Y,
G�	g�ny��*�Ej��E4��~�e;�V6�s9
��g��͚������w8���F���T��	��v��M樅|&�=��.��	im���	ϏrQ�kv��l�`Y;��x�ʊ�Oh�D����*�韍��3o��#������T������Ξ*�C������۪\.���r�z*bp�Q�N��%�����0�S��SB��;X�6�j���ߪ��#4�T=>�fs�tTV�=��㸷�]O	�l�'	HdQ{����f{.���?�h6=��}�[���z���G�H����@u߉��A
�P��KK��^4���=��P��<h[�
Hl!�Ps���,{�vQQ^4Tt,kzbb�kGц]��� �@�'�e�����e��%��G\�j)�A/[�������pg�B��z������}E
Y�� �W�6z}O=%T�\���X"�P$P �>Lom�u���,�H�t��B)���ȋ\'�-(�N��xQ#��B޳��R��Q�� �l+ �{�C ���n�`�d2����z���˥�n�i���r����x�x�:��kw������������:U---�w������?|������h4�ʵ���7���@����� �*�J��7=�[���7#���rvL�����c�^��(h����@_3��։s6����B!��7PZ���_������;���ѯQ�:U����7���/����i�nll��vx�ʕ�E\���;88�.]�t�����@���Z�CRf��`6� ��c �QM���иyp�\q�c\b�J;�L��8��\7����;<y����fNz"9��C�v���7�^�����V������0�,�/[7��\��h����V�}c}�c;^c�r����[׮^���흃����D�Z=��J�D#��a=(!qc���
]��K�!\��R��x%�Pb7H^��r>-v�H�q
�7xD��4UD��kW&o޼=��뱱�?�������Թ+����'�N�_�<���������WCժ7�������o��_����4I�4G���Vk�����3�<��˸\��9qscK���R�*���M8�&/?��@�1��\���Kއ��f �{g�������M2z`,R��M8�c����W_}�l�U������p�������g�6���g&�쓫_��v���>�[�OE(�)���9�����Wn���c[�776ǯ\�:x��̈́:t�;��*z EJ[�p/���رcjttT���3������ڪ� �
���\^Lᶾ��d�&��J< �&L���;�0��kjcs��#��@X<~/--���-ڔ��Eu��A584���pOChl���x�����Α.������t��ӓ�O��oB=x������_ܹ{�Ϣ8>��~���裏���,�R��P#C�jrrR<8ɄYYY�_R��E��ׇ����gZ
@��*,>/My�J�h��p.�; 8�O����V������Bth���d",,�)�E��tC-]�{����k�}��y��Q�c��s���|/���}wrj�wn��#W������k������+W���>�ş��7����߾}[]�|��x��{�/_����� s���8?(\FM"��!�pp'i��x��a {���'���d!�=!8O3ga��~��u��>&��@��<8����y�l��_~�����AD�P��3�92/�ݻw������?~\8t����︕��[[��샇����W/��C/\��q��Z���E�kw�������[��i��x�$�E�/��Ļ�����n^< 8	�����޽ǻ=��!��ϋ�(X^^�ED���x&ԐM�~;�Y�Z5�
Ko=|^��#���̀9s����⒚8@���H�U��V>�'Y��J:m�3J�r��	��7n�R$���6���E���v�*K��G�3[I�0R[~p|g{�����[gW��jag���{rq�ĄڮV߾~��_�"�{��:w�E�kY9C|@ǜ:q�9J? n~nnN����B1�.WL(A&Ù3\�t��b���ݿІ[�+���b��p�эTNp��Q�2���ApẐ�8p�l��)ұ}�oHp#8�5�\7n��!5�76��i�K��8I��_ax����y��髿B�g׶7�������r��a�"5H����#�K���+�̙3�3��p[������qc�]�8/��ax����h�E����!HL_��JHB߳Ş�4�	�I�B�!��=�5y��F�1A��-u�����2�;�U*5�'��W$�I��0q@�H�F^`k�aJ���v�����l��_]���^x���<�`�ޞ~�_6��~qe����/��֦���e��!���=���!���E"����X,��J&
!��W�5��Eù��C�p5�!�C�s/H�Rv��8Y,�*�f�ek�X0��T��k t�炘�ٮ�w^�L���B���ł:D����f�Ty���e�f3*���p�s�j~q�;��o����W'�N��7��ξKr���;�w�q�fff�gF����M|��'�浫�\+�m5P�S�|!1>�Hn�B�5�_7b�Ħ���&P��L*�5�l�Q"dHXD�D<S]t�WdD#E�:��U0.�NB��-�r���!���KO-(8�oݼC6Y����o���u�Д�|�<��Ŝ�+x|�F����f��z��n�A�]	uccp�έs�֭}���f�J��whQPUWV��zg����SDv%�71y�9��2/ޛ��g.c22�:Ds��'E�-����0ZE�iN���8u^�u�骜������m��"%]��6	�7�f~�ZVWh�>��e���\��6�*h��ɽjE�LG����S�N������O����	��_\X|�ٟW��Eehae�I��g�-�� �.%ѥ�nԊI��m��w�v+DT.g%���1�������{k���������7�-w-��8j4Q��p '�SC��e;k��!�0��3���s������M��3g�WSG�,I�
<,�������C��`}�o����o��޾U��IΎ�f���h@;
���آ���m�������U�ʣ�6}~P�odl�v�6��Y<�W7X�'6���0lAv!>ǪJD,��M�PsM�z�.;[A���߀M����,`�h�5�k*I����x�*mTӚ��W�d��#��s�ՙ^ �q@M���s`�d������
����_x83��r����[�;t%T�V;A7� U hh�;G���i�$��|����믱����e�X����D���s��Ő�!�f�[��qՆ���b�<'��8�yeY/a��a�B�����+���������9��hw�#��퓸�씁'U&�E}���l�5	��+�wY��t~��'o���z� ��������"��D��6	)C�C�?xx��j�p",�_��	�G�~:$�;�o�x�E�G�����,0�1v`B:t��W������,�8P���k��ɜ_K�q}r�Fы��E{ѣ�3�b9fI�p�e�%��R��N���*���
x�����a{�d�;�,�e2�㦲�����5������+���ϝU��c��f�xc�^��b	Ql50<�F't����������V������q���N� �k��H�u����h���E|�w��]Q��%b����`����=��� m2�l!�D���:?8��h&NT2��g�\MЦ@|�3��6���CWs�O� �E%���k�?����X�g�0BǎW�^<�N�yNy�q Η��R� }df�y�HM@�ɦ���'�q���%���48p�D�e�ߵ~��Ф��B|g8����,v ~V3ˬk ���.-�A�F�N;?��ZHAm��d��:�Lp"�a�8�~]���F¥b��w�.sIo��y��á��M��Hԑxκd����A�7���u��HRL�B�������0�����'0qo桺v�:{mN��1m�E����蹧?��쿐Ε�I:�>�\>���5w���Bo�4B��V}�Tq��*�"�B��a��`}L[�%v'�nm�.ih�)�-��SM�5 
DX���bD$B�j����=3���I���P7ݤ_ :�.T�5i�����(�MPtNp]�!R�y����/k���a	9to>��$
r�LϝQ}�O���mu����uWI筭���k���Y��Ͽ��z�uu`d�A�*׍P1��PPT*c4Q�"�hi϶ev3�׈.����n��\$�C�#G؆�xDas{����-؝@�a��}��7w���=p�Av��^�o��I�q#L�ok�W,�1��%΀�p��u��	����F}��|���a��Hӿ!aJ`sTh�D�)����	���Ç�p�J�. ��¢BF���p��(�6u&��"��5	�}4V���8 n��x_Ėx�����g\M�q��; J���)�m��<�q�C��S&n���]�z�	n���.��$0���$�KB(�Z(A���̨�V��\s�������j|b��3@ܺ}G?�����LԳϟc������>�1�sP�vc�\Ӣ~Ko������Ј���~��}�E5�p�1<�5�#��ʸx�u���������������z״^�!>7ǲSW��Ɂ���AH
烛
�����Ͽt����w��S�O��(��\@$q�����q�:�� j���� 3�,���f��3d��l��F��"���׮]c�r嚺K��o>f�~�{�Sg��0�n@:�4�@��8@�+&�&h�Yo�Hu� �3�٧~�Z�T��
G�ͬ"���f�h�E���L�N!�X��L6 �DfE�I����`T/,-�=-p�����C� (
��.��|@2�֭[l4������'O�K_^�H�vz�\a�}mcC=���� *�&D�n���f�����^V^y�Dڐ�r�=�K��eB����/� qa�Zc���{�Y��������)�?ٚ��F�M��H��:�I�d3�{e�v%��y�!5:iQ8Et��b���]3�VnJBx�4Gb�y�q����â���y�]|�GO��c��G������꧅�̢��Ԋ�d��΁ ��q=��{��"D�_���q�:uJ�;wN���?�◾�	�����jxlT=�?�>��oP��z�L@I$� ���� N�w�>��\6w]�qt�(۞'W��,Jn�p�p�0X�e����6D� ���2�q8?$Y�<?���'5*"��0�as�@8���/#I'̑�v�l��/�HGT���/���YK�M؋�U�����{�Ν;��O?E(m�q� �o��o��a �^x��'�'���?gn��~1G:gC��o~�D>E�ݾyS}���L ��jYg<�����3��:P ��\�Dn!���(�j_��^-�
�����I�<�= ��;�Ƨ��4�RVY�Y�b�}��/���$���9 �Xf���C��l|�@"R��h��u02�I����G@m0b�-�%8�6�����#�3`�g�X�bs\�rE!z��������^�$���L�M��`T��&P�!zޣ�O0��V(�@f&w3wc��b'r�P�2���E(4�-�.�r��T�bb�
�3�MGJ�[�>��g�)]��j�C�1��)cN�X -t�\������^
���X-���go\�0ǳx6b���W_e"� ��~�Z&}έ}�su��֩��X�:4��7JFn��yY��b�Й{�lH%C,
�����L��|�yaz7�|�Uկҳ���l.�<.U�+��&+����(���ϑ�/�$=��,��x%��%y/�iM?A~Xh8De�I�KbAM�%�{"2$��?���g��ay���� ��Q�l[A����/^d1���������������0r��E�v6��@����x=v�(��0��78��P�~��p�:�ts��L)�~�s����+~N�F2�IO��K��T�'aH8�?�	
�5[�!
�)�dWl�Z�1����Ֆ���˧B�9_&�h`�P��//]�����S+k�|}D�(�RS[�#�c�"�s9R�!� Ȕ��)�bro XQaK����Fh�}�d���O�����"�[p�����Nh��M�0�.�b��Y�I��������o�y&V���Ky=}^ܗ$[JDB'Y���4ͧأB�s���3 ������CɎǀ8��lN	��%����s��R���bo���r�b�Q���0�N��g��i}���J��|rز۹lOBM�&V�ǫ? ��Z&G��M��s�T��D����ɢ��&�š<N�^�{,[,��rmw����N��xmx U�a��.�8j]�8����7���H�LO�[6�k�"HH ������ܪ�"��	"бc'8�������/���tN%���1�8�V�d��s�k�	�=	����?�N��iGI/Fפ�z�d���NG>�>G� �t�=�0ViT����MM2�=[J��t��|�8�����vvݫ�?�|��������qn̾�L�C�Nc�gn�l��S��W�����0�ח��&_!�4�g�"�ŸM;k�ôR�ډ�^(i��..ۿ�Z��=ٺ��ѝ""�ϒ�
�A���O_[ϒ��<,*[����3�ׄ�6:2�F�9�^�E{ˍ��ʯ{^��'j��XB�
����R�g�p�8�8SKbR�"�(!�,dz�;�jh%����οb��'�{�j�s�{j�=��i �2ɝ*L� #�ޑ$�(�ŤGb�X�c��+55�����k!뉛���ɼ:�c�9IJ|��XB�E�nܘ����3�Lb�,�,\��:-l�E��]w׏����:ǝ"��V��:�9�?���~vs,���D^r������gH�qBi>��	��u��j�Bi�(����&iQ�z���'8�(���}����_���[�^�xG��vp����m����)ݑ�ND��t]?�\D�ٜ<�g��̚+�Q>B}��6�v�я��pq��PLu3�B�*F"�N����P��A+w�������gA�:�J&����,kw�d����R-}��i�)ߑ��tK��')J��+�1�}�m��Mƺu����J���*()P��D�τi%�J�QL�ضkq_���p<�HNGiB�Ŕ .��ҋ�N\ym��ܖ��"\7ni+�k�ŝD��g��X�d�(q�""�4G�r!rjd|�9H���k9�\�%�M#��є�xM�R�OB�'/���JɃ�)�[����󨳘ڋ�v�Ƹ�������
ג�g��%�,�\��zُ�����,46 |~[�NL	�k<v��ń�Ԛ�	�8�{-�jW��I�T���(F0�4���f����*��l{�����F��Ig2ɱ��J����J��#)�?����U+��3�"ɤ<�f��]�/	��/�i4#��U&�a��-��$RC\M���l�g�P�) �ڑYPo��#�ϫ'8��>���ʕ�t!JZ�	a���M��T���-b���ծ��"�jC~�(h���[�	�
;�yv�خ�M"��%��yN�uS0��ix��{�4�XJ�l?����	-B�ttOhR�VV����:qB{�]:/G,�)6��N5���P}��?�+�8�9i�J�@�#�]���x�a�Z-ŏ�F|��Sg���;����vy}��� �$��s��S��8��<�c��Na�<��ĵ��m�������L�<��F���+Ľ�j�����'8K�F#���"���&�ҋ�~�ݖ�?����;�99:BuC��p�t���0d�L������~�#�����w�]&��;��|u؀��0�%�C��1%������BK�l��:���o���Mv��黵��676�8��"�M�u-5���
��k[ߦN�<�h�<i�ۋ�҈�a�M��&�~n7��<h���B����2������:����{�ҥ/�]"��1 ���չZ�&b�~W�"� A�8a�g��9UADd�~�*ǭ�~ k�t�F���z�cOB���ܛ��Sܬ�����J/v7�����{j7H��;)!H�=X(pPl�}�X���0J3d��"}uL5Q��C.��tϋ���
�}���4k�?�M���/SC;]m�;	�n�g=<��dp�w��-N�F�e7�8��W���P;՝��;�oH�4�@�64��t;�4��p�Kʲ�G�q{�N����k�?�����:.b�����k�#�2�~�}����.3H��'����0�s����Y�әsH˦���dPA܋�ٝ[�����A~�H�vL�bΘȀ���T�͒<T�#=����_�i#��y�	9$Qk��ђ���~B0)�R��O/->��M�r��NdDƭm*
�@i��v������<��q4k��ՋNR��Y'}1;7�v����$�+���E�[��P��ב-46q@�k�,�]u�'8t�m��N�����z�'��X�NyC�F���Ї�I���7����z�Re�L(Y��<F��/Bݻw�T���n��(@ki��#��t�Q,6�. �kE�=�FTm�ƤT�����zC 8p���~;�Gr	�7ZP��+#�><4J��O�?^%]��m�)f�~�+.2c<����\%HHm#Ψ"����wWy��ݓM��A��A�t��Fp�a�{g��?���S�����qi{Jz9��thG{�"P>+edt��Ah��݈����� .�!�q�5B�@w`5�Ğ�pm�x��B=��s�߀ti  �����3T�g�E�x��֮M�8X�Z�pܮ��t�;$K����/����%�B$u���kr���|�B^��%�kY"����P�`A�\�E�	��hG��Q�h)}�@2yq�Y@d!A�C�`ǲş�iX1�b����U��i�]��D�X˴8���i�tėP�����`�=F�����X'�}��M���EZ����o����m���I(n�,���gI$}饗�=��7���ӫJ���k���	�Q�!�䶋�vCW8"��K�4TOsR�4��[�V���A���~��j�\e�y�뫜���Sf���>�8����@ON�kts��¼��/�\�
 �8Qdp"�7���U�%���;�}/�s*з�@i2������z<.��ɀ�@(l�F�g�ͪz��YK�*��YZ3�NZ���R���q�%h��4���!{ӻ*)*k��ڎ�B�W�t�͇��@�юFi��ϩSgN�N�}뎺C�h���JE��ydð'`CZ=�T�q&N��:$ γC�R�(e��kg3�N���Ç���55G\���Ρ�c#�D ݍ���z�.C�&
bv�@!�������H�>v�X:��bu���	e�6)�Ӏ ��k�7-�q�_��H��.�l�B�Ǟ)h�`}�������3�,�䄣 ��7��t���E�wY�`sT�a�42���v|m����L ��cǎp[ 	�\p;ٞΨE-/��c�ܸI����I��uk[mml���lH	���)C#LD��:q/82�@�͇�m0�]G�;��aN�qt%T�Dnl����@��DI������m�w�&{	jY�i�H2���P��K���jxl�A �|�8�8>�&N���ja�����X[a�jV+*gR��T"\K���I�Ǐ��!�q�u�Ψe7�gӢ����悙-��A������{U*�A,QذE�~�ƛ)������{�24q|
d��&�_+�5�Ъ�݅#]��kC������7@�K���<T�}��*�pe�-
�.��2�^]F��5����{�c�fY#=G�s5j��8��QR��\�൹;[w*��<�.� ��"���_f�gԋ/����l_;�J�Ǐ|uR�[������C�_C�� qj�kٍ��w2�z�#��LٴW�=E�p �
�3��;8� XH@o�qum�w{�t����&�||��k����T�ϜT�#��"������@ݺvC�2�t3�dq��>�捶i��(k�Ӛΐ���_�K����O��ӧ�/~�3W�f�#v����p;ӆɣGA�l�&ط����+��s�(�P��>J��|�r�Gwτ^ɨ�H����P���msvu�L�$a�.���Q�+�L.��+�D�a��p������y8�puu9�7�M�,�?4M�gl\�^ׅ�Љ(�p;T�gXGIḘ$ܚ.�]�6i���	z
�6����RC���n�	é���� L+��{�7FD&	q������J���L�ι�:n 7��i�F����N ��Cp��Yu��Q��@Y(��pz���
�����nݼN6V���RGg�R���Gu%g=ݼ�]Q�菝8N`�('��u�/d�>�G��������d{�=n�z�2��u��8�&�kqN��(/�Hp:E�R ��F�#��7���2n��P����q��&���,0\�3	�w�	�L� 5P�����gN�9�� ��6��w��f�{w��̼�������=p���E6
�*tc��G��<�^zE���k\MQ1�i�R���(?{����/����d��=p]�&��$ez���ZE9�=��ɺ�J����`����5�!�]؉�KWq�Xөb*iq�$ai@%�HO�	���
�P �M��WbyuEݹw�헍�5���B�n�&����$�����MB��� �i��;�z��ak.��kH�8@�� �Ңބd��޸�쑭'��~`4�\��P=�9�`}��ܘ����T�;�1���nHb�%G�T5F��W�û�B�K�)	����Ђ ������H���?�][hq')X�A��s�����+�{������p�B���J�n�4����d�������=ml��1��G��~֣	;y�ys~-Z����
�����	�/\�F�~���X��I�G��籖wq�X���C	�a���]�)�y���t@Ow��U�z!�y�}����9��Y��-��CPe������3$�$�Y�d�\9�9�p�8_�#�-"��n#4:ԅ&��@f�r�t��K�M=��)�i��&�|���N+du�\�Td�oaa�7�.(�$Bc�S²\%φC���'%T�<�H&���ѕ�l��-��n^�MEJۣ��dD7Sl$� 9^kDZ�ɰ����'/��ې�}�=-�A�;��+1i �r%�7�� ����	�(#��_������ك����F��8�9�Şc� L�C6!8����<��%��̏��C�]�%7��b����`7k��(�f;)a���0=VOg����������Fs�$��L�R�ĠƖ�"e�eR���P�L$��xF��D�:��I�v�>�@?'�(�6]�ŬXA��ŕ���L�	��n
2�%?ϊ�%l��b�z���ͱ��Y�f�iGi�J5M��2[��vh��M���BͥD��	��p⚂[(��f��-�S���Z���F2��s�$��MSlJP�6>7�K�}�`!q��j���-n��@�	�C,Gi�m��hw�~nq�� �b[�|�9:Tl�A�,�Svȉ�� ��ݰM.��N����v�ʿ!^��pB�g�J�숨�L�k����x"�������ѓ�w�D�ko|K�9���ƣ�!
����y��ǈ�Q/��9+5���#�#ݬ���Ֆ�������>[��lhn�&�ur�#��U*��;qG�x���DJo ��3&�u���. g@�h"0ᤚ0��xrޕ2N�r�-��#����d���ܽ��^�y�]w��i3�4��H!C���s�����ŋ_h�	�f}�*c��:0l���56#�	��JՏ�i�
Y�(ܧ�c����H�\,IX�@�v1��^J����D2�AmD|����c��� �?��#����qs��f�X����x�9����P#&��<F�'O��
:�d��c]��nb�7W����(.�\|K�J1��}������$��.��4w_CYI rhd���m�����5���/�f�{N��넦�ؒ.���-�S=dc�}t��ް�G�+M�@|x�e2��[�����b�"��k������X�3j���`K$A���8�����#��M#���qD�ݘ+�8�����f]��h݆nRưƿnXZ^P�/}�Y��A�JR�j6�>������6�M�8��[�gY������2+
1�{wn���6�u�'LZ���}-��+bY)w�(�����Y"��e��۾��bM�Ҩ'}Ӓ�'��`k|�7��!�<3s�
[�8��c�o��m��/��^y�e����j�>�+*t2gю��f�]�������֝��fȆv!�b����y����9Ҍ�bH���^�;uey�m׉9��a���8��-����1󳊉�m��?E�Ý�G�S�#!v2|�}��N{�Z�O�'�|Bp<�ؔ��{�!��29y���K/���6h�1՗�)	t���@K�? �:B�;��߈�J�VU}���ru���w��m5;7�]S�9��6�j�<Pro�� ��~��=߲��8RO�&���G�sP�a�Vb��_ҷ�.�`gB���7���l�k�v�_���z\��쬚S��]HĿ���d�FeM�L��-�L�����S�E���d��^��f	@bHe�} RL�cR�E�
�1�"������1��,_��/0|��ibaB`:���Qu���Hol�]����9R�G�>�5�)�w��=c����┡�C�J"%�0��TȆһ��F��M�i��H�!¦�w��ٸ�B���9GS�t�ֹ4���C��j��x��.���jG���i��2�����v���}�;��4�˛!���C�ح�7��G���?�N�_\��"k{G��F����HO!�;3����x�0a�)4p-!�]������w��r��jq�E6M����0fO�g�*�5���� A+���-c8����E��S�������X�E�{��6���\m�������������8�8z�8��#�[�
����.���:G^9H��g�h��p'i��w+�`�bq���=&��B5��HE`�_��7�d3Y�LM��ҝk��.N E�v�R��bq�9
�9\����Ƨ"�2юv�Q�#�I�D�n�Kǳ�t����L��S�y�N�҉ ��lr����77�9���͛<�A�;��,�נ������~>��(�&�����n�%2�6�&�ӫg�E�QY��D��ۜ9�>u�h�B�>L��g��cE�P|]���K����OP����N�'9XN;��y��<����y�2�BGf� �$q?2�[%��#���.�n@�Z��N=I6�UE'e� j�gz̾��K�4P�\��n��N���XP<�)N�ośf�EzS&khŜO���c̹�?���ܒ��~��8���7	5�KPj'�G�Br"�w��O���ruK���	WR�^�g�X[Ovq�� ;g駐�9	�OY������Y56:�N�z��؂����;b�5�;vL�����0����>��7�_��Z'�aV@�@cr�	$����|�^��8����!�_��N ���� 'Έg�W6�癐�OvI�nQ��N�N�$}}W4ز� @��H�7���X��iB'� ]Z�Dm��$$Q���Q��烓u�}��Un��֨�B��j/n�����7�őW�3��S�:¼��&^|���H�h��總���2&�9��}>�1-����A���	�psKb=ϳvO��Z�j�����kCm���3_	��m��k�Q[�%��@{&L�L���H��6
������1��� ߃{ ���cA�Fo���̧��A��?�>�Ն��gt�+����.>?��q����&~?�c��{��뾅�y1Iw�}�h6���J���{���`y��S���}��WT�.��3Ӵ��@�� ���@kX.[��Xt�@pd2����B�f���4O���^{�U9������B}y�3�F�8E���d�����sϫ������$���7�ɰ�@�j];��`�����d%����J�d�t�XPn!�Ȏ�}zϣf�{����鬿�먘sPf��Lz�K�K���ϩɩCj�8NP��G�hI"�	�f��.��R�n߹���HX(�u!yz�e$j"�ٯ�~��Z^\�vd���m�uBNh��j�Y3Y�I�s��߫�J���y�2r6��`�!�eqeY����"߫ǎڳ�bw�'}7��I�����>=0�}�M~�x���/ �_"NC���"��)O7x�s>a����:�� �e����ʢ�䓏����B�^T�c�3�!L�"����]_Y�q؇M�������j�sHjbC�F�U#��ᾀN!� @4��}��?=7;�R� �$r-���8���Y�u���:髽���h�_�(�Y@p.!Ė�����v�U_|�%s�q�a,��s_~���h ����Ϝ
{Sl~���O�`.e�Aׂ/SjW��"�<�,߾qS�"��ib��\�AQ­�Q6���T��-"ȘP B���y����I_����+g��Y_�̄���{��~�V�{�t�N��M�I-�$e"��I~ @�_&x�:���	qWD�
���}���;�v6��wr���h���
ܲ�y�҇�1��b��Qe9\���!f��D��mEq5�������/�bQX /Ov3����[�"�Rީ�����2]���I���k��k����؋@i��p8-,�� �@ 4"�qQ���h
�����0jh��}����Q��̜��ӡ~ I4��3�w���š�-���ąL��hcm�6N9��
ad�|v�yNܙ�陎腔e��AN�#N�h�f��#Gս;�%�;�����y'��Q��'��c���ҥKZ�;�I�N���ex�91?�Y(e,��1�y�z�lN\�����P�S珞dOD�������_dor+?�9����o�E���>��/[�.�y9��j�/]����H��t�V�a]��Q�Ց������_݈���o�Cl�O?��kk�pL�rځÃ�̩�j��T�O�T�O�T�ü8�z�+<d�%�%|t�o�N�x9u� �;��MC0��[�9�3�z�ӓI7b�$����#�S�+-Y�zM�)sl�a�@�, ��W�Wt#`��%��A/��" �����{�#T��W$w�ﴇGv}?FF���߽}�E��$v�9G�n�r�e<����
�
M���/L�Y\��S�܈b�9ǪHQ�������3A*�;�8��T��_z�ꙙ9��ո�H��H[C:t���a=�ml�C%��T�9��>��:��`
�O2l�bc
���:=���y�a�����M���8��^G{Qr�(E�'�4���b����Y5?7�C��+�;�����/?d;mP��\n�;�SJ?�#t��A4����Ou���fC������z�[���HM?�Q��,�͊��e3�(�N�Y7`L��Е��ͻ�����aɇ���m:�`O����zjw!��� �+9�_�P���U�&B'�ޞ/�X�DR�(���(}(`�4׀�z���7�=\����؜�� �����Y=E���ڪ���I/ˋ+�-2H��<����܆��c�)�fӥ��l�$/�5{�9�5@7��+�F)�y�����q���S������;�RJ��+��l���A�d@l�fŐ�7�j��	��T�{'�9Bq�����_t�zcs��M����[�\c��ya��짫׮��ȓ�z]!��9��h��6)o������V p1�!��{�~DB	�"];�K��j�=���L�i��'�x��Ǌ�n���YyCd�v��H�_##�3-�3ԲU����a��-kZ�a�%;D�8v�kq���;�K���K�P�49�Q	j<�n`A��!C�jtd�ŤT� }��'�i=6P�ů.��Mݓ�����q\��f&2������������r�ȍ���(^d��E�A���t����Hv�
�#�鈧�?Z"@�{��z%+!�|��tp����� z\G+sĲ 2��1����m;�/?'�XR���Ν=�~��$>�H��q�E���eu��-����ν�z��o��5x�k�PU�`Ͳ��B������|_�:����@0�F�(8��d��a��s���H=^&���Ҋ�&�,Ǽ���������n�k//}�:�n?:�[������%��/~��� �C��V�27�,����aޯ,-�VVى�W,��֬W�no�����6u�g����0� gcX�J���=nI�Xlm��#���(˶w�@�0�^���X��"�4؁؏#^�܎��pI2#���o3�A2Y��B/$x��Ra��hѤ��H�3�#���B��	��,̀����K���[g�ؼ��ﺗ��ΎjGz����s�Q��Չ����h�u)�{�D�����$1};���R�$��Х�I� �7����,�$�{��Y.�RD�]�a:�xn�����٠��I?F�o���z�v��iџƧ���-OFi}_������~Y��L��ح��rMFu���Ju��+`�0�W�w4�<u���"�,���y��p�C/�j �z�t�5>_3���.�d��آ�x���u�X{]���^E��9�J_S2�Ѓ�{
��p��vW���~`ϡ�Z�y��J%Tx� ~��^[�}y߶���4�G��Æe�w��,��B�G7��M$v�{q�.����/����ifL����-�I|q�7<��_�9P�J0tޞF��&C���r�}��X�ýpm㉀3c�Jj��Z�
�ㄣ�8ܿg{���0;Uu�N�Ծ����������p��L�[���J.x�Mp�s�,�(5�K�6L����*�f�ܤ�x���A�9=א�Tjҏ8�H�}Z'b�=�����8q{#�4�Hj�2]#%���Hn�vsQu��]fB�/1Y��zt��9KbF���|B;uY2,��f�xRAe��B�C�!+����ʆ.Z���N�=x���栿�G>�ը��ػ}�bNo=�'��w��������u"bG0�R�i�.!.����.u�:��Z��&M�AW��p֘x��g��~���Q�d�������T�`��a�󦏽l�]�i�߽�~�5+~$%�t��d�IM�1���'�Z��R�]x��dV3zJ��#_���%]����N�w[��gWb�G	�p�GJ''����LI���I�g��]n�`�����I��x���O�Q�(��Z�nvP�H{���vr!��n�A�s�\�>P���nI���I�|��ۜ[��N�tju�m�V�/������37F�B�8�SH=��#:K���k{�vLvib����|��G�˦����ڿ��^�÷��şC��R�0�n���6��!�:]'��ҩ�V���MFv]헣KX��-�X�?�<�EN�q�����:��i���&�ef J}O%E_�{�摆v�LU�E�Ȍu�QG8���ޢ �A�:T��)���2� e�D��?��(��1m�ǋ���rS��G:�L��>W:��n۔���Z��`²3���E8>�gۮs)�y���̰���j�%��]�^6w]�u���]][fO<��U��_Ҩ��P���5�~E��Zv�I��X)��>�+���t�>f}T�[vF�2� S���8"Z��Z��PQ�.�q@;��5P;K��\x"�l
�@������B�g���ѩi�
��h�c�X�a��͆oF���F��%��{�g&!rxj�E���y�n�����`���k��[��~R��N��}�u<��]CƸ_D��$
Ӑ����h��/A�wy__I���r������"9Do��`�9:�l��d�8� G��Ԣ��V�kj~iI]��"����/ ���\embV1�#T���]G'��;���i都ږ\H@K�a�8���	��X���@U_ vP{%=�������sh�~���p�\�0Q"�"!�<+}P+H�*L��͘�˸�����n�ߓa*Ȥŏn��qЄ�kO�,����~�v��;�����fI��+y?�J��S��h1	�|��K_�(���B ̄�g:��;���o���@��'��"lr�J�#Ʃ�Z�q_A��R��-GWs@\�P �YI��A�!F&*�����|?�����ǰ��,��\Z̵t`�OJ̙Ik=�$����*�^������آE\[�dNì�,�:,��Bal;[`ɖr����ɺj��*��غ+'����z�x�h���vp� v8Ļg�Ǟ��V�cE'C����ͺ�Z��'84�Մj��V��t�8��� 	�L�)�tǒP��܇��R��0ՊwYmau�(�&< Jj��ڠ*=lfi╶��o����0G��bl�g;(}t3�#cHp�&M$����v����)�j����C`w�P�E����"�.��('E\�,%/���9nh�������Y@b:��Mk�;<�E�� �ѕ>�<g�%,�az�i�,��?G����o'��8��o�H�>�0��/�bs��p+JsطF U </����v9r�q���YN�F~�������`"l�P6w�l����:i.j[�ز���	訴;��X��eH;c�N�e6&��MD�Y"�X�����ǐe�x�pf�6�x  ��s~�`���$g�㓓��LSa�./��/��{�{�� �<�������V�b1k�H�l���gC�#��<�I5��c�ݐ[�Ʊ�f��QRȶ���8����.�y���Pc]P��������>�tI��E舸��'[6z<`�޿�N�9˺btt��� P�d�Bdޢ�r���0D�.�9:�l�(�G�ѫ�kSs�u��k��K�o$�<<o_�v�^�M�����Hw]�ױ㐳}U�33z����_��N(����/�q�A3�>�X�E�canN��?�����~���d�������^����g�XE��J��;���{����`���GTtrf�fdIo�ݙ���?tu�,�S������n\��N�QX�B�#ǎ���y�M�lT]�����2µ��I�8��:=����=�[,���0*ȏ�����b�Md���c�Tl_'.g�F=ic�ӳ���&�cwk ��N�����c//yW�kOD;1���n߾�lz �� ��g�'Qu@���h�Q�E_���d�z�g�&T]���6�DR��4��5C��I�6�NDa���d
D!
��"V�w�w(I1��k� ����#�"�4!ypK
T�q�kz��E�]^��ӿ����}msC��'Os���F����C�>,z�Q�a�.���G�i���fak&.��I'��s�Q��>nmP�Vb��ej5Ҽn^��Er�_ᆽ��۱��\lq4�\O2DY&���.]]����Q��J����gĦ����g:�V�� H耍�-���'�|�&�@���λ��G����;j��u��5u��=.jr�!qӘW�ǌ';4
������g�|(r�${g�Q�Gs�8�a��]7i�\����$�0U<ц�����Oa�ڬi,���N���ڻ�임��!B�C��"��ὀE'?_��3�b [�ݙ�+Q ��l_]��vБ�����	�����έ����+���S��nEf�ݠF$��Iya����0���!���yp�DL�獌�m���j=���.��msi����н�����%о�
���nGO��b�%�&T�<�L� �HG3m�ډ$��=�����f#�z۝�
.��^�꿥Ŭ��
�ÏLV��>WQ`߾yC�I���f8�K^]�����8�֬��sU8� �n�#�8�1��믲~�&�� �B��s�Ë�R�����W������#�<�1C��(����~�O�n=n!��tN�t-����ݙ�&�^�݄�"
���#TR}��L�b����{CÃ���i@D��c4��u/�����Ut�i6+Z�l�܈-�(�mӶgD����I�#��YV#Y��;��Bl���窅��='�`̟�\�3�\��2��5Sp1��i�����G9���#M�ǁ��,U�N�a�5��B4��,�c�TR��� o�!�E���SD�Yќ��\3g
��:8�g���`���h����#��O/�Qh �`v}�mL�H?� 	�.:��|ҕ���v����vT�xT��Оd�������K/�����'�m҂�c���֧�S07������hL�����,�)AmOW�=�-F�r��I�ê������qq�]�w�Q�uO�qQM]�~��P��54���@c��p{e����0O��:b&�%
N7�?�xң��y�����|yyI}�ѯ���ayi�!5�HH��(��!�-�;�9K�"rܖ1)�K`�q���&ۨ�ۑb�{��R��y��.����w�pu"1�gX�l���.R���#V�,�2:�MH$Z�D(�����í���T�6t*f�{��I�tߊ��t讣�zU�Q�.�mWL�{
X�!����{؃�l�@Wȣ7s�gB��-�yވt���h�?��`�J�L�c�P��#���B�M���CD<�/InWkɸZK��x�S3J	�p.�U9���� Qgx|v����~�gÐ��].���n��݉��뤯��7o�$�����
2pL,g�ƚ@����C$���F:���, \�i��΋��j~q5Q�;�H	�H��j�)l���I�i�ϳ5��m2��=*�syz�����^��gXB��?t���D�NfD��Z!�)P���v�j'�pigl�#͉�sI|�7-?m�8�vd�pG���#�I�76M�z�̡�E��xe��Ô�ƢK�q��*�g,7�/�#� ���qq��s��	�8�פ|�0�/8yem���:xx*��$́����q��sȮ����D���]���i�����ЈK�~L�cKg -�kȊ�$T..��$���9�����Į��������R^Oɶ��(��NBR��ֆ��d����Ď�k0��L>�N[gؖ㑲��_K�*~��ooB��Q;Xh�n�M��9�;����!7AF\��kG,��Qi�؞���VR!ч&#�J����E���j�T�'��'R�@_L|����F"뱡j-�!8A�e����Ɂ�lI�pk��~^+]h��	E7���vw2j�	�Io�,$ '� 1�vM�А�2[���Y����$�5�!��a����g�!�ͫ69`�'�
B---���!�.\��7���2Ľ�ɫ�W&@
��or&-G�Ø99<.�T]����S�cr�lX�'�*:�ku�N�S'@����Jg��SB<��o���bf� �P�)�1��*���8�G*��ՙ�ΪW^{�r��Ok{L:��#�	�ʃ@[��Q��B�7���� :M�`SGl�`p�n� ��R���#2�d�t=|B��{d,Qz�g�+Ml���Ń���ʬpz;L@�zU�:��\g�����w�<v\H��:X(x�F'�����o~�a�!�w�[s!D�c��+^�T�U�:`%"+L=�k�$_�Ir9�h���0l��Ңl�����IOL(�0{�����F����8hM��o}K�Ew.�sQ��$E���4�� $�0��O&Q����ߘ��	\/|z/��ym�zS�upfp�T圮YN=��1Kq��+6�M� ��h B��S�I��D±g�C�Q{Ǣ$���h/�"��������Wo��������626��.�eN�y1����s+6�`yv���]�w�	�ġB����>P��	4���Xp�wET����WΟS���k}e5��d5-3�׈�tb����h��Y�l��d�uh%�Lh=*;�ӆ����ϡ��A�!�
��Xч~��Kǌ  k��7��[̰��C���2}oR]����u�
�h�M-]�����;:u��3���j}s3�Ԙ��A��v����_�>��S4u�?'�a:%L�e�Ԉ%^��L��3r�X��aq�i����@��=��	:S��;j�M�,v�@+p�&%ʍ�?~��f���{D7���*ു�����s�E
�ʘІo�#����>n��G�}u��a�l}��~x��JCw,<���Wձ�Ձ�	}�B �T]YYfW��ʚz�ྚ��c��,*e�^�@�!���l`�����2eްHo�)�+�W#«\�
��*W'ʊ�P�#�p!�f���o�h*W�'��@C�p,z���F_��1�e�ðk؍�} u�r)����/�xXd��h2��V]�<�V+˫ܲ.�J���	1zcll��F����༁�~�%dPऺ�HY��q���J��
18I�vZ��H��ņ�kj�Lt�*�5�{����?��o;o���7�i!�s�c�� 7o��e��q�����_M������@_��Uv�taˈ$�A,K�h�奋I��rĖj�,V,\>���ۑ'^��u��l��f���bY�k|�fT��WE��,'Ru����H��I+����ߝs�x��vv��|����A^�cE�̳xi��HG!�
�n�3Q��t�q��-0\�>��.��8*Z�7݇|��A����Zޡ�2�%��;~�&h�Rl���$t����6��,q+L��紾0x
;J�}��m#Ƭ�:��>���U�f���B-�.�'N%Ę:4�G� QY��[��y�ʥ�_��R�+��H\�=4F�	67L��`<$���
�=�" 9�E:~�z��wԇ�q�]���.���r���,x`죐E>cA�r�$��F�!q*`�Ls+}޽���I���}])�5ӯ}�;QZ�#LX_�PC��Ȩ-�lS����h|���6�%�
�D,�a��p�:x�o$��2<�� �L�OC�.�����f:6��qz��n�Q-ƭZ:�P����%��IR�`�a�%̄����u-�u(����?��^E�1�?��(�%�M��v��!�����[���͟�H* l�c�b�T��}�9���7�PgΞe�s���픣Mq��)u��Q��|p% �V�����C&���b�k�s:���1m"�
�pk,�?��ݽ{���x�����N�I	��Q�����V��u
�J����~z!�41$�	��Q�!1#]٧ �\�D�$1t��<���i~���>a��eŸ�w�yG���k:nĥ3��-�9�m���F��=Z0���fף�hZ,��W�6>·ȭT�yvb��>��<E� 8ʶZ�7ivO#]R¯�7y�/��H�6V�s�Fص�Ȧ/�����]Yl\�u��2g�n�E���EQK\�V��Pe4I��(4�C��S�`������'?��@Ѡ-��~膠M�M�cˁ-ʋ*Y������e�{o�w���s�r��H�M���pf�����쨫E���I������U�TpQ%���f �֡t��ڰY��T$�hvzF��λ�έ���g��N�$�S��|��(ӐE��*��r3�W��[�
=�!��z�� �P���n������vu��i�.}��9����{�N��_J��y�lZ�X��qP�h�	�[^����r�#$8-�Z"��&��yr>|�U���Z�0}��h�_��5��?�W�ۦL���[���P.���G}�j�M� �z"�<���)�8���k��YDMU����]B�Ԇ}�ǜ�s��ҁk߭6ح��_P�O�hb���B�qc�7�)&pO�?<���� ����{D��BPP#�T!��ۣ���������0��;��2�w&wn�����m�a�5�e�!�v�B/2����	���e!��/��'�0�\$����-�`���L��I{�pܶ	�G�6���z�_O���^Zd ��H��1:&�$
Q���'Dgw&j�U{@N�?Pٍk�ʤQ����b��_�p��a�`�WV��) G�b���D�O>���F���ZY�Ĩ��u�P��j:��{9ЦD�d�� ��ۂ�C>M�i��r�qٶV5P
;]ٙE7d0<u�z��M$\�o�B8�롂��S�P��>�C���i�W�^�遅/�Mk�^�8�����j�!��x��}�6s॑/8Ekmu�]Mܔ�0da�gq}��[l�ւ�A��%=���Bw S`�A�9��9���LD�!�8��^ ����Q���Gq9)1��6�
��A�������&�{���a�67(�oɴʹ�$�ϝ;���3oA�~���;�bmu9G����Y���f��	Fm�Z��ߐ�#N������s���6����¢�s R�����F�R�"s	���]&�=�O]� p��{0u��G:�F��B���S�T�F�zӞ���c$����з����kŒ�'��#.(���U���r�[��F:�bejrs���*�+<�u��]Pk+��L ��7	���i������Dy�u�Au���g�s�CYe�B�P��|�Dٿ�(餬jDb��k쒂�e-/şit��dȰ}0aɆ	
L�y֖$�&T��A�z�%ԄV4���smn_x�(g�5��M�w��>ڋ*9 �8�"XsK��{�I7h^��"<hoS����L�l����sq �"�n���ҍ��H�m���a{���s}���K�<�aѬG�ZV���P\c����Y��m�,���&[���t�-�Q#��D��ste�������]ny��j������hCӬ|�����[d���2���sS���%13>y�sd�y ���f�[YGtЦA�$���9S��֭11;3�i�1��Ј�����7���*�J܄QN(S:]���D:��-�g���Þ>|�k��'�o��(F���8�Æ�����Hj��+���KސPtl�|�����j$Þ���"L����f�LLN���#�$�׈X��/bc?m������N\6��g\��=8�0��2'�?��3b��1�	�)t�����d�^��B�U�&�`4��.��,ä���6��ϖW�l����>�I�	6����c�A�9B��;��W�q=���,���+�*��s�c1��pǖ0���abh8$8���	�M�,�2�Z�@�d3�&�����~�l䢸v�:���씋\��1����ʏ����Sb���x���#CC���26��+_q�x@��2QqrC�B�2:t��^|�q@�ӧOsJ5l(D�5aT�:��=�d\��0rw)�F���aoB=��	$d���� �#O�"�@��ݑ��,��nzܽ}G��?�3��Γ�_�1SlG�Rry(��k�H�`�� ;)Bbs~�	��p�Ϝ9C"2#.]��u��`n9�iӶS���	�T���q�l9�N�Z{���'ѪG���0���>�pw��)�i�b;
��	����&D��j�ɶi(�4m��8�`�}P�����c��C&WV��w"���"Q�E��pG/�ƨ/A����+�W��#����S�4�bB;ѲJ�f�×�t&�B�em��	�ԋ�:���!�̊*v G�\.�фWÿL��.0".6]	U����� ��Q9�*
>����/�ز}��ܐ
{�\V�r8<���ڣ���x��U7�^!O�����2I�8 ��[�#�.���i�V:^�!��"Y���s@y��{��02D�&@���a�u�[0�C�5�
H���*�q��~ћ^P��\=�VCd@d�b�3'�Gdw�t�s�뭳��pi2q��-y�����0#~b��7���{��"�9C:᭷��ĕ<�,����-���#��ƛ=���!;���Io�,c�!Q��$��;���'�di���2
m(�gTu=s��E1��
�~ч"�cҿ�cn$����
�A>�6��L9�Q�(�,�t7&I��$������r� ��.A�"�����sp��G#��)�)b���|��y1�`�= �_1u�Ó�5(Lq��䄘��d~��1��[m�qT:���s'0�%>*O���;z�]��tF�ᚨ0$o&���<���)�Ce�^%B\����"aY�����!��*�3?;#���?�e�q�&
 I�$=��V�I�7�EnaQ����\�I�;�)a����BԍOM�_c�
t��BT�,"�1Cfߺt�5���nS�kc_�������wlw��V�w�s:�[g79*T|��q.?D��^����6)�v^���i%?�[��Ns�(�8n�H<)�;:���A���Tj�iTgFi0�.Չ�3,ݝ�/�<4���66[���D�Ͻ�������L�B}SБ*'���*������E�X�4�;;U�Nt%�{��q��b���-=LUp�{f |�wS的t�a��MQbmPl����A5"P���hinү�V����@��1���P�jڗ.�DD�Ϯ�0���t�?6j���_%Czמ�qsHt��9�9J��ɬ{�����Wcx�L�z\U�X;�j^^�s���?�+�����-TB��Gq	 ��]��,u�/���_��uQ�����g�8p���ςm-|sd9���(2��1j�l޻�z(����TW5�6�L���ح�]�*�낺���JAC2(�bRO��^o���.�,(��fZNY,�$��3��m��^���|@ &��'�tȮ�GM� j8QM����k�th=�dF�j�D�z]6�� b���Mz� ļ�zEރdkV�3]93֐@"�ٚP,ZM3���P�}�RI� ����ȜzD�h=���!��&��/�T1��$�}�A���Zg�g���Pp�����k��zo� �fB�)^����ʶy�:�:�f�lp����k����l�Pt-b{8A��`(
���J�OYYoNЖ
��
�gz�0�����kzn�Q"*Ǝ]Y$��˞�4�%%z�
�ޟm�`��.v!	4�rE<�z2|���_m1'�� �֔~J����-3�*,��:[:эu�米��D��.����\�w9*| ��^CI7��]�+���F��wՔ׭�s�������S!<$}�4�� +��Iݤz%��@��[R�%��"���kqj���Ϸ"mET?+|qg�5hb3�q��<����`������z ��ZB��~��.�:UY�qk8ٮ�C$N��϶����]F�J�$�VV��I��;��D����z ��h�.t��|�:a��&NČ��z�2�n�pZ5o�������s�]�����+�+۫Emr�`�#T��������BB�M��:@;��L�,��Ujڔ�*T7l=|�p�z�7�#���"r%� .�,:��G�˞J��J�IW��:�w=��R��\K�>����^ĨX7y�:��W��U�6�]ɜ2m��̊S挱�����2�H��l#���f����O�9��oD� '�W]>���H��Y��J4�aBۃ�����,K6��b��9r��Fn �>.n���8������h4^�<�����R�9̸G䦈-��/�$�۲�jm���������H��?G�I�0P�j�B��nNC&J6˕���P.�?W�M�eI����G*Mn�Sf�Ok+��,md3+!f�e�w_L<ӳ3�� mN%)B�!ďX�feG��.�k�e�Eʾz�X���&y>	���].*gp���O�x�I�PB�U�9�.$�`3!��!2�@�����m>p��(�A�[DƧ*��(�"N�ԜL�Ņq��r}p:N�k"��$��-����8��,����(�B�Q;�5���Zth#Q�%!�2:�%�K�� $�������v�X�Dpg��O]��X�G,,�ʾ�6���W��&J�K����� �8�ey����"�Е�rπ�,��F\��$��VR~(��s��p�w�����ݻ�;���������m"�_e[ʒ���
��m�P(�����Jw��ꉼ��6�W���[��~���f���#��� <�ٴ��稄G}��?����@:*�!.c�$�e��,�	�ۈ��<6h�~B��=��2B���W���Q�h��={���� �}y�,��%�z���,�Ų7��ېPX�L�'�d�^�P�3M�z�^�5����aT�f 锭z��9 Bz���U�]B����F&,�xmJ5��*��Ŝ�FU�X6�������T <���t�,����<��i�	�z��Aq��A�O��YG�B��`��HinJ��~�^��G�������1]dP�L7[q�MQYi������0���-���w��������ҽ�36�sX�Lpt�ΰmJ��t��#��V���)k~<N8ը�'��q:��06�����E�J5��P�s�<!�j6%�G5�X��4�ySBg�+}���'羿�X�?kE���}m$V�I�o�z��k�&b�����QD�=���u�����nJ��B�W+/%fg�� e������y�;JYWg@J?�7{���	`0=�@N.��)��
��:��/ȁ��&ϲ���j]�K(�T"�a"���J����^zJf=K뇰�Ҡ�е�Z�0�&��V�{!q�fWiUGՑ���1�Ι���޾}����$�ĸ�fL$�������� ����f	����dB���FDH\"gH�$�U!6�� �!�	\�j��h9O�����ǏO���_[XZ�Gx�_��a���	� a����?���FP��<��gꮔ\�g)W|o��($c?���k "����v���"2-�2M�އ�[虲J3�&��'³��t^��lK�;~�H����� M˥��u�n[X[��c�u�X���0/�͝$Bq� D�ί�_(̓�饟�D4�OC�#|f<��N27���q\�RO��>@/�\~�`�S.[�ް1�K����ؓ��e�K�5�L�1��A��4�g�x|6�<�0��p�s�`v��H��@�~*��X���5C�� "�`�B?e��Mfe��]�/2��?�{d�:s���?��Ϯ]���O����[���v�s3�t�+|�Cd���#��V"D9:!{�'S���1�2H�R�����wH�_��MjW�=Bz�B
x���#>��#�C�ufq,!��T��ݖЊ[U���=n_��������hN�X�A��cq�� z�c��A�O��9��,�-+�1�%�b҉ؿ�����3��w��Cu{�O�����_�/.�dyr��mm}�R�L�L�UP�\�$�&�nB?csP����s���G��'O�.�!]x��7���<��B�GI̡K��	ls�eH7R��^~Uz#���+��˘P����_�ϑ?1$�a��S�H�#�1-;����x�L!Á3����d]�j�N0��p�|$����ή�s������Ж��Є�z�F���7�|��L=�~�����6{�M��� yqg-�p=����
F�Ai�ǉ�.|$f�z�1�RN�t7�f���Ԑ�k$ZP���Қ��mX�����v��<����d*ɳ10*��8�UbT�	��N�Zޱ�7���s\�@����Q�/ax����2g�������@\�Ez����r��������w'���$�vD(�?=M��{v�~�����������f����?H��e�e<�JP�5�#����䕽��1/^��w��fk>��-�;F�f/���[\��4��uɷI����@���� �uuf� ��b��H�n8�j��g Q��ׁ>!��܇��ʃh���ȓ}�X  �<��P�_$�����方����~��o���������^z��o�����\����\��ح��tcC�(��&d�OTN� ��4���7B\���A���s�+�N��"b8p@����2����f�-��4��zAǁ
HU.����(�*�㎁a�-��0�9{��90�q^D���|��6Ў����,���y.q��f~��+:���v�w����~���w��;�u��Y��+x��������O���?�8�æahJ�;#�����`8�"�bnEvq!�k�AYd0��߻�����H�8q�=���CFk��l2|^5�Y��!Aq�o.\��PY@&7\�O��ǟxB��!�G�#�~�&� �Ӟ�nvE͐X���!�.��|ANe���.a�wv�_jmk�Ş���9qbV<��cB�+��2F?�^��7��r������wr���B����LmN�6 Χ�6-N��NF�с#L�R��RK�:Ć�9l(zF@aOL<��Z��zC�d�F(����.բJ�ŤSu&sy�i��%�$�pmm��z��� ��؋�9&+��PC�^��dƳ]�_f�������spp�����x��J�^xn�;x���k��o�{w�gjj����������0:i#S�x,���h�7%R�):��A�����E����ΈE}1��x��6'_b��ioc��u���	��"��	��6PAHn$��-�#Q�����s��LK�e*ٔ�ߞI��;�}��-9AfLA|C�!Tp��⋀O��1B:���^j�?7ז���'�$�|rfvz���u=��6>%<3J�d'Dh�,�H�����@#G�����WU�$$�C4�'��e}!�+z���X��d.
�d"�iIϷd2��'���lWW�]2�G�������sϝؒC�Q�o�P�tڲz��~M��gf
MS��:�V{k��=�B��Np+�^�Sv�{��WF�T,�2�H�KX��l˳툧�Qxr^�T,����]Dw�J��Q)��%k�P������b��x�i���T���&ى3{���e�����vB�[�!��}q���N�36O8���Eʳ��B�-�	�9�Ѽ��<� �K˶]��Ŵ,��J��.r�����a�K���$��J��L���#DY�����[A�͖�[���_]�+��K���t�`��6�    IEND�B`�PK   Ŧ�X���j_  `_  /   images/43e0edf9-5f24-49a3-b78d-83485af402b6.png [@���PNG

   IHDR   J   �   q�   sRGB ���    IDATx^�wx��7~g���^��m��^\��$����$��-	��o�|!		-T�)6��n������}���{��^�W��}��_���ciwv4�S>��s�ߗ"EG�� �_�
���/P
Px�%�������\.W�^-j\�{P�rϹ\���`p:�Z�ˢ�h�N���ʡ҉:ѭu��N���	q��ΐ���`p̏�G����^�5.�[��B*�Jp�T�(�A�V+�"�?�NE��t:Մ� �QԉZ���k�n7����o!��������)��,9�%�+�(]�v�6�T��Tj�Q�p8\�cF��[BBB����'�V�6��w�ѸL�&�J�r�/�ifg�����`
0���wt��Wxh�S��;4Z�j~nN�t�Tn�[-�.!*�R	D�ֈD�":����]�FT��*��Ѩ��F$D AN��h_XXp�Lơ�ʪ����>�y.��3P�ox7>.v:&6�ob|4��L�J����r���� ���Z-�7;;K�v;��V�TD
�t:��fs�N�K�պ��Z��p*�J%j4�V����H����A܂�h�jA�ӊz�^��'���p��zT���.��.
�h�������:t����8""¼�@��h -��_����z�N����Qj�Z�r; .^z=wb0��Ą<�I ���@���yx��v�po�Z������ ��A�v�J�H�=�#22�8�vz=a�!�I�I/��������y�`��D��/���Ё#WE�Z%�������A)@ H�
���<@��V�=R �{����w,0z�*��\��RQi��-,�Q����$d|bt^P����s���1�+
���h��1�����njh�l��դ���tvv�'���������<7�  �KJ�*���F��=���M��^�Fg�.������I�{:m�A�{�{�FW��ٱ�3�Q[�>�UT���a���K�Z�(�(x  �7���z�j��K�b>�N�" ��TZ��t�,<<�$%%���b���j��m�o���{r3�!ˮ���^�_SS�M����ܹ3��@���������@��E`Py P��j�_$�(�=��Y �M�4�O�n�t�{N����d������:�Ѩ>_����M�ٝ��B@��f�����T�®ήo��ϗ�@�����Y��<6% CB/�OA��y[��S�����ޑ����=�(���O�L��ד5kS@�{���+~���� D-(�&v���D񨶧�t�[%d454����^�^MZ[[���	�a��`�7��@�T���Z������d�s0�T��>h��Inn6IO_C�&C_Ey���ܨ�DT��@�Y��\��g;Qw�=��di�:���L�vbw�����:/Q�/c̃��H����Nn�x�AiB'���F���@ge�?��.����
���3afa.���������� ���N���_$N���N�<��-<H�=[N�x�$^��=��R�ז��Krss���?X^^�pvv�k� ����Ewuu��8fz��}��7n���������AP���(�zH�(�*��
ԙ<"����UjF�G�Y����/����׮��X��V���ڞ����ݏ>�u�J�Q��G���,Y\����!�pq��B��%W'� ��%�[b��w��y铫��j[�t�����]���l�ɬ��dff��z��FEJ�1�.^U[�w�s�ӳsiikHgk7���!�[��� r�&gپ�R����o��	Hx���tJ8��v�����_�tM�Ʒ!dT�"c.�%<��}��;{6���&�'���Y�X<L]>�Jot�裄ɥ�W�r��xPѠ��C�9���a��@���[�ܞ�UP�$z>������~��=rmNvill%C�a237CO�O�5��
]�rj� �R�,��r�ץ�3�����deeA���l��m�ُBCC����� �}��?��[�ޒ��G��?H&'��(�<�D���3��<y��y�ǳq�J��̛?�/��:�DP����۽�G�6�?l�| ����y��}��HZ[۩D-Z���Z��/x��/���?9�Q�q*��}�HEE�(�F��������/�wŁ����?�ӿ>����5�������Ä́�W9��u1�Nh�����Of�`��ǃ��U/55�����DY,˱�}�-i	i����^cc�nll���_�Mkk{EFz��3���J|d^���ST#�s���a��Er;%WK���>Đ��z055�h�ۏ|�_z�Ƙ�W,{ l�޽������?y`��KM�@usK����Rv�pS� �?�帔8_ �@��!X<E�も(�INN$���$,,d$77��ioDF�w(&&J����l�'>�裫C4�ݤ����y����Qrc͟�+��;�+��V�A��ˡ<��v\q���ee�(��e+x)JEUWWK�ɓ'�����i�I_� E�@2��⍽�Fy{şo��R�&�������H\T�A�
�պ���=�c�s�(����N���+�ݠ��u�M�da�Bff�<@�Ҁ?�]�/c�ߓ{�3�(�k�@3������"z�v��������W<�Ž�����G����������H]��2>>I��(P˽x��1H�&��r�̓$'�,:�D�]��������ྜ��'��S^��9Z��F�{�j&�&��jm���^��h4�::�H� �G�nV~�o�/����>�3�r;���_6
%St���ei�N"�K�eeeP�U]S�`vv�NA	T�Rj�4��IG�<y�����F??]gG/-0`.J��"x�*�a�JN,y{�p9O��-1�R
��~_Ra�^K��gVV��h�k߰n��̜�]� X`t%�ꮮ���Ύ�_��w�Z	H��1�S���Ln�y��?��|���B�����$��񜼺���Mdaa����ʜ�A�e�����ql�(v�6}���a??��������%?-_�O\n����7����'U9��UU���uj!AAAd͚4����2��[_swnn�W=������Gܻ����j4:C_�2���H^5xіmx�+B�P}��3�{N�KJ��[EF:��?.���L&���D	gPp�9>!�����wCO���(�S�l\����y��?��Y�EGǒɉ���O��fOSs�xp0�ؠ'H�'��c���CP5*Vq��������Nk[[k�w���߿����2��N)jnn.��'�����͉��BwO?�(�Ԙ�K�<<�x(Y&T�||L�D�D���������y4_/� � (��3��R�92:d����r�=�gg4)U?�@AG�s�=���o︲����������D�=Q>W���{��� @|�G�o7a-D ƍ�X�J�H<K��]WIQ!)**"=�]����O<��m��I �ʔԽ^f,�w�{�_��jbB����AK�v+��7S�s�j�CG��x�Uxp,J �R	@�zB� ��1p���R�(����S��{P�+(��z�}||����|�δ��c� 0#y�׹H�z��}�.+((�N6����0�%�|x������7l���ru��Ҏ"R@ ���R��y�{�p0	(��JtLL�bY������ӛc���v�)
b��顸?�ṿ8xtsQQ��T}"V���%_���Sp�p��ox	D��*I{�B���R@ �l�)�X��OV�{���FJ�덎;�mW_}�*+��R�������~V��ϛ[:֧��V��h�6z�v����TU���EON3()� P �s,��cA_��n�Pi�*�6�e�f��ZW�|ƚ�SSS�Z%��ft�?����ڷ�~����i������'�ԕ�s9�AJ���A;��d���vy�9�6Ƈ��ǂ|�J��IA�JOO'a���e[R��|"(��\�͈IR!��w�>u���w�~�.B�@�0���m?��z�?#���y�ÎP1hoDc*����%��  p~���6�Jק��.j�!��Tp`��m���MOφ�:#q
^J�RMN���:�����x�&��O���C{�,֥ޕ�®8^"�<���S[��qx
���g�a�
zE|�0�;4�wҥ4KPP@gIIٶ����+�%I�zx�cmGk׏_{�͛A���� ���0|8���O��w�@�G�� �z|:�	m$��@��nRb<)//��***y8**��d8��z�477����~<?��"���da�J��<\A�xu����$��"��>s
��P�@�����p��?�z555$88����x{^^޻�#͢2��W��C����ߣV��<`dMddi{3z;��c���̝��h��-�޴�j�R�۲�z �gee��h�k[��z[zz���%�233�t�x�u��x�~�S�Cfzf����Q���7�Rg�(_1!/M<PrG!��'M�b9s`敕�.�VӲ~}������·D	#��I����������̛:;{��������"�M�xy�����X�GPxI���GҶ����N�i���~��� R��#�ٜb�9.��o~�k??�qxh�ttt�{����V����z-����灒S *,,��dgg�������*����ޯ4s@�
A��>97��Xt}��7ߺ�bqG�����8�����O�L�WET�z����/r{��:>F�C�%��BCc=��0  pgIE����V���ݻ?�~�O�>=7�P��[H&'�ICC#�9g��������v���9_�k�S:��.O����z,���-��x���K�v��*�+�(����#���7���T����LLL��E�@I��}�1�$
��׍/���$�I?���9���AG)@���Q���t��-w߶fMV�Rϧ(�p������Oj�YZZNZ[�I[[;1�h4kNx")�Q�I�&r��3�V��A���Ͽ'��*(�#999��=�G�l��qq݂ �v����'�z���w}|EAA	�7�������^��tʯ���3ly��Ր�����z��^d@�ff��f��~���OIIoS�P��m}{��K�!��(�z��b9�Z�w_��7*Wk�d��`�@Ch$�J��i���O4������D����ju�ɞ�ԯ~���PeNN�����(4�&�Ln|��"^�������E�xlT~~>����t�t���+)��0""b�ljGϧ䠣G�����o�۷ykyRb�jpp������ �����z�o��v�l��P|!��>H�/��FML���"�_��򥢢򷕮ZW\���lx__��x��'�gCFF�HwO�{CÃ��>����y/M����}����L6��r�|TZZ
�p��7]p��׮�ܳ�.lx�'���|�k��v��.�`acSK3�Z�4{p&[�ˆ!PhOPbx־e�����Wm�Fi5*�e URRB��������ͅfewp�����;{���c�u��*��0&�3�(�%�a̙�;�9���Й��<|�����"P�INN&�����j��,ߖ�I�4���(Q��������{�~����&���Q20`��K�|�^��x��E+�C-����ӛi���Po��(,�f|�CB�zJK˷�:��]]!���pzSC�O>���f��4���Y��X^�1��K�|˫"���M^-���ߗv�iT*륭��-=��E��q>�R��mki�ɧ�~��ؤ���Hf�-�Q�&r��̙W/�t�L��r'p�7�L���M�yb��K���Q^U��0�����sQ=�3��6���?�~zzVj7<4�d���y����0*J^<��o���9R�BRr��,w�������m��E`��gQD�R9󱑱�_~�??��Z菂���$�?��<O�I%��K�䡍/�� c�ܞ���;=c�p�Ɔ��=����@Q�w.����Y3;;}�o��ea�����#��r	���'�_����������J��FQp��_fV:�u���5TW�l��M�vzs�2OV�D�w���ݻ���T*�axh���������g�zr~����A�c��'o�P��[.�.�t'�JM�EC�����]�k�UTT퉊�J1Puu_f��������sCFz���p���zI����r�|q�%��=��T�ȾX������G6o��tww�OL��_��k~v�P�7W�Y}����er�j��f��d���j�<IJ$���u\�.����/��^OK�|��j�o`��G9�������z�k�fC#�"�~.@����~��K/�ZPP�3��'N��[��U�/��o��9_A-��~��Z���FALF�Z��i�٬�#G�o{�������9��*=PE�SO=�;�]VV���Yff���,��x �s�Sn{xi������������JES�����[�{����RO��U��x��^[{evv��~@��u�g�b�B^�%g���KU�D:q�~�a����`�K�i���Z�'�[�����'7+�H����v�\ҟ�}֎uQQ1�!����iFC�1��S˽ ��Og�^�����w�X���o��'&6�lذ���fKKkC�E^��W�z���^��h�"�� �����Ç߹`����4���F2a��$O���m����xIC��E�z8��R���x$*44�����F��1�*:|皵��I�Iݟ��w QaaI#�#?y��������?�N�j$��3�蓖��/�+
A�K/�yE^��F����ǭ^�Jǎ7VV�ݓ���w��,��8??3���g�˯�z�¼���Γ��f��7��i��9v��7��:��	���!�P/f��)I�`���m�99Y���o��P�`Ia9t�(���J�[j������~����	���Of������Sȥ�l���\�x���<><���LLL��Ln����ks!�[q�Tfso�������x���c��bq��SMd�a|�v%����4 sr��c��E�R�p��թ��.$4����t[ff��(Z�p.�2����N�<��o^����Er��)▬����������.�OޝM�x�)���i�b@��y]M����RH��t*x�fh(>����}�_|sb|Z ��ob�-N�ž��Ao�����9���zSy6����
��qq0r�V?4mذ~{vv�{�A��j��V��ut>���ګ���ԝ�ݴ}��`�\�C	:S�Mn��(����1n7[J�'��Jk��nb0��H�K/�:����������hv�9��^�ٜ�:::z���?����� Z��������� 6i �r6�K�|99sG���yg�1	��{x�V���Қ��鴷�_��g��Q�
B�w��f��ᑫ?�h׽��&0�'�N�����K��n�1f����9r�����&��z*���qka��cɺu눿�_Wqq���̜����0J\�K=�356�����Oԝ��444\?;��<_�K�(-�<���_��n!P|��P=�;8���6>��A�%%E�Ok���7_��6���l�N���ɿ:t���ZX<^WWG\"�-~y��c�pp����UHp�?��<��I�wb,[u���	)* 
�b�Ͷ�������ޓ�_rT)EP,Q@:��׿>����q~^����inn����Ş*o�Q�+�"������E����	��X �L�W�|޵�𻟞5�A�����,.����Ǝo�z�mII���
PQ�s��m���37l
eN7H�*9Px���yiA������y�|�4z?[���š�����"����0���	��������!99��<���gϮ+�灿l�pA������Pz|����}�8<�>R��ǅ���
�ǎ?xP�r� W�    IDAT���o@*���z�upp���m?�9!!�RԨq.����+/���������B��梫ԧg��x=9��Y�p#8�D�?�9�����>D�a���x~u�Px��A3� ������{���]ii�JKV��������{>ٳ���/7���QC�Ta`.��$�WG95�Y5�����!��� ]i�I�^���#M~$66�TUU��!��Ȩ��_�ڳ6\�sE�jll4�v����컷��u�V��.,���cu��|�(����T��Bi�
��ދP� ����9�4(�}-�\3��{ �����e�]Ke�#��_(.,x)3�`e��b�nd$p�������ޏ��s����K�v�	'o��F�FQExW�^��R=J���e���㝆F�%3J#$��3�ʅ��r�g�w�[W�5/���ƍ��VBK��gl�=wpt�O>��FsS�zq�I��ۉ�9���s�n���Y@�7��w�
t� �5��������I���w��Se�' Q U���tυ��2�]VU�����YV�?jl�#opp⑏?��jsS��;�׳��Kt,Ym�/X8�%�,7�@2��B4���PH,��r.
���\�	�f
%�����INJ %e��h
�-�.y����|�n�C��桱_|��˚;�m�E:Z;�[����;��h[x5 b#I��*�l�@��@���](`q����&	O�N���V��?#�d+�z�����ёG>����-͝�iq��f(��-���%
n�o������F�?�D!�|���#���G7qK�'5v(K��^k�$-9�S�������EE��9�wT;4d���|x�G�|������n�
��ܞ5�K�xf�x�ī��Ѷ8h�q+&��d��B� �ۢ��x�4��
[X�S��INJ"ťE$ ��SUU�pqq��hM�B���Ƕ}�ᮯuP�;�@l`d�~}�Hx֎j$�� *�uCh���g�� �����5a����&�쐗b!ӝ��L�+Ja�AgEE��K��u�Uott0kbbl��;?������v79��H���e�B�,��(M�˵�`�@!�h�S���N�ZVW�'ÿ� �+-%�TVV���ť��H_��x��9у��쉉�?|w��]����`e(��ڈ�bc?�����
�	U
�����w�#=�����eA�%n�I�T2lKT0��͙������2��iz�rҟ���zkժ�N%��\�R�wvf|���O}���W$����"1��\8H�?���v��F�j5���;��H�����<F�J@U�n�&�r�>-�؝N�*Ņdafz�i_<���]����M�H�rA1΁Y�w�{?��~RUQA\v9y�$�-,.).����n
?n�8�_a�w��XRqA$ ��E��!Z���m��W^QB�NM���'����RSSa~���3���Dԟj���[n��������F2�^�Y��?q��Fw�7���/��c���^U��6*�R׌Jt�B� qs�&�CUj�3���z0�fbttVC�����;�"#{W<54713:��~���s�s������&�Ņ���rNŧZ���@�ǩ?0t�b��$2�',p�Q�T��p� �tz��3�n����vV����Ķ�wŧ�B>JQ%FQ�5??�����[�_��`�3��75���-hx�p��r۲�2�<ú0s���v!s�i����[ q�$�[�@����S�Ewr�@A�fjJq-Z��;Z۞x����;�Vb6�j�&�zg睏��ѻ7\���NN�,n]b��� ��,�Jz3����ÀY9�+�	0
 ��%* �_ J-h������K�&��a$55���EbwLu�4����k��.(ؓ���h�
E@������ګ�����C��ܴ&+��L����Nb] �Z:!�'��T�.�G]��f9(�?#���d�wA� H$�v���4p��	(�D���VQB�*���2�sqa����RS\��_�����̕\*{Tk2��F�����ޫ�����z9z��,�h����9F�]�D��Il����&j7c�ni4�`*]�J��<��n��0�gNiM���A�ճ�Hqb�AM3	���,:�$*&��F�"��D%�:�W��&3=飨�$󊖫�����������ko�x�d��Z�G����H���u8��@�j-�ON�����8a���A�rjԔ�E7шrh��2��)�A!at����4���%&#�[�Ġ��6 L���&.����=��.�`�&�\�Z�TV���_��de��ئ�[���}�9���"C~.�S541�vlh�]�|~mk{����"ihj!��.�#�[TDBU�9>I�μFG9���H��N� 1�������b�C?K���������zp"D���.'-�A���f;����۹DB�� *��1u�� ��g ��1����8��Tee��S��w)�|.@�����Z�۶�;p��޾A�yd���O����A�0IC�"��Ut��kz��=�7-��U�LTtn7�	��	�_\ �1��$8 �,�/���iH좋���(�Z�@�;qX	�� N�m��FR5��R�-ml��ШHښBj�*�űВ�����䗲�����!�Ql�M���'~�����a���)219I���n#��9��DA�-�����v�L@�A���r�D�����t���9j�"BB�9����8A�T,3@ǰA��� nh Z����i�T� �3�?�������R�Sp��PRT�l��a��%�@�������-��r�X�ƞ�23�J���z
�(u@5�j(�Hܦ "�.✙�mU�h8R���̆hDo ��H`���h���"8$�5�-Z�R��$�w	�.,R)3���حj�U-86~7��H�)�@Da0�T�Tm���R�+ۚx��I���y`p���S�==�&�>r�8�HZ��A�CK��A�-��'�	gj�8C�j�g�vԇ�s���p,V�����ề� �X)�����T��@#�&���U�����P����\� T1	�x삒�WWܘ8��
�����<]�!���� ����F��V��71��/�VP�"���Pzs���5W=�CS���}C�1�[����ggg���*��� Lq8�a�D�i_����":=_EV�(�͠� �/�D��		%�E$(<���������_�*�^��䶵v��ԩS��Z�₍t��ЭN`๩)�D��R�R�X�/�F[��@JT����:OU# (�J�"Z �j��Z��� �r�K�ń�HlNQ�b ���5��I����퀭q�Ep�{��S��HvV1�+*+���&�j��Xr���;E�fki�8|��G�[;.ѻ]]S<==K/Db�f�8 ���4�8��N�Zq]BD�^\�o"�V�`��[��.�k���q�&PM���N�Y���3��1�v&�N6�R�:]@�hfTA���EF�թ��H"##[�c^���� *̯A�6�J�Rw�>�����]=))�QC����-W��
3�ƖUn���(�$0P�E����p�?�HTn�h�[>HX8d.�Vh�\��.'���zV`��T��j ��� Rε&!�N�_�۬��';���_\aͿ�Vrڏ�P?���~�UU�N=3�@��h6HE���E-���	b`�G�`Q�J  7��Y�M���[�w�n6��S�C�N T�݄8�RA,5����M�h�0VE�Htz-I���ö�Vptuw6>�u���9iG��P+�(	(��?����۷?SZRi�_���'OQ�M�kt�:����u�.�
j;�%J���}D.-��w;`�
3�n�L�S{w�6O�h�p�Do�)𺠢 ���F˲�NH��D�������nJKKlUZ�9����}ս������J?��M�����@ᦩD�R�TvVJwK@Q��DpI����B�j���
��{ ��E ��r����4Z+9�|��@��w� �\N��<�w���6�|��DR^RJ좃t�u�m�r�M��ٰ�l�jJ��(�[o�|��O=���r�~jj���w���I�;K�sQKD�HD��E�����UPvw�[�>���� 7�n� �@�6�3�fp�5(�
�VH��`�4E�t��J���	�FEO���fgA�!���?���k����@�����3�{��G�y��˳��u6�HZ�;�ua��mE���[K\� ؙmrk��V�^�`�Y�T�Ŕ
p�����R���W���w��W��!m�*:�����d���S��"�HQA��������[oy<7�����xE�"���]���ǎ�mkhj�6��uz���JKr����j��č+��RO�z lS{:PT���� ����w�<%m�e�h�����	� P�t;�ƭ"`�v��ӓ��hRVZ
��pڏ�?W���3"=]�{����,��ӷ~�w���=�p�����=`��.ǲ� ܼ��ҁlJ����C���a�'GoTZ�a3�@@!�$[(�j�����O�.���EIRBm�V�sUu��5���+��\��Do����=�}�ŷ�9 �lXj�3��e$̉c�h���ϰ�E���eD��LTGL)��cok�*�'�g.k=1SI� �n;M�[_I��=�5��*J3��H6�V�K�D�yFF�s����۷o�7�;�@��b��w�Z 
g��a]�J
�>�j<U�E�Gp���0��6Jڡ���&J��1��G�a�����ƒ���`�fy��4�����hw�����}���v��	�W Q�uI/��u=�Z|%{h��Vy�g(��b�2
��º!KC�L��X)��cwؠ�����=�!!A}�5����8/@��v�ON�޳��}�:��1?�{������/+'؏ ��Q�=|����rJA-����P���ëz�F�EUWr
��!�@A�thH`oeE��;A��z�yFGr��&���}W=R�@�NCts
n��LS����f�y��4O$��qڤ�d=ؐ���PX�cR��܅EQ�(f�X�+UG��H���tK�kʡH1XZR�����*{N@������T��7=R ����Ff�fe��e����U{��� x�ao9��໨zhgQ�(��uR�f��(o���`�YȪU���7�ѯ�������W΋������/N_�žw9r,�j�H]<�%�� �.���%�f$�6���G�`�û�.�3�kIz�����L<���u�n����
�ZPu��>�n]��+��<��Is�����8�����J��'�N5�Ͳ�!�n:8(�N�����C	
��U^'�b�0 T;l���9�$����f���eꏶ6I�5�q����8��L��\z�OccjW\� ��޶��k��������ёq:��.u̡T��ƦU�AA~@���J��B�Ǡ]�����'�����*n8�Y����D��j�����55?[�xrr2��������Ʒss������nd�̐��,��Q�z�@z�u`�,M86��w(T=8 ���.)����Cj!�����XL�*:W�,�}��W�����򯾥���p��?���{����� #m$�28M�xz��G�J@p���c�	;T�(����tP�Ӆ�'OD)����(ޣ��1���Ј�#q1�$/?�M�斆�-w�ukna�I�������v�[�<���`���5.7NEՂ�9�(��v��X�xB�F�W��t��7��A��h�&��u�x��:KMR��Inn&	�uu��=p��'��A#���޹ �ߵ��>��C���-
��P���aY
����u	�ý>af/�2uJt��T/�+z0�(�h�0<M� 
�R5`#;m�����l�Ã����u�)�~A�W�pH1P0���7������ܒ��l4�ȉ'ɂ�y0sL(Q�9 j���`�w1���A��cCޘ�t�ĵ��L�92�;��H� Cl�v�z`�E��2>>�p�M�ݕ��������G�j'&�s�����X_�y]ll��d�Cl�F���W=�!h��5.��!%T�����po�i���|�x��(,�e��`.(}`"��Ҍ!Q���E���b�&�#C��^r�KYk��*��6�u��Id8�Ğ>��s[{ۥ���p�JG�O6���yGc�.T�	n�f�M�����4XeA� ,l�ƖEx^�;~��oTl�#:PJ�8��,��u��8���M}_VV��e/����WtK&���ŉ������v}�ľ}_�Í�@I}�%���ax.@ ��Wrb� Cl���ѽ�ic��������,GdHTuu%��������ZQ���R��TZ��l�J\�Z�����=r<�G�#j�3���!�;m��@a�'��5�"P =|�9p8�8#_:�;����2>��TLS~Q�#�հte�G�ō���L������>������1uu��{(����x��%�r�aL�F��:�gĵ�x.�ЎE���	�����z��c�1�o�/�{t}�o*��%
�,��]�.�������O,�� s�Kw�����a�#��j�@�{��H��4�6
� �w�E���.�C8%˲2JC'�GEEu�?RV\	�Q+�é��i[m�X��D�����/���2���Q^�)�'��	V@k�7�"~4޼$"P45��fx��N���K���'C�.tD���J ��[X\�DeyͿ���s�(���`����7���b˗���B⮩��z=|ɟ( 6
��c���p"P�$�dHm�R�	����ׂ-�@x����p������r����8@	���).���O�|����V�n�^ofn���:@21e��)�*���Q����>釱";S[^���̘�sP�Ņ$<<�����W55@�VV��u'���o:z��/>�����#'O��N9�1袙��VEХ#�Df�|>q1#J! `���:�wO���C�ו�*�����܃��bgdddS^^�/��ׯ�1�4��	��(۽���w�� 10 �455�T0���zc>������`��N����u�Ui-��c6P*�:��x�Y.����U�z��������'7l�S��c@|���G����{睝�<�|���)dnv���Q���1�X�����'�U��
@ 7Ți54
�BƎ}SP���'�<I���S��v�1��� �n?�a|lt�qӅ��|��+%���E��O��=�ӟ�-�/	���5qlb�u�Jq/Q��E�-7��>�m�0+lx��g��+(�Л�?(ګ%$22���v����M]7�|�S_|PE��\�
ؽ���?�٣/��͎0�Hm�~O�<�f�h�����-��.`\�!����U5f��&AO^����Up���(:IC���{����ߝ����W<���^���ǟ�uQaY�N�'Ǐ���r�1gZ�H�� ���� ��ю��<�N3	*֜~n��Z��FE����\�uֆ���-[���y�s�(Ë/�㾧���֊�# U_�@&�'<��(�z(!|ЌO��q��ta��e^*Q��3x_�e���m����ƍ��q���$�:8��x���ܵ*.�>""b��~���#���_y�׬]� ���NҺ��ȣ<�q�9c�7���>��Ǡ�ϹC��K�ډ3�C�7�yT,�J�:�6�S'�~t��X]]�ΪU)#gqxLZ���l�?���{�F�k��!᤹���ͳ� �����||�vn���xgo��=,�:@��� P�c��"����
1)**"V��LoOOwZj��o}�?��T5(�@P�H��ߑ4<<|��:x0�fu���&�vA�K�  IDAT�R{�@����B�����9PH\Q�>�p��llr~N��&!!!$$8�N�_�UV^<�� �+���R<;;�ս��>X[[J�<@��.ߧ
��or��8:;E�����7�<h<-A������q;X/iRb<����B�[
�ذaL�Qd��811簹~�����{��H?C ��d�/ɃR��L@���[^�=�דy�&�\.}��@d2R�&���b|\lgFzƯ/؜���>m6w&�,��<|��ݻC ��֖%%�u�(qx �6fiy�?c<f���#zGz^X��s������T��@��Ą�����kjj^[���ᩩ�����[�;v���Ga'������*Q�� 2�«,oԽR���v	��K���ԇ-?���uÆĠ�����>s�9?/�,cc�kgffn8x�Ѝ���Ch�Ag��x���L�w�Tb[4�)y�B~�4��`/
(�����Q-2<���Z�۴y��կ���C����\X�|w�n�ݷ?w$P�淈�9�4�$ϥx�x���m;�R���c�˶����T�"�B�e�]&���޲���+J_V�P��k�������~���W��ɑ��Y>\Z��{/�N�G���Ͼ��(���X�E�"8v	��4[�bÄ�r��*���L�ݕW|���f�r���������ＳJդ��I������%�
���������9�/;�)��FU��1&�����ꮪ�|��,�%A��;��~WD8������]� Q�8������N6��w9M@ �$s�1Gu��	�c����߾7CcΤ�M���d���{3''�����A1P���!}����^z��:�!<<<�?q�7���nS��%��x��NX��u�����zrIB>����oܸ�,��.tnܸ��/��oqqq�6�P�(���ڽ_����ϚL�ё�Q������z�B�x WTO
�|˫���?x��$ƻ�OPeV�z�䢋.�es�޾ޮ믿��͛/v���Q���SU�_{ӋiikB������o�� 9�6/���{��4zՓU[x�F���nY�%�А RYY	}����������-�������GAkbGGG���^�#>>1�~�ם �W�PZxZ��Fɍ����vr⾀���У���{Q��e�1jI�\0�-ͭw�y�}%�k���sP����ơ�o�����Ā� r���3��	om�����y��B`�s��� &�n��^���{0?q��F���,hzu�����������r[[��4w&����/��ϟ��%D��T}#�����y�cɧ����p9�U�;х��M�L��N���)���&�N��P���K.��?������ZI4�54����/o���]��j�BB"<{W�!/M��^J�������Y޸��	k��(gZ5kن�TEe	,�����-'#���kSު��|PI�APpif�9�f�+oi�x��ߎ#DC�?N�2ܼD�Z�q�rR���0�T)�Z<�VRU���4t���udUD�pqq�3�����dW�б������8��G}�h4�cǎ��YoI����f}�K���J.Q��I'2�`;�!9�$!.ޜ���M�J�G�f�<*�J�����������/޻wo�ۭ"mmmdxd���A�/��K�/�+�Ug�>�z0i�Z%���(�����$'&�Y���E}�YAV����x���ãG�~��g���\�qWG��Y��r�%�Q�19)��T�0VD��M�1}��1*BbbbH~A6����+��˦�%�9/9s��qá_ޱ{��P�Ο����+}%7ؾl�ټ�� õ58��[ps�rB�_aQ.���/.-����E�����������ٵkW�������>]>�t&�B/'�2^e���tUd)bX쁪G%\2�z���K�IRB��ڌ��m�/��vl4��������[kkkW����H6=Æ�-w��$��Wt ��b��`����b��{���/-0��`9Yy�����x���~'ʪ��d�a��Z�������;vD�1�=@Q����f�&����#�@^v��f~@8P@hTQq	4��K�a����>����u���󒖖�'�{��0�Q�����4rD������m�/�(g��I�o��� �� �K+Fa�) 	cGj�U���sII�o��s��j�*E��s�������ƺ�������������������ȁ���[�w}��yS9�'Y�o)P���ڂ�HuM%�X���4���Y/����Cl���������O��_�����s8ј�f���g˗�y��H�rBY�P0{��f�Ҳb~c��h�쒋���+��G����(������7�x�)))q Q@f�X$^����UЗ=����M�FCǟ	(�(���;h$���56��暫����+^8�;���.�?���5k�$P�>(�i\jOXnI����
8����=����^$-$$���eC�g��;1p��7>��"Z�l��9ITK˩��}����'���%�C���(_ގ�zri�BF�ǣ4y�����<S]�Fy��Qc��0�RG=�^��H[��c���|��Y��GF*������Ѩ�{���O�������АH�����������Z�"0�k�]���?�'g�x��$��a�ebb<�,544����m���+�.//� ::�_ɖ'������~���w�y�/l���Q�����40�!J �}(e4������|�(_l�W��;ƻ	>�%SSt�y��c4�Y�<��Dye��l��ƚ��a�Y7�Q�n��h�d�kff����9@P���� �+7�x�x� ��(����w:`ɹ��͌�J[�9����`���;������=..�DRRz�ʩ(����VT?jmi���_	Pkt�TH��5/Q(q�ұ�.��rf�#��.N�<���ӆ�Rl4��-���ssr���g�K3>ޓaYt�^_���w��b�3���&2h�d-��A7��+r0����������L��NU��f-�@**ʈޠ������͗�*((H��D�@��3:ڿ�j��z�x�u{�|��aЖyh�����i����������ۼ3yT��|Q�0�깥�zLL�&�Xܱ���^���_��X�4A�α�'��ڵ;����V����/,K�@�b9��k�i�\����y���q(s �����2����Byy�S�E����b,����'w�|?ya�B�[��n�] /��1~���$C�/瀪��P���x�3��zP)�<���3����*Y_�d�1B��9�zCCC.�b���߾�Ύ5��&r����'��]B������(��%��J�����~�J;�`ΰ��&��Q���K�y��\�i��G�������[���O��hX�N�Q\�O:QϦFH*坾�񐛡��<�oz�b�1��p������ 44x*;;�Ś����d���b��fs�(:
Z[Z��;;2a&r}C�`s��A|�:�Q�l��k��;O+���$�*��RP=S�?jժ�ɼ���>�4spN�����h�[�P���'{�f��������z��B\��K���_n�y�?#QE�/���ǣ������H�jU�Tdd�7n�}RR�)%U�sJ���\��g~����DjiQ)�ol �!��Y4���+����	nH>���c�8S
���F��`�TE���� �{`4�Y�fs�w��?��⫫�'�w���w��s�H���d����Ϝ�NΑx�w𞜰"X�+�J�/Jb��[�y.�����D��doii��[ݴi�nS�W�b%]��[߸���5?-9�4�����!Oo��'��hr�P-qI,Ox�F�4�����,�2Y��%���<b��
�i���@��l���[����}�t=̹e��5?�;11]�:mM����p�|��\B|o�۳�m���$A����8��r���U�_��| 
��&�u�a�������n�VZZ�x��b�`�^RR����.?�V�r�hffn��������c��?|�R�S�p�F ?�K`��ha�"lh)�]ֹ���J����܋��q���NB������F�ux��s�M7m������"(
@"�$�l�{�}��͑����466���i�RU( n�>� J>q8G����O���%�9Y X�	����1y�	(���dS�`p*�U,�+���/��9�&&���;�JuE@5v7Fu�7_��������7���&'�&MMMd|�u��<>a������*�������R
)-�@�(Ps������s9<ll��@#���!&������PNNΗ���/UWoأdoE@uwwG-.Ζ�l�M�������0�ם�����w＋�8;�M�݀�	�%�C�a�X8�)�5�:�Z��ԏ�]���,ˊ@9lv�w(s�͒�7����f~~�#���^P
�A�%�*��ͮ_}�?t"lw�?`>-q'�K<���A����HZZ9���y��7�$�����A�1���d7�m��f�EC&�?ac������_,+����d����Y_����@�������������|�GA��r^��k�j7�3X`Xn�2Ж��ԨK3�qRx@pK���x��?C�nV/��'P)		J�X��6>c2E�!� �@�G���TC�3;w��v�����qcܖ{yK�,�$hL�����?�3�7��� �N~�|���>�flNdEEK�U���2��:�_�k.|"88��8q�5:�hZt�r;Z���޻;�a�e{[7M܁�C�Ğn�+�k�(Hx ���ZB(q�9R��e�p/tw4���CR?�3t{4i��o��B^~IMM�X�����5��L�I*1~~���ށ�_��aE����B�ٻC�ܘ�,��C��JP��s��6a� �=_/DI���,��q8��K�&Ⱥ���B\\�Tff�/����|$�K�"M�'�|vǻ;��p�����0@o����X�F-�Cq2�碠p1���g�%wIȤ��v��`A�
xx�������ת�+���[q@���G���ϮZXX�O6�fW
����	\��(H���� ��{*�c�wp�%�4�.��
웚�Y``iTT�TNN���5�����҇�QP=�V�28�w��;w�41>�����sޣ�M��,_�u��
��d$�AR	<��i��z�(p��Ġ� 煺^eU9����}gs������9'�@���.��b�����:�N��A6o-'I��8M�$��i��K�e؈�����*����0	 JĊ�g�Y�FE�
�h5��W~���22>]��0?�X����=��o6��0==����N_@Ɂ��1���t�4��@�E�/P�%/�(�*I�fi$/��-**��0���6������_��5k2a���.l��Iu�7���������������%�N<X>m7X��)�(t���ݦn�L8^�N䆭���Xր͕r;Yvb�@��2992��η�����S���1������Ȏ����iii��O���V\�E���>��v�岜b���e���
WMI�/g�\:�����Mcׁ�*��b=P���U6�^w�o�			 �w���bc�G�?����:|YJr�����LOO3�q�m'�A:h<&5��s�ԶP 0�==��ɣ熥�N�w�Y��M����Za䈖J�
���������뮏���Yq�kn>�t��7�87�X�������%��,m��v�3c�DC�D�μ�I$�+������y����L*�eh� �GX�.{�׿����z�S���\\\t�mSgE�`x�?����7_�ǿ�����*�����I��+_�@Q������.�Eۅ�C��v�	YV��.a��	�ˑ������@��f髪�ةRk��k^����u{g�]VPcc-�N�W�45}grr����!M��i���Ą��x���
%��&�����2�|N5�� j�t�L��u؛>g�E��z M�EF�����啥�2��b�S>�&+H�ݾ������W^��M�ӳ���A208�s�
�{_l��~�1w8ρ�!P�}��ɘ-�c���;ײ���@�
z���l�qQlذ񞨨����M\\��l}��$
z8;;;���tG�<���w\�r�A]t�\��1��Y9c�=�\��d$=�	8&�n����a $8'lti>�f��ρu{�����/���;���zzz����g�(��XO��!Dwuu_�ګ���aw�����4˒2���xă�n����-��F0{ÑJ�nb�?Ý���w��L�ဂ�}H����XKbR��6m�_�h�s�Q����:	����ƞO>����T� �-�|�aز��~O��t�����t�� H��w�+%��@� �A1�Tpll�-1)�͋/�������3P����!����l��_x�)��kaff�N�#x> �ri@[�=	�f�l�=L��3�)ߒ
��9~އm�,�*yo���m���VGmliPP�G��R�q�o^z�ƻ��9'�jllԍ�����olmi��fuD@*x~q���� 
����D �aU�IP�D���>�U��
����:e�j�6�F{H��\:��P�.���@���It�*�ZC�U�U�zMfΞ��(E3��(	 ���ڒ{��"��׮�����&��Q�|v�3�^Z2�6� ;��l�4N�Ap@�p�.<��HY�@������>����&�� 
���v�?M��CI�U�hU��V�"bՓk�$(�$^�ɳ����x��(^
z�Z��A����4�b����|��4U�-�E��,&��͛��|��<la��8Xw=�9759�r6s�aO��HYw��j�e��\x%|258x�DUY,�%g�R�db��'x�큒'j��mY�����=�,%&�\�F�)mU �oA(`�r8�&�C�#5��@%����ڇܥ+�d27��I�P3׮����??4�� Rn�KˏB�MnR���F Q���>����#��(��2�G:�y� �`��	�G.��n�B�ŽH8wܵ�\'����t:��I��������''V��j?����OWޯ^J%6664�X<_�KIzD%@&��DT�9�R����i�T���%��pha&�O���<>����r qP=.t]wJ��27w������_�J=������7���ҽ���=��ƹ'8�}
#��I&Rp����E)���q��s.TU�\�s]�3�8������TQo�U۶��i�Z�2J�p]��:�,��A������[�nxg�N����G�M�=�uٶ}Y=)Q�o�G�/.�:�ۛ,����m�D��@���Th��F%T`��(1#Fj�:�-����P�T(>H_a��N�0�UF1$+�Jʕ��6\�0��w���|Ϭ7\�)Qf�p�0�'��!<A�T���2�2���'l�K�+���'ݰ��ӧ�EU�-/�զ{��8�Z�iB��eY��
�١]��ٻ�0��/�0��<�'Նs���q��h/����y�T�c��)u���U�a�'�o�}ȃ! Ÿg�OL��0ٗ��/��S�P{�T��Dl֑��@� ��߷û6�    IEND�B`�PK   �<�X'(�5W �@ /   images/4737cce6-ef6b-4e79-82eb-dab57378d86e.png��?���?��*�N�Y�"<)�J�q)��+�9/9�ͩ*������i��"����ls�a�9nc���~=���O�].��?���t�^o�wL�=  ��߿� 80 �<t�w'�#ĕ�c��]}�C�O�!�������[� ?v�{Z���n���<�{q�>}��B�
n���O�;+@^�?�5D� ���~Y"}�~J٤��@\�,�m��g�;�o��]Q|z� EC�J���2q�D,�۬>�Xk���i�_TO�h������T,��@7A�}½���_ؓx[+��3<�������9�X��,v'�W�K���R��2���W���&��0� ��ِ���MA��+@]A�3JY�`���=Ɲ][h�Fq�M�p	@�3�Y���>j{~����;D�oy��s��-��y�����'���������߷��o���۾�-' �o�����������Y�w���9� ��2H*T8jfVtðKݠm�촿�h�X$��p�Y}���03a�H910�aUv�;�bg�"�gC��wf;21�m�1��m��K���0vTss���t�bbf쒻����|��F��C_���\7�.�2�%+���Q���}�Ȫ��dVO���7Kj-ڲ�v�S�o �>� 6{H��@��|��k̰���D���Y�>%QO�Kߚ��;9�ܠ��ܯ:�E��g��"�4TfIW����^�m"�ck6?[��;���qz��Z򧹤w��� :(z��P�F�:�G[\�'#�vg�#jKKʸ��Z���W`zb��+A�쫯1�\~(�J>�T%c،��&��ݐ�N8����_�h�l~��}�BU6�2���|!�`�u�OЭ]mz�V��"�����"��ձߪ\nC#�M��E�`�,��OV��H<���dP��)�����t�ӕ����E����O�.9a�q���:�bug���(�B�xg	������T_1c`T���Wcɟ��jܺɉs4�7k@$W,y��.�h��<^R�Wo�!����|(��/]�{o5Hn7�ǔA����4�//�蜿���%��6̋�)�J�6��7�a�/(N�˻@��wмiL�~�[�SLi�$S��q.�b7�_*-���j��Z]8Dj�'�^����cRe8��_�=+ZS�N����X[��MuF$���I/`b���=�nboZ�A�z�����n����42�����3��9��5�^CQriJ�>t�֖�q崽�j����֞EsV��,�(��>�u�w�8�$1�L�sd_�s�3R0Ոn���������r�bZ� ]߅�3�i�w�?��,oީ�����R�Tb��4)�@�{��u�GvލZ��GL���^>~ڥ�|u��,���Oٜ��W��Ij�̈L/|^7)��d�̰^��҈�	���y���	��v`�_o4�}��;[zoå�\B��fk�4N.������s����Ы^k��nH~�p��"�!gb��T\�{�O�L��t�K�Iw�����Rdl�d��B�oR���e�m����D�����h�qC�����Ҽ1.�*�>Q�>��c�8�
9�#��DVB���o3�mI+��5
mT� �hR�2��a�L&|Bn��^;���nM��}hq�W�΍��s��*Ʊm^A��xy�ڐ���ã�_u}Syk7q�	KeΜ���mC1*"Sw�&���(VT��-��>E��EW�t��ԫ�M�ce�.6{I�H]�sl���9�עQH3Y���KϦ��*��.Vj��g:rb$f�~��	m�'9���S�Z�Բ�(��2�s�,����_l���I綧:�J�B(ra�����l�.��ɬ�h�������H�v��/	��´"�8
�u�O��A��3V��3� {����|i!A��WNp�Ah��0�"�����yC�Pʾ���U���.���ه1�9IU�-�v�_��|�ɑTwƥ�0���۸��Rh��љ�±g�ckt9��OE��Uֻ}c��M46#5�2�����s���3�wNp�d���}-g�'�w ~��+�_{���UZ���\�m�XiI�7�r�'b����d������Z��'�t����5B�:Q������ti�-ܧӔ��0 ����!�ݎ��#G��ǧQ��5$�KO.�/��ԣ�P#�Ẅ���1z��]�C�>Z� �c���	��J-�ʺiZ2�xT�����@�>��Ӫ@��$�Gكg��on.���;y���Օ|p\W���E7�R���>9&��j����)�ѩ}5�$^xF��J��
�P/H�����a�w���ͪ)�q���Ie�G�
�dq�]��2�CBv�f��?"������U_I8�ڳ���4�R��� �}A�;-4S��j��:��t��<H93�O~|�A���M*�&�s�@����"jq_E/��1+�_x8���T�S"L#�I*_Џf���;��T�d�MSҦѩc���I��hj&�#�~��L����C`tk�� >`db�7�x�2CE� n@�Eq!�@�`�8W�׻'�w%��Z��<�������vw�>�,ͷYd��P��}�hy���qSǐ7-IXg����� ������R$g���l�^�|�j�6"�Mi�$,d�å��r���\�ۻ+~F�B��M#����͉l�����,d�B�k�G�^�ɂh���]���Z����q�Hx�C������ګ��f��nC�?#�d�<s)N�2U�RX�g�lWz=!.��H�^a�ח��@O2�,�����:�6���\g~�	ix?��z���\b���6��.rRU�u��Y�t"s����ya�4�����H5O�)`m'��x�e���n��fF���%ڪ�������(�{�7���}�L󻠫�)
䘱��9J d徵ΦtNr:)�=�S��xBN�[�9��S���
B�L�6�٭���'3@fKe�0����?��_�1V��L�����j�!��#�b6�>!��9�i��������XO��c����/�~З���eb�nj�.�������ey�F.���_���+���H�8�-!~.��%�C������9]6lt1ьh��-��B�D�݇;u�\d��]��C`JN�Q������AY�X��q���S�Ry��֑=���$ ����#�o����T���F�T"��9������i̦r�5�uٱ�}7�}T*ВM�q�Șy����ـ����!\�S^��&�)p�´E�<�_8)�3�i��m���8\��{i18W�u�Ɓ�M�5M5/f�Y�a��~wr���;�s �Ҙ%��|��REټ�#9�W��㼪�?3+�2��z�d��#�-'�"^��������Ra�}Ϯ�j�>�w�hI���lB7����;�V��/$wv��=�>rRK�
s�3�	�宮�œE��,��k��x|����,�w&$�]�W2Z�׵dD���ywEwN��w�DX�aN)��F �*Tca��m�.�Y������]��I��$�}���=¬ _,�F����s��Yj�W�n�>R��LMϋW���=��MYP�B�|ٜp
�I&�I�z����039pp4b��2]o<��d�`�؞Тg~n~�����C�����j�Um�<��pk��;I-��͈ȹϱ���."��/�o,}�X��-���z��;��M��sQ�zl����T���I���m�by�hz��kqv�����<���e���%�0�'�^��BN��� ���5���@,�v��n.C����hf��Х���	a]a���Iޟ	e,EO9�b�`��)#b�]���7
f�.���}Fl�H))t�)2�.]���9櫻v1W��m)D�2��[dow �Yx|�vw>��^�>f_��]�ߙ^��s7>�va�'s�ŝ��{1�1�4�ЏuW*���$��L]�>J�@�~A|��)ז
׵��A�~�[�\� ��?)'5�̗�{4{h`!�1��^����m�	�{��AeX}1"�Š/�����[ooA)����}r��Ŝ�}p�i&A]�P�Ik�F�F�`k�����RXx�T���X�i�X���]�^д��k�1���s�����3�5�u%�T��u+B����a�V�x�m|*^�^�g%�_��K���vֽ_��aR������h�����y~$6 @����k��{�~�%^�xb�o�����V2c�����9�6M+tc̦,3���M�ww9����.���m+n̥��B`=Y��bĶN�[$��o��%s/���a-\HqJ���sS���(Xg��	q�F`.e�x�������@�"wܬB�m��|�.�Bv-�_,���~�z(�_���b�������č�Kގ-��:��'�C��P�J��D;�Y�ON��)}/@o�xQX��t5ؔ�P0��u�Y-8;�EN8�*�F������n�>��ó	��x��ƌ��srZ
uHX*WJ��:z6���K�g��ɵ#�V�ZI��喱
1
�ea�e��j���c���!߮ ��Q�����AD��!�����_ת
�G��R7�6��O��,����L>�i����^d)O�s.ډ��MJo�����gh�U���;"G��bi<��$*�2�E�N��ԤS��}��@��`Rv��%͑nR����9��chU-�5���{GWt�-�$'�=��"����ǜ�k=��Ij�ɢ� ��J�ވ�y�~��IY�[	��/2��R!|��4a��?�����+éO��x���Z�G��_^^ܣ��M� O;�r�Ơ�$�X��c�{ �N��M흌Ɋwhi����<��s��7��1o��~�����'��S����!���:���ئ��'�6�7YM�!�
 �F��F
��4���o��"x�Y3�"U�r����i�݉�oOن"u�c7��m�����H���*�A]SN��<�1vh�����)�=1�Tb�������������Y����v�֮�m�/��ɀk�������m����FП�c>+{		��UjV;/��sx�<�8v�V�
��d���/�Gl�*Z�C�|wがQT""�ioTMء�^��Q�;<<Ί������X���s�~�ǜ*y�~'7��N�d����Awm\��D��+周�e�ɉ��P�z��C�k�I���\U�V�Lu�~5$�K#Ex(�g�%.s�o����S���\�F�{|�cv�����n�^\�69Q᳦�54s�����1ƣ�9v�o�ho�ՔL��Ȕ��|TYZKl��Kd��J�WC�%wY����c<��ؐQ��;6�����o@GK�[ܩ��߉Lr��h�(J�!usD3�����s��?8~#yg��t���~��Z�̫49$��`��KŅ]X~�O��q���.�<L�V���,��ǹ�J�.�-���cvn|���������ƞD�����>W�E�YQ	�ח��y@�ƪ��D�����p^N.�z1Sbu���*���İ�U��:�K4��h�ac>���m�۟0�W���ZbGޯ �_�ym�#qÉ����X#�=wnb������e��M/���v	?h9�N�!���j�i���=�7_��cby�#7�5�џz�g�gy�95�dw��'����CJ�S�/ic�Ãe�� �]���8y0 б;ڄ��S���t��A�icK��O���V�*9]��曖0��q³��;uY��3f/�1!o ��V\�:�z�^S$���)x��Q����
�UL������|J��Y�����/��sVY5G����i�^��*sL�J�q+�f�\«�X�P�v�6D֯G*���!kI���\�Nl�SŖ�zΦ+�_%0�~����R7�&#�7�y�oN��t�n�=tp�x7[�N�C���h�j����F��Iק?�)ğ3b#��܁����W4����O���d�Tս~�2�s�g�p�7f��˱IY���f�^�N~�݃����./*�:44�)T���#�/�<�/y�'ܰԢ�� _y���i��#.�n�^�9;�F,{ȩ4�=�����.{I)������r�4��(CY���v��_�<(���/s���'F� ��ޟ?N�~��=8w���r�z����I׈�'X�6u�~�,%m|���sҜ�y;{w�X`��O_��bҁ��VY��>t�
��skŨ�f��tR�T�e����|���`���49��9���2�^�~�l���ˍՋ���ٷ�q����%/���w��R�~��Ϲ�z�T/mp�@��w�5j�~�y�%9���H�O�f���Q��و�P��T>r�7�����>0x��8�:?����r�&4Z}lI(��$6I��$��2р�|4�;��'mt6����'2�op��+Msg)��jՂ M|����	 ,|OS�1R8!@8�-/y�ߺt�7�'���-����I�;�.�OK�C�a�jw`R���vSM�DH�$ԑ'�o�vQ	�CN<�_��h�A{��A��XU�BsG�B��bHY�9�rh��.�����.G�b}��)�M����S�x.y��^1���*y���3�D�ڜ��9ިj��f۟g��鬻%�,�1 F�|��Xp�b�u����s�2���� t�������hB��8+�좀����y%�Z���.󿑀=�^�Cb��0�#"ě͋W	9���OT����� ݗR�{��")J1&�T]j�J�aþ�l�)?�?����V�i�ɦ�y<����'D�*�<a�d4���GAD����r�w��-Th(:�"����"���)�uu�ʁ��[��fM೔ӥ0����]?52��-�� x�u���������}��5_ͷ�hx(�����q��;�
�Q�\��	h%ۤ�(��m�����3՝���T���s������H��+��Nq��M����ˣ	m���G���(jE�gy;���7���'`�� D8z��)��cw*C*�5]Y0�|��r��-�9$��Ϙn�i�.2�
Q)��uv�(���\�Gh�紨l���o뀦�)4)�\�o]�r�@U�Nb��eZkr�(�{������!�?1|�{P���d������)���kdF���6.�H�lZ�����W	�����	9x��. ŴD���?�봀��T%א�,ƆX�����ZC��4R��}冑���ť5,��Su:97!
B�hA-nQSיMAs�ugjlO���:h>�<�*���à��C~c�X�錄�X���O��X/���_]�L�3U|���|R����Dt��Ӱ� ��g���������˲m-���f�u_�=�i�ꋖ.���
Q�	+B����s��J��~�n�-���;��r�p�m;1�'��D;3��jEt.n�� �����/_��_�������3'���(���EK��$��í,�����@��z���fQ0�_��>���?��0*��<"z�� <[�'Q��^h��w�c�~(�L�����\T��{����~�a��N�f�Z�2DO�֗�RXJ���N4�R6x��"�e��Զь_+�9�,/���}����E�Ǽ��m?�n�q�ո=��!�a�}��6 ��=���fч'�M��j+�P+O�j/)4�|��`�4��U�!C�����6�C���ôl��LCO�h��]������Ԝ4����6Zo��L�b"K,�/�k����Ł���
3���_d5t���fD�(��6q� �+�`���ol�^U����~�>O &�/y�ϵ�w�V�u�y�t�nο�ؖs�Mg�T^�Rӌ�NR�����BBdiZ��Ρ�$�q׳�[M�'���C�ۦg�����Aҏ �ҋܗZ����K,�*y�f�syM]�
\������R{(�{U�ȅ��Ë+B�R��*=�ۀ�O�A��'�(q�z'z,3��!u�Q&Xp����c�����$��s��n¾t��O?�_Ij��p���`�v�j8���1#�bWL�}�oK�7L*:.O �o�׬������$t����7$L{y�=86}�v�bb[�RK�KK���+����];��sssWh �����;
�Zv�Q[_��_Nj7����R[���7:p�*�#	�I�k��&��]S^��2���:%��9��[��J��H2�^�iVONd��1����u٣�FB6}NU�Fmp�!YKTmbQ�1T,����iX���%*�Ol�_W9�an'S��A�4�P)��7��Zx�1O;3�G+4ޠ�?�ɹ��H9��s�1��2~jkl{Z95j\�O)���p{qj���
]
Ny^��d��*����z,��9���?��~����{�Wݥc����8#���Ps��՚߽&:q �jwz<R ��Y�qW������˷]q]gQ	���9&O ��o6�5R��|���Q۩k�/>E�e_��'2'��}΢�<��8S���7�f_�,��sW�Lb�F�ȥ�z��MHc�#�:"=� �����q1�����X`@�&hǩe�V�Qҽ�钷j�K"�fI/���� O����hT5T����>�9��^O
e��r��K )ó�ьMqz�EP�v� G� S3�(�q#�̞+U���9
��}j[Om�7��Y�(3�v�{��ot^��;9*�q��C���G��������ĕ=B�z)?e6,��X�Z����JS�[I�M(�`�J�ɭ��^����DU6II���0����w���_�c.:��Q� ��L�"пbc���ȑ5�w��>�1�X�*����c�ڃ���WEed����ࣗ3NO(=�F+��\q�bV�d�~܃�e���RѠyc��H��L��V��P�^�wi^#�����m��̻~�@!G��PO�٢�N��{�~6yY*?)P<V�Ut�va|*a-v�S��a�
;m��i��3x���}�n3CX�Y.mX}�Zoc��/kd��Z�|8��􇴯�s	M;w��?�W~�����������Ww�v��%����Ň���|
?Q{miz���'�Ow�o�y!6�t^�|6_���lߧr=���B�����9o?��g�8ROդ9M��I����Q���g� 3M�֏p��� ���A���s�7�m�0m��L�0T��CA?�rp�|�d����)iTg�Ͻ�	���r@��슢��SMXN��<B#,>Q�ˆKp��\�L�-K���G��d�1�$���q���ieaj% ��]j�o�-�Q[���K ���
�9^$�h��2ΌF��������_O;t�6������� ����	�>�*����6~pD�܇`�`�=��ƕƅ��28�J�p�!G� CI�������s��ǐ�zY�?�<n
�A���:�z���|,_��Ӽ-��#�@���>��@�m��o�.:rH�G=F_]���p:g돐�+x##|�a�^˖�X6W�
nFo'o���[9�ƭa�u1�vWX~ڰ��  �k]	���r����mz�79_����N�k�j�	w�� #mTO��ZȜLH��(N|V�Q��dr�����9�~�����AaxM%-��[B~t�A��y<l�P!����Ƀxл?n�  ��yc��!,�!��ȩ�N�����I��_���RW>g�8�*��K	=���>�8�㈱�i5Gٟ�dv.�n�2�Ȟ*��zO�G���\`��W�K!��[6m����,��K�v`���]Qȣ'd�yq)G*��.��.Łjұ���A�)X������'bku'�"�c�2؝
�o@����[$���Ƭ�7�-�+���.s���"<�u�����XI~�v�mI�1Dn
,��^���^H�{��]Q�D� �����
$�{���݅�K\ V����BqRp���i���B��5�	�s�!F`+�{]��	�7�(�{4���H��7���Xb�����xf̽�yfο^��OAV
H�ʁ�a���P�0]�z*�=��2�""�}}�8�Z��㴑J퐐�E*���e*�֟}aegg'�{�.~����V�ڿH����+��7S�,��5s��@S'U��L��ը�0ݸ���o�?����$�
4Ʋ���С�'hz:c�����C���Y�RifT�b�v�Ȧú�~"��<�ӊ��b=�D��B6�1Q��Ŏ4{��I��	�����E��>>���M�M��V� �W�\��O}�r����/�>(�RW{�3�����x+*!141�e�����7fR���5�^��kuL\\xlͮ�LN R͗|��N9\X�`�#µ	���Ek��THQi��=)�8�6_9y7��f��r�>�g#����?g��3;��i<ox�ܮ�������XH�����cu��H�������� �-��_��}�j0�q k߲L����9�\\��^��?G�6�zL@`(�%uV$C�>z�Q:���Ij�=A��DƆ���"3EJ\p^]g���^_�'5A_�Uu"�-Жg�·�@�;��>��<$s+y�	t������sg2Uй8���=F�m���|#��ǎ��rV���My��|�i/��	@�����^��,l;�A0_�Ryg��v@ߡ~��u~��8�u�b��%���/�}�.6c���{X\]�X�K�����U��\Ͽ����?�)f�1�����^��NR� qE��G�����<Xg����].���N=R���!ja��o*�e�R*L��������[�rj�=�P�[TT�)x�|?Ԑ�^�?D���(��Sg`�ǉ?��j� ��ʨ�!���[m��m��_��׻!�O��ǧg�C=��3�(��o�m��l��
�I&&�H�#�i<t���'��Ŵ�0	�W��c"�$H!.��<v��|��0v��6!�����������.�E��}o����g`Y��i5غ+�G��0�e{��?X��Բe銃��a	����x#gA8�%��0)��#�dO����S �p>&�恄���	�-0c>n~��� �[Ӂx��7���&߅��Co�m��,���#�2��)2�ou����l�qy�m�Ѕ���O�<�-��Β���+�ˌ ��EQ�#4x}�|E>ux�D�s�'em��F���:���*��l~�Kl���P��(����ɪOOW�>*�<�(��'#�/xIQ?߈"��G+9�_�}=�j���-����
^�����ȼ6��f�bx1,�J:�(��[�S���h��X���Ƚ�F�_��7Cu�	��̧�����e�}^�����JjRUb#�'��� =�Xz�v�,)�Bح��s7{&�W�C�}*Z��aצ��2$j��ޱ7�E���� �����p_H�v]�ZcN� 7`d���!z�{����8�޷@s����k�?Y������������|�ʤ�o�|�?u�W^8���O4����3�o9_��h��,%��j~A��s�G4YF�,;���[�_d�7P���
�.����PRR��N��Ø��/_��j�?HB{���BK���!��:%iQk�W�^w��.f�ܲ�Bim^ck�{�?v��*dD��|Hn�A{rkg��TÀ3�"&
�S�3oV�4�4�`�XX����ٶ�Q,��C$��8mg���$���؍!� P�7q
.�eK}�񣖢��$	$(��'}0|�7�����{��l�o1�q����j��#�;}��"PT1�)ͱR d���A�f�N�ɰK�=�G����Ğ�P�5"�:��=YS\]=�^5Ը��˕c�!��b0Z��*¤��7�)u�Ch�<j^Jr�-��C���T7�����Kd�(��Z룇�������ۿϩ���զ�g�\�ޭ�%��g8͊��#�M|U����&p?�wu���CZSէ�,Ｖ8�.~�r�i� �дy��эO��?���R[*�=�	�/�l�]F���m����z�`���ʶ
p���5�fW9������'������*���ڍ��~�0Z"�A������JG����Ɲ�rj�ֶ�|�/y�Jiٚ��*�0�2i���
tS�92*�Zz���ohŴ`mxI�,�=J���mQ%+d��L�^��#
��N.��.w&80ŲyU��ɘ�G4��W�@�e�h�T�?�O3�WN�;W=X�|�.���)_hX��,7w�H۰�!%����H�tC���ߢџ��ME�q��S��gK,�4n�K��v�D�[IcJ'��={e߳Ί���Y���r2�0�|����E�?Q�,|h�l������G<��SF�+�D`x��	�*�&�0���4��+Ф#���h��D/{�x�	o��>4S�w�{�<��v6������7=����&<*.*�}*�Φ��20RL6_�x�Wɇ�_��.bP�uV�Fj͸�k�`�SJ�g����[}}�f[����t�U�������r�2�v���O/��
`桩��'	7��S�h�J�GD)�L���K�e��g�1%|w�mN��u0��l�i�y
�V���t<~e�˛�
n/�vJBRC�I$R�o$`19�^]���o�T4��d~x}��ώӻ�< @c& ����%�BXt(:��7�T%/k�2k�a	��@��J�
�]���!���AK�Ű����\�B[z�!��o
WUSU(������zT�TИ��� ;���UL�"�jb2,��ШQ0k�\���)�m�e?��6�a��I��B����ꋇ�R���J�}��НL�����+��ywd^>l�	��~?��uJ	Ainv�ܝ�.2� �x��t�t�uɍ!oւY�!�<�
�X���PB���*�K�V��"���^m�i���'y udȢ�0L%�Q�^����Ⱨ�6[��عǨռ8��3|�3c��zN4:�
�ߘ=`��h�D��܆tSW��{Wc�s�!Ý���ȗ� *����h�I=鬋���dK�%��~��{ı��%��www������(��z��n�&J}���Fh��l]p��uʕ�w�Ԟ��T&I�����?��v=�}�iYf�>xB���se��To�/Y��Z��ļ�dMZ1�-��p;Y�?�A�1�k�I^n�ɕ�vW=�[��*P��wX#:An����.�t�Ʋ�<7cE���wynv6�_�E�FZw������?�e�p�p݂Ka��)S:�gF�r��ᓘp{R��=�6��u?w����.���i?G�{��{N��)�����FM�������_���\�Ǝ4�Dߔ*�:~e&�0M�K,i��y�m�du���só���>Z=$}�lKy�ְ��N��6p���6�w���J[037�#��s�civ���(qK�U�A�ST�.����*X$�P)�7o�{��n�eh6OĮW趒�+ӌ��oT?����U+�nL�~���$I�Q��鷀����;�s�?���\��lY�49xk�W��---[�`���U�-c�8��F���3>�tujsR���ր��Xy)�	��Ϡ=G��ո cy�Q�שd����R<o��ϽR#=�����t����[�Gm5��VVZ�ɗ�Y��P��;���`j�����;���(��g���&�h�3NM-s{�f-,\P3r�LQYi??)˦	N<z�P��tg D����
!f+��fR�O����)��pc��EK�k�Xf��&��1Fx��Hoↆ�V�4�@ �G{�2|_�n��ȥ#K�&��+ޮ"�ޮ���R�����Z:O�ڂ4�Z�:�[��roI������{�n��v�`r��m�����PR��vwX	�@y\���9�k�4

"���l�ձ���ּ�6`�K��-����
S�U8�2A�9�7e�sH�q5���p��@J�Y?� J�F��e�իW����`F���S?H��t���$�ݾ�ߴ�:0��ѵ��C�nD���ɐ�kw�����o�q���J�@�_*�����U̱+���Z�A���4\�K�(U�"��=hg�%a<��>M��@Q%���U��'�$�XϮN:'�hΏ��>�2�kg����}�e`3B?��]���Z�b�����GWA-�U����BK^)
m�z�~��)�2f-"���x��<N��	��|}}Kȡ<&:Dg�y=�
\�����q�����~l�}�Q�V�^o�a�j��� ]���jJIf����f��������pf�17�pV���F4����w��CPڹf��:�HJ3A��`s2%���X;5���h���C�vGs���FDR���@�֗^E�g�
W��w���4X;[.��wp�&���lc]����a�YF���,����XҌF��Dť�p@��}�ۢ�dd6��M��I2k�~ސ�B%��3B��4\�.�]e���
\~_�XF:�P��#����YV�)z�%��k�a޼�U�ߣ�04z9n�wG+���+�����%���rؗ|O�?�r����Pl}�})�BC�zZJ˺�q�R�dg�Zw������c+�R��|���f/���U��C�yn�`Q���Kz��@��H�MH�OQ����3�P�{j�X�������b�:��߃���nR=:8ܴ�2-F�����Ԩ�W�"�E�"��]�/!U�y/�\���U}����'�u�X�Z�\�|@Y�vh-~�_�x���
0�-|
��qJ�o���E�w$Q��i����R�ȯu��M�_Y�ʭ6ɽ;Oge�۶�B��RQM�5SʴvN�ph���!��vm���_c;�/C��j������8�G`�<
�򱃧ԑd�6iL��,uYb��B'��\�VZ����T�@x83�b�jkj>� ,�a��~Vc�f�7/�a[�WK�|�����V���=������TC��iÏ#G�ի�"#�q�+���9��C*����>��}@�J����!S�%7b�̾2A��S�];�Py�~��|V �gY�~�Q�S-��� ܢ���ȑ�{�4}޲�I����Qr�Қ�?L�9����̀
�%�;�e,�_|�N�2X��߻ #���6��pP��}(B��4@�������h�VeS���h����z'�i^��`��v�O����*�H��Kaas_RC��SZ[�9��.���Y��:wR��T_�L��E[��C� ��A�X���@4�a�
���`n���U�6�=O�=-1W?����î��^��6=
f�حK����-..?�i�eA�;�"�7(�ÊA�*��Wx��� 5��8;�t���{�qur�9-}�q�_ݧ��N	ol:*~k�􇰡-|�"�ţ���� ؃W�Y���rj���j e8�o�˧_s�Q�ي����n��+l�	�n�ƹb�F������'k��Ƥ�W�s:$�I��'��l`�`U�Vvl1��6�^��"$R��az���CXicꈦ�j|/{��#x?1�4��l%Y�eETh�eʳ�,��n
�y������uK�H`h���cjf����l�#�9X��J0�3;����KS�3��Ōeo���e�k-g(g�,@Qd�c6C��.��0Wp���P8X
^ t�5� Q�'?_��q��q��]p/��N~���}�y���z3k�AB��e�gw9Ws�|��g`aI��MtD�m�fj�� 3n�F��:�Q�m�`��5s���t�cu�'��?���q-|��W����͝����VI4fH�$�������St{Rl.GC�o�(p�QP0���4�Ԥ�w/u�YPūqovӑ�-��ձ�N�X;0TJ��X���0Ib>�`�a:�d�����-�N�����L���H�fM�����9�/J3�a��`^�I�=�N��y��P�����;�i�Z��2jӱ�H�O������`-�S�؆<�Q<�z'��q�~�~�wƏךT�֡�O��K-r��e���3�z]�� 㼈�O�ѩ/0�O���ơ���U�]J��!���ٗ�N�U�!A�?F�+Qs��=��j�8q�/���	~1�v��l��QZ;�[�Sc��L~�# �>�LK,\�0����A��TIH4H��&V�����S�3!���j@�W�����kN������G�/V_�?iK"���[��غ���}m;��c�c�)� 7}��ф�kRhƏ��%���@E��M�cZB��b�A�j#������-����j�
:ʚ�YL��O�$���ǖ�j�ۅw�mvH9�٥��v���%�}����*y���)*��r�q��[|��"�8���ݏa���h��s�	}���N�Ci�{�]�Z3�K5��mz���L���d*��]���ׂw;�������#Fd�7����g��,�=.<���+ok�j
ߴV;�`S�dV�V�6�.��z�x��[����`������*�n櫶L��>����<�����/濎j���RX�
Y�Ⱦ�w���m�
kZ㦻�C�ST��9���H���K�k���e��Q����N�<�}
Y$����S]��J?�NO��t�PԷL)[�Y��L����1��qM���8)��%R��))"�"���0:�Q�K@0�FKI�1F7�a0ꋯ���x���������{��~�$��"]im��H]#Rj�~���^��mk�2L�I3���q�G�T�L��=��CD����hM*��>_[>(`����Ŋ��HCOc<��F�7��Wu�Wq9h)IGj��:�Y�)�!Ă�rS���MvV�~��Q��tM�%�=W�Rg�����������5�V�x}�{XMܞ���B�z\2æj`���=�;%����IxV�[@5+��Kj�K? �\/8����I��!z�1���M������}�=Ǝ=����bjS͋샺mD�T������38��P���/뻳qR^�k��L���tS��p'��P���/� �޹�7b�~oi�"��/'&\���0 Ǖ�G���%���շ����ʗX�^j4�4`���ĻV��f��ӇWJ&��z@���1�G�1Q��t!�Vg��>sV�����k�D;Ƕ���]�MYh{N��)_q��6|r�E(w	�k�'%�*���v����N:��\�dLg�g�O��>ϗYLQ-�V��%�œ��8��e�͢���.���{n���;eʻt���m�= j*�cfw��SH氛�几�����.-ޔ\Ej�"M�Z}�R,��5��nsX�$V�$˷4����yz*PO��L�X-��{-�&�x_e�QB�@�ȇ�f	��m���;�h'�:�)�X��=�=R��|��gH���C���7��/�F)u�2M?cbZti�\»��m���e����ˀ�I��ȫ�|� -�6��׾�R =����1��ߜ3v��mB�ކ���\���3�i�Fm��n��=��7"� ����8��y>�Ɓ��Y4��t*�{x��8�����c�g����4��U�"��j��iT��s6�R�8
�q]�	��U-�.A�����5���C�r���=�}dI��zP�������U�͍�`�ۦY}-�j�G��7rO6�{plνl�}y�� �:)X��sr-�r-A*� T�rf<� ����!k��U�-� �>��I�G$8��s7�)�ڎ�+vi�g�w��Q�����Q?�R�?�;�Î��4�*;/�>�}zt�n{�%�tySFEBok˗�l�e
d�^aI���y����(��Aӯ]�b߷��2�>�`���7�?9�OӶ��l+�Z5X���خ��m7}�S�TMX�v]7�,[���b�ٯ�w�R��)�����n����ڟ�#*�,
IIМz�����U�$q:u��,�F�Ļ b��5I�'��:��!���v���4�3\ϷZ\m�I�Ȭ���I��q\�]���U|�r�Lw��J�?9T�!~��a�;�׉��	Nr&{Df�d���.��v;!��{�	=�f63�c�P��(�kDy3,��G�1���m�d��)�j�X�̛h7�?`B�[��&��.zze��~˷%!Yf򋷐i�8 C�{���U�E��K�7����W'��]�^lPFz����q��d���H�+�A9ی�w�5Y�-��]n�P��m<��W��-#L����2F7��#s�o"�+ey�x0Q��7i ������m	g����״�8�6�ac�؅��yn��S������7�V�n#�$Gv��|���s�.Ur�3�9��QUԀm����T�z���z�"��(cN���,�.6�yߧ�+��z��9γ��N����w�T�qZ̊��)�j��Cۡ�̯@���*s q�
f�7"�~=�6�O[��˻�^�{��*������@$l�~[m=�L�/�Z��M��}_	��_��4'o�P^	��`� &��(+Y�6��Mf�D�y?%O�n�ch�_t�@�-�
�%�;_=u�X�%��b�7F����?�ݖ�O�a���F�2D���\k�O��ϕ�k��^��y��{X�x�r�b��|d_�mM�9���G^5H\+���\/7]\�4�f�~ ,��e�3{n&���*���j4�ֹ*i��)�;�Q�c��ۘ緋��_]��C�8W�st����}���A:b-�|i[s��Y�ޟ��B6DL{K�}^Q�.	��r�����+;�;@���=�����4�L�m��D����M���.�Oze�y� c����6격3�)3���z(;�'''�J1<�<����bX!��||�&�[҆&�#h.?7W*�����g�pX��B�w?T�8��rrdI��X�̨������W�+�q�,IO�"�(��������T�_��1��2y?���7撑N;u�:���u�p,r)���)AP~�_f*H'���zUWLw"ڤ�� A�w�; �^��Ҿ�j/�J�z'���r��1���4ei4`_�*O�����LN�?-��ѷ��Iy&Y���#P�� C>c�6��I$����/#�Yȟy/���!���Y����R�|n�B!ϲ���k�0�l��R�9�ِ�{��X�s���m�iJ���̏����Cn5�9�*����)��y��Y���T�FoY0��Ol�A�!����ا���a���>����Ͱ�:\�" ��~����w��=����cYx�Z�1�M�H�6�ߵ6�����c\�.��HF��/���?�{mVz�Yfg�{�z����(�mZr!�y>�(QǼ��L���1+$_O@��p2h�@��.g�CS���{�w�H�!>aT�.<z�'��%Zuq���J;kx"���b�XeH8>���@�5��3ļ�/ۜ+��G��ݻvxw�c���:���阷&'{nfO��t�(e�����n�u֘IQ���y��z ����^�RCuu>_�I����;��[��I�A�5x��y/�ֆa�e�?�����<g�_�R c1u�U<ţ|t~��ɘ#�*,�u>�˗�a�}��s�n3�2tINǅ��!�k�m���M�I����F��-R��с��W�u��D��u���F�������-��xMR.��YUP��>�S&.����o�L� �oW�a�뵬
��0�z��E�m���4��3�xG�ti�|*N�e/5�Iǅ�����6�1���T�����Nh�uq�\b�|���Ad�5t����:b��itd�^�y�3���e�aT�2��B�o��w��.���ר�c3pBd\85��&��U���"�2!q$�� ����u�_�}!$E��`s�~ Yu;����*����g3���lU����x�HY�7���1#q��{�^��Y����חQH)��uV��!�&�6�lZ��M���&��2M����+G����c��H�與fn�Pa��C����u^�_z9�]��Q�W�I�Ǵ�E��>�ң���3&Gh\
�H_o�6;|�_�0�uq��y�%+��O�ڢ38R5�s��jcndM��-l�,zCP6�VF��.���e�`f���p9�Z,����>��vk
�YЍ'�J������f�J�Ϛa��ڑA�7�2�h��K��z__ΐo�e3��xL�h�|�[RRBc�5ӧx��ڕqQ�S==��y����CgO��M�m�H��MB�k�6���s��'�D�L,Dj�e�W�иԠ��9N����~5C_�����7/]�e�0�5:�����I����3��%�_�s��%��pq�z����w
~ʛ�M.*�1d$+�lRvx�Ej�C��U�Ł��^�s� g�&+]��Q����Q�R�%�т�ҭ$6��QB���x�dVG��5����^Wb�ti��oy},����. Kf#C���^��g�č�N�;-���5i���s27G�����y_�^�{���k��߁���eQ;Nz8�S	.R���$ᤍ�Żv�=n�L0��-��;����ׅ��g�!�a��J��^ ����	!v���Yl��0/}HV$i�`��8�y:ZKЅ?�q�!�5����{��� ��:�h]��1�f�������u�[L���9�]0yF�ޛ_��YP�@�-��S�(�&�v��E�3bݖ���~@��nm /�Z�N5 �b}��ثS�3i9�r�}~��ڗ����xjF�V�ϻ��N��SuEmaO���RvP���ݖTS S;,�^�H>heۜ|L�<��~5�(�7�>�G���Ʀ���h���P8Wya���	��I��;���YL@0"�j)\�6�+mn.j,��� ��0{G	��H�����/�EÃ� �l�?�[�k���������4�^)�V�"� Z��L4�����I�̬�s�3���9���d��)��>3fz���"��ȇ���4���&��)b�%�S�yp��%;#Z���V#���k��Z@�Q;'|x�s2qkV`=�ǪU�Q��!-N�7�S)�2&Zk�w��1O�C��#ɻ���=���4k;͏���o9�$�:j;r�N��q��$��'��i*h׻��O��(i(:Ư~~2"��v2�`r�C�~�_FKyܿI\"�y��v�+}&c	�ҋ�>WJ�-���S�#�������
S��9oS��{'�����(5s|0(�S���i���{�K|@H$2_�sz8��ڨ��D:�����w�xٛh;����i����Ww���"���M�ڹO��;��&��;���)U��E�2�Βl�&:z0����z�K��lu-�!�#m�ô�z�#��]�o�Y}]OWS�8��kK��2<9��穹��,8s&�6}TЬ8��W�p����Wk~
�wQ��N=��8o��oI0�g�
Z���E��>�rs���
��P��s��"��=�P6��zZ���c0f52�@5�pJX�@����	Lh�N�Ɍ���-�s�>�8�"P1��������� ��7Mƻ��
�� ?��5<���΅��NY�F��l�MP�̭y��5��y
vx�7Kɂ��s˒�,�?���y�i�Y��b'�Y��>��и
���<��y��{V�w�:ۥ�x8Y�^)�K���dn[��z- D^Jj#g�J���"`1\h|���U�&�U���n�b�c�3��V�K���%�P�mv�ٹ��|�v�tZ�c��HXR���%l�W{Wo��4u#&C�0D0� SL^��/;��-;���E���\%�vĨ���lD������f����6�7�*�q�i������ў��D"q{e���lB� .���3B��nd.�!yNQo+�6�N� �b���ڇʭ�X�Z	@Ri�E�Oz�'m��h��5�2�Eb���sT�I$\����C�_��9���3r�{�Ag�������!JH$>�=�c� ǚ��.�q��EH���K�Ѽ�vv�������s��"c[���E0cx��<=�������-�Yi]�/D��f��S�[����gIjO	0�$��)�+�iî����m�n�U�3C��f�� q]�U��l������S��g[!���كW��5>¦���b��-���U�=O�|��Xy)i�+�st�٦�D[��{�{!���I㠣m��|䳑�Y��sS+!1�z;���c���ov��I�B+��z�~������G��:eu�A�1���/93i�^|��>Y��d����� ����.:�����N�=9�Y�ď��`���m��ϔR�:D?���}
�0�\�r�/��'�x�[�����VK�&�/߃Bo�>`�8�*��0|N����P�4�m~Ox��j���D�M��dKhS%�6��
�O:�K��D��_Q�����A+�:IDHasE(��p5�f�f���8���}�r��)��'����ŕvAn:���"a+>��ig��4,\ml�]�W�J�{�0r�����%������ϟ���á�S�<�5�+�s��٦�H�8��QT�����3��^X%�XE'�r*�B���t�h�7O�e������:�SL��|��d�b�e�������D���#�Y�R��pM�������7F��_ɅDoE��1HT?)l�� �~�l����-̢��Ha`w�IC핡��39k?�tn�Ok|���<�V�O��ҩ���{��qW2$Ș$������0�Ձݒ�,<Tԝa5en/U%�P+9�m��Wdf9zӞ��T�� �ۣ)3�.z.f���cgc0(L�mFy������w��z\�oU�蚹*[&�7Җd�v�,/� 	��M���%��^ p|u��a����Bj���9$�]ԤQ�9iS�.�M��H%�}�p<S�rᑝ�\��G����9�%�E��%nխ� c68� ��n�����N��&���$o���U�C��ڣ�/¨���*"�W�ߴ�J��]�6��쾛�}�&�$�*�Ϲ�yk45�f����lx&qv�
)��%~��zG�h���H�G�ܢQ�9ܡYq��޳i��N�g�րm��Ja_���V,��.ز�6P@���7=���T��^��ɾ��런�ݝ�.��:G럏��
��*ͯ?�f۔����z������ŞLz�*�sP�Z�ZD��*����+���S�!�n�HIoFZ�}%��t����w �x֒�r�/��3Q���݈��l��ɠ�'p�'��a#/���x�x#m1�ZHz�����k�7y��w���Pk��ů���Zo�S4O�����(����b���o�R�vTq�"�d=�;��Mu�.5,T����O?Z��i٩_fǗ)h3���A����J�d��������F���B6	���PH���֌)�q����%C����?s
V%<M	�R�4M�	(�L�2R�W�E8����Np��>�6�|ʖ�b�W��P�$�nb���bVD?�5����W�<�#��N�G�҂���R�=�VFF��A�{!>�V��	�x�3Pϴ�zv?�z����l��bY�e��e���3r��@��*��]ϤM��w>�Ƃ]��NSS�5;y������G9W�G]�ȸ��=����(KWAA��Ӆ�;�iaq,�@�rL#�7yS�|�����۹�� �!����M�����$;��Ë�E���Lo�������_�f�av~�[w��4.���4��U��,Z���'r"�"�څ�8�d/���+y�ȩ6a�l�|�<b���a���+?��Tv���p�W�1�2b������.�li��6,�󋜄LU��@g�Kk�=���h�]z4�}&3�� A�FC�.�"�oV�aȽ�#�,�ܽ}j����]h�E�>�(��>��J뜜[{�L| �c��>@=CV̹��Lc��|6���_�c����I���lǧ�u�2g���b4�"�Ԙ<�1>���a
���cC@�d���XL�GO�7�+2Wg�%�n��c� �Ii�dN�.B�F�_5EO�L)- �9Ae�LP�W~k<Rd��PU��:���	�W�[&���
���'�x�?Ak~�������A�7~"ծI@!�V�s��@�9��y�s־���ҫ������;��� ��Q�V
[��8/A�5o>M�V6�2�bڐ]���x	��n������O���ގ>���Z����M����T2H�|�ۑv��L�8���i�y������ylz$`:���	D��/�mя\k��~6Y&�A��c�}&!jQ�r,�뙴�H��rز�V�����h[�N���	?�_���Q��EȑH��Ǥ�p	�Z�4��A��>�tc9R�g��맛����*��n{:�-���*�?,������� 8����<Y룢���(���"i�5nQ�7��)�n�2���>]�@�O�\������Ԃ�����踳><�ʴ6�JUԗ-.�)v�`/'�[���'w�&��fd��~�<�^]6��4;|��^fJ�>���Y�')�33�����b���<)�U���~ŷ9Q��93ɗ�y+��+6�_��̾�1Q��6~��_]����U��2�m:C<���r�|8h�*��0�7�%0���w��(���0���Ű*���{ &\'��Z3�����ui��+��!]�&R�E먀�ϸbg����ՉpK���*����@���ŀj������I����.�#�����,�ǯl�=��϶��zc��B6��0	X��;��o��yt�i�;����b\h(:�I���>�K�Up����[��n�LJBY�?kq@������|�On[����A��"��,�-1J2%;*&�0�rY!_rs>�.hG��Ӄh�w�Y��.����vo���3j#XM�x����12�/�oX=�Q5�ߙfO�'�@tk���}�)r��#�铟u�{Jm�0�����l�v&��q%@j�/�˚��*�mL��Zu��E|y�Q�9�(	�Se�tK�~-.y��&s��kf�5���Ռ�'�uJA_�\�����˺��O�9C�Rs�*��|��qئm)h�on��h0�zz�y�d��\w�sl���}7?��F��� �r�H�ix/�rd0D��=/�\�Z?�!h����v(2xL0�з��H��~E�~����p�NiΫ��2�����%Y�ۚm���^�&<�C�ACC�������/��N��Ϗ:d�$�nI�5�_��[�������!011�k,�gAfI���+L�i44������@2ᓍ'�O�Gjk��G�Jn�u��|�q�Glb��b���)�7ɥh��W�=�f`�:;+����37/�t�M�{���XK�M��H��[�7W��Wi"�m��[�A�X����WI,���O�H����6������;���⃚$A���?=
Ꝯ��\0?w�Rڄ��~�ԉBƑ��wXE�J�{_ס������N��y���6J�E�`a4>Ʒ�e��?:�)�҄�� �R'�4�g:�TA9�|*�^ �r��Ls���zK�j��	 ))���3�g��^�(Aw�L���؟R�۶ʵh�l�+Y����H�T"���Ѽ�� �Js{�\�#ONN�Y0l��qԵ��ǭo���Z2�AR�,e�ǮH'��T5����������م�X�Y������Ϙ��s]�WX�W�pc7t�>���N�"�׫u��X�h����/���G�E0�K�骈��;Y��c�T�Nn߼uk��S_��<ޓ����n0``��|idC�i�Ѵ.�?��9�̷c\\_e���e*�������*�P�ޤ���}O1�Â9�����%�y����»��@s��J)H3�({]�r�qBD;��Y/e91
>�Կ�n���q�|ً������&�_�8E�ggh0�u�߭��
�R�+q^��E���w��L��p*n��+�<]��!×�&��B}�����M\�Aں/2c�f�m!Wl��Ni1�>���c�vT�z�o\*'��Os�(�����IK�8Xl=�h�\�Q��β�W��]��+��![�Y�W�D���4].��R�]����U���l�V��=va�GT��&�	��C���T�]���kpaƠ�-�U�V������B�υST�&	T��O�O�L��"@`�s�fx��F�l��U�
i�4IJyi&*n*�D������M��FKV��μk�Y�,u���33,�)آ�'<"�¨~�c���T ���M��V��'�?y���g��-�h�!e�^����SƏy�8b�������;z��D�oF5{�<v݁���fˢ�w��=��;���X���?4Uh�N"���{�Uvzf�[G�sR��Z����Q�,���B?��D~�iJ7�mɥ�x�ѯCt���ă��re�Ptu�b���)�ǅ�~���SƁ�:MQ���������젡�z�Pp�tt�|rڟ�m��\�Y����wл:_��:)��xF��!����Nx�g>BN,{��C�л�L���J�0��)�H��	�[՞��~��4�١�9T��Q^[�d�Y��j|�|8��n�� ��E �?G��<7,b��c܄dM�gLOw��u���ӆ��ג�f	���Gj��g��һ��Ţ�]�(��]���5��TQ���F'�caC< �΄@+�{�I97��H��ޠ�>k�ڠ�56g���XN&�^��ˁ���Q��x���rR0{���Ѥـ{ò=��>b#�@-ǆ	�z ��K��=��\���������:�(�,۠�������'aE���ܼ�:���]dß�� �k���'b�/�x\@���
�֬ճ�������,��O%8X�	�z�����W��&Y1��Y�����î�H+�����^�8���]wQ���;�(��/��4{<�Z�J൙5���H�]]HQD+��1�T缷ک����!��g,0wW�T��v��o^�ރ�v8?�0��5O���`��������z'���1k6)|��-����������i��I��2"{�5�V�_�ޫ�bYȨ7���6�M�2��m�l���<�pRٯ�-�f�#�D����@����k%{�\K��n�N��7����힥IjR1�}�6�at�j��V�����P��N��`w��t���P�ʿ�Ʌ����n�f�B�����bg�O���_�J�t%��[���R���x�ػ�q�����}_tM.��jh2K���ėe���}6��xp��L�q7�xЭ�f�x�#����&`oD�ۚ���Y]n�F�&1Sā_Z:��`���Y!���n�ǭ!�Y��'����Jׇ�R��Ҽ��ge���f7L"�.u���$������}������I��m�k��� ś��)v�����A��!� Tmɕ��ə�����+��,ꏓ�����%e}e�zo)�������Juvg py(����+�QVsS�d@`�g��io"i#��}(�XPk�;�U"t{��R���W_m(�ݽ����v�eх'm�b� t��qҜ�k�N(�K�t �`��=|�@~����J%ʁl+�Wj%�+�(�~��<o�6s��Nˑ�3 ��t��~�S	_-Z`ɻ��"��Y|ڄ���#�=���-���@����C�C�9�����2�qsȟh���o̾G�H׽V�n�� �5����V��H9..ߎ.����@�)z�?z��`5���ɡ��z麟#�$9�7��dJ���쓊���S�n�	�\H����D���Q��9�6L�jR�ν0o���s�es�8���{�7�Ǽ-H�"�@����c2ls�q��<���̣�C�y֚�.�Z� w��~�:V�iB�k�+�ř	��u����wq_�_��ij�R��d��6�_�q���b`W轿�Wb��}ŧ|��hm���H~QY4��Q��҄p?|�����W��m��<@�+�>v%_99�Z��uҘ�+2g�B�ā֨7x������p[s���2msю�,}����dQ�{��Z�`�E��Ϗ<���T�`����s�wR/Zeھ��1���]D�5D����=��B�(-���[��Y��=�����Gr����;Y��K,_9�C��[q��PQ��ܶɐZ0��q_޳�1�$����󛃡~�	����
�J"%���9D,G��Jǃo�?8hIHb��0�ha�s�&}?���}�n��Qz4�����G�]�X�*��@:�9���]��ځ�����iv���'�j����'���1P�d����	�K�+AUI��7�����}�t��5'0�r�%��7�'���M��5�^�8�l!���5,@?���������޲��f���f"4m��nŮ��VZ�
�R��K�uI��Q�bd�I��ݻٜ,�F�3�\��e��0x[L
����l@+�M'@%�����Sg��6X�Y41��'���h��s�O�����pL�@B+�\� ��z������ۍ4ȥ���������%ϴE�5{�'֯:��Ka�^0Y���/_&�a�n���aެc�~X� ���ʗV8!���R|o�״_+�.�7!�a�w���P��b�_B�*COK֬-��5��y�K�@ɑ�/L SEoJsY?��'B�r|ʔ�MB����՛%�?�<R��[Y��)���!+B�tk�2\)���~�1�r�����G���&_��[�7�n��]���
���%��s1b��A:е{�J���'��#���0�6>���#+Õ��Y��e^�AiZ)i��Q�A7�wTbc#ˁ�),ݭ^��6��@������jm�(!-=}_S�b��Y�����ϧyS�e�x#Ekང��Ox�X�繿���=uD��-��d�o�Zg/�Ĕ��Mu���mut�����e�潆�l*� ���N��ȵV�4<�����7i����b�$?u�i����c���Ƨ(���,x�6Yi*ΨL��Nȿ���%���b��rt�/��v�I}��b��fM��1Dv��J�~^����U8c�KtR�Nq޾���&8/Wu��W�~�/Q,I
�O�M�(ǎ��>�I����?=���h>�E�'ᩡ+"\����c�Բ����[�����U�՞����w�_���H��I�8�X�E_�r����eܟ@5���EÚ���w�>trAt&&&TTT�ד<����;'/eo����clp� �����U|��r�^�`�bo/���r��
����fX�{��B�Eg�\��QRQK�^�Q%����(A�[���v`߬ѓ�}�/�:�Z�M'�\�jX�-ʺ1׉Z�aP�	I������dZ�_�bēy�P�&����+o͓��`���2`�����*�jy�@/#��*����	���_���Fq��)72$�(����L��$h�h���*�}!.Z��4;�� g�tz���/=��b�ł��n(r��H��bC��i�k{�����xؗ$��Ό�����Zz1[RR�/�Ӊ����N��j<w?�76�����m}O�(iM�$c�4lv��xa:99]��u�nmm��T�Z�w������PL�	�ϕq�5gI�_7���m�}���ƴW���e��ܕ=��K���c����Cw�,�aq| ߧ�`���2�y��+��i�䜈t��t���t�&�� �~ɱ�Lw���I�'�(q�{-0�Ν�d����oWI��B��p��w�6GֆB~�<9�Ώ�C!�X��o�DҢ4��B�s������X�wAHC��{�v���+t�>��,Új���r&uglܺw']���G����\}��ި=!�&/� D>A���ߧJi�*U�a���/�8�D�ar�ÿA	_��K�<ل�P���K��
X�yNN������l�靏�+U�t���U]w���\�^*o�¿a��/z0�'8�Z%Қ-�%��y��2�߽�]-�ekC��Ȣ��ȗ��!�!$97���gg�H�e5E
_��tϵ�~���]f�-R������`��O7��e�ɥ�4�T���9�ס<�����Ofv���e>�fs���>�5�10o!��{��\1I�&ݸ�a�3�3����3M�I�������y}��*���4x��h��bg�5��y���!�鋼�P�����1*��ôP�z2Cզ�JԦ��$~l�䉳�k��z��s�M5P`9�����;���U��n,+��w��k?'%�����e�6��5�eS����i}�;���������-��B�@�-:�***��I�P�I�2�<�28��r�>F��M]�w.��k��Ƥ���+�'�T�Dh��l����UT�s��.�z�i�b�ҕZ�����9�;�:��\�N_|5>�AV�Qύ�?�{\�q�o��f��UD@bY�-͟v4=re�U��p����?��c-n`���A�[�/�7�l����DԮ��KJW�A�U����L�� =��U�����/�Uf�M�$�q���'�X�;!��u�.}���;g�.����Aŷ�:{�N�L�7�1�=�4�*��h��m�x7�,IÚ���7x��(_��O0�=;�xѴ���#��m���LV��Օ�_f�؇���o�!l�3�ey����ϴ<6��p�[�G����=������dct���%�vҩ]ME~�l�x��d&"H��6��f/�\�0O��"H�r��(����oN���qa;�Fe3�����فi3zΨS�Cam�c�[o;#�$)�;oK���{�rk� �E��B�_��.]%#�Ր����op�b������w���`F�XUz,d�d=Y�MA��U9,Y��
�i*����[��
?nE٣����l�&
Hgt�X���dzr?���YT�}5��$�,�jK�q� �X�0����9�յ
ʊ﵍�z��#,8������[�}A��M2��Rx������a����h��8�����t4+(-�N�q�TkQ6���t'I�(��V��u�o�۟@����	�����1���%IIII�38Jc:����6?��}������S��=�$��}���>% ��|{a��OK�ge�
�!ڃ��Q�:�pw�(��+�����6��6"�)��(�/��;�ے��urPn����D��)�Dn�����b��z��B�Sb�VDe2?u~�+���J����!����$\"\�Q���ř�ր^��j�B����Ʈ���ꃜb<�ޠ���XK�}E���Jc?�cW�}�$��#E�=��]ߛ�n��K�MK�"�	��nO�E6E�'���
���h�Oag��s��穤T�>�y�ƒ��JCkJH>�����$䭇�"��Ի��Yn�>�.�r�/8�V'
����;����3��[�t���w&F��[�?�/��e�öb.�ޤ�[��>�[�-�
� ���I��.���	M�,B-6_^o���L�#���kЙ$!#9oiE}��'.��-��g�$* P���m�z��  ���/�!~���ET��M�:������F�� �ae�@B�ٻn�/�Zo�ԏ����cL�M��Z�;M��P�/;LS�@�F�*q&N۫��S��s�߄��b�M�6��7�\_mG��?}���.ķ<��̌;b{�c|"E���%���1��	?w��k3���@:��}��v��[ca���rK���1Vq�3R�D3V!��y|8v_��q�pm(R��;�!'��_i�h�`Ӊ��u��6��!p���VVB|�
e�v"�\�Pw��>Q_U�4ɖ�����4#�����ᓖq��
&8��Y��4Uz�p	^�����U��*<�u�᜚e;t����C����
�����j�$�~�F��T*�+Z�֮�J��ܷ�N�o� N�ԏ��eY^�]�Ԛ~�ؘR���`ȜS5�/����FXklf�S�������Ӏ��Ml�/�Ы��>=��oMT��l����r�s6�Hh�(Y_�թ����"�?�5�h]m�?���\�Z����o�Ŗ�����*�lU���ϐ�W������,��� ��4��.7��)�)�1/�ƠUtQ�
����C*�#���=%�K�P�'G�,��/a�M�Y ����lj�~�l9&�l��MV��&5:�N�ѡ=_�}$��Nﴣ1���_��7��Y�F�x���|O�J��:�k;�R���������`;����66���>���`7˝O(^{��<�ۓ�����U�௓��*�B�^�q��9�����N����I73��u ��s���|"���NM�c�ۨN����/~�P����f6��ÛR�LC��A�Y��*����G�A�s�f�����e�G�䌱�h:�?����9�5c���5g���%�W_$d��N$c#2��h�
�DX\���;�>�rĚ>A��Uq����:���
�頝|� J����Paf�����'���*�*��c �ٜ�	�`>���f�F��憟Љ�����g��·J�����@��瞥�l���Y��dț�D�;�d	ݼ{���� ����o\��4^[�S���?Try--�4>�����ƵFAmm���{F�?��F�vvw˼2a/3eھ���'��.­?$�Ey�r��±�x2�_�;�]��Ѝ�/L�h�~��[�����f�z�>f0:ϩ��L�]���my^�a�s�,vg��}=�"±���A)&����#�jP���uv���Ez�p�Y���'��:[s/���.=�p�E��=
�q SRhQp38�3�I�͑SZ�q���%�9�h�Xô4�'��up*^�R=��"��r҄P��^W��h{�e/�F�b���Ks��*�o#�HRE�s{o7N=��~ؖ���I��	���‛-��������8QkzN��٭	��d6tz^v&�`ܹ��e~p@�X[1gX׿= �����ޞ���?����oq^�%f���V�լ�W�߿������]���������S���1��Qm���8�)�R�w
����wEw/�)��]�C�νg�/��/�w��=��y�0��1Z���u,������a3X�����:٨��O�^k��솒��y�����<�>���&�d�A�m�C5�nOş������J��T�B��CP�_-f�CvZ��'Ũ���I.[|P�Ķ1v�����d��#�#bC<� ��t�	ۓ*�<^�Z���M�ԌZ�����g�$檌'{����{�`�����D��,�k�?�F]M�eFw�.d'DC�I����@O?̠RG:+�T�
)���h��|�w9��}����h��u�umr����>�CJP��J[F���[}����Vp~��l�{��ٶ-�����]�!��Z�������_Ҧ5����/f�m|÷�u�� ��Q����A χzs�|��z�*�O�ը��,7R�����D�[М�`���\^�D�Ed�Zzѭ|����/}�����������i�8X,��>t٪Ǘ����4��%���m���	���Ĉ�]�8�$6G:xLXn�xPE[�J���b����Y�|2����Ss�Z#6���ݩ$�+ڕ%LW j]�0k���S�~-{����'f8�mE�f;UDw;�:�[��F��`3�N_$\3�@���Jwu����2��y0dc���p?�����,//�Ɗ��2��Ӂ?��l��5�[�뿔u���]f�T�, �OA��>���v�d��&@w��O1�C������WU�w2wJ�Jc�gTy�<gưEf��g���%��=T1�{ԑN��\,�9��B6r�Ǟ���q��ݷ�5�_���(1�V��W<E��ր�k8!c-a�h�	�oa��0R�nK��=�%>�M�w�f�lV��S�Y�]9�f�#�`����{�ScW��(��+֗vq'���у_c�\@^����h��"]2:16���
�F.�'1yr�HZ��;:�^��VOT-!O��JY�{��\�Q-XB��/6���	9�����m��[�6����<?Y����r���-m��Ym;.#����Ûy��f�|rjJ��C3���F��;<?�I&}1���)|ZT�	����X&����VA��=#b�W#�Q�;D�4�k�ċO�R�P䲼�:�6::�ҙ���`�&��bm�ɇ���VvW��v�7�Lȴ^´+��f�ؾ��C��]���G3�"��n�Z_�>�uu~�: �M�$�o�=ɆP-�ʙ�C��j�Q�C�Y��5;0��6�� �h�ƈƇ���xH
�t�����D��� �.1s�H/ �\~ρ�L�03KGܵō��xiGƦ3kU(��w�#wf�s�u}��\�)Z_$0ͬ�Ӿ��\"a�8�����mxv�̿�b���x�ҍ�Ņ�������k+���^��Uo��7�9��_E� ��`�������/��8;c#�>i�ֽAt��^�U�E���i����l	��6��=#Fsd$>�RS,�_I��gV��h��m͢]�G,1���z�!���l����lܮ���9�3�~��fn���z|�����&I��X�F��^3�Q�.��I���N�|R�c9=�i����V',�@� ����PG������n��g@��y�K��u�����8��z;3g3�����-�\��0����׹�k�;":��cv���b�D�Dp��(;-D�
l��]�0��ҰG��9�S��xƌ���r�ۭ&V )�c� ?)��U󲽜�IEbO�*���6v��������7_���������J�}��{��Q$<�2~�

�kO��зv�r�� �]���/A�Zo���{U<w2����=���E�@������%�Yh�����z�����B�x0�3�J'���:&~�ݥ؎c�������+�@z�p��f�Pn/��l���%fr��	����l��}���0;q���Ϛ4�e�Cx���Lc�LB4C5��c1Dv-�5��j#R2~�m���ɡ����?�;�4ֿ$�k��O�h��s�Y�����:Z�}���'�uGO��>��x���jmsh-G�]#��uz�+v����sO��ylw�ܨ���u=X�v{�5�B����H�������|qc;��?���tg=-dm����� �WPzŞ�{+[۾��o�K��U���	�"�*	�B�w�xb�����Ȱ�ȭb�Ö\q1'����b��9���Kو��XTn�@	�]n�w�L�;�Yg��q��1-&���ӗ���]��p^�S��kw�Bn�u:��\����F��]&Jt���׷���qWVr��ul$�u�d%��sI����Qb~kw㘗�Q�:��L�'�Pg�=��i@Z2�v�O�����ǏbL��	��m����w1SM�A�����G�ߩ�Z{|j	�p��"pm�|�}t���I��G3x}�C�V�T��QV�Ħ&��NX����
���������WB?|낕̎�E�J�v�Ը�M�3G�̓r���,}�j̽�a�Y+������uFGGk������wܶ�n<ݮ�93��l������]��f���kLGGw>�r'����v��#�/����:"7�K6g3�(l�6��s���OZQS�"*H/�c�Rk�nP�|�1�XK�-|Z�O�� �9X�Er�i/.����m`�~����7�|��y�el�I!�����A��웋�2�����cy�-�r(�o6��8a�Zқ��՚�M��ԛ#����Kc�},L�bs�ab�y8D��ƕ�r��%��r#���>�L���ݩ���gPt���s#��gvBpi�t��r,\z?����K�}�ݎ��Tk�DgH�ߠ
�2���ʫ�fbN�½����P���Ԯ���������mB���v���e2|��`���s�*���ƞZ���)`_�j��A�J=�Hʱ��&��ˣz��ëX����WNN�k�f=�%���B�=�`����k�����:�?����1~������쏡x����ZL+�-F䙗�c�=:��d��d)��^��sdt�Y���Q��]����ٲ�ak^O��G�Tp�PP;6���o>��@PB��C~��=���U>[C4��p-�+Щ���kl��|��$���~g�%��~�d�T�#��1hD����)�t�s��m@��*IY�9���\����cF��jS�7�]F^�tur��b��KS/����~b���c<�b���)2?ÿ�5�`0�M���zYR<H施6}���*�9>��ǲ���(v<��"�P�S�润k��C!�v�����FJv*2�"�R�^Tajcm��S�+l�U��}�/.z�jQ�#�_�M�+S��b�]�߰y����y�8���6ⵇ�hq��Nq{�tJ�>˗o���U+�e7��/2׷ �)d
�^W>�e���+ͼ�玦�l��S���<h��⯬���B7By�n���K�!]/�NV���t������@
T�frIgl�3�����>�Y3���!*&�Y��[���?��cf]�06�����9u�pf������� �Z�ԃ�^�Y8���1K
e>A����Lx&!�7�b5�E��KGh^.�ƍp<�{7յ�@+)�6tϲZ�=��h��"B�Y������qoX��WOk��щ ��!A�=D.X/����¬����3��!��z�Dwr��+w%��rqg�`�������-8��oQ��ɤἝ�>�`W4A���e��x�q��S�O�MT�LA�iY�� ji������Zy9���:%�Z�f+���w���������u�DSItEm��$���j��6����
$�rk
d�6�N{f˵'gg�\���1��8/)�/�V�W�%F6~�\X����rN�-]���b	褗��A�Tb�}PEM�]��A����g`X�Y5<�nCC�&���A�C�WA��V}?�z���%H�m��%$"���X��U����\A���|Ꜯ#B̒v�|Wzʠ޳�e��^S�� t�#�U��٧9R[��[��0D6�e�>d&��a�ha|�x\X�x��n��sb,��7��ǆs>;�U����)���+fC`\��V��B③a+~��=J<;�����p�u�6�F����E�>�����6�d-��� �α}���˴��4{	��y�)�)���IݼQ��B�l���ej��w��.M�6��ZS�΃n7AK��[Tv�@��2����ȶx\�|kp��tC�>x�6��Lɻ�kΨ�=�]"���v���"�5�
��#�T֤�5��HuW�ˆp�(����J��������B#`Ygҿ�y6,q����r=�j��M�b���w\F��ǋb1\�/V.:[vE��3.�*��*Cqy�F/�m""Y�����MY�����
�f�!
�y�Xu��,��ˋ>�V�o��z�=�	9~H������a�h��$Ѣ��p]�k�|�6��v���}ؒ��?a��J�`8x�c>L(���Ɯ�.
��9ݹ|���S=���5wM�U�5���PY���ExV(��/=����~�m�n1�$h/��0���I�c����B�c����.�ZZ���1'T~�3�*�5��V/�u�>fp��K��) �a�m��a�ƙ�&ۛ�68�a�`�ה��M����� �E�*`PC�ɒZh~���;)���`mԥ���H�\���qn%��4�>��y��S ��t�<
r��=�Bba9�?s�t�)����EO�0+>�F+�����n�����|�u��4��3a�௥�q>�1��c����Iݦ�>����F렙���lF�nn�F@�^�)v(
���T1��sv����i�����2=QGG�(�ޜ`ͯ�bg8�D //?_m���}!�|y�?=��薎[_���;������Ӓ8�m�8��!2!�d=f|T[s��VR?k�eӓ[1:��'�i�xqs�8��(8��7�\����F�\���L!iNO�=�s���VH�s�2��~�U�������(,�8:�݂�z�SO�s@a�����/b�e��~��tˣ��mi�i�K� ���,h��r�4���CTe���W���1�ќ���-:���4|�#��㳌�zZ��ŀ��#�0�_�dG�j�?EݼR��ѓ�����y�b�ع�"�h0�L�b����a|2Sr��|:y���>��������`��*����1�_�0Q�w����tކ���_g����P�ڱ�1e�X�&z�r����X��MS�]g�nW�曝�1W���� ��j��w�_��.�-###WۭuX���L����wd�d)��q�WZ���/���n!%ǣ�77��k���'����Sē@!���1��'j��j���+a`��;j�瞾�P��q�6����"��Q���r�Iq<K^��0uw��n ��
>1�Y�NvY1�R"�,�Y��zu�@S'3��
�/ܼ:�x�~V��J��[ƞR?�$[3�1|�@��Q}�{�Q��;M����V-�iq�����ؑ<mU�, �DHxcܻ�I���ϕ��ޗ?�Tvo�k�Q7O𡒟WO&7F�\�A�̳*4�j�ko�a���2�\��ۯy�b���t$h���Z3�=�sV1�x���f�x*i�[E\�ϲ�M@�;�CW��Ӻ��z���B� KΣ���_�Ɇi�P�I�o%�;pR?�]�5R�^z�uT��Bjj��k>�2���O��d7_�� Uo�$��Ap�
��	�\�v���Ԋ�Z���X��[�r����imKM�W�rMBY
����L��}�8��QX�U+�v��=j~��C�!68�ĸ�������vY§��^�������)���/>v�A2W(�,����>�tA�iv_����AxR�U&opL?;�p��M�5!K-_�Dk�8]����zr�b��G]�<�r�6��19.���~��q $c��FOE��peQa���iC�`[��N�>��}���n|��A�F�,\��of�����ӆWU������G��	�,�f�k��[���n����-���(E����
S^�-�
9�����B.��f��������Ɉ-�Y2]^T�rvd9^9�D�1�}�v�#\��;�$V�>;����j;���I�^�O=�� ��cc
�WE"���_hj�}��Jk��t�k�q���C���wGR$�6��?v\�n䄒�)**��\�	�2� �4�i��!/�ȿ?�Ujc�j2#�������Q�_�hj��W��'1T�d�;����A����y��y�PS]Y�\ۑ����+zk�+��+����R��|C����Ib���~�����(�Bw�Xyj�BTհ��ş�D����͒/B�!�E�C=��^q@��J�Œ?'��VYқjxEQa�F��7?J*��_%�ɉԆ��y�z#o�-������7���(��a�`��g���Rz+��W����l}5����u���0�E��{e{sȋ733I�),��e�kb1����A�U�����/�}�����@%�>%�c^6�bT������b��>�Vi��%���hRx"Щ
�Z�����q�}�x��)��v Y���I>���'d��S�X�pg(�8��u����~^�n�)33���?�6���rr�5~X"�U����K/;�7=�HX:|Q�(���U���qBN�:���w�+�RdWX�3?��'�Z���ua�?� X����Q�7=
.�hP�tH��E��nK|��� �H�
Y�Kq�&y�����^y���~����ѫ��A�A������
?<>(���m�c3)������
�'NzPMa)"¢���n$m9�/¯����}cm��4h���G���[�r!��~nN�[�a�͡cS��g��;��I!AZ��W�w�6B�950;��\��;�=ŝ۱r�z��~����y�xo���)�ԆQW�7X��N5�%t��HZBlؕu�+��\�<e�!��VY<8�{�+�5��ܙh�q�x���K^��Am��F(E_W�h��^���&�@����ci_�s�I����/��F,燅3͛{zɮf_��x����a�2 ��T�$8\�R's+�;;K�^���	l%�-> �U�;�j���0PxU��p�(Ѱ����7u��$�k���k�R���}�bB�L��������O&�sx%����R�^�b�#��(��x�{L�k����/�>�BN�[��w�z�'kvWB�+x���Бm&�z�L�,���<�hI#����ŋ��c9���
Z��c'V���oS�93b� �B�ho�hٵ2�4+`"�<%�V��B��P�M�C^��B�{��6�ЦE9<��X*���/v> ���A�3�|�YKm!�J�
y�o0�'�95=`�����}n��PL�d����/���2�'ÒN��sٻ�bn~�p�5o�ג8z�\��� �EQ!U��Q��K��]F��O����f����3��G�	����� [y��g�_?/��xu���x�wJ�R�z�?I�)���UhRps,e�Rc�S��)1u�8Bmĸ�ټ����Ä�&m�nOs�&R9�C�hQ�&�>a��v���_M���ry��{��.x`iw��ls�w��W�|���ؙT���{.p4�.�[�����s�'c�����Ly�'�8�{]=tT�b5�k��l�n��)��G�xŴ��a���8k6�]���cz]�o�h)���v�Dz[oTVD�j��5Q(�-8�o�ں$��)Eˢ�턎������&\@�Gqa�/a*�N�#Z8��c��]���ʩ��Nz&���)���K�.�z������� �����1�RQQA�+��1*�����gR����A���;����ۭ~�g��a���3��{p��B��+�y#���BK/Y��ͥQ��p��"{���!5��0�2�4|4$,�-�Mâp�|Sp���(�Y2�>Uk��P��]�ݝ�%�_I�qL�c����R�w-�2��?0��o����W'*J�Z��cM`�H�(�
>otlm�V���[$�$uM��T*���ě��$�՚���n�����[1b��F��&c���d���oȄf�7��ʦ�x�;:�EI��ѓ�j�Ӽ&e#�7}�<���wg�Wh���;k%�ύٝ�=vw��3K�h�k�81<r��0�\('�Gɻ�Ab��Ko�3a�9�r�P;Iu�9�BT���#j�V;��B�S"�k��uL�}&O��~�?��s�&_o�5��m$�&��hr��v���b�8pMu5�+����|<���?�JD���75e�ե7��y/95�ʙ����ֻ<���}��в���bC�_՟��g�\���#�o�&&9rKgHj�qo#Ҡ;`��c�0��Z�T�����D���,"��ē��>�g+���n�	��QՇ���BDwS�R��p�H�> �����v#�{����[/ªKO��<&ˢ��:��p*Vy�k]V�~��Q�`��3�U&M����j�0�v��9��$b�8q�`��X2�6lL��FsU_t�Z�R[U�g�8�Q�	0PQ����P=~kR�[���+#�N���OY_�z�f�=WQ���6ml<K���ey�����K����D:Y���è+><O��h��~W��%����>f3���\���k7�4T����>����a�E�ٱ,���gB������.�-��]��X���'%��I,������q��c�|���{�$�7\o���]�j��ɤO�� �4:�ǆ_��.�=�%O`Y[Qs�J��J���攕����AB�L0�
H��Mа�4�T�G�W��С!EcK�,<� ������N�y���oZF��9��IRqµ���c$A�E����^Bg��b�U|�ZpNI���}�Ksr��j�P���5gn"����_s�Y���}Q��1��D&�gm�gjI�}���ؕA�zsE�Xѕ_`N����8m2�g$?@w%��X��Mvdg=�w�lKQg�� ��%9��C?7_���I��-qJ�C�Xj�~;'O��/�W�n�O��l�5�C��D=dEA�k�l�v�����E�B{���H�\�?~�*���"���n^�Nb����6���.����z��+���5h�o�����W=ł�JD�ՎGdff��lQ�>P���'t����B_SJrKE0��}Q%��^^�T�5�5u�W�UrC�������p̢0>슏|Hߏ��^�����q���Ý���Xn �݂��%��ZF.���.�=�wR��[�<k�^Y��=��[���^k��ph�2�{[�8Wo�q�K��fl��P9�Ԩ<S����U]ƫV���@��!�8�ĘE<d��w(s|�/�;x�d���n��U٦>�T!���R�lƁ�q_V�l/��qTB���O6�ؽ��L�nU�^p�?�u��	�LZ�\n��P���yY����J�9��$#[N{�i���<�� uE�$�PeL��ӆ�}"򞅤�.9�g�ڸ��Y7�$\��n��g'��yB����B�b=�0Wa%3���	E{�b����_#�[1"�G"0&����s�,�c�g�	/C��X���&���y�&�D�{�V�_�2{��_�VlR���}3�C�P�s+�za�6�	�G{��V7]:^�4��#Å��D��{5� �ʄ'T_bHqB�����h��#.k��JY�����������������?|ĢT�q�Y�Y��{�Y�̬�T�.����*�g'#�Ã�`)ʳ�9�P&hw�%�����}�L6�w��]�ID����Ҡ���ZVғ�*�/��r�ݞ�s��T��E��#��;L�4p����50k�إ������!C�dQ^�a�?� ��S��f��6xX��$�sz���ɭ��)9H���>&�fTK��h޼$K����;27�m?���s�Jִ�d3�`��E�W@&�^�A�8;b��$�I�������~��Fxµ�_��c�;��8*O�K������Я"�p��UH�=~�l�U���K5!�q�>S�v���jpN�I���,ڊ��]�՜l�n<�ϻ�Ӎj(=�9]�p)l)���\i"��Տ��-�H��w��`���ZgC�_:X��Cu��L��!^"4џ�/U�Ju3��˵�Zwq6�c׌��?���,n�3Q:!��t�)<?#鷥W{Z��+9@���M���<���_ް�?5��i~_�W̏�?����q���H��8�n�k��(+8�
�V!<�ŵv��3{�$�+���ր�v}���$�x��]�����1��J%��>�HL �լ�^�0�E:]����Vp�--X�����4=�,�?��֮�y��{��~;S�K�N��`��ER��wz�(Bcm�O��D�]��]�ZJ�8[�������4y �sq�M���|��Ō���o����(�b����L_�H��{Pn�~�W|Q���.;�B���"�E<���4�=��w2e�*@�`�0�'{�!�3�t��ki/�'z�N���?�)���&|d��A���ܾ�L��8%Q0ti����5�5N3'r� �Lf�Q�`������L����R�_��$���y�E�����?Ʉ���\�J��O���"�Eíp�ȵ;b�|�U�	t�Շ�hw�!ֆ�׶�o㥗�B#� �p*ڌ��{����)�Q�{1Pu����R���9I��q=�g�3��4C�ckVh�2����2���C�i]�����?rn�|�3a޸����͕e�e�	lcdg���i9b��f:���I!SP����~�ӞB�vc�kYz+k+���z�>>>����@!���xe���4B;D�"6T�E�N�U2���U��C��<�{e�l֩J�h|v��g�L�~E겿���>>$�T�)��y��u�l[�<��f����^�"�~���]��:N8�3��r�_�^E0�v����d����ѣyHVh���e�8I�b|tkݨY��j���gϪ��*R��0�"]t�;G�E�#�>U<��|c���;77��{�L���(��7�,�]�Jf�?7�;�M	��w�;BGr�3m��1v�.ܽyL��9k>ܠ�(����O1����f����]�d�C�xg��� ��扠ѕҪV7�����Z��'�����5� �i�~��/�������v�	�+7�T~��&G(z�YJ���"���y�嘀�Sl-x�c��T��l����&>ׇ`�t���n`���eZȎ~������ D�ү s5���L9y��8���5�̔E��߃��+9�Zo$2Ђ�%��u�$���
�3�ӟ�����ۡ��d��VRD-)8Ṵ[F�᢭��ߏ�
�k������v�,��L1����:�z2���5Va�f�8lF�J1	����d�[��MSq
�y�z6�x؆��*�{�_6�}���Ղܡd<�u	[.@�;���c��x���ƍ�dY�|�������)���ћ�Z���-)��,7�#*j��j�d��8ݢ��g9MD�[�mK�VO�� 3�ls�~hx�o���I��m٩Vț	<x���q-��2p�$��!��W���B2�cO��������?���j��&�}�a�:���f"nkg���*�'3�/�E�t���I���p���̀�����~vv*�Y;����|l������	!ږ$k5�;@��(,[��14����J������:�(�M�)G�#�АV�B���8���	oE���y�\����g�Sq"j|JG�	�@3RYo�:�g	fEUeO�)OW�ʃkʱ�DS��Њ�����Ӑ�GG �%WER>���^/�pK��h�LWfY�e�%���?�b����-}���A�a�����zAe�h����! 6��ݍ`s�s��Ƕ�̦�����n�Y��p^<�B��'6�:7yt�)α�GGq��}ٶf��z���fg�*��!%����X��/:̾�R���̢��f�t0��r�V�����&�I�:����z�dN�0.>&_g���O{)��c�Ip�l�ަ�B�1T��R9~���8:�'T��wf�,o��F�M�߫��'��A�֩�tl,���1��{MGnn, y^^�`����#}�׏�`��y����l�.W�khJF48l�����\\�?.�b9o����A�;�����	8n�^�����j��)�4/��R�^��Xji���U�	H�y��>����,P(S�����><��{e��}���wv��N�6���f�5�ݮ���O!�}B�)s o�R�o���n�o��i�]��JM�
����Y����U���'�`۱��gqO�u�m%��>���5�Z�� EC`x�v���ό2䴱����:��{�h�d�ٰ,?��)`��r	����A�G��em���#�\<N��#�<?Cl=~=���4� �uDy�s�}|&����1�l�W���Z���'��/槣��[�@k���5eqV��u�b���O��բh�w�����&�:����j��+đIغ"d<M�/�c�!��P���:l2DN:��,�j�L���v��|o9)��T5C��������i�y��4Ij����v����x% �Y���sf�ݵd�Ð��Ѯ����`��Sl���{N׍���PR~'�F���C����cC�W!Hh-Q�~����x����`��鬾n,��ťF��P��<ֆ,B,��E���ڗ/��8�k��{��1W@��F�X�Z{��������4��l����[�Z9��X�~M�b^�}-��<��'�;�7�:��O�<��k}��B8��m:%e�����\��Qj���o��� 5łw4��f����4�P�}��|���]��GT��{1Le%��X��X<UNx�5���!A����/����(J��y����|�"�5�2鸆�n]���$/�s54�o�Z{��ۺ�.���G�o�Y�c�X[-�\��py��ZX��c �0�mR���o�`ܦ�ϻA5I��u��9lOj��O��v$���/ݑ0�g��1���!v.��������k�h4��p������L�(�L�]Q��CE��}M��k(�=�cwX�n��:���}W\�_I�,���R����Mm��I�v�&��@8�Ҟ:�`�&27k�>H:6�XB̈́>Q�ZE�lգ-W"��|��Պ�x��&�Q������G����vޙO�鈙��ښ�%p�%�I�p�~�}��<ex�����-���ک����	;S'���s�C2��S���@�����]�։:Y���^�;�A�<��s@oݝ�����@2�g�4���\����]��]u�kL��l�v^�A"8{P��1��R�⣰�|w�_���/ޜ;e�{�f�1E�v1{U�Yp���Ô����ddLR��{[�t�3�\�Y���)�*%�����O^ݠ���X*�F6���	R���5±2�e )�LJnM��3{�+�6O"_�xj���zs��{��Q��t�7׌���^��oq:�ͼq��W�E�~���O\ތ�ǂ�����-����6���d�PV�%� z�z3�1�b�����	�kk+��~�-w^��2a�?��wE���v�"�����(G�4c�I=i2~���d4���1K�l��Xk�m˱q���ON�xh�2O0�_C�?U���bw�k\e٠�����o����'�
r]R��dx���bA�
VO��G2����N	���� ��ss3�=r�V$Q?���w���/��W�c&!���;�eFjFB_b��P\�K4�z~P��w�^����;�	,k��M�0�m�B�0���-�e����I��4"�b����xu��֮b�~T;B�o�n��F������3^��]��ݛ'�ڿ4�ԓF�≙n�oYF�lH_��r�nrp��՟N7S�Y�!..e�Y��_��Ζ��[w;>1���%�%@!I��ve�B�9P���}ߠ���Kn�L�3�=��FԸ����=o|W����[�Ҧ2���g�_�t6�@� "B�K�����y�����{��{��M��m߈�ea`7њ$TOL ��5|����}���B�:�Z�.y�a�t�>"�ʕ��
��>>Rͥ��XS�߬r0=��И�T������[)V�j_��o$z�Q���q�����oH� '<fF���d�w4�V�CŐx�qJ_;|oV?��y�\yo�λ����@���L¿��+$��tZX�����d�CZ�u�3h���*W;Q���T<@�4�o�z�M��VU�`ef�q��
��'v�X����.r��z�A}�.W*\�c��Ј��۶�(:�Y�v����h��;�_��ɆN8)0���d/
�thyt<�O^ؔ]Ԡ�so��m(htU�J�*j�T�%��K�YQ�T��E+n�/�V�Xq�]}�f�)���� H���5~�xh�4	�ǧ�h0�ģ�8�P���Jf�T
�J�Α�Gk>gpdC�����	ŕ9����G�u̾�<-OHBB�g�v�V �pӲ����5�'�歕�E����i���-,�v�*��qm�Vc)��YF��u*�Pjݷ��&�V��(�()�%���(x���iF���Wʷ�߶Q%���N�Q�۰)V�]�9j�O�%��R�Y�=~��2��)r����"����B�72l|���s^���\<�{HZ��&TZ8 ?�H����v���6��}�#w�i� &pO��,-�ߦB\��;A܊��k/l,y��'��:Y���[2��Tq�<�7�=�e1�0k�뛲vBd/bT/�ǮV}!��O�uԏN������yp�rձ�$�=�r> ��3��ȼ���Hjw��h%t�G�vt��KLo>N^�L�����8���{�a0�L�+#Kp�;b��a��sU��Φ���7tP�����Wm���Uj�� �?O¤)Mg�9,�4��F'�u��[\���0TS�/W�O���a[�0ػ(�z��|��\�Ŵ���5�(���`��r����ژ[!z�����bp,��zI�P�J1qLM���r��u�귣�Yw�Φ��1�yO��  �.x��g���A��q2�o�u��&������B���=̷������#�+�+�S�wK�t�{�e������b=ac�	323��/� �S)��нt���{��y�1I]!8.��^Tc�<E�)��|�ꊻaz�5.vP�A��cp��L����g;.�tܶw�?�mL��v�R�����:�����{�����$v����Q䢪�;-�v��Fz�%��|��Of��.�V%�V�/���0t��P��*^��h_+*'T�8ˏ�qu��.����x1_ΨW�8�߳HA|�x\��mĜ�Ɋ����fW�.GGk/�g��8�j��{I�~@"�d߱�C���.$ҹ��q{���bZN�;�/쉼x�8�r�Z��%����YS��V�����&��<v܏����Zt���ܷ[��	�DPk$n
��D��.�� z3��Y��%���J)h��֣�K�K�ŋhy�n^�������|�c����w�2՟K�g!�f��ЧD8�;��be�����I���x�����CO�2�|��^�Ѧti^��a.A6�2�:��US���^ɖ ��S�hG����龜��O�/�~����Pb1��I��8^���z³Iwß���-�l2S��.�$�$�)����6�����n��R2��'n�;�z[_y~/�<��Ėe�=��׻h��/���yf+a�O�\�U�+L�P��T�
ʻ�?FYHkwk�m��It�g[������t�!is��R����M�<��[}�3�Y�O<�;�����X��C��7��KK����c۶��fcӐ�L�Դ��~Y� �/%���Y�-�v�]q3������z��/���^��	A�4���;v��owq=q`�aht^�n�gygɀ�qٹ����'�&�����ީb�H؋K�ÚG-�
־�1${Yi�Oe���Y�^38&Ѣ���zVń���=�{�t���fS�iT�hO~�H�e���J�aQ<�*	u�}ы��O��4���	$*�3��]��M棌�'�tj}�3ro�ɊG�ݩ�I!}�b;�֌�,�?��S.�X���B^Hg �ubZ��QC�4V����
�,P��q�i��d0�nh�����}���GU<�MB�^i6��%B5/��9�Y�����^��.����}<[����q�A:&D�m5�cJ1޾�V�6B�I� �P��;fc#ҥUOL��/����2Ƣ��ǋ��:��p}��5��SS�#������q�ˑ y���Vȿ���G���nY]L���#%~F��+�C�0�n���'�j�S$��Q��C��*6�^�}�0D�3��۫WP�6�ar/���}�f�$���%����	~L@�ג�B�Ĉ���;�;�[����w��E�"�D�ѣw!"���{�=z'��[��F/c�}��������-���Y{���>�L�z�	ŭ{6��.?��R͐f3j�(�4�\�����XtP
2������q+30p�"R���,=��R����LѮ�ZY�T��ʿV.{��8Y���_������d�n=��[�f\��ֿ�l� ��צ���Ƒ�9�ƽ2�h�NW���ȹ���n��JW�,>)<oǛ?�{m��feK<+cb�nB�_�38���m1,�Y~��Gn�a�{KⰐRF�'曞������3v�'���&�JmseS?����r��ɏU��Ķp}/&d�[JԸ#[�=5�dzWfF�=>��42(���ڨUd��9�����ӻD�M�K��ۂ$C�he�N�g�L�`U�=�ȏ���끠�ga��~�EY�E�݊���`���ۯ��t[�����d\ĉtoe��K��/=�B^n�7��� O4�O�Nh`{����B������%Ո�3��J�Q��La��Jg��o�L���|M/�}�\�G5����NNƒ�� ���t�*�|U�μ�1;&�uM���Vs�l�g����N5����1`���B�z4 <8^��\$o,.�z���wk&��z�'�_�[���P�z�R{�<����u���[n��U��ˏGl�v����I}�i�y�t^g�lp�Jz,��Ĩ�����Ϟ5��=�nsv��|���x�CJ7�Z�%$�"�ȁU5��4T�g����@��[�H��p�PH( ]�!0�E#�l���eY9�b����m���WX�ԩ� n�������7�z]�#4v����~��4Tuass�ig|VE˟Dl�_���n�����]�r\��n�����t<���BC;7pGS�4���|݈�S�N�HĂ#�#68�)�ڐWSE�E���b�J��K������c ��
��������6��d��H�9�B�Ĩ-�q��.���tI��kf"2l�te�G�A���"��i�Uj����29�V0�+C���!��&���&R�gMLLp!|H��D�68<.��z�iCd����Q��Y�h?�/o�n�9��{��$��(L ���3b�\֢7\Hf���ڦvE��e8��G<�� y�ҋ�ǻ��SX�eH�d-IA��yeͬ��2,����#WS">C�v�Uho;�}H�bUC�T	�e�h�拴��Ԛ�.փJ�U�4�o�+u�=�pk��@�^�%n�)c�5�pl�n�"(�n@�%���sj�(,�tu\)���
��[i�����������3��y�j�W�b
�P��op�8�m�"�r���v0�*����T��?�p��\���|�}��P=O���c�����D���^1+f�����}�?�v���4������ٵ��}ruРi�BE�cD���rSx�db�k%zsY[i���^��6õ��4KϠ���V��sł�ym4��D��v���H�T,��E�(�V�4�Z��ش46���s�~3F�,k*��^s< ��'�&!!��keOeUdx���eW��\�rQ�]I�?=y�?��b��o	
n/��t�fT���7^{��T�T�jN�Q'�4@��q�����`rH�1�_f�����Lv*3�- 0�឵)�q�@��֓\�1��q��ZV�M�����eVsᔑÔ��՚��X�v�DĜ�y��gdv�n?�*�I��d|�vv�~9�lXx�s@L���ͤ'9$�M�5��Hз�])U��uA�6#���Mo$q��,�;��sʇ�.�ί�ƀ��O_7��`��6����@�h�6��g���[��T#��>��x�]�vx#
���߼@w�K�Wgu��7��K�vu(*�f�_�7�o��?`�b�%m��%�C�W_��-^�gs���胏t�-u���o��rB��T��sƋ�qUʋ�}����Y�����e�O�@��H,3�՘o9�����Q����+jM���=��v¸U�V�N#�O1E�qw�w����}�	��-=<���r��n+6I���^�s���W��I���&��H�lOd�?���Y�9R)*`�艸�b�*��P�=�i��l�LN���B��I�)�YM��[�]�I�-����ڦq�Ux�e�z�|�'+%p��P������4����\��oД��lLc�Ot1(��CI�X,`�x]�.�ۺ�?��+	��4�?����TE���s勵�0d�D�[r�`�����o=tv!�Jm�Z�~�~gE*婏5��j>�|
�]yj;ln�_`8Ϙ��;����n�F"�W�t��(�-i�1��l�jBU?Ł��l��3t�}_���h�*�����R�$��ɐ�-�z��+4����|H?���mD��n-���Ǣ�%����31*���6�vb;�kb�Lۈ�-�����e�������\_Z�촗�c[��I	�����&K��@���C�3�\_�i��dҜ����:[m��uI���50�6v�( y.�h�rٵ��A����ӥG w�	��I��V�_u��|��  ���h��(ea�#�C�ɱ��)C��F�Tz��Һ����ֽ@�h����
�'~�/e*{k?ҡ2�B���S/[@=��~܏~��2)�^������4c��,Z���#M&�d�ճ��A��HNw(��c��J"�}��r�����A�FC[[�j1�`�F-g;�8����?Ɂ=�_��nZ�����҅$�F����r��d(?�Y��ډn�֩gA��ԇ�䷌�;=�J��S�'���:v���0-JSo����~���������������I9�2�cC�u��G:q�}n�Is�nO�l����5�J#�Ȅ��F|8gɇs>\�*�~>��&p]klo�"����I�Gƺ]�q=�ʃ�����vC�D���s��Ƶ� $ �S�� ����B�B'�bj32P��F)�eD�ì�g-�wv���>F7�U��G �Y-zn6�<����0��[��#{�>���Z/V�A���o�B�:�Z��鿹��R՘���:�)�m�P����5�����O��5�����^��I���a�,��VJ8ո��
�b��J,(�y�������J�V�����ż��6�)F��H߄��4x��J�$��?��o�y�(=m���f`�^w�>:���b�BwD|~ ��A]P_���, y����V9SkGA/������0�Ӽ���È�Qw�+>P澠��� �8]�U��x���T�L�����i�oX�N-����������`�.��0���k[���'��O���.=�~5��������=�md���Q�U-��y�_�ʵ�h
BJ�6�=n)D�G�Yq7		�ns�}y$�I994�x��)e" ݝ����q�����ɱ�ѭA�#���gjb�uE�M���ۺ.�dBP�#�[��S�:����h�fO9;�$�w�]&No�ѹs�:�9�?�j3�I���[Ѽ�����C������&w|���X��4�w�ݳ�i{%WIwoN����[��}n	�?
�Xl��iOt�4�>�{_���f��؜��������24��a�5���|��e2����pL���!�)9ws~�M$QJ�VO<�@���q#�d�'=��X��bΚN��Y5H�����I1F~Ό�x�K��Y��-sX�8�KD[\p�G�X?�i��NH�/��uH�ʿp5*���{k����ZZ�l2"�Q��s��$��|�g&~x^�W��5���SXID��]6��7��� ��㒹�D	>�P_�|Z�0�|��^���E�8u��X�]@k@v\�l�ȗ�:����U u�2�Xw_9ġk6N
S��`��Ñ7�wwv�l�S�k�'��3³�s�k����+g{p���qk�N�ұ|���B����U���f&��蝧�~Qق��p�&�&h�p�
ם"]�����0��!f��'��d���5����Qː!�՞���9c��'OwQ<:�:o���z����ٹ�(9� h���K�ګ/~k��%c_H��+�?�\L$��%�Ӹ�`֍-mb�"#.3��f��;��ll-�Pb���~!�>�3���È3o&\�㗸V�X�-�o���eLvr��.F � ��IO������B2�7ݡ���";��|���z��
l7��򚵂6p���}���V��?)��D< b�\��:}4ҨdN?��	�*���L�K~��h�o��	61.v�4 ��� X"Q[��n}��K�:�?��^��zR�\��D����6O^B�AM5U�)�,P��)�T�Q�劜�NJ�n�Ϡ��`i��������4/���啨��]z��a��� D
�;��IQ�P�a��%h\��Iۈ�o��� �4�n=���y9x��kva�u�M�� �Q�އw����+�r��X����e�l�:�`���~�a��AV���	H6�he.@���>stw�^���o#FE��K+a����;�&�_HW�[�ܪ*�����2"�W�P&	LT2/�/kg�N����L������H�������D��T4�v,)��B��Ue<�+=�����޹��%��^HMd`d��S�0�?�ʂ6��h��y��T��ʝtk������uQ�c�v`$�-ٟ�O`�fP	)���(���Y�|)������!"�dp�F5>���]� �m�K��߄'ʰ�v�����a5P����`O5����/ҷs�S5��M�r;d�+6H�(���v�0Qx�]3v*]�Ov��SUX���+�En���c�%B���}Vh�rb��ڭ<�' �T���⁛�ҵw�AF�M=g߳7�.��y���D\�}*A�##������/��O�V����-��z�E�E)9��m1�+�1��`�v�F7������+�Mcc.�,N�rDY��
:��5Ʀ���8�x�,�7�̒�9�|���,�OǍ�EEE뼳�+�m9( ���-<��Tm�`6�~�:sN	�Q��ڵe���r�Ly��pm�c)�E>�lr?'�=�o4_��H��a�ʜ��l#�)�*d �7ӵ�Y)e�Z�v_p�i:�rH"�.kH��~���]1WX�|g��NI�	�̢w��S�Wr���oc'e)�x�[�*;B�6�,�y���DH��mIm���#�{������T�k���T�>'��Y�4�{��15PۤE��ҷ�~_�������Q�+Sg��fS�L!U-OC����1�D2(曢�L��7�����iL��u?<��i��6�R���:�hJ�Jګ�0^���AH�6�
�C�`JCkHx^t�Z��OM�b���Ѭm�C}�/ck5F[���3�t+�<��}
[�5��Wn���_��ZO0��H$��W�l]爹p������b�񢹟msmV�n,ck}�,c��ײ�<���Q"�O���ta�"�c|�/��(�D���Ϟ"z��x9�[�o�!�iu�wXX-��Ӑ�����e�k�oCεr���{������dܳ�?���B��P�sT'�:i[zQ0�տs�\��*e��9J�A֦N���GY9�S/R�>h���w��qx�j�M�dC�
�n�������qe�$|S�Y�5���_�So��	6}��{5��䰖�br�ӝZ��?� �_FD�3g׾�]4瘜�Cש,mE]DR&��8%-��j�܊�m�����sp��CW,
5�J�Z�)'�ͭ~tP�/�k��;Bޝ�����-�)+�z��T�����-Z5����#/M��K�JWf`������g�z��K���_췮K~���4�i�9ih�������# ������8���ZK��#}���}��CB�>O�v!(|�(e
�@Шe}[��)�y}ޤϠ�"�?�d�\��Ǭ�)�'�p[_z�@�X����;5|+��ʜU�W��y�M���'�e0��{�>�j�(�?v���&����֪E�R�R}���T@�t��R�B����e2.%J��A�2��,�XJ��,�Z�.�o4MR2�������R�!���G��]��M�Wj=�Jl���6�]$�7}�'H�4bԖXR�[a�X{Nh:	L���AW�4G�4x{xE/fS���Z�ڣ��ipØwPYڮ�*~���l�M��c$~�D�XO�;ZKÄ�9&���z�J��q�	_��.܉h���0���а�j��-"A�!vqܹ�q�P}��|�+�<�s#�_M�}
>�9nɉ�2�^4�Q���,g�G�����H�ո����.x~8�o?�k��4�JE�
�R�2>'���u������0?��$| ��R�_2a�BU0������.vZ/�u}Єe8@�O���O;k��G��?=�}�w��	�h3ř�w>�	h1�KC���4�7��-��q|t1�!���w��[u�����ཟ�%������2f��(�{��b'X��N�˵�-�x�b+c̸��H��,�\t�6P/>.��W�kf�>�3���|\s$��g�g:(�0v$I���@Ov��5I%TfՆ�Oz���^���xws@�'�|���e�W�B���P���X�� ��$���]s��?SUIJ�.1��%���X�,Z�\���x �y(��F�`�WVz�|W�Ÿy�7+�/9�n��j)i>��t�݄h�w�TZ~Ͻ��Ѧ�w���?�Ȍ��ޚ�i�&�-Ɯ}�'�ݠ}Y~+��z%k����_��B+�I�R�+	|ph	�9�䋌C�l�@�N^�\>�X�p8�o�z��D@�ƝT��T�������0�`!u4rβekC�6�P��w�	�L���ս͸���Ƞ%��y-�OB� ��`�ѡ�-��n��2��v�V�克��xc��ϔ��=S�?\��B���61��V�zvQ�q¹x��oL����tG�I��-^r�����F��H�e�G+N��Vw!I�YzϷ��76���S���� �(DQ<_�圁��Ӌ�bf�P[�D:Y� Qo;;���FcR>�һ�
�njA��f�fK3S���84t�>s+���$�<�������w*�n8/�~��b� _���K`�*T��=+D��$�tm�HC���x�\�;��F���~ya�B�,����-v��Y/�r��z	��{�9��׈E���q�Df�=���B�Ɛ ;Na��B0����kA;	\��?Xm�]>�� �2<�]��ą���c�LI���H��ľ^�����r!a��W�.��$k�8��AiY����x��d�.�TDeV�!�����율�o��S!;�� �_�|ꆚeJ
�+�ѱZ9l�_x�b�����S}'��<�����B�H|��u�G9�����;��X�?]�*���jy�'Z#��s��F|MzS���y,�.�j�Ԩ�r��C>'��Yb��0���ۏ�闏�/�����~�
Z�J���+|���������	!f�J��q��=[�.��#���!�����A�|�> �8��C��f2�gZU��$W���-�7U�.[S��з�k�N��t�����" lkT=����cM����~� ���AHh_���F��,��ZzN����c���ٚ�:���_�ݖC���xX/QG���������n��EE�����F�ꑿ�:�'��I��+:��.�|��=�����/��Z �h|���ى,���|�Z��7��7Ue�}��4�<��N��}�z��_���E���9d8� ݍХM2x���#&W,������Ai�?>�Q�ώ�=��&6���
�V�._��_b4v���d��k��5��S�"�޹{�d߀ف��d�
`��)Fj�i~zr4Ƹ
�1�ݷSƙ(������O�Bd�s��nB�c��"�X�O�lTE{���+i�*IV�\�����_�7�ͧ!�� ϸh�/n�X���͗G��u���Z:!2{��Ih�@���A��������D�o�vç��� �6.c��?q�'�Xtp>����Zε�(��M�X��J��V�QZ����r��&%X�)ɕĸ3f��~�/����������d�N��wך �y�+;*vb�r�2�M	�|v��Q�|����R�^p?Y-�P�6F��JY���!~\Ր6�>HÕ`��l���4uJ���Fv�'�r'5���nz�a�O�ō��R[��������W�L�3�ZV#8R�$�ָh�j�T���:�q���{Թ�y�r���K���_3���礦vLh��y��Vt��.SJ�� �4��"�DЅ��a?���2LJVS��W'V�p|�z~oA/4A�S$J)��h��.0V�Yh䊟�Wq�dO�F;��8W:�a��=/�`���\s秢,�fW�v�	�e�{��@19�ZE�Jc���Q�i<xV���띶wvQl����/�^����\Hy�@^��V�Q���j߼W��㧳�M���V�oSh��T�/#\ͼ˘Z�E����c\}�׈h�����ݻ��UN��0��Y��� ��Xl疷q�X��o��;�	��s� +RtǠő;�D�z�(�hs��b$&i���XY$����T��}��ئ6��O�Μg0M�5�}$��N.���0��ߘ!�j�)G�������������j�ڶ�LeMW�E�ܾ��鍾TP��f+��;I����E�>�Є���-�E�a�������W<��gs:t�-�%r@[4g����' ��ʙQ�qk�'k��Wj��������b�m"Z�j�b������f�p_���{.�	]5�v$ǣZuv u�)�-�*~�����ܚ韜v�'W�M�w�4_���d#Vl ���B-d�-��6A�}���n�������ߢ�)㼖�Q�k��}�^WEQ���h��c� '���Á�6�j�����~Z�+rN�Y�W�Qywv��-��w�)� �֗^7��3j�C����52 �^!5�
qG�	����������{M�3�²�7S�K�$E,U�Γ��{�0EHn������N,�W���c>�~�my�Uل��7UvZT1��у����jRy�9� � ����0��ΦCZ+X��B�\.�+/�k�E\�$/;��Sq�_A��O�h����f�tX�bmYo,�Cx�qgj��+f�</��p�ĘZȧ3����h#���Yw���gZ<�q�����)���Os*�g�)������֜���5�ף�P☰R-'�h��7�d���s#�؊z���)�u��1`���k7#w����g}��K�f�Q�'M�3c�b+MՅ�H���.�R��o��3�����0��V~�7aK0#�P!��Jd6�$cPj�ġ�P"ɩz����?���{�+�E0�z���a{�-�!�pI��Q<�%�?�m��U��+("�+�����|6��"�����:�����U�9\�6��ߦ��b=l�t�a�ә����8E��\1��#�$0vp>m/��~[{m�I�d���g,ݝ�}���p���ݭ��U~����vۯ��H)��;ۦ��[��F�+�k���:v��N��2-Rƛ�����+�j8�ό����Zdה�G���>��0�Z�'�ɝup��V��{�$�B�?�ep~rx�,cb1jюr��W!#{��=�jd��xM�,{B?~��D�tFW���g���co~���m�vmp_���Ђ�u|�o{�^	_���4 ��m���l'�2..�Z�U���W<{������y�Y�-c�oa�Y���q1�j]z�#��.��ƙνJ(�͟,!Ͼ�[��>�:SDW�h&���<�^���X����/����r�̡0>�������Dم�ڃ�=[ �<k�?$wS߾�Ly<�\�t_�>�#�}����gC�4���ю�,B-l���� ���MG���)�D��9��?�-S/X<��n��& �S|ۺ��6�����
433����N��<���vq*&eH�B������G)��!I�]Q�er�ڨ&J^�M���3�7�ewL�ٚ��t�1��w&1��-�$��{
�5ބ�ym��f��	���S.s� �yY>�xOu-��=+쇳��]�Ęï�tE=X��/i�#���U]�gJ���g��{�~�k]X{�Q��sYa�iJ��^�&�B:蚦g��k��!�F[X���K��q�<�aܪ�A�^f�g�5���G�������i�6��"U%`��'��u��蹵�+I�I�s
�����@�y�F5��-�T�t������k�rO@?���qyM�U���e���F��P8�S,�h�52��MzAc�5]����(˻@����BӅ�dh���D��6���y#r����)������(�*�>�vs�!bV��w����Bu�p����`Z��"�kf�9dx�D�Q$y$u*7��f΋����E�k+(�x�8�t�h�*��V��h�?Y���c�;����$yeV��B��j�i���Y�^�;�h�j�o�n�V�liޮ1q})��
ʇ�zm&�]����Ō{�y��+q��N�-�=Fz�)/�q����k���ȍ��>�q-#UK$}����|�fNkk?�֜匼=�O<�vU��۾RbwP�Wl<�HE�PG��ߏ�S~Q�#cףtLf�1���F-�\�7��K
�sU*�F�{j=Ł�ؔ��.1������G��$?&����'�b�o'�Z���z��6�����[Ѩ��~�n�@4�ܱf&��Ѧ`��?�0��wNEoyq�әU���v�[<\O!��q�7�U�(���p��_�#9t\�#�VR��r0��⨻����З�)������s���S��������uQo�������Ep�6�wm�2�v1�R� Tf<�q�k����9l񳫆�RJx6E8��s�ra���b�\H9L�y�cQT�u~��N�݉������*�9p�
l�I!�K�-S��q�hق��et�4l�Ҏ�����>��4�Mcщ�~�����R�G�ti��ݼ����u�V���_ż���A3�oe���Y%�5�5���i;�\�j�7E�G�";�����Rߝ�����v���\��֓?np��;��dv��k��B/߂�&_Yu��y.Gql;���߶�Qʳ�/�g�OEhS\���F�N��\M�1�e~;���2�g�k��#JJ_G-Cjʱ�4�/��~.�;J"�g1�hz��$c��J}L�:�o�a�b��NTYy�qL5*_#��� �c���Q9Yq'y�ǢhV�,�ϰ��S�� ��g�oy�(#3��w�9���v���E�s����=ǉ_h��N4E��D������yF>�����.��$Ei�Ntv��E �K���{4~� 0�T2�k��x�C��[�ĩM�0N�ߡn�3���3�;��e ���� >å�#�_}��dr�ᮖ��He�FEDR�)]�����޺�)��-�	B�+[��hֲ�̿ �Z��T,�����e�b�.�0�-)ꥃ�fk�ʜ6t8�9���*33��������`�H/YmW�Q�y_���n!�KϚ�~SJێPR}!k�O��MU��s�+r4��待��5���:��i���͡���t��^��W���\|y�u<�'4-��Xu��gF�ݲ�?����?XZ�C�`	�kC@.�w�4��s�%%��������8J���߬�žMp��hԶ/���ۆPh�;��V�I	pb��Y"l��k����|ƨ�<�pe���5��cDX~^�����!'��3����l��:@"���rؑ�|
�D˟jg��5��oXI�ڏ�38=}�W���%6�%�n��d޴7΅���ϞL�j��������,�mV��,N�lj�a�g�g�b@���3�M��Lj�K��Tm�>�\PO�0Y<I��[g�b5�pC��l����W��γ�Y�EQ�����o���/���9�2������������	
�Ʀ�
d����M�������:����5����$��� �/�>R�T�ʬ΃s������`K՞����a�0����}_�N�i��#��q��J��j&���`!����?`nF��l��
��N�4n)A*�@�,#X$7r����y-��;ڼm��Ͽ�Qn�|�4C�D��q��>C�R������Y1%���{=��NQ��=�&�G��Hs/e�oCD�"���t��dY�@�����o���q�L��!ô�&)�d��$��Z��O>J;���j�%?�V�2���WK�G}��39U�$b���7��J�K;��3�*J���0���d���0����ѧ���ҔUɣ�|3��Qӧk�=�J1�a����b��kM�>Nۣt�35@�*��a%4���R�?�j��o�b��қL#ۓ��"��\��Xr����
���=n>O��?Ua�[~z��������A���?&�����"v�5.Q���iGgaL��9B�֣��������������ڙ� 9��ICߢǜ�A��u�;�{9�[A�����%��_S��l�Q`�~��<��~@ŐP^������ރ�|�>�-���0]j�V":J�>�1�D=�����zcWi��J*ɢ�?ev8��x�Ȟ� �܋��~7��CţTv]w��ǼBufrR�3݊$�:�{ު���%\V�Hx��>�O��`�W� �Fy��3�t�+v�r���^1�V�X�=�������K3��ip����9BNhJWo��<�
��̇)����;�\��~�I��ʇ����)�,�S�F<oob���T?{~�B.#�r���U�d�͎	G��y.궸F��IR��C���e}�nt�T�y�b^�̪�I���x�H!�u����+�U�t��h>I��5Z������U3}kQ�"�r�*@VL������4x�-��v�ٳkK�*Z��F'5��g�~ɟ�UZ}�B�%��lKx��^ϒ'T�k����%nDK-��:��X�4NK�#5{%2���J����D��-3/�{N
�g茒�s(��Z^qMv�;����Wq�7f���r�V�27��ˤ�_�뙮����<��Ԫ���<BR�H>�w��VP�����L���{�.���e���f�'������a;-��+�}���|s�
�AVwg,�4�
���b���bn�*�m�)�~AՅ�2)�\��1�61�޺���z0CE)'����X<��>���`/��i=.ģ��tSn����8w�t���Dx�'���%��*�շ�n�i����2��8�Ü���V��D�
��n]1��V"6��i�om�!/�[��.�JI�)yn��v�2��iQX�?��mV��L��G��J���p3iS�c����xw2H姄D6��Y��]#��KVB�Ҡ^LSxrày�uD��.�L�������ݫ�ے��MLx�!�k%��%Էy�)�ft��bFxChVƪHG�K��dr����8�Q�a�K�J+��2 ��_sq���;d��gޙ���r<W����eO���pEI��>�b�آp�ĉ�mW���(K^���Yݴbҵ+1~pL�c^�{ʫZ>c�'��?n������v�=��4�DHJ�֐�a��Ji+��nZK�_�g��������BAm��_����~7�F���)m�>M��+0GNӨ$�����VN�.4/������oWV������kCj=#����E�.�!T-N�{�Z��E�Z':��������.���ǅ���%gh�%H����,*��D��8�}�����K���� ��S|�o@�B�ʔ�c���i&0e
й;�1~��;.�&�*��^��}s$�;	�P3wr)+�0]�g��IZ4�s�Tkxz���ϭN��������c�[����p�8w߷�
Y���]h���4����I�J���hգNك��i�I�������G"�6��2�ߵ��=��7��e�����W�B��0�9��7;�x!J���QH3a�K�	�NR���G�P������o/��D��$�)��=�L/,Z1ʕ��(Kۈ��(C�7����HD�=«P��85���9���VU)�j̮��&1� ��j����FCo[~
n0>s��������v�dq�ܻu�Q�N�AP��7��
������ybب!��[�8�&*h�d7�5�ػ5�!�gL��z)�ϸfx�#�]��5lԪ>���W�[y��M^�-/�������\\��y������-V�v����>D����,'^Y�omܦ��UzVa�~$R�Plf�DA�$p��#��k@��}3!|���#�>n@���S�Z$'ٷV��(z���TJ��@����]�	r�w�gM�*#�`2���~���B)�Ce��5V��nZҢouY/��t
�gn��>���Q����������G�Pأ)���vz:\�M-�Vs�u�;����N�j��a�ۈڅ����A�V_�M����V�cة�hZ �o9��݂�H��RXg��$(�41���rz�Q��C� ��~��G�KK7�2_��9��sLN��7)�y�H��c��7��wC������yao�خ���$k��y(Ę�Zߏ�M��g ³�#7�=c���o	��5#�͎��a���5�6L7�hk�k��WX~�����Y�3qgm2>�0�ؙ���!y����u�83֌68��o��{���6,D�L��r$��|�< U�|���
Q�!�>�7�G:����į�>;��,y֤ăX��r���j��4��ΰ�����TV0�~#��^�+���k=]�hoԋG���f@&���J���eԔ�h�=����~5��O.��ᐼe��1^��y#m�H�{���N��Ѐ	�P�����	�U���B����\�3L��Z)>,���眏W��%�Q^+��X��������k�V���̄����$NX�q-��_�g�S�&-=*1è����%Q�ä��z{x�x1r��Q�w�l�����芡ꮌZ�y04ؗ���;��^9{�k������[����&�H`[T"9]n���\�K�o�,Q;�t��M�iY��¨�n/&��������"E�z�����;c몿 ��.H.N0��C;lM6;���Eo"�e�����|ޓ�l����o9��
�����, ;R�H�vl�[����2��;�9��g�Տ�������3�X��CCN��Q��)����5W�f�>��ǩ�	�Fi�$YG_��C��s��BQ�,�v>�w��)g�_s*U ���aΝ��:�/�S/��^^�NY�;4���g�,;���
�m.NR�K[O#�� ���>KO�Y�];�Ӟ0�l&ȹ�g
���Y:P��<��^E<�H9i5���4����������~�E���[wQ2��7љg���n�υ��͸L`M��7�-��?���&8+���o/�0�d3r��3��̓K�_���'�y�ˠ���x��v���rl��s��O����ވb%�!�B���w�CPB˲��/U�q���܈.�dTS��RWbՠ��._�u��9w�͵d=�J�i>��p=��4��4�<Oȹ5�G���$`�<�$zjl�gQ�����q{9���ʉ��M�3���!VG�t%�Jԋ�K�%�7"�o�ká�'��֯�*Q�~`��[���[�p�H
bU�_?���\+Iu�Y!����4}굶�<� r����z�8吤爋U ��3���ڍ9O�#�6�>F���A� �=1�`�^�cxV�0�ү�մ�QD��ȑ��P� ɢ��.��o��vL��0ߓC7�J?5�BC:��x��>$��c�|��>��Cβ���?c�U5!p�N���B��ܜ�[$�W�W��?��ۢy��I��;r��̆8��k�7�uD������}1Z���"��9�1�O��sMa�� ��zz�&\4=%�A�H��1O����������^�z��߄[�k�2ȿT�C$G�N����֋�J1W%�qՇ���*�FvP�Q#'�r��
~Y~,R�#��;�C֍Σ�sR���H%����=��`)h�Qf�,N?�Z��_'{�/2�냝��̂o��f�O����q��Ak��"}���/6���X���R�}�"�of�Gz�����S6�I@#�\��K˽~�I헕6b�=�/G��JpTX��וk_WnI<�,�+�o��$�sYQK=����,�F%���u�x\��s���� ;kB����ny�em���^\ y�!�Z���U+c��z=��P����~��Kh$����֒Әf��%L��?Ը8�i�6�o���w#�	c|8�Xw)�'��7yE���H���&��w�%)��,�N���2��!\w��P�]Kv�����%���͍%NK��l#vQV�Q-�N��0����p�\�T~���z뇦��{X�iF���[�n�Na�]#JH��tw��1P����F7_�����/�p�s�s���3�"�� N�{.���nP��G D|��I��4MX��k��~�F�vo�<ϧ$y_���Ud�ԦX��V�М���4���5�>eE��Q�u=�H�f�Ņy��k@��f���I��T)Ѱ��{��X���ё�M|u�Y���M��	ay�è�/�˙#���=[���X�.�h�K���j�U"V_��.?��;jE|�X�,�0c�!�Ph̑��t�Z����#�B����<��Ӓ��>x!@�ae ��ý��%6�È����t�\��4'�7c��d�}���_����q�+A�jUU-�Vs��8G��T&���7�(j������h�|������χɹ��Zvx��ɺ�O�t��Z���� \tZ؂7�D��ᲁ/�-�����p��I겳�lJ�u{(�n}?�z��K��=��'�DbUٌ�XE
��&���p;I���P	�;$���>�R���޻��V��Ǹ��Ʀ.9
i+֌�����l&
��C���-a�u�xD�Ԣp��J9�u8�J�p���˴��W���ᷧ-Nˑ��ǣ[V=e������&`� �IkT9�yBC��*s'*j�ĝ�^�-,��*�P�I]qss�:�gu^��s���G����G���.�(ށʴ�����;�*tm�p�#o��w��P�N�ԋ�bG�)� S.e���MI;���CT�oqor���uj�15&�ɚ�]'��a𴆜&�`����`J���#4���v����������a�j���Id$W���(��"	/��½hg��>���������=zdS2��̨D��O��BBy�_|��FZ�&O�T-�x�E���=�����Df��L�&e6qStf}]��"�2�ʎ[��%�j�v\#�[�/.4�G	���TGG	{���V���FP���ӭ��1>+h�)d�e�۽���S��pt�=�`�k��&����*y��7��E��r�}����ӥX̦⅟����F���˦Di���&){ևlO�hO�QY��v��i�HP��ti}GA���	�HnM�T%� 1�9oE��0U��u%WjjZS���O���c��]M�ȳx�ߌ�����ᴌh�	c���#�v�}��/�?R��.�(I7��RQ�����2�5��*a�t�P�lL���ш�lQ��i~.�Y�c�N�l�j�U*k�ekwD����.�sc���O�:���" �[�g+�XU��沞}[���B+�י��F�p�����g���Q�;�D.��&��~i�1�����~�%����i�z�"�C(�]�[/�[>q�������	�my���)�G�<C+�:QݞYgI���y�}r� �z��3齥J���0�x��=2�u��x�wH5�8��F�><P2���w�����Q���a���!�?6�.i���b�5Ϊ�+��#�nM����`T�4�e-ί�����E^_����II8%C�E/�no�
Wj|�E#y{9{�J;�C����]��/��ݹ�21>@��tV�����8{W�/\�:÷e_��c��
? \yz��)"Q���ۣZ^I�1�7A�TO�=:��\�2��E�^���O����6�Z#',?�=4�L<�C��w?h�m�/���+���?3�f�Z�D����?/y��`;(Ҷ��w�\p��Ti �w9=M˶J��Ѽ
hȴ��U��S��L�)�'ҁ5MQ۸ah�^���Aoې��I���\dY����o�s� �W�5�!3��#�U�E�5���π��cEɜy��1_�'�m�ތ���P�����YU(`%��/�$vn�d�>���{�����[B���m��Up���������]�LϽ��/�Z�����:������B9g
�������aa9�l�U�a�+����v�)�ܲf�{�*�@����Kbާ��Y�S�4���V�EY�[�
��$^�'������36GP����n/q�7+����<J�R3�?Jҭ����v��/�}z�a�k��GV���1��|��n����Rv�^���D���a��7��lRҰ�6��z�z7�a&��q!��,��qd�N��k�2�j�//��d���*��$�������j���9���cY�z�5 �M0�f�cRE�����s�2~���t�Ƃ�X�`- Q���?��w�z�.;?��v~��v0�*6�!Z,/{&c���E,�&�c�*���F
wClT̿�²�x�n(*�,�a���F�(XC��l�nK~}�+P+�筨S�Kb^k����	h�#@�W���Ϗ��Qŵ���Y�r���SN6&�/I�S��J����h��/qT^���_��BH�����̋?�	�;k)����'zߧn��jN�x7��6�����3�]�M�v��V�X��Xݤj�l}nt�"�PN}�u4k��ELj��Cg�	�����j�#���/>(K�v��ɥOX�;<����u�j���N�cƦݪc+Y#��Y>5ya��>.隣;!���#�j̦E��H�/���v��&S
i/�����CG��<�K��L^� l�l䣞�lb&�͍狳^�~ֳ��/�̬�
\�Ȟs.:]O��G�Vn�(��ݤg��P���;��N���pj9�-ь2>�h���[׷���07=n8��@ƭ'�)Q�]D��������XOM�S�X>�q�L�M�:ڞ
��JS%����Ex����^���!���{.,���ф:ٟm��X�ퟍ�Vͺ$��-ϥ ��<s���mD�T���T r:d�_�U�Ԫ�T���+7C9d<>U
bCĞ����(���\�R��h*|z"g_��d����O���,��^O_�g�d�<1�bE�S7xL4q�U�;�׵_n�M�-^�m�lUH.L[�Oư�����O^�'P�'(���Q5��%��ίA���'ޕU���yb�s��3�Y��F~,�֓V�ew�P���n�ef��s#�>�m��m�~��tƫ��L�--6�K>nj߯��Q�܁�p�h�z{��O	B·�,q����#�?��73�+&s�n咓�]���i#F�܁dR6��t�\{��Hb>���viw���a��J�^�i��A���?-����;�/�Q(�0xs.���Z�ME��j�Ir�s ��d�Qv����~d"O�CYce/9�f(�GH���d�S�C���V�>>8^��[��n�'�b�ύl�Nz��)�n��=4�K�h�	l�~k�
�-��&�/j`�B1V��`�hn�IH��Ȯ�TvPw �
y�T�M������'Y���jw������ɷ��O�<�����]�-��r�v�9����rJB4'a�`M�����p����k�Y/�M��S�|�[=<��Fp�8�ɪ���	5�A��f��

ݢ�N�[�S�,�/V��~&�a��H$Q4�P)�7�H��4[wǬƤR�Rߵ�w�ິ�s�����xi};��VN^���K��.�eJ����~�`hl�����>�烵6��ù{����i�~�4&eX��Nl�ǂ����m��'���Z��磢a]T�ĝ�����Lə ���6��!�`h}�r����7�?JުG�Co�<���������/����J��p2�#�t}m��_0"?�-M!�;_hz~gˣ'z�Lj������E6����&�,��F9 =�*��O_��c��l~�K�N�A�J�6�1�-�V���78T�%/�ڍ4+A~��Ga�t��s�O���aFYY�z��憘ם��E:`�k�K��>:�[Ll�
#l������������i�C��{�sk����c����)��TF���0\������C�^�#�loRɛ� �xy3Yg�����ES�uÒ���^���-գ�WG��{�^���τ-`��%������f��L�Q����
���8�yK���2Lm�e��`�朾'Q�1�ֺ)�ɇ��{����95B)5�͕����;����iw�Q��Y����� `�B8��[?���Ft'�w��s��K{����[\ҕ}��D>��!�"�����S�i�}Sx�M����e�3��9�
�Ҿ��<�=�Q�;0�<Vߡ� ܚ���sa�6���m=H����n%ڄ?��a7��BS�(�
� �7MS�b��;Ӻ�i��d6��>7��̪&	9��O)}���8�zE+%},P-��\:�W,�P"Z �:�#�'M���t.�Gf�)�9�Sy� )ׇMK4c�6�����q﷟1�Y?.��lP�|"�m�\P��d��y����m�Szf{P�U���L�4����C~KF��3�(և���zH�u#0�\�{�7�v���3������2UW�)�A	��?��)V�\^������T -����f~�'���Z?5���l�|:�x�9��r��}$8f[�����G G|g��xW�BfJͯa'�޲Pd�m,+�אꖳ���u� �瘬k�W�� ���{�YF���[���!g��6�ȋҀ��]o��ω��|��:�wx������v���d�~.�O#2Yt����;�	����TU�}���r9��&�1�h�z*��M�y�n��(6k�Ղ�L��"er�iM�?8����{�S�lT��r����g?n�(���*�i�䗅%T}���e=���~.eS#[?RB�w�!�L��*G��Ӏ�S7}��d���"���e̽ ��s�)X��u΄�u��r+3�Eji-~ދr�Z ��^Bb�A�}^����B��)2�D����Y�^S**�ܒ�X���4������yT������8�Ph���+j���X;���_���L>��oc�qW������Kr�+�c_J��"5[o�j�db��7b�q��ug�6m��x�n@p

�Rv�a��ס;&�<�:n������~�xN�I	?)$�I�8޸�N�:)�'����E�úz�|m�uI�),G�ܗ�J�i�=��`�,��V��6z-;Iv��ANj�Fh�(���J��@�y(B�?f�h���p	�H��&�
P,�N>�_�ݏ��h�k��u�-=����9�7�Ϝ��5�^�x��Z��Pˇ?v/!��9�C'�s���o�d���"���y*��v&� ���i�^/V}����^��\P�k<��j�"~tC}�7&�v0�RQ2���J��t�Ni�x��K�7��[	�����ד=��8C���:�}���vKҪ� ӯG'x�Gk���# ��o��1�̸��TE.�>�:NYo�3>WN��'@�����G4���d��:��}.�>d����
������� "����1��2
���k*g�li��_C�:�� ��`��5"��c�<�%�A'���k���DI��jҥ�؇D���%�c�v��t.�c��-J�N)�e�i"�*6G\�T)�y���Yj��ѡ�HQ5�{�CϝIm-�l�sQvι��`k�Pk�P�]�b�ޡ}c���������(����)-d�$xj�����u�W��8/��&���/�ҜC��g�:�F�n�~�뎣�Ѷ������H2I����!�6��� ���`C#*0~*gq>��0ʨ�?�hg�m<N�x[��<~�eOOE�k�����?sOfϷ�K�H���E�SJbe^��m����d/�`U!���6�{ gZM���~�0��Ȉ�js����=�����'r\�i$�M����Mst+��b��"�!�WR���5l�ٻ`���3]E���PR�#�����:nD֩�O�MQ�HL]�1E���,Lk:�m{��N{Zm;�7#[7�����S*��>RDǦaeZ�}��vRrl��Sb�'7�Ah �Б�u ��%��4�ca��kD�i����6̖��g������*�`.���v6�i��غ���!5���W�<L��̏�{���s7N�&ӯ���wA5�d�`QTW��.���
����4���M�o-)��3&N~bm�{�&:��x%�'q�Bwq���);ƫh����_(M�a������Y�ȧ�3��_�?�����ԵFI��{�W���#�2]ƹ�����e֎��i���*&�-�ءFʸ�(�a꣄b�͠�_���"��[^ i��}uwƴ�鬻�'����eRo�|�O�o7tq�6�$����Ø"�j�cL�T�Ŏ�T�_��;mؙ�WA�����-!� �����N�����ǛO��5ǜ7ַ�+?����#����W��g��D�^<����uzV1�
��؍E�F>��:�&bRĖ��A���^ܟ����}/�n�@R����[��X���U�IQv�jX�I!��~���Z-��Laۚ9֗|O�෼?�E+�NM�>xpA�3�:������{ϨV��c��;�	n���-��9 V�.���wD�Vn\�.�P[I`~����ڼ\��L�j-LE�P��`z��c=;����W���X�������&���q��v��ֈ�5�jS�(c�`+�)�{�䒺�����c�����[����┝��-�͢wr ���Jȩ�4��	��. �COj�Q��P�dL��UuP��DW!R"^��8\�lŨo�Mϥ9�$����_ITCg2)�����9�ʴ��K�S�Lj�"�Oo�9�0�o�G�8�tw���B�9���y�^!?c-��b�s���"	;��l8YыF��ĢLn �a)��O�:�s!�t��!|�p��mr|�Rx&n��2��R��(	�z�<&H0~m��b$�$u��x��j�����'%�B��'{>n�������R5t^o���I	؁���{�QK��n�ϬVz{�9V*	iL����c��G!����e���t��᧍D�1/�����P3�k��k��ws���O#�4�<^���(�A��.�a�\��g���:�m��"�
9�Yh-]�=��0���pԦ�烨�6[���5���x :6s����k��o]�F��H n�6y����z&���-[`0qe��+y�S�3sO6R���������)R��H�<��-��yk��sGp��٠�֋쵘ssy�O�ή���d��^DƢ'u���ig���-�շ���Nj��уtn|o�e׿~F�j*t}1Wi/��؈a㛴��t��!�a3��>ݗ��@Xu5�*|���m/Fps���!��ٗ����E�Vf"ݯ��dgI1�6����+<Z6��Ao�̵��6oN��r��IFw���e&����t�T����W�KN���^�Ī�lX�RFDY�'�u`�lq��ܐg�*�Ų��������o��0���}M���'��l��ct%<�����a�e�uȘc]Ĺ�m�R�*u^��7�j&_�ꕎ.��5RU7+��`�<�ײ�D8��L2~P|���tw�,w����r�5Qҙ�8�pq��½|d��{[}��z���zAR�5�xTWr�R�ۉ�6��+.�f����{(���,�,6>:V����v��ԝ}k�Af���v�U�t���9'iΒ�>��ue�tN\xJ
e��`���6�ng&��s��w�CJ<Y��rZ���3�\�YZIx��A1ˉ�n�qO��R�m�_k�p��)�&�{p�������Ւ�.�|�����q9��V�ttlVx��Ma�����R;;���R�����l�;4�㎣�	�'�b�t��NSn�=�@��`i�^�7�0No�
mD�%֍ ~�x�L&�g�}�I=��{��(�� ��L�CXPL!���iw �;5W�b'������B?���N������Q�j	𖱵T��I�6��{œk�Np��/ׯ:1i�40�Ϥx�%$�x,�E��g��&��1Yy�'�Ӫ�O�g��7B^7B�Ŧ]���7=�D�:�5��w�f=<E�Pĕ�k��Dٷ��$�5E��\y����[e�65ktW@ŀ��#B�w"Ap�O�����n{~wی܅ŗh��[���D�{�Zwb���Ix_y�cpWJ2�G�"���Y��|#$�'o����;�L�\�!�<��Iൖ����w����Xs�-i���2����庫����Fƴ!���˚+�.O2�ڼ3�o�����E��P�]k$T����*����n�
�G<z�ώ��ٝ!�cWR��즧hfZ���&���6���[�Z�
�*����.��%o���ihK�b�����'?�����v(��ڳ|�uf�Gq�F]�ϝ@7�{m�����vL����<(���H�i��gJ�0f1�3�l62�X)=t�Ƙ�e��g-햡���B!�v�@?'���-�������H�>���w���V�[�[��Ŭ�J6^b.t��M�X�B;��Vuڜ�,��<;��1�c�+˯�b�%j��kC~�Tx��0D޹;�|�:%����d�\�0uP^L�MV�.�8=���l������5�.:[^y㠻J'=�aջ�y����rRŌ��SI�ւP�������fzA"3e_�'k̈5Om��]�j�h/�V��)P\Ȅe�:�/������ᙔ��hG`�1ﭸcۑAu~R|��90Nt��p1w��y�n�5�R]�mZj�z�����P�1��F�\�Gab��/���Z.��Yf��� I��
�{X���n޴(�I��[|A��>v�9��1v��
ˢ�mA����첤�M��)�2�2nχ7\7��]�����P%�fI�-���t>��м����@�CE�"~t�r�0��,Y{��v�d�yN^�6��f��V5mG�z�&�Q�'E�����v�Ā�]ҋ�%�����m_��rj|<�7W:d��>;F�}���9����1-*�[L�O�*"��a�����s�Us����JVz�Y�d���H��&��m��Ơ����k �m X���:������:K�In+�߬�>9���I@�{p�3s>_�_i��"4:RoW�VfV�L��h�4���7�)X%}��W�c�����-��3��i�kG��]E秧?DFL�����g��獐� �U����X�L�.�jp'/�
)s��;� 8|�Ѹ8
�J���2槹%bcnL�
p���U5V6�kra�}�W����/d���i����]�����%a[B���W՟��ߓZN#�4-4�!�Y�~����G�c�f�,x� ?
��F`��[�gqb���K�O�vD)��-��yS��f�^U:��ڽ��4���K+��݁om18��XӒ�"�:��.fЌ\bׄ\⇸�W��n�	h5�3Z֞�������b2�Qg��E����"b@)9Q{���f�C7���ּ��KiI&�3
�����Iu��u͊�%���<�M|t�Ա��� ��H.`|,�����b������e�˻�2��olB�����+b7�<���YĖ�[�	j��z6֜C����U=E5`���|�mmTjN��.���4W�0$������j�ܔ�Y;b\!�z��H*@1�p�*J��l�ʌY�^�m�J���J�u&��������߉$Z�rz�Q�B}�����)��i���Vn���te<�h���+��~���
���t^O�#���7��kH�����~̍�_'��3;�ڄ�?N��ʹ8��CeJ�^Ϲ߬=j��i&׵0��
3�+�+@`�63�����NyHw�k���nmk&-��D"t�ђ�� �@����0!C:�^��~��J�KP���w��1�k}�[.��10��PX#ǉ�=z&����Q�L���'o�T��a0����:�i��\Vʆϸ��0s�Z<�u�S���|6���_���I�pWk�$+`�ͯ1�#1?]~��BA@�F9O	�q s����࿬8?����Ӱ.��T�:$��NL3�w��e������� �Ǚߺ������1��l�ؑz�ws��N3�<Mhw~��{Q��LSI���B���j�d$xd�_�̉{�>�$�5�3-���uK2/zQޠ�z��(��ϏC��B�	�� ��*KhT�Z���mf&��}�����x%		c�C�F� N�O��*��#{Gќ��uTecpfb��_v|��fpK�����.u�Ht���M�ī>�q��a���6	��jA��~�-?���A�,�]Yt73����K-Jz`��{�c�rJԚ!�m;K3wD�<*�z�&ޔ��[g��&�Imc�yٝ��qw�ʟ�����J ��Φ��p�U݌^���U�v�Z[o�g�I
�����k�����X�1�v�/~�K��n���l�t���`��Y
ث �p BN���%�P���ߵ?�U+ ��������ȅ�߶_�X������$��\
Z��~0��A�Z�s�"�0^jߓ��L���])�GV�P�;b�\�c�~�^^P���u����q��Z�D����3&���=v`}.�i��B�&�U\P�3V�~�i�QU�*r����hV}c~#��Zw��k%i��k�.�#�t�[�^2�p6n�S|zr%��;����rA�f�`�+`�Lz. (.�Hfr��~�6Iy����jAVǒ�Li�CN��.ߛr@w�
�Uϴ���9>@�-����׆nVO� +;���LwP�0d{���ܡ;}�]�zb-�$�^ۡƊ�����-�?J=�YB8�BЁltF�Et�G��j�v��^�I��%lĉR�-6��K��󛑸q�z!��!ֈ��t�	X@>E�i8��kGg�Ɵ_G�Z�].`�q�M�1���F��>�~�jކ�6��=ܟ�f'�޶�WN�&��2�� Rޒv&��u�L]NB���e]p�J7�_J�`��]o�.vB5^�W=,�w'�z�Ten�Z�Cȧm=[��o뙟�}q6�n���E�Xԛ����Wcz���5�÷|3�qj��G�R�K��k�^�	�|�.Nk�K'	�Q=v�t�42�X�*~մ��gz?ߞ�q����TH\E�R6�DH�h[�ϧ.o����(�&�|���b��ǡ�t��P#�{�1�5ް�\���K�� z>�+����K�h���] S#v�Q4�I��bv��"��Ɇ�O�ë�_H�::� �q+$�!�Mh�WW�c��mh�TD�J��|PG���u�~N��w��Z����ڜ��S��"�y<�'��y=SSdrUʅs�1�4��5����8;����-u��HSAt�eU��՝��j���Zk�>\\�X�Qؤх�����Av��-@�!糳�Y���+N���S$1�e\W�W�%��"/�^�����+Q��Ҙ.P�Z��#�e�iUv�B���I�V�
�#�(鸃���.r����{�Ws�ɗ"��ݡ3� ���43��t!��֦S�z㮵���/`�9�&>���C�;��@o/�!��n�[�6)Wm*+�,̷488a�[e����O������|�XD��mw�s�VI�ʜ�e�����m��#�U�֒0��1@����`)�vW��s�i{�n'� �s�Z�����oR�W2k���J�,̐9��x��^�N7�͆�o�@���oug���m�����I�}kռt������>�֬��[��A�R���K����0��{ȏ�w��UK9D�&�+Ҏ.�*o��c��u˶�zT������0Plz�"l�C\�|��Zb��U�z�p�qIR���ŵ��i i����@՜���n��8~���닰��N�y1wW�r��P��9��Z#�U#y�L�Y���޻������V)�����G�L>q℗K�_���Q��gHF��,��Џ�ԭ�=ϦE�����`�����������_�
����:|��r�sw+/�\�l�+��9��7�3okp
|+L_�t'�����]�Q�����ɾ5TK*L�
�]U V�:F�^7�CV��a���$V�6��s�g`��q.ě+0
ś��*R�\������z�Qj^���;'��+v)�8򵐼�s(��E��������'���ʕ~Wa�����]#7s�t�me�4D@�����WY�6��2������>��CB�S�/�e����B��ۑ��;&����n��x�ݏg�/]I�	�#;�ӡ�JO@6�Xi\0��:@�N�7�Cyzc�1��n4�8友�J��O	��-Ox[C0��=!��cj����e|s}v-��M�`I)W&R���p���gחr��g���v��y4}o��T�GP���HQX8�FK��^�~��Obk�J>#�aM�y!���Z�A�,!�N�F>�Dg�;�8��e���=]��J�-���ϊ��<#�Ꮎ��r~:�������2n�e"��x}%2ʶ(%�-�?����V�����9�׳�s��\3.�po�u7��s�v�Y���8��fN	�n:�=s����4��l��F�!p|�J/���7f�y���h5Т���p(���{j<ͫ����PNRvt���@
7W~Q����2���$b���J����k 퍕���вd���_Y��V����x�X�Ulڍ(e�w͗?�3�&(�3�%9��?�}�|�E�2S��K�X�nX�C�`� 	~�'}d�N7օxz�~�n���b鄹]�S��*��e���'=�����u�-��.o6�fx՗F( �Fz��(FC�'��Oq3?�����} �Ӡ�6��"�+�/���ç��ѧ.YLLR�^hxD��D}��Ԙ��@9x_?���7�p|�ȋ����fUJ%.X���]N@O�F�.-y�E��Z�2��ʞ�-��N���Z��xh�����(vx-�7�9V�FM�>�!O�|�^�� :;o�S��-��A�O�L�~/Y﴿_�XO��YL;�^G�� ������LuJ T`K�3	P��C���OSL(˫��Mq� �0���>��4�2f����Y�)@�}-��g�+�X�(6q�u���8�*�z�
�"��n�0χM��*`��6�z1���>����ƿ��q���)s��U�2�f1���pO�d$�����<�3�2%���A쌑GX� �_X���4wk��@_�홐?H%�hfu�!�v��p�l6T���[ �z�_��}'�R/���@�[�ݹ�{�����?B�� 5�.����Kے��`��㋣׏!����24�wr#�~J^t5��R��_+}[l��]u�,����c�L�G|�޽$kB�vg�|>�K�2�G�Ӝ�+b9^U��nk:��T���C+��.����Y�O?OZt���2��v[������ ݷ^߸K��['�)ֺ�*&�����)6M�Y=#� /2��Z#}M��GU�.��F�>Y�l��-]�y"�1�y������.3�Ȱ�^@�<�>���P�r��(���V�j60���a�{:Lu�'h�~r~/�$]3���M�m+0��ڂb�M�*]�����e��bQq�8o�� �z��q�޼jy1+�Y��/��S1�N����+,T(�Nki����~��n��uIx~�q�����>�**��f�ވ�d~S7��ï�#���n���%]�۔3mAya��#�33��,��P�%,WId��E)���	���S�a�6k��=�E+~���Іgyٶئ3x�ئ��'���n�1��d��"p����v.0���x���`�����(����FYF`s)^i�P���F�(I{!%`b�W��7`�"e���L#�>�S9DI���e�,��o����p�.�*|�+a�9q��:itSd>Aϥ�Γ�2�Y|��M��<����ݥ�\*ڧ�cl_��?	�����Y.�������^o?6�M�W�"A��>��v�+�W\>#vV���=aY����^�xy&:�:s��F�wDE�Kӡ1���wl���U�9j��GaG���_H����2�p�F�q��ۅ���|N�1;+��o*��#]6��A��B���^3������M1�<��%{���f�^��������ٛG��M����(���6�=;��'�;t��9H�c�o���K�w��\���.K����d��j��jU3����v �"�4AF��;:�;�\�s�1��� ��O4�T4�`��F�V�\�և�ZUz2��o��l�	��0u���ei��I���b�;�Wgk��n�3%ϷW����ߌ9܂%�ދ�d�+���no��r� ���K����^O��=�ɲ&�؜ry�`�o���I��w_)��u6���}z{7�Q�s�1�����������n�ă|���0��D�+d]Z���A��er�Cg�����lֺ�Eb��˙�ms
�.�:���g.z�<պhG�����eG7hxv������I�+݇���O��Aj���$\��'O�3��"|��S�3_�vk��۝7m���Q�r x�o@����k���ޞ�x��s�����,�2��NzF�~�t�~t��j���M,�}���X�ӜX;�|t������~�(�^�`lA�
+�����"^�\��5"���F���E:j��X�s]]�띥���؉暑��7"F���!7~��L�;�m�K�1�)�K�\�T��*Y{��\��G�(>�Th*�#={���`t�j�=s�ڋ�%��4�d)�h���u9�o�Y<�3<F �1u)���1����>�;֕66 �	�V;�H#9�ڸq�v��Z[զC��JL�%�Ua{lI��w�20~��NOO;��̖���.}T�T`�>s�Ve�+��ɳ�.4IǗ��ߘ��mй�M�Ð�"j2"�[�jHȁ���9,υT���iE�7v�X�}EC�V,����B�.=��������#p�0�)��4��k;�vi�C@����|���o��}}o�%HY�0���xLp�n��̰���Έ���ȭ��CmF��q"�R*pp��p��`�r�Ή���*@K�?��[�����fk��r�����1Y�^�.�+�)�A���g��J����܀�+{�!��r[�?O"���mg�cL�Z�d{EW_�`�{�Y�͝�z��,-��wgd�D�!�o��9�I�9kOV���?��C�h�G��}�Az��QDK���]O�h0 }�S�Jc�V~;�!I�]�y  ��_��ʼ����@�����7���(`�Q��ɭ��PDa	c���Q�"��c-Wi����k�s�b�ؘ7�Ŧ�W^U/���qM�	�2$���9/��v%}7�����<��N���)#5��;��,��o���-�����~2#��I��c���"-�MNp{9���k�ZG&�3瘩�Up��؊�F �.�o��U�ŵ8º�,�*�|�ڱ���a-_��t|3_�ð�J%���%�����7_�J%�ta|[3~�h+;O�9YmVl�w��|������H�P!�oF��9J ]ٷ?��vU8?��'����Z��N!I�e*,�e4 B���ʤ��|��g!�6�t��=�RO'E���z�w�:6�B�b����@�Fg��tmR������u7����P��[t"W	q�u%݄PCNd�8O~.���d�I�Qb4û��b7^��&��t<4��24��Id�]I���<�;�&�l~5<�G�Xj��{�f��QLV�(�C�me�_�۩�و�ȯ_p�[X�Y����y�K��A�P�;�����%وhwu�Ne%:�[n�����A|�B��`���{�?���y�T�`[@*�j5�]�w��������`��Q猹�����ob�,jEW�hL��ĠoԨj/��Őj硎���j�4]�T��Ydv�z�E*CLaZan�Z��<;I�*]�%hL���;F��|�"l�����BK{{�Ո�8�hȟt�iQ���\��k�'}����R������̏1�R��5c�#3����C�{�GZNX߫A��y�Yĝ��*�µ��҇\)��{F'S;��Ck�GE\�e)ӵM����!IT�Ӆ1��̺c���3�m�y��
�<xk��P�~��?
�̜aV?�'f���Z
�1��7�Eg��('dr�g�&�p���`���/%�J���C.�	�5���D-L޵�op�?�EC�͕E��[��t��m'�7�T4�u���)����'�d&�Wv�ں�ԮP�zĕ.R`X��V��-~�d�C����3EbWi$C8(:O�5~��O�K-�p͏�J���f��]/{�
ʶ�h`�(����"~V<C�]A�cre��Te��"-���
�G,��̸H�2�m�z��P�<���DLT��W�nZ+�%�(�IP�%�FA�aH� ��V(�T�:�#QS-9����B��s��5����z<����4�@j���lL����-��8N��L҃*jȎ�$ *��3I�ɃW�ޠ>'u_;<�!�K�I�j�.�>E{"����Wp��u�ցR�Kqw� ��;w���R܋C�(�N��� ����\z����1���kMYk?9<�G��i��)i�3�m%_�l�������g༈*Q�[��³�O)��R/B�&���3;��`|?W`�>��>~���ō��L���oܞ�+��N1�D��[i������8�S��x[f�Xc�i���W�͗��`�G>���Rj�QJ����.�^�<`'�����Kj�r�|'&������5m$DA y^�x+2�J�ʚ�(�5�r#�� s��P��R�b�WGܽ�a�����ߪB��Bu�R+��o��
TZm|�eC2���l�T<�r�b�xlU��-�����&�b�����R�b�ҔF���}�~�k0���`���0����l�-�}�>��l{4�*M	D�i������nUx\
߲�\�=I'e��A2}�{�a���@وlˏH���f��e�$*1����A���܃�[��zi��,��3�Hލ$��X�ܯ"�鿯�)�/a�|��rH���,Ɓ�?��K�k��יO:�?r�-���L+�NGݚ���W���,"��1&�	ω�O�q�ZPM�`g�R����3yV�E�la�O�T���I�a��6�ҟ��e�ߦ4�>�	~�/O���l>T~j��D*�C��T�5�4��V�Z��;��|�>IY�;�q���Ç|î��ϜC���WI�i���x����J�}���i|�{�V�T]��'C���s���l��+�<�Wd
��<��=�%Τ6>b�酁)���g�C��Ul�JC!n�$([	x|sh:!��j!}	v��"g�T�΅�i�B̍O�2ظ��]�M铘��EX�'dڂ��!�ʣ���l�g�m�1&����^p�M��#���v5;јfڠ�tR��a�'��u�ģ--5�U��_�]�,m��<SZ��"�vx
��uj5�qWM[�f�c�zt��\ۭR���/�c�3wN�_4 �u��ōo��_S^`/{^�4mUb�y��.��Y���d��ڙv�<���e�e+��f�M���
�2O$j��/�_,�����q�N3�N6�?��/o��+RO�d)Er�y����2���_���3���gv�+;��y�����]y��	ח���6f|��j6�$�o��K�Dt̜,=��Y[�+��K�IG���J�rJ�w�(z�c�b�\���Sۍul�J���R,����ns�ӻr\#���jP�6"��|��}���&���veYY �6�!B��I���ڻ	��f��3[��kR�W������ɖ��D�㘈<2f�1�c~�6֩%�ݺ̜_N�ƻ�s�lE_���Y������:�T���m���.s�ki�m��U��� ��v�*��3�r��>c�D|:��� հ³)Kuѷ,�4h�5�/�L>{
wC�����ޣe���D<�ށCG�S��9������o]���:�ƙ��MPS�%�ca�{z
�x��*����3o����
���[&��!��	K
�MCH��rK���@iu?=������ۿ�-t��L�+��F��Աz�՛�����A�wG�ʳ����k�E��ޔX��R�����Tx"O�s�����O�6T���8���vaOU���0t{��I8N�	�g��6셔�����y��|P�ۢ�j�zQ��f4O��rlh�v��ʃ-�����嫧魊�{Ζ��b�K�����/e��&��v*���;�6S�Y��7jk.ϸ]2�x�I�?7)~�I;#!y	rx@�|*�?~���Tc��
,��F9���/	�c,+T�uW���B��l��U�����k�Z&��TtN �^Ó���E;'ص�z�r68��,4�	�R�x��x&&x�0|;h1���/���w��1��bH�P��o�x����̋#"�db�Y����>�V;��c��>���W�ţk�Ä9}����ƣulC�}����Փy�$��Y����^wVFc�bHt��F��󦂌����f����^�\�$e��G/P�Oid�H�9Z��ڙ�'H `����"e7`���'�
��
/}����e���8�^f���br��e�?�������2y]c��x�PS�7>�Pi(�W%,�PG����R��.�lq����D�	�}5.K�� C��=c��>��ll �t)ܙ�`�k�`���	�U�B����I�y���)v�G���v�ǝ:vV�M��H�ú��!  xU�������
˙����Ej�"&���n=�RR�zLMmѷ9�<�P�PV��
*�8��B#c�\Z^�>o�Uޗ�J<g%x*|��P.&��:��=n�V�v���S��%o��o�7��٧*��С����!n99�a�t�,76-�&�o0�R��l���&d���|�T���������N�Xﱭ�{c��9���A��؃�k��ʙ���X�j�Izoc�^s5$�V0f�׋���:�+��sޢ��X�e�[#w�m(Lv��Z�|�}�/�Da�'9�a���ѭ�ˀˌ�Kd�H@�ޡk
��,)�t�J;�O�#$��%�<�8DJTk��Y�����#�:���Պ`���5Cս9��V�稔])l.�����=x�6��%v�Kְ�8��۟q�7�b6EX�p�|s�� K���ߣd�qOJ��_�Bd��_�����C�u�X�/2V�|�V?n�r��;P�]�Q�TVI3��-���)�o�+����o`� �.�����f3�y!��3�XBқ�W]�]���i�����_���/эB�qY�~����[�dڠҎ�A�9���tK��hls�������������?�ō������!���*��y\�C����q���=,�����66B����M��$��7��:��9MOf��JV^n5�R����æ���MX�A�v�#ں��k6�z�/�f�bZ#���AU���)L�j��s~b�)����v�z��x�Y�h�������&�ٱ�;u�����$�'	;�-�-�n��Ɖ����
Y�Z��׍#�u���}ɇ��Ly��ɱ�@���M���̋��YCk�qca��������qQ��
r��D�x�CY�%�V�_.��[5
�Z��<eB!����O4�g�����Ű�� ���
]�x�Fs~��u~��)��B�-f��Ձ�ƿ
q�?0��7��MW�����'�x�'�کň�.���Z^=�d@�_�>#1ԉq���%+�� o�1���n�S��`&^4��A���G��w�J
�>s�CWn��ԁ���σ��b���(��a�uNf��R�s�[�-��،Mѥ^0%�%�8Ǔ�\��ϻ�<Zˁj�~�c{��Nes�N��ϲ6�n٘���ZV��&����E�Qnb�N�&�ao[�ӂ�+@����*�l��E f;���Fz�	���@>ĲI��Wؔե5��f�3����	����1�ê���ʛL:L�2"��r���
\�K�3י^�^$XU�,���Ef�z�'�Ҩ�A��~&g�5Z���i��QI,�ߩJB�O������1F-�Y���}��w�l5[
����p$�M@{�p�&(-���[_�Z�:##\�SV.َr�?اfӴ5C#,�磴��ԛ0��ͱ?v���D$<��nost��RO% jSA������dy���>ȝv�*+)�(®��.r4|�2I�󧘈z���	����2���Ջ���A�U"l'���"���~ǐ���,�d��SA�:
���\sl�Q�`�D�����)��Lv9|W�p/���>���h6o�����,P^������4O5;���l�{�߰%��bm�sW/W�ה����y������]ZU8S��	�g;��) �=���[���1�df���XI��A�X�y��[������>����2ݛ��S�6	�pB������D>�Z�I,�5�~��L�F�#�xш{�^��"�k���z��.6�a�������!�1Tռ�(��y�b:�-k���E�4e_#r��;��-�r"jM8�Hۑ~?)�@����}=F��g�p�y])�-��ɼ���''8$=��W�cDC�Ѕ�2�۽�m�&&��w��-LPC�a�d���O�&���1W���ʝ2P�VoK�Z.�\��"���!�Co0D(�Q�o��� �)~��H�b-,��U���9؃lK�V��}�/I�b�4j`�jL:��Gnt�E	��Mߊ��mA�K�K�+�2����&����CJ�s��w[����[Q-ȂB�.Qi;?��Z�(���sJ�F��KR�̏{d�}V�����#�y٥#x��n�q�,�hzC���xn=Jc|1a�AR}�Nߴȍ�zv�O�6���>���.�7J�@c'��N��>w&x���[�7�\��GQÒ��|�zĂ�/�c��\N������Xu���7�����T����!� �}�N�'�r�g�W�z�.=��d��D�(}m�Zh�x�k��>e<=0�5��U�uIZ,������:������Ki��S���I�Ȋ`Y��p�~��%�.^?����T��]�,�����[�G�Fw&���j�5Dng��S��J���V�����+�5�i.��!̂Ѡ��V Z�yO����j�Q��pZV��(+1�g�|�+�OϑM�N&�5�/�w�;/�s�c )�t�6��'���O��ח
��ٮ�%O�?�τ$��J"�㦅�BQ��;�`q� �0oEU_��YM�z%�#�s�o�-^�@f���v�6?;���IަGJ�iG���Mo��Tu���r	��ݝ�v��ְNK�O��,�Cm	^n=��D
~�<����w�W���\Dtp�6¨��r�i[�{9�*��z�eaf9�=:�c���t�WR岞��[P��z��
WIzqi��#���C�̥I
����|6Œ1�(��!�ޭ۵������W�C�����Կ�tm�?��j����Nĩ�]�x:9��mO�<>��jS��V����2�T\�nC�TG�`�}+�7ʉ�,�^(��nI����H+�/�	I�����%��0�cȿ�h&�M�`'����wLUS�ő���ڂ����R�5�]�mk����<�OA{��'�f��e"N���v�(���ͮdT+2+@~���
�k�ժH����;�}��C�;3�_����2����Pa���/DI�N��!��f���43���������DaZ����[��F ���
�?8[��/��q�|j�V�^���X(��r�S����K�$��r�`�dVL#�!�0���2�DFKO_��0��/�a�x�X���R�f�m�/�_.��f*�-���oԳ@1φ�I.53;=3����y���-7\|�pr��+�=+���l���|S.lcƠGa� ��@16V�0C�6	g{���c�8���1��~{d�L�[8����T�fl��O�̈́A2]�Kz�{%$,JMz�p�PW䉴<�5님������;ZO��	�p��rx�/21�F�=�9��t�e�yr�h���yO���}��V��>c仞�-,;�7NhEO<+�fUyU����i�͢�ߙ�6^��jΦB�~�z�O5�:�k�m��̴�e��5"��ѐH0n�4�Z������[��σ'`��(1�ɟLR�Q��aW��g��g^�F���B�*>��ŦW�
�a�G�z��$Mٝ8v��Z�^�8��6"l<|���Y-ەb<�`�[��\���u6�ny,��TA�W1�Y,�o�w1��>�w�y���"<YL��T������ �J�#�kC��O�n�>!`lqf2m�z�Pb�r�mf��ݒ�x+��5�`PJ����Z����gh�X)ڌuye��ȣ��c���.
�Q���u2�RHV��k�2;ү�lr�A���ɷ�n%��䋿tt*!Ie�6���ws�e������v��j�O!��9�L���"V��K��1~��H��	o�������?�_��2�V��hƛʘF%���J�W��D�1�Y�Y��$��F���x�DP��,[&x&k���׳����_�cօ���H���.��a

@�S)�h゜�A�~範I	Le��� ��a��S���"8������S�Bo␅�@?�����s�:�w?�.*V<����i�6��s{9T��b��wqU���5o�h���q$�v��Х;mV�S���N��:�E�۾�?�x2�=	���Ebڗ ���W7����B��4��n���t� '��(a<�Fz��Z�%�D�z��o�x��@O��ZU����gļ�tw�E��v�^�>2����	ARcU�G0�n�p-dcPz��M)��g�c����	�wG.j��f���.F�o�Fb.$11l�$-��f�$12�H�:�f0�	K����ޝY?8��P�X��ԌZٶ#�U����;l�mC�z��I�݉[��|��J�d��qK��p��%(J���p�S���/'��#�3)7����֥������v�^o�TqhD�����wJ|l|�6����qUS�Cݦ�3a���>��J��|hm��c���Da��u�/�<�zk��Sf�]�I�պ,����;B�욌�R��E�1�-�� ������h�}��Ej�����H+8dmow��-�$rs����!� �mA$:�`�0+Z؋[�|��� �H[�ئƚD�Kg:�>�
O��-�n��(�Ѓ;d�7��*�����~��r�^�"9Ɵ �w��G�4�� �G��&�:w�:="��c�<@s�5�/�o�ot"��7��c:�r���X�oW�����hf)�?�P������yJ�L�@�q<Y��m��R�����6,�r��1Շ����?�Q��6�4�f[(��u�lhR�����`y�h��(;�=��b,
�.v�u>]�a��t��ٝò�|�hN��s��n��Ds��%�ێ�(�\B{f~��wP�;O]�q�e:��|:��ñaX�<�jfJ�!�ߪʝ�&�#�~q�QA���nT͝�ݻt�7$���(��3��꥖��GM?
��@QR�_�2��g17�͑aR�SB��0�"S�r��_��oP8-�p�u�{K���^�_��䕄M~MCCH�$8f�]c���n�;yɑB��{���.�����b\�Y{c��`h���	���<['��t������V[h�����Fhpu�AҾ�O,��������Xt��K��O���1D
*���6@q��^9{W��xd�`�B��5�fݬ����D�N)�$:�,,j:�����C���w-2|K�J	�(��yA!���WS��NV+l�5 �$H��'�(�c���_L�~��~�JF~�����m"x�vw�������(2qW���F�U��8b�+80^e̼�Z��c�c��J{�$҃o���[82�y6�8��\�f)�ѝ�恎�wK���=������^�형�ƚ���}8z{Qw�阀��A�|��nj��O^�b��[��l����i����#�@uAS��v�lk܍ƌ��RY�iS%�@����7�:�nH�jxO�q"3	�h�-r��h� �H'گ��=�C��o�H���^57cb��p��(��Fٻ`꿃G����_W�(M��~�U����2ic�ǖҖ�}|�+��E�~��[7�?��Ǻ�����a������!�)���w��}�����m�����!G֯�>�v%}�|�H���A���Ͽ�+�S�X�M�/���H,7;�p��.D�G���=��q�W|u_�L �r=1
?�b�-s��8?�;�k"Ra��D�)~�F�F��N26+���=�K�6Y��E�w��+����k�D\9���N���`?|l�k����)�����O����S�:RUO�=�N�]K�0�����@Y��y!�J쵱��������%�ٍ�9WA�*x���R�����R��[6νmϨ�K�� ���m>��w��˧p0��t��4t����tۭ*(�͢����O��� վjs� \���lP8]�!]�c	/4���j��X�6V�7�YYPOC�b6�M���b��h��. $}B^@!�Kv�g�d�X~���`�}q��!���z�NE&紦�ad Ҍ�z�Rd�Щ�������3�%�Y��\�>�4�z��NP��D�-�x���$���ͿZ5*� k$����b^Tբݔ�P^�x+�nt�߄>$��g�k��0.��q^�.�Xi����)��VQ��3ܩmV��"�)�D;���3�O�/z T�ن9�5{Ĩ0�V�M��C7�ZA4x���T���Gh���2feb�or
�p����G��|�Y��j[&8K���_1��	�RG����\*7�+b����e~4yqud�HZ4������a��$���=R��֧���l��*�6٤Q�#���e��Y��~�-��Emn�I��'!摾%*V��w���	�4F�Ҹn��r���	D�o1~��PeB�?.H� �<3����h��?�Gy���K~�����u��'�U�n����'+�[���c^�k[7U����Ǜ�>�BH�Q��b(�~ +����k��y�t�[=�.�Coˣ�t]�"��F}@NF=����T�� d�9f7������4���ףb��'9�Qt�8:RgE���KEUn����lϫ���=JkH L��7��d���>��)�t�y�<~����e��R���曾ֆ�3��&�,�_]W����	m��%=/}!�aZ_�s�~�xs�
I���gj!�5�+���<��Y�<i1���=�Q9K��"gD�6�mS�%Rh��q�ӧV�@�-�^�w�"Z����G?��<�j� Y_71^�1� lM��]R��I�+��/V�#Q�١�YB�����_�ں����<k���ũ�11=��� �*pO�t�ů��N�?�+Kl��j�>��x��#�qm8�_YQ3�ӻ?�m�,%v�0JN�����B����(����^㆒�>ip6��+o%u����֣��3�]���|j�������&�1]�F0�UϞ�|��I�[刦^�]鑢�fEt�W���e���Rq�^�T�w ���P6�z`�e��N=&��/��5�z�?Y	��j�_~ ��2�W�r�⏱��鵔���G"��a�|���B(��G�})�Vъ�!k�B�M��/�'%i�[tޱ��ݵ��T��;u�/|�y���\��Y��{��0d�%���fL������Vd���m�;H�E������$�q��W�'%�ua����ĥ͎W�Ǚ��~\��o��U�Ͻ�2Г[᪞���~��s�S{�2G#��WGǷ�;��|UY���&D�S�g"���&:/Z`!�(ף�Cn<��{S�J�b�w~�����!�4��:ʱ��!Z�[�ِ�m>����ͫ�A����QL��X�����R��m�^g�s��;��3c�v�C��{O��$�X�H�Ť�f^y-�ϦV�;�E���Z5�2����"��Ī��f뚢|�r���W ��L����6υC�l�"�?��6CN��Hl��[��e�����ٿ�<��xMeR�C�����Fѿ�n�C�:p�����Q�+
��eT,�?�f�&�������O/>.۫��Sc�����a6=s+Z�o;׶�p�b��Ѽ��Mv��`~S�=@*��-�bͷ"� �~m=[sW�g�n|4O�B�����h�1fmQ�P�U�á�L� ���F�]�l��yt����I��yQ�qk!�j�7�Gf�S�]���B��V� 9�b`��x��QH�[�^9�1��gw���%6H�z"���Sf�w�q����o˙>��H���Z�i���<�0��w��<	9���+���,L=����N=>3���2�!���+Mչ1�3� �F����L�~��^:g7YWS[�S�{S��_��oߎ]��^B$v ={����Y�gz®���ql"?vz�	U��"��.��K�2D�E'�'~+.�Z9���gט�wI��D{�v�L�QM� G�viŅoh�����k�S��֝]�8	OAWܖ_7��Ki����6i��5��Cb��-Ò����s��Y"}�pT�6O_ U�.`E�K*/y��^8���/0��y�L؍�)E����~gI����T�ޝ|=�mM?��X �<�]�����+>����Σ�8�mDMs��$�n^�����"t����o�6�v0��9�o���r_�17�����گ�QwG9��-
�:M����a���chGM�m�Φa ����⺃r,3���^zH��?ߠF�]��ax�j�s�2^C`d��u݆~A#}�{��V�Di��}@ �D����s��uފV��@����,~���r�l��*)��������T!ƅK�7:�o��nq��i�����,�P����}�!��\\X����R"��Wg�R#!1}X��������@6|A��d�ݬ�����{�b�M;Ь�h�n�tϤm�=��ӛ���Q/�5۾P�0��_T��P����5�.��J����b���xt>MM���6�-	��i����?����qT�(���3�渊.7�:�5���eo|��f\vMq�i�:�3��vz���Q��Tz5ch�/�0�t��7$��Q��������g�+r>"Y��8��Te.%;�7�
��߉���ڮ����؊��׼��쯺`R2�U_�3��O]�:?����*����/��HS�h�'6luf�P�	�@�Md�I�t��\��WZ/Z1#<0�]�_�6�P�j�J�Br�����كP#����is�#�I%��sD��1\���U����� ��SS={�_C�3�J�7���	0>�L�e)�U�j�b9�?���]��"4�顃Kv#'�4а�wl	�aO�J�L,�<�E�u�n���޽-�����Yq�&"(a��t�8��n]�'h�����0	��٣*�Me�j��]�(kEP�/o�F�6�t�(��<Y:���EWv�ޤ����t��$;pӦW���x\�'\	r�&���nN���w%�{wG�S��v\)f����x?;p�e瀲;�.%�f����t:�@x�q�r�:�a=6���2x��v�%*���ʎ!e�]�tM׼yn��.y��)�M\"7�rC4�-
�v��筥�C�V@�ge����X�m~�D��;�m��bG���`6��A����Ҫ�zO��̛��P��.^h��<�Y�_c�Ux�d��3�?��j����b�Mf�h�)��W�v���>4f�S�z�6M���֢��i�̔�7�vj�#_��կ�_
}�4 ������\�~���#����5��ýz��p�!��u��Vo|����[�h��Kb���^�̡.l(�`f���t���O�x9]K�^}��h�B8{���95��nߛ�߇���\��Ů_����A�'s}Ju����X{�qtF�����jUh�r�;6�o�	E�ڤD��#[/7�\��r6��ϻ��<�9�(��i��-'�!�x��L��S�h�!.���6u���N��3*-�X�O�]Hz�������KX��Rb	g���i������z��#�Wm�k�;��-��0 �L�������z"�|�}�ɀx4��Fu�5'��ʋ���MҤ�Y��љ������6f���|YF��A�[7�щ�#ӑ���^�����9o^�6E��zA"�D�U3�;�f���ؚ�T#�c.Uמ%K����VʀAH�J��^D�X�!�����mK��d��G��ݜ��`�$���\T�ǅ�N�o?��j57]z\{������j�8�$�� ײV9��Ѫj���@z�ht�����ݬ�Ӄ���һ�n�-{)�w����������5��Vܧ���0�&�f��Ԥ:�I�Z�Ë�3b��8x<E9+E!Q�[=���1فl�+�20Ə��7�Z����[�tϛ/n�8���X���Пl�S���6��Ӳ M	�H/:���z|��PB�aMb&���
��v�δMK_�h�nkJZ����6��� )���]hד�Ǝv y�K�*Bq�l��mRT�!s$i)�M����e��Y}~[�H*ߠÏ��d ��ޏr�7y�6
rO�"�F����2���,�����C�n�v�� X�U�ڞ%V����A(�*�=z��"����(%�rx�_)�������lNU2�f����WBd�'�r5�x����@�b�6��4q����o�4�R���������>]o����+$H�r��?oH���ϡvPK�5o/�S�=��u�[�Mf[�R�/p��)�v�@"�|7�**�#�B��8ţ�wh���ՙ��]�G�����(��]t)�I���ln��+�;mS ]6a����5��]Ҧ��ͣT,E�et~ɇ{�/�drW�6�����|hymR��G�\�B?�x4�B�>�2�'L���&~�KҴ��tV��<�J6i��b:��'O�����m8ylA%��<;����J$�����&1��PD�P|��}�&F��F0�E�\w������b�Ae�:��o!Ӥ��-��h�$F����a��I�����K�^p��� �b�\�r�O��6z���g�&�K6���<����q�m�ǽ4�Y�ލ��M�]�.��\gQ��yֆ�%5�^k�"u��)aS-鵳K��*�ϟ	���r�{�e�>BL��k����E9���6�^o����Ҟ���yb���Qe��A]���*'���i�0=�@���R��	{���G݃�����j8*�^��������{&��%�6_�\��n+�Y���9�򺯒g������eo�>�*����f(��`i�<k�AΜ����Q~o[�0��=���ۧ�<u�n��m��~��#Y�PWL�nD��7�}p%����j���ȇ������s�_�"i�fr<��[��Zty<^��~Pd6�ߴ�h��2{�ȏ����Q
!����GO���E�h:m��S��V\�d�n�i9Ϙ�������맘�~�z ��Օ��A&@�`J�	UϘ{�B;U7�ڬ����K"ot�m�rtm�&m �g)�3si�[ep{��%��:���6�ݠ��'Ꭰ\8d����;�������6��df�V�섩�c59Y(��,�8�Z�н#��ӧ�2�1� ��l���gl2�����A�s2����嚤kX�Y����0�:=?Kc5��2��T<��{!f���{�'��ޕ�����}BtR�{\a�w^����&��W����%B���^u�͓���8��i�;
�U�	���8�p0�`�d�Ɇ�}c��$v��"��I�p�:�]��<RE��j�u%�f�%h���Q�]t�l{;8��q�݉^D�R	��Gw�mB��]�L����jpЛm�O8���K�"���+cp�e-~���ag��W�=��_��	HިȒג2#w8'<����}&�m�連<`�ED:����&sg�">����^���.{�㚚�i��5"V$=B��"����N{����6�W������l����0�H�	��>(��W��b�Ju~6P4N�(,t���w5���w��+!p�cB�L��W��H����nw���=:8���t8˱a��@�l?>ἔ[��zڹɀ�n�L�G�����p�<BNƃ�"ۼ���8~����i���~D,66R��è
�B*��9K$�V}ّ�,�&鯗 :�kK~Q.3f�ӆ%��yK<���e����D�����Ň�\�?�b@;Z����.�[Fw�,�]�^bP6���Cj�,uI�$��o�;1Wv��4�3�S���|�k�5z�A�>U�Uiē7&�a<�����#v?/�q�G����7��xwO�n�[�M��ٴ��>�=o����2�ل�E2��u��W�U;��U�.G%��� ����i0��	IWVK2��Q�Ń�/��N�op��EPVŕ�̻�1�D��x	�lyg�$"yC�&u�K����������p_=�l|�@kA��!���p�D�t)]�)�Kv���̆Y��R���a��NZ2�Ê;��G���G{��k1���<ˉޓ";�� \J�߬�=�7�Nx�����2H���<)���=^����ϖ������O�S\�fU�:��L	G�e���#���{���\a��8W&�g���L������U�e|]7|�8 �$����[ڲ���D(&Rw��t��FN��f����v�ʗ�}����M�6��.�?�.��1���'��^�O�$N�"\�v����(�dpCO�ԯ���6�{�L�X$��W=@
G6��oRw/W�~���`�y;2�>h�h&+��0�l���RWJ;�R��X��`�04p}O�? 0l��S��Dߔ]K��n�k�b�\,ŝ�m�N����w���6�"�0#�$ٖY��1D�
Ǚ�V�0�?2R��04�����S�O�>��.�n�FsT B��33���.W�t{�[N^]�d�RF�|��\�:n_�]i�L7�Z�ٶ�Sl�*�w��hvPʇ�<��|7��s�\�?d�0������{��@�{aYsp�ba��.b�tr�C�+��"��~C3ÞnK3L�eo�b��pd�1��l�2;���T�����CI��/E�_�	tsF��8+�j�e%�}��ƃ�>��M_Q�y%�Ǿ�l2U���Rw��*rpjӻ��4�b�B$LS� &\�՟����N���}����f�jr�%��-Y-�{�c�Ę֮+��L�XCTi~ګ��+��_��9va��W\��G�A1�l�
N*�2_N&�:��#���w�����/�_���]��*W�E�h5�K�`��:���j�m�����dc�s̗�0+c�[�����]��ʥ��B@��|��m5��bp��A�F�K������~[�� ��N�K�d*�Ae:��ڠ�Z��l*��}�v����R5Zs�\a��]�v�K2����|�³!1���L�!���F]-7e��0��1-;�./���I��׉�T ?��]틕�7,>�d��4������9����Hv/m�h�%.x8oct |Z�%/�H(�-Oށ��D�:֝����.ZW��
.Mo��=�n�M�,d$��nwb_X"|
��:��=�����X`BhQy8	m��.�D*l��ˠ6Uc��I����uQ�m��+��M�|]x��!�cj�/E������AHR��6��������ແA�(s�NŐ T�s��U�]����^�i��4����m'��w��OV���A#���K�f�'T`���m�!��1��5-�<CY狤���)���W毿%����R7h�ViH�Hd�������L)Ju�D{���R MI`g5]��\A7�?����o�s���v��<�~_�[<��qи���_Nr+��;w ��߶u	%����ѴTZ�_�p�n`�Y�-�N�ն�{���dz��н,�d͐V��D�O�4��R�eU_� �����1�b���U�Eۤ	�!9�% }�������a��o��]��i�i^Z������Ǆ�yK�����P	�g�Y"C�{9d��^�GG8E!E��]�|,��Θ�$���ܒ@(A�N��y��X����QX8l2�?Qӿ���%bܳ�_9xqK��$������q�~��,���VʃU:���vnޱ�2�����Ӎ�y�q�g�*$ӽG���.�${F"nsO�"�D�_��$.A�/\w8p��!�\��A��
�1T J��m��	i�zτ��_�jG�}ݗ�|���-��Y������w-�;�.�g
y��S����a��HE�4~���_x�Y:e,_�"�د�c����Yf�ļ�m��inY�|T�m�����"�S\�;.��uŮ���zy�g��$���n��%���ʱ�}�z�-9����� ���Vk�kܔ��Gr=�?�)��-�pP�e$�����R�O�%j��(|��ޣY�@E�F�Ry;�Z]5�5p1�y�-����j�4n�v�?o��[�Xf�t;>������]��=u(���!�] ��ޮf�"��?��ծH�2kI-6[(�t�urNӺ)D�����v9�b0vLU��X��N9�T�;�@/��5Ț��G�����f7���29˿BD�ՀГ��6����I��n�U8l�x�6��Ye�ƬَE��w�G���\�>�%I�ߕ|�����e���5
;�<�����^j�ﳒr�៙�pڼ��.?ZB\H��5�,�I���)�u�J��l��6���ɽfR���r�Zb�� ��2V�)�΢�ͤj�Z濦�V�|�Ii�����y�2H�am~9ГT��j����:*�FJ�n6�9���P��[���O����
����� �#]�H)H	�-͐*��1�9 54#���9t� ~x�����9`����}��*SO���gYcU�w�$ݗí����gՆF�$K�)�eO��=�ϳ�+4TNPF��e�;�h�v�<'��(̳��|���e/�H�yJ�=?�牄Ξ͊s����fp[��(�\}�gWXK�y.�+UC����u���P��q�=b�ߣϴfH-�>#kni/o��"�!��$��g�+C�])��E�*��չ�T�R�K�������|�������h���[���r���b^��;��H�3+�e�a5K	���M�]�����K�'l�Nl�E�L�6>����.���֐����ШǾ@�C��'g�;F��u�^�i��+��
T 
m�WQ��SR��v��lB�2�=ШoP{�]5�]s�V��V�FW&mz;�<�Jް�կk�wG�p�ˑ�������α1�^���� cĩ_g'���l|�!��/�k���I�{K��Zv0�[��|Ǿ�;�FYV�|�E�� �⮒��N/s�2�]��6r�173e�b�̭&%6��:�
~r��b{T����ݢP����y��52Oڭ"�ʆSz�t�R�V u�w�yS\���*����nT�C�B��Dς��ԃ�L�k�Ȋ*���0/�䱧��]��>��_-�������?�u��"䐤%h�r��L雷r��;s�$E�ݍI�)P���,u���������o��M�)	��*NÆ[�)�/ַv�r����]�[�/�$x߇�N����<���h�hS�Ǘ"���41�|R�7������&P�/�a�g�z����7��_VF:����j�ƥ�i/�W`�+�r9���?�����_l<� �dR���Y��ȕ�`�v=U��=��/��:�S����9��Qbrja�ݠ����<ǢX�e���Z{o�Jo%�G�I�ͯ�Ԥ�ά�x�j��b&ƻ���|�a�y�Q�5 �_N�S��>w��L?9� �K�;�$���h����pI���?C����:�QA��N�ǿ����]�y�7�M���O-ɜ�w�&d�
��%5�x	�+��.b_�ZC�.�u����ʕ��
���gG{ڗGY�=����g-t���'���������+Eͺ/7)��/�MHt���c;*�!��t�ˮ�zmO?�f�����13?q%��Q�X��`��,�rY\��)h�}2���F�}:Y�Rݥ�gg��g�ۨ#`Peτ(brD.S,����w���1��܏��ؤ��ہdM�NGk��l�P9�Խ���-�ja���Y7s��6��e��V�G�v�����x�Uc�nDc���;���+j�E�U+Ͻ^�ˍ��7����'���L�qX�.��|r��1@�e��o(~���	�ߓQq@�ʈ.�L�5�p�~��,�3o��´�.���T��ଭ�X(C�Ң��[�¯�.�ݴ�;j3U&	�q
H�|���ڧH������veЭ���"��
�_7��̲&_^
 eK��F�OW}H0�[����2ۦ�%���!}�A\u3Z���Lb���B��-�z7���Iu�WJR�	���ax�
q��z�8q�~7TO�)��3s�84�X�ҫ�8�\y-^c��˯*n���l5Hn�&Ȗ\;Q���G%kl-�tG�&,���1�1����ͼĘE �`�ڼ &�4��M��)����Pk&�E�󜃦��=p����rϼNh�����9���!#���dE����$����V����X��;��_�]Јx(�\_O~I֋�qZ�]�L��*���X�R�~l\�(R�H�B!�d�)Q/�����cJŮ��k��q�z*�fN�IM�*�Ӣ����8\�l�lbz���X�����0��?J��u�&����E��=�L6
�|Q��'$9A�:P<�,1���/���7!��OZ&�-�΂�`�Z����<��ɚC�|�`�=/v��M޵�JHc�Y%9�Y� ������3Y�1��!)�#�h9���
�{�*,H:g�A���u	���ZY�g`��Ok�\��c�>�N��g5�Ѳ �0�.��s[��rW���"]��W�3����e���X񙮺"��CrIL{8�>q���[�P����k�߿l���K��+D����]T]	�eSm��g��J�u���`�1��I8��,y���T&Up���I�	�hm�G�^��Wfĝ`�JIe%��ð��X�}RBC5�x�D���=ӻ��}��<P�Y^����p-�W�f���3�����jJnv  ��f��h{���y���מ����<n����,(;���G���ۥ�O��ݩqIw)�=�NY%��c;�؋L{���Ky���f�� �5El=�9dR�B�&�A5rŀ�3غ^�۽~@a�ݻ��`�"s������xԌ;*��~�4@�)�G4�`�{�nC��M����'�2��0 XX��i����/4��c*�ڳi:A�,��f�ޖ����:��=\���D�ގ�w�kN^�x=��qq�1(���W��ѓ�V�4���y�s0�e�W�a�S���Xx+�y0uK�uu��w%�v�wӉ�Q߈�l�2׃;�?��+�8St��-����|��GTf�_�.�B}}y8E�طEm�U=�D8��2k��|/%6�{N�FM,ڱ�<a?&�24w�ٴ�������&��|4���8<��掕���
8|����K�8�;�.������!_wMm�&��c]0(3�(��y{�Ҵ�PPJ�.���Ş�F&�ր��<\X�R���Lbd��L�C*��/��\?������k$���Y�VHϿ�4Y�o$u�F��a��Dr�z]�2���*$�6+�UU[���_�B��U��9Lo��D'���_n9���[1Ðg1�� ���W�{e.m�+�����W�J���4c����O*0� 4�y�=���!�Xz����9��'Q��#�Z]W�ʏ�|�% (�Z=O�&f5k�����vO�_v�tZi(x뤫�_i�����9E=W��r8$���\ďg�ب�u�h���8��\�bS;��������&z_�����������l����ԯ�L�v�L?
�FUu]v�P���͒S�Q���(ǿQ!K�<�����g:|�ܓ(��F������ &��}꾘�	YD������X1�����p?�R��y�9��&�����'P����A����lۯܡZĚ$6%H�ƾ�<�nrn�Wӯ��la/�u��ݜQӄ����6��3ҎG֜�n��mԟ������ݣv+e�BvV��!��6�ė&)о��D'�S��AŌ��(�V�b�U�1P�(~p(IG:]�Qc��v����Y9���b���?�
e�﹯�
��	X#IQH����nVpx3��L�ԉ㺊��w���$�Z|* ���򭥒+4��d���I�ؙ�ȥ��M�Ji M�r����.��Gk=�q�ȕ�MN@�5��Tu~�I�+�e�SK�"���)6�*�P��Y���3�;J_�/$ A���j�H
s��Re���eV��F��F8A�q���yغ��ȵ,�#ŉ&Z���V�������h3�4��R'�v�Ϥ1zVޅ�0A����~�<$Ic�y�[���f�@��x6�8�|n�#�(�$`�f����\t��w�{/,�(���mE��bUXL�:W 򸴻J�+Sg�YH9Ʋdw�N���]M}������2L0E�^�;�
Y};�}�`d��Fl0�9K�x��,��L�gz�m,���nJb�F��]��)��{�B&��7
��+��k��.�x_��,���$^�5����@�����_m���/�t�)�?�U��iہ��U�L����$%�����
0)�
匹�=�؉��țٗ�su�)�˥ֹP���?*G���[���fzaԄ�4�BN���q��cp����=���|��%�e�Y(��"��M���s�ˊ�&.�#\�}ܻ � (�6�-z��;$2��������i�%���'�Y����|��f����n7��v3�����Vx��e��3��pӵ��_0��3,|��}?lg�z�>n�5��~z(~�����N�Z�q)��\r�\?vim��a�lN��E�H��Vn�܄;��:s���Y�֗{b?�\��z�q��<,KĭC�-��p�9{i�f�%y�<��ǡ;��]q.�1�[�M�q8\+-��7�p����ܴ�z�����(�`{�*,gx�
b}��|H�^�s�h�����I�z4<�}��f�8�ޞu���_6�Z8 ~�/DWY�W�[�Z/�ʥOJv�w���,$R|�K� �C����fe%EK^ָ%��؊5F�b �����qA�cARIH��eR >���-V�樏������</c�����u>��J
�>�v[C�_c�y��m�����L���Lo�;96�U�ҝ�@
���ϵ�!�hy�ÑϹv��gK>�>ы���vi3�*fX�m�Ng�А���xmj'�z�t�?_�ΞQt��7�w�������m=C^7��o�M:�@h!��^�བ�L-7�'��J딫����~K�
��*3�F%!Jٟ+<b_�$�ₐ�C��N n�i�����If��{���|��8T�&` ��k���M��er�U�;T���$��v��U-���c�Ǌ`��Y��|�ǦС��{��x�?���,��Q�MP��2�'?-�܏S�7nڶӨy����N�u�quoxe���XF;��!��������3,���W٢pܩT�tj9�E����gc(����QX-Fe��dm#D�#pҦC��,��>�l{EN=ն�P�ym۟�/�I\��Zzd�è�:Pw�U�{�ST*O����B@s��)�%+��CG��hy?~Y�-�K�v��~P��S�yϻ� ��y����M���y����빅�G���o^h��J�^ fn>�҈wh�.�}k�2����rQ�w9Cd.�=��e
i��#:�Τ���Y�'�Ӟ��>~2=սt��y�l�QWt��R@p��#��=_5�_O�F����^]�p�S��t�d�]���D������]��g���K�˝v���7�zx����X�w�.���U�L?)%�\|L����l�Y(�79��ž�սSq貄��6�F N���c��&��h&UD��r�s���W��6���ݾ�%�Л"�o���(�(�}�e=,U|r����b<�Q7 _�u���>l���B�	�;j3l�|"��@I��������l8r��<���_��E.����H����E�57u	<䀃.xe�*8IaG��G��߹�IR�u7�E��Nq�K��m�d(����P�b���滋�U -�9})�Ϯw��+w���z-��zQv���"0�U�]����*O�/���������9�Bb�^�h29���6׀^3&cD�tZ��?����NA.�%j=��&8�f�՞��̀8Fx8��n�$����o��{c��<e$Io���\+��-R_F��7���R��R��Ey�mR,��2�:]a�9^D��<T	~"��ƻ�Q���Vύ6��1������ڊ�S��z��e�]�N�D�usS�{�mz~����fҗ�-Q�d��7�-��&8�^��wB����$gI��5�[֧�&7��K��RnΑ�G���#�y���Ɂ8��D����Y�/z*���5� ����
�x�7�r��L���Z��r��"vXj�NЙ�Ij�*�'V0p�=7B��:������k�wg�����x�M=?�{���굆��H,Q��E/�F�W���@��N�SvjLGߥiʶ9���8���Z��(���c7��T�zU��gk�u�</�O�����&�(�k4���:i�IR��MM��xy����q#Jk�:����ɟRr㹁��*<Wb�b��@���M�j*��*~q���}�}��se�dY5��k銍<Q�םwr4���}��(�,��@ܓ�=�K�H9-`Ok��@T_������IUۦ�%����N�e��(���{��~{�_x b����p��f�P���F W�%��	�q�U' �UI/'��}�Y�ѓ�&���&qB�ii�����0`2
��% YDocc"ܭ���h�c=��6���#���å��4������W�Y�K����1"R� �M��֐��<���s��	.��?؟�:?4�����o�p%69�^yo3�4i���,�����s�m���e�Z�#<5Lv���^/�M����8TF�(��0�!�5WM�����aױ�D��D�׹���`�"4u���>:�v����oI=/�X'�J�D�h��]*�Ρ����g�	c�f�8����-�_�����G�o�-I_s(im`��y\��U�ə^q,�'�p�|{�n>�"
�(8~4��m��<�yd�sp�r��(�6A�ueb��!����U����Ў~��'	�!�T���a%3�����0a^u9��$ҥ�B�ܟ=� Mv�ȷR;�S?�� �JFC*N��6�B����:�-��9�#�	�X���5�()ť$McA��&�Z�b��|�K@��3{1}_^n�s�;��S8�$�/�ܙ��K����!i�>���1ڢ��Bt����&���x
hR �zˉ�����~_]�c�򽾠�ڼكݔ�]���G��4S���vs�����H�-3o��(5�H�c(*�'����8+�^x� ��O��~7�U��:�����n2�:�d��^��GM�=��>��3|g��_ܺ�bp����[s=�Xdr�t��zOZ�P֬�:�R֋����Q,����uW���������Q���#�]���h�T"���Q�_Yb����:��J�p{fQa��@�.����0�����@Y#��n���������y�N����o���kgM{����c]/Z=I�ydO4�R����/5��q 6�L�b���4r��A���t�J�Z]��3����o��f��v�����  �>U�ʆT��� ?�</����|��}s��2'G#_��x���|�ݚ�gd?�^��#Th�2��W[2�d���1��f�c�]hb^?��[M�� �����v��}��E'O�������ǩ'Iu������.�0/�6EL�팝��7���.7(dzY+��.�O����-טzrif*�o�ҍ�C��P��O@��}0��;Eй�w�.e�>���͵�1����>�7�:���ӗ?n?������9����.��D���c��,<���^����X�
J�˿��J�4c�Iг�+�$h,V����/+F#��5�j�%T/r^K���â��@��r���B��t1 4�,0dw��$�.VGؽW"�ksQ#���j���~��sn�_�Nd�4�f~$��r? ��O�m�#����=�b$�W��5<wٮc�I���Vq�R|� GƯ&5�X�X�;B�L�Š�w;W���P���G����0If���� =��n�D<�d����G�/����տ�:!�� 83�M�olx<w�֯�2Հ���y��=rt@��y�_�^u�H��Jm����a����زCR�Jț��z����J���~�ez��ΆH�k(���X�4P�;�/��:�͓	�*�;����Y�(Te��K}���Қ8
�@�8����ea�[`Re9$�D-�VLr�����+Z���Ѝ�?�Q/�b�%w��0�,�^mg.�J'g�O�0�a����e���ة��ϭ)pF��S�&&���T�Σ��sY3��1g��J��g���?Eu��B��3_���3�j�؅��54ׂ�P�t:���.n���E��t�6�;�c��G*��װ/��Yc �87���CM��Y"���}���Mu���<Sf΂��o�0Q�l�*��Ֆ��d�������%�ۀ�!���j\�=1�䗋��U��[�`�IfM��VVD�⡰xv"�v�8��zi���^�!mB��mtqj��W��r����/����%ޕAxZ���f:�p"���Xz�M8��Ld�xz2�:ņ�v��
"|{�3��q��|����(��d���2Q��Dh޸5ڿ�	=04�,�Rj��/�s�Y+MU3z����~=z�$���Ȑ|�<Q�j06%A���U�b�Nm�lS�t�(ea�����)2k�$�A�HM�ͫ�1�{�$��A�����t���� �0{��9�h^����e\��SG[;��9�2Z[��X}�"�,6���>9�Ͷ9<Ј�m��bYL���*��C+��;�>{�;�L�nikC[�+_K����M����U w��1��gQ@�`J�����:�����z�dMW��G.vq���,��COaX+�Gg���vt��b'R��rd? �ܺ�����S�w�s.�T�Ki�~�,���\g𖥲"Λ���	�'�Yֺpi����iBR˽
���
ə�c���_W�d3��&Hxy���"]�2R�@�G�4K��*���mM7����p�S���H��a�Q�����wh��kB���B;�]^E����Jc,�8Cy����PVi��F��?��O���jm˯XAd���{t}� ��E��{��m�u�/ ��K\6�uo}K��3(^m�FF��~&��@�K#g}G����F����;kQN�V�k�0F>�2����2M�x������q��g����?��R���fV<"�X`R�C�%��x�x�XQ�xN�c��hu�6�Z���}=	��6�צ��+��)��G��ɇ4(t��A�,�Q�q�8���Ԏ�6����g�7޴�NG�ƞx��������ăQ{$�L�y(�S�;Nc�r�e�+��ix��[:Ys����Q@��%�{b��DWeʴs�G����-�ϙ�͹MX)� ���x|=w��ʴ��'��;�q�B�9��v6�������I��1Z�������&��܀�Q�
��VS�H9�#�:8�*���H&ګxdRP��`�ĆJ���ܹuevE`MH^p����a�����ɇT�~J��c��6�4v��Z�"��d�n�[���E�<�3� �=7�zr��䵏IH�� K}��R����R� U!L'6i��'e�ʬ_Ub��HdbY�����[ϸ���J}_��vw4��r�@��^L��!L�]bV�y��;�[f�5�_C��OX)\�%K�Tg5��Ʃ5؀;�j�/;����Ǉ��\�5���l$��\��(�mY�}q��@���yf��k�9����Ԯ�[q�/H��g�	p�@;}o���I�'}��)1��>_�Uڄ)�$�W*�^)<�^��J�P�$d%'�������(Pȇ1��K��"�P�p�R�	P4	t��n��nT��O'f �H4��B��SF�z��G��Gm��T��Bd��pt�N'�C�8m��0� �;���zG�'��cJ��J���N'��H�`��S�\VX�o�C4�6E+��L�
?,7KdֆV�N�v^�b~	��'�iق�<�E4��~�%dVN�qx�[�b�i�[�Z�zY�n��[�X��#`��׭����-��p��O!��n/Q�_�P��u��&��(�;r�_��w�U-_V��f�n���X�^�8#���ݪ$�l�*�l�=�;S�U��C�SUWM+���)�z�L��_�cAK�ba�ڋ �^�	?��87}��h���w��f��G�"�:e{��zY=��un���kv����	�����9ˬ���؂��2����>!��A'�Ͱ���gѳ僻�Ľ��{ͤ|�[�Ξ P#M�$��{,?�af�G�F��:��+��3)p���,c�R�B��>&r\�)ׁK�J`)��7���]l��Q����h7��Ua��r�O���:-�Hn����:��e'�R�PH_: dP�QI%LU-�vTQQ���SCl�I��H
���(ۋB�;��=�2��v\:]�o�������^��Q��hX��@]/�S��ryl������8�>Q?� _��@����!c�ӳ���A	�������S�2߻��w�����>p��S���,T����p~��6y�;Tx�ԇ�[���c"��Ù[�w�PU0��N�(/½x���Hz��:io��$����&|���M`�|ec]Z�I��5�����L�ǚ�Wy`<LQ"�_8h%=ݪ��%�X�и�hsS�ƻϖd�F� 9U-�3xh�no>_�y�%� ͬ���(L�r���VH�L�����)���{5�.`�7xè��j���H��[>��~��n��u��D:��O9~ct#���yU��V;/�~�~�b����$õHi�;�&�	�H^9�n�v���Ean"�k7Dn�[�+���ơ#J?�鶥9{V t$�&�r���{�?_}��1��1�J�t?5�m�s<�ɍ� ��_�u?O��&�/�8f��9�O�P�G�|������[w-�>�M*S��D��T�7'������%'X͚��2�F/z��w~����m�|a�n���?�����>���,Dk�uJ5�qO*�gz߹�ѹ��W��#��ɇi,k�:��[D�Kj<�)OLEx�"�㤤F4��Bc��1�0[Q5��4L��e�^7���_����?mg�REbER>�w�bDz�Ė[�Wr�Z��C�$���>��J�+���٬?�oIq^��v:%�7?(#��lh���|PU�2,m�����c��T��G����Ѣ�C�akD�Y�p��ܾ��8af�hH&� �7c�u��$�޾��迗��z�j!�!��^�`����:�и�tC$�mY�d��CqT5�$�u1�_d%Y n�䝎IdN���&�ex�M߱�rk~��A�lŜ~Ts��&�GgFd=I�&E�'HBg�����(r�-�[���K̔�=���65��JR��;�k5yAϝ�=]�A$�f�X��rk�z`ͼ�R�I�ME�)~�l�<�I��d�.�LV��#3_D���Jy�&V�[�m|� �y�����C�����"F���C��;�N+u�Z��Q�H�ᄷ18
� =���hk�  �3X�^���f-LǷ��L��p�E+���H��l�p9>ǡ7|՛P�ȁ���ਢ�:���}
���o��WW4�.Jp���ߕe�i���xO�8	*�n�./k��jH�1lt�������D�CG%��Bn�C�ꅉ����/�=f:�<$]��Q�2;.�|.��] �i���z�de{A���X��4�E�}������y�T/H��p�P�I���4/��q�Iݭq�%m$T�GT��^)s��{�:����L���#Y�0��Y>�(�ON�<�ۺWU�ĥק	��90m+�]̚�}-}�=��������!����O:�V��k�鄼�&Ȍ�o!��Kl�4IF�0�,��y�+�ZȖ��Y]U�������!����o�.��g������.=��b�%-R�B����n����͡���*A �� ��@��Ѥ+\Ƕ��+q��M�RB�0Rl�W������n` ���'�?��mݪ�@�+m���i���P�bf������TQn�ͯ0��֯w����*Q�,h����_�}`|�ۼ�7�H��i�	���Q��wj��F&����g?g���2��]~�.�p����z8��y{Y�VEH���H�P�����s�Ǘ-��w�Ӭ���vV���`��d� ��.�Eby��n8jeZ�~JX�M�	��UU��QQ���N�i��C��!����*hWA����$S��ʲ���G�BJ:P#c�Xaj��[%2Ux\�Aɝ��l)8���bO�
4�� �DY/4O����=��I*���F��f�+�����Ī�#м�θ���]���*}���[+t�R^
��Q�(�a��b��o{ �璽��J�	��57��	�2݀�$M� �:��[=u%�����Ý!�����(j��9�6��X�R�/�D#CDǗOr�),Q�WnN����*|\�zK����qlڡ�Oş2d�S<]������B_��'��	�AM��?�� ,J�w�0�p�B�{3����|�jt��B-WG1�s��ys����K>!�!+ݒ�' QQ,���Z^�:�c*A5�g�����s�k;d��Þ��n�?9�����.L��2��ܱ!2�l��ǹ5�ҚX��.�S:fD���1`੮<����
EZ�_-�hF�j��Z�z���yO,�M�o�4�d@/<@��-:�磬��W�MA_�SӚ��מB��Gb��<���<���3��սj��r熫��L�d�y���ɬe2T=�W웲���ސO=F�����m�(u1?�i�U��:����	h{�YN�.R�lS�K�^��9�{[4�?�qHѦʔ��2�LYl��l2#���u��~�]��|����m;}�nyߘ��0��OQ�Gq׃{C�dmN��;HGW�]g�w������|�9��=5te��[�Ht66R�O⓶4��/��D�ۤM�����Q�5~�V��4 1�'t����57�R���_�fo*H�<��Kf2����h_ȇ�h@j��$	��j�*�r0�f��z�Ki��2��:ʍy��7��!j��nT�KpP�[��N)����tV4!�-+��l ?�e�M�Xl�;�ܣQ��K�f��#9��?��I�q���F[��7FB*���h��w�h�l|�gO5[��c9������WQ������n�?�iD!����u��'v��A�v�G܊�����S*ߎ�WիU@=�;*�)JJZ���'sς�"�z4'��G��:�^xz��7��D�n� "��t	/�!Q8SBCf���D�o�L<΁�m���=�\��.}5�\l{��n��J�Ʊ����ľ�㇍L@!V�S�:���bI���Lfx2M��)�"B�#�@i��# ���i"��PO�3 �0^0~���u���&��"����'��[���mu��?�x�u.�z�m�vE�N�K�_�<ƵL�uj+�Q~��#(��"������#?��p�8_�[^L挆�{HJ���J�p5��d�hri�{ͯ'���~�Z����S����4T�P*S�AIJ���?�;�,����4=fvԮ3�.�LS�����{�"�1Y,{�&m�M��N�j��1o~���U�Ӎw�k�Uag���l�0S ���)8�Q���o�>��!��v��UvZ��$��{�U���u{��{c�;�	�oά˫*��v�UU/�9�qP$͋HpZ*f���/��W�|�F?;��ZM��z������*]�K��Ft��5�U:'Hc{m~��O���T��e�^�}��c�2/�������֌�He�o��
k&�A�]yʔ��R4����Bd�:��Nm�U:O_ҙ`��E��7lE&�>�}�"�(�V �g璆��m����5g<�2
���>/]�B "���aE�#%xqq��>�U�t��(�92:7>�;3ه�`�)i��ﰬ'�T��^ż0쯯�Yw�d�U�r\�M����g���aqKdb{3ܪ�31��Zk���	��O�o������@Ҷ����æ��҃��T�m����#���?��c�Ne�������C9�:|09fG9�Cx��Ή�d�bL��x��ɘ��h��劒�������RN\Ö���M�5�B��ek�����f�E���h��ƻ���=T���&pQ�O���^��E`�ڒ�Dhb�6���;!�L��]㩟�;�:c�n�H�����rc-z�O����R5��X����d)�E���UY��!MT�~���~�����
�O�	62���%��T�[!���t�c�$�21�w-^nl�=�]-�y�`� 	ȩ�%��8L��s�����������q^9\�(�<l�]VH��ĝbc�7�����V�Z0ϙZf"�s����&�����������5���D"r�����@�˯�FO�Q;�%� ��|����\n�����`�{~�h�y�_	C-ĺ�D��掠�>���.�Q���3��4����!/��]N9ɡMB�]�����M��N����e���پfQty����� �]j@pk��k�ջj���%��)�m��{I�����	v��U���S%�޸��`�?��_��
�4ˉ5�	)���t.R�U��\l��zp�0��d�o7,������ ��[�u���/ ���u�-���X��o'w���^db������OЬg�G®L/�D��T��N���J�,-��4m��}�pYȭX+A�$pb��[S�t)i��]�UV�^?D�"�\��]}��*��ChV�Rh�M��eo����_��Omڐ��ꅈ�B%����:�<[oߝ�?GF(��X�U��9\���M�%.�.=$�3�����4Z�j�H^���}z��>i�����sJ7.
}\�gJTi&��V�
4�ڑ}�P��G'D�9��f���7#c����|�3a����0J�I����A����esO�"��H��g�Õ�<��OV�0>�3��5�����#țҚ}��(;�3^B[�Vsb`Io%a�Y`�.|��X�4��j,��5�h4t3<t��ݲJ�2��
._4��i6�ȴ"�?<oJ�|%��p��s�hzl8Hտ�9��o%��aRC/�'*�a��L{�I�~������8��o+����4��D��b�3��2�[����N_�̣�('����#kO��w$�Qi}���Pt�@�6
8�EN@��ۮ�2D��n�����2�EH��V�f�r��՛�D0O��1�5��0�W�1�ڌ﷨|Q��y���^����R[�L�o����t���a�=fVP}@CT��Q����}���n��h��y��$�	�b�Z�ٸ�p���k��3�j�=�%$�2�^�~�_�r��۝��8����i��A08���k'��M,c�����R�G�`�~�b����Źq��~,nO�?���)s�;Y���*�L=k�K��s0�bD:�d���g�-^|x拤?��)k�s�<3X[V�^��Z?[eչ+��fo#�pE���eb=���im�,j ����*�o��r�i���E-��>Sߘϼ��SZ�ƪd��9aVg�Mc��М�\�h��GvWg��.x���O��螚ޟFJ>r��4��o���'�۰}��r���!�͋p[�#�t��KIS+��=��8&�ٲa��ϻ)Bx��u&m�d�\�/u��=;!>��Ρ��iO�_��a	PW����9��G��/��/6���������~�9lM��B#�&o5�b�ϻ���j�,ɍ
`y�kub���f-g�x�JX��=6�7"�Ԋ�yk�/4��H�8��^t�ׂ?H�5������G��<�d���f-'������1�$7	�l��P�/ĎxܟRM���A_*�5��.'��Gջu����t���8a�	����q�C��4�x�"m�;�i���u39	�=S��2L*ʷ�E��j�WB�̱Ӌ�"�PI��o4����wG�IsqG��?Ma;����u�8~x�+�Q���*�/S�Ž���`�CcOʦ�ʍ����`Y	�Sm��ۘ�۟޺���WD:���1vJ�)�E�^ ݶ$�	w�������������j��ɟp���� �Q�v�Q�J؂8;����2#�
�s3�G"2Ű�`|x���F��kx9xe�����ޛ����#��r�{�K�Q9�}_D��Q�`Y<A��J��"�+Ê�;3���ts7�.gT�'�Ҏ�q>-����fW���䕻��ѷ����Rۅ��t����n7_r�~��>p~�>"�'^�rO��{���oB`�:*+�9v8�m�e�k0�gk�0�t
F��J�����!�v;�<ԩ��(e�؎���z5z�y��Hߤ���멩%�����	y==�N��e�a���c���31�0Ƴ]խT�A~d�f���KR\W�[�����-��lӂ��_^'aa `�-	��X�oW��ah2�R���`9������E���������We�_�O�^���M�x蝹���\SB�a��ހ���O���Gϣ�W���g	�������Y�N�W&@ϹZo'@�����s������#lr�|��fpB�� 0FZ�q�p���V��`d�'KX TI� �ztu]E�"�_D��է�|�[J#��!����<�c�f�=�W5<z}T�fK�j>��C"L�7^Ōʫ@�k�gN5����`�y�V�(�B+���
Ԍ���uT
�>�o�j��0�z`"�9>�OP��9��d��8�?&��!����(�HI�t��t���tJww��%� ݃tww73�0����~z�_��Y߷�����@g.0��z����@L^i��r1�p5�,�F�a(�[:
�E��U�´P�Ie3h����Ͷt��8yKbS34�w[7������S���R�j6�ay�^[�����ۄ�:��2J?(�$b��������t����em�й����8sm/l��Kf�l�\[�1���0x+��������.ئN�+�b����jO#"3�$���e��[}gU�4@Wi��Cx��)R#�W�
h?��I8E��xJH��Ă�X>�;������!3��?bX,w�Z�.-y���������!�[LW������i8�A�	��C���;-��B�n�#���X��&]�f��|�*G����9�Qi`!C���C��|���ROϕ�L��c_�7�?�>��}�PR�{,g���z�}^�F��X��x­�qn��^.5��)��ӽ�Ī
��$��eI4.�[E��a�	�rA���
{�D6��E�p���������.�iH������ޗ{ |��s�C�b��P�v�9 M錅w�3��;�x�T�ti�r�\tj�*����j	�����h/(G�D,�Gi����R�v`�XrZ�Z��˚˃�z�\�{-��-v����$����>�֞/a���C�M��/���ærl�8n�}�08oM^b�ꝥ�ּ'�#���d�R�'���}%���؏%`To��LƋ/�w�Q��&��4󶣯v��0����ks��Y�o�&��*~��,h���� ����$��lg�*�)�{RD��mU�S���r�ޛ,a�R����??�w�Z��)�GPy���$��-3��lV���X���w?�%M�bi�7�Sl|/�-��X�����	��K�2�B�,�꺆���vzl�p)`	mD�r��nG�L,r�?��g�y�Q_��N���R\w�EVP@�Wm��"� ��Xߦ�)��Qg��/�o.*|�z����6��g�'^�\��_��8G��\n���O	A��Y�E�ȯb���l0��R޻��R*4��22|t�s��Aq{�&1/L$r�:i��g����L��]�j�cYjU1�A�0��7L�(���!K�s�l&��f�sY�t(\'g�M�B4�_�"�6]Up7»��&��\�s��e�lK3����S�N*�R)m��Q����ǧ���B߫�ʵH5��������ܾK=DJ
�O��`b��͌:}Q<��zm ������ߴ���`z����ۏ���8�:y�'�H���N5��G�'{9�Tg@亀��3��R�����hD�37/]��N��MM�/����S�.��*��X/t�#~ɣ���3����y����0oEO�[fx=�C	�ޓ/����"g9��M)���7)G��*���>,���"`8������<ym��I�������e=�����eF0v�ҙѻ��wt�Z]�Q��=$#v��s����`\�r��ۿ"LOz��s;;�ޭ٬_.�� �HW�E4�zE k��m1��4��!8U���7����J�����Ao煗;
�nv'�<�tJՕ�$�0C�ԃ�;��^y��w��Xi[�2]�!ю�/ƭɍ7�C��x����̸��B)0����z%}h�:T!z�m�L�ƒ��g�/�����u� %_��0�K���[Gыw�4:���0WN����G����h�j��k:��7Mn������ee=���ֵ򪭟��v:]�{P�P�Y�gi(�w���v-Ckr�3h�{���}��^w�n�9�����SRTY/��/rCq�J�mE��Q"?;Q<L�d���$��GzUۛq�r�Jۤw,��K{ד3sF�G!��x�E��øuu�B����gvo�u�f�"���Ӳ
п�>{vETt��*"%�դ�;��0��M���t�a�D�<�_�Sr��zGoڃ��ЋF9���Ani�����q5�,qQ��m���igV�h׭��[�/6O߇��.G-� �=�8c�;i�U"B{���R�1mq�r1wнIp<��8��z��̇MhD�$�E{��M�T=�$n�r�K}����mI2u�DM��;��n�����ĉ��1�BY0�\{Ǉ�:���^7'���hG۷��3��~۰�X����M�(���<_�d�ό��V�ilK�W��	�a�z�<ob;�_䂟P#H�s�`��m��j�u�v]�K:R�qj�E}�.�D��U>b�QG�&�xI��4�c���Z���|!�Ȭm�ٳ��$�lA3.�̎��ig]�3kGܾ2F`vO�Bi�Ϸ�K�H�墡e���i��I<���'^���O�.sr�sJ�"�#s;��g�%3��g���5~�8x�@7ý���3�Ł��=mi�T���i��7����V��OT�A�fږ�L�������K�D��䎩�e�$��Gp�AtcT}�(���c�Ÿ���җ�ѯ��ufSh�&=�Y�aOx.q:ɘ�.�m�˿��v]("�Hs�Kh��&���q��[��ۇm|h�t[�pn9j/V8�7U7�>~螵8����������I�y���WX�L����7�3�k��g��B�>_��)��YU���W���W.�y��4낼.��l����
�����vQH����<,ꌿˉ����Y�y������"��w�e��ٶ�x<����F�_M �јh�g����xKN����^J�ӥ��u"=�\�[ �8B�þU�[+|������x����:�b!����d�Lo)r���N��*	�km��B�G,��sU$�쒐~��]IB��[72}�E��Hp�}��+�c`agpv��H姭�0�a���Q��������-��ӧ�Z��%�M~�.���������؄W�.���m_;+�/keWV�Z1_��y}c������	�c߳=�Pv����-���l/Hβn�o9)<yRB��M̧?�@,��������x���R�4���==�4�=���ys,�����Ĭ���1�A���k,��wr�(G4͟jjۛ�J.>��jX�On��o 	ew)�2�l�����(] H*H1tk�}�*����.�2Z6�ğ74� f���������ط�w���3Uo�!lS�8r��	�T5��w������w��lI����k)Q����KB�3�0����U�º`��q�z>E�夷o=��@���F�9k�Ϣ��]X65���J�~�$�-�3~n4����b����XY>���֩�O��@����d�6=s�;Y�8ߓ�q��|%�	��H~��C#WȮ"'̆ZY��1�x}��,�I�=b�P��^Y��$z�O
��ү1냪�et�����fD��������P5����<�S�~���V����0�}N�S���~�$�_UQ�P�MXl�0��&?/D��7���'�E��L��jyQw�~��]�޳�&<8����r�fG�<�P�9ц9�GgOj�}&����L�8����V�%�Dg�%��/��̹!7��H	��+W'j�9��吠�RO�省/�o/C��_��9����v���9:���\��[��l�nx���f�Km�Ұ��θ�J�윽�Zps6���~�0�z/.mX���B-��P��K8��w�����J����{�@"�e��k�D���'±��۵�V�<c?�W���t����-?��|a/'f0�)��>�F3SxAf'����4zzC#�U~�r���������&��[��d��\bnU��:�N�0y�Z'ᘓ�?�M��|�|�a��È7ݧɞi*:����>odE0������y:�~��L=a��<�a��4 eC(;:O�k-
�_��L?�Z��[X���W���j1��ʝ�|�]͡Q��h�
�߂p���` ������/�J��!��C��u�������9&����kJ�>�s��X��:��+��T�-�3W�&�0���7ǥ�K-`��7���R�y�����|j����f�V݁��'���;]��͐����
w�� �#��������GWh�m"�u$xŜ �<(��>ҎGM���\����]#*�vQ>���J%ƌ�r�Q��d�^	U��� ����H�un�{�^�$��yE���gE�o�m�7A~^˶ߵ"�;����ON���%M��_��\=T	=�R(�i��x�����N���f���,����IX}�@�s���y�"�͑��X���vS�h�q�}}�ɼi2�}$�#��y7� �}8���������6��5�o6����+b�RF%�7�GE�uَ̅�?b=�:8Ē4B)`�[`�z�������-�3[(�*V��z���b�������ͦr#�!<�����L�<�`�K_���f�V7̙۬Gg��/s�o2��TȲ��-P���_�&^u����=��P�!��Q��D���Ʃ��K�N7��0N`���k���E���숉����Pr���w����.5����Ұ2�:�#��ʳ_d0�1-�����ph�S,^�ԉ�s�M���"R]B���3t�e��<��V�Z��U���R�cmj�Y=~<5b��B�xl81�N	��G	8d[>}N�ݮ;���6f?ա\.e�~��&N6�&v���54��%�j���,{_ɿE8�b_q>�pb�8Bh�k�j������u��F�d����P��������/K嚱aJq��3]�m��݆�=�bu�6oyn~I�Yt�J1g��pr#͏�)]b�3w��Q��X����0C,�^H3�gN.��ؓ�6s@��J�h�<��OO�=
��)�v��B֏���ּ������X��-��z��}͓p\(�g]E�;��$��L�u�|3��P��穲�SR���i��C�K $�׼�3��h���u$�E�s1�{�����q��0�dF�Z���1��Ѝ��5�Cǻᦒ�ض��ű�/�-!^���M�S4Ţ	I�H|�ƛ5{O��C5W��yg6R!M���]k�%B�N����)z/{����C�w��)�*m�Yc��w�g��hv�io�����A��g1�����$�o��
�5��=��-��Z��!�|���7}������-µ��M,����lG�n2�r�.����S)GxW����g8�B�Au�:w&N*C�=j�3�Ju�;�uZTx���4��%���t�M��4}��xÞ�ܷ�( ��M �����%�ݖ�~Y���|�+�)�ꓫ7�Q��G�a�Iy��5�����5���}+eR�x3��Y>R�D�p?�M-�^��YNUO���z6�%+��''#6�[�WW>�4�4Y�,Y�e�)sYC��3�ظ�K��i��X/�Ev�f��c@�P�������O�{Ϸ���'�Y�4����qsd~N6Oܘ�|ˣ]@�{U���\����e�]*��745�?���K��n�.�ѡ�|"��������rH�I
��?�z���	��O�Tv��Kx��hO���0���nI�,�Sj~���m��bd�'{�sx��i����5���0�9e�3d��L�%,�>ug�Ӥ��β	�<��@h����^���$<d�{!H﫭Vq�����ل��Ek���}N�"/#����{�Λ��P�7�F�X��_��&�QV2�������'�z�܃x/=�{�#�7d��x�gaΉ��7+j�C4љ��|��~[�u�a����F	#9~�4���ul�{Yguf���#l3q�X�x����K؋�5��id����#/u�H(⟯�V��7RW�$q>m��
|��`�E�c5�W����ջ�6�}��`�����z�W�=>k�1���p.H�R��y>3�IO�VՋ#!�s0=ش�j�}Ӻϖ���r[��&�z���[�Z�+���k���v2��왳o�l�� \Wi{��i�y��D\7�:G���'��d�:Ud�|"�	���SQ�ýoӬطx5�%aZ�M��q�I*c�?��!�e}ڹnHӱ��n�פ Hp�N����v;Z�]+2����Q�Z� Ȟ*�x)��`λ���)j,�q�hj���Id%q�-���_5��\�'���^�(Sԕ�?��^Z�m�Zq��_A=8Z3�J�����kH���[ʥ�~�yF�j�o	"���N1����r}F��;��-S�Q��d^>yu3�	io��[x���9h��������r1�s�z��eMOO���Y�VI�aj�b�!�6�jkJ��@��'0y��H��3zZz�|2pM������$}�k��~OPh�u9K��J!���˘�ߦ�B?~\�b l�YEJ�N���|xo�W����"\����82U�[�[*2�Q�΃^�F5A�Y�U䠵�"��~_g���������S����Kt^�ٗ�N��d�w�#?+����@}�����8:4�h�ѕ �������o"H�$�h����.,��5;���,֒�q#�����>��E�멑}�$��������gg�_���ࢄo9��ަIsp�\��]�[��UT�qx�KAb*
�8>F| ���:�4�l�J�}Y�TgB|��8j�����Zu~�r:��s-0۾\K��������ۜ�㫫m.N�C�!�Z$�����~�}*�{j�෍��|ͳ��V��9;l� *GMW�y��=H"_UC50�tl%nK���{0{�^��sOƼʥet�nɕLr4p�?�: �c5��+�Aۜ d��*˓vh��VNI.n`�jae�����5�Xc��.�nO�c�">D�G=���e�\�i�>����������a�\�g��Gk��Ⱄ�}EA*��p[Q�=]u#�.j˧+���5�2�\�@F�F��՜M{���v��"_;�K���$���n�N ˎUQ��!�l����Se�����D�����P� �!����ye/n��S诣��7cK�a���#c�- I�_��{�ر�cnf���VCI�]��F����K������tB�;��[�/=�H��VW.��ܫR_�yxu� �V[�]X���5��_�>��'�MU�??G�nd�-����~�8d{R�_�����S1���:cph	�W�G2���Ԭ��A��g;Tѫz|��l����Ys�I�O��|������?"+�j�}����-\�5����{�����s�n���A�%��VT���-J;��F�A|;Q�,x�X��|7%�8h����^[G�LZΞ�p�EZ��Ȉ�<�H &)9z/�{����f� �#+�'%ʃ}l3����}�JK ������(-�tOi}哏�Q��+�ő9�@>ވ)Uś9�ĿW���`�����<� `�Xgi��x��?Wn6�X��3&�}zN�+xr	��^�׵(�sσ{\t鉳ʞV��hkz;�)��d�.-&��:�N|�*�>�K�=B2��lj���N�uTֶ֙@�+���|﷢�c�O&����Ȼt�F㑑����SZ��/tVY�~8_�BSj��Ν�5�w�L��J�G�;�u۴<��3���:ϳ��֮x�z����>�OzQ��=U�����1�����F[�N���{�?	�|ׅ�J�"��(cϚ�I�&?���xᡠ[ue�x��������$��:���C���b+s`��R8T��u���"�*��n��@�T�ˀ�+mgֶ?�xp̥�j"3Ŗ��+��w�b�ˍ>�Kce�V��,&�f���C�l)lx�V٫���l'!7B�����5��	Y�F��"b��K}/"&0�|b�`:�KVj��"(��J�]��k[��D(�R�$���'����I+�P��߳��Y���`�M�P/�l��H�2����y��)�����Kz���B��:�6�L mݵ6��2m~}��oJ��0y޿�+����r4!M,�`�u�q�XB�V.��u�e�u�l>+��z~�\B�����qMc�3{���h��E�����
��p���'f9�ʅw���q�A4���-x��^n;�,�y{��@aQ�#�h[�%�O�pn�iP�T�և����x�����sF�������'�W]݊�^�z]�J	b�&xE� Ѧgʳ��[�8���5��4Z��$�G��ק�99����Z7����}@ΐ�)%"�Sa�+��>��N��0�d���0�(���s��CϬ4��e�B�����4�+�$M'u9�x%~�R�i>�=�U~,��鋐��Yn������,CN�����{I�rX
�y�&^�X���~Bo����FPl�D)������}cm�sS���t|GS�����p��M};&�����R��s����I�#��)���qn���s� .쉤�v��4$^T�����+�Z�^z�0 w�j:5�gk�sd��<��{�!l�(E�m�p�Hv����Y_�l����Snjog^�^<�z�c���%��D�\f~��"�@�ֆZ���P(�_a!����9�U9'��&��${FFU 8��\7]ז�p�t¡*=���1Zg��ko��jK�s�\�u�Poz!ۢ�ǍO�c_�z�5���n�	z�*~���,G�֎H}�>ť�3b|��{'�M/�xo`������f9xRe��N�����qt�+�b�*7*�2�$}�T$�b�k�	 ��=�YE���e���[Y�e���+}3�=��'�8�ٌ�ѧ��E��>�9������X{[�d�5����z���U���'���T'魟W�4l�ږ�dZ,�\	X*I��Aj�����3�G*ޟ�NXXT�_��*&
���X�ca�P/��(�}m��ڥKS�5�>�jY�م�f%bo���ܽQ����+ 7��i�hM?x�V$�`r��Cq|�p���h���Q�m*�����]A8�����Q�dz,p�n��k���@�#ă6}�_i����ZXKGxgF$'�mɠ(Ϸ�Z�2��A�f���]�{!u*"͙�`
�*��G+�������ic���WW"�G�o�L�L�|؆��M924��TKY���3�����(���+�a�\S�r��Xhi� }���a����<��*������;�Ǯ�b����?<E���f���z:7њ�߿e�ƍ�<@��O47�r�A	�"�>ș�`�����Q%Q�u��֍'Pj0-�4�]�m�iC�����r���'�J�!m�,ȁ=1trM�ʯ��K���xop�TR�x.#�m�Z͘	���vn��gY�}����zw���} ��z�\i�f�QU����0�b�\��w�5�1�����O�]��0�kA<s�&i��щ+��P>��#�s��#�m�Pdr�;�.�-��5k_>K=ܩ��f�p�ds�z���A<!5��_�?E�(�,�4_�:)���LE��8�6^v�P�Hh���H-KR'q��%����ha�&�pOj����rf˱Y�hr6�줿�7��}��R���J!6Ŋ_�_�?�qGO�S����� ]'z��X-��	�Y�<ċ�#��p\�a�o6���)�m��e��K�Z3{"�}RB����Đ3
�seH�fe��gY��կ�E������5��0=�bX��I��@/�����,��!�����C�5Z+6�4}8�� 	�{�������N��䁑&�z�I�"�K5#�eS*1��d7��z�2.��8���\��/Hb��3h��f�"��d��{�Q��=�ũy��&T�vx3Ǒ�]_�`�����;h �g_
�
I���cU��rª�oZ_��0��yŢu�&vm�k ��n�]q ���a@?Q.\s���Y�W�+���+��{_�w��:&��x�-:nEs�"����f!OI�����ʆ�S���zRd��R�������+�Ʃ��Ɔ��׼�[/7�rg}�'�(�f�n����(C�4�,��Ϣ=1߆�V�Vt�-�΂�u�Qi��V�T(��w*��ͯ���@K�����Bx��sv�t'����aN�ݤG3f=��bv^�!>}��[*����o3��Yd�(�K��WS�睷'��`����
!��r/N^��s�DU��!� �1�����u�sJ}�����'_o2*r�ͺS,\
�j��f%wGQ���3�'(F8Xd����&M��M�AK��}(�ᛩ����]��z�ɺ$s~�k_H+���ly'�#3\�r�*y�.�:�T�ԕf��+T�㉅�瑘��h��c�m�24s\4�<~s�5F��T��S��`Jl%�2ZI���gR��x�����x����Nmu=3����0���~<�X#���,ph��XX5�T%�m��f!̚����C�}f������
����~qOe��zdݒW?�|�N���s��;SUe�r���D�ٛ)���;Ko)�h9�e�DD��0��lޖ����2�mQ��1~�'�s��[}�Ň�����pm��>��+sWCp�w�'b)�#TQ%��w���DM~⯂r�8�X���6���ơ��D�J��w�>�H��� wI�����ϟ����R���Y�ܮ=��L>p���:���xGWdudT�dl�E����u�itHBb�qX?��<�GRs��Sv��	����9�Yx7F{�G�F�9X��3=rH�zk$���;�����\X ��k�jܴB�f��ɶ�X|�#�w��p�'�p�y�G�.�GC�9X�u3��_Ge��Wk	�lֳ"�=T���c�2�)s#[�ݎ,�z�ξH��e�V�4�2��#�"��$���_�Ԙ�@��U�!�j�8I�p;хi��7v`����&����n�-��[���7g'$6���!o�Z�D�M?�$�y�<}ivI�+:#�[kklÄ#v�g���[M�1?����s�y�{�����hWt
�
��Y<�v7�r�������.���-	�,Gmnjs����|�6`>DHUhJ�5��&@����[T��0�8(�W�Y7����g	�IR!Hv�.m��]�;s)�W�6�.��g�\[dD�D,w���b�N!�,oPe�V�j�'�\m�;�l^�=��������^�޸t��!��Ɠi�~�g]�M*$�x3��Ñ1X~A�LPF�kO^^~|5CO�B�AFv��G첦qTL��
�>���:��U;�T�e��
 ���'�DA�s�7媪�.<��	]�4\N��m쭒��82
ګ^OW����S
��,0%M~HHd��x��[K�,����S�1�Vy�̌��-����Uw��E`S��|m��U��S�J�Tn�d��7>b�Ga1���5��/��Zt�û���m��]�M\$�Z٨o�<�LK�;������T�cR�嘊�z�����]�L(��!UW�l���(-��?`��4�=ۜ|yuumQB^pi �v
��j�Δ�\Ս�3)\>4��^��������v�����,������t��hQ��N(�OG�#e3�r���z"�D��� ��J�q�n����h�x� �pl�z���i5�vZ�qt?uHEO��U�].�-�LZ�U�숄%/�K���D�]�����JmN���I�:��E���6��,��/�w���M3 �F|�ytT氄~IV*hX�\HJ��u�N�̃i���}�]��T����y�Z��?����9w�D���Ќ���w̌�@'/O��\�7e��ŀ��V�$S.JU4W��S  ���'/���Q(���)#�j��3d#l��%��1�tu9�j5X��ȍV�o��8��y�.��A47Hh��J&#�"Q9�!^Yf��MV�$��oj	�]�3|��>���C�0����Y�.�D8p�n���}���Nq���;?~0�!�H��2�[���ǧ��\`Sr��U�������̏q����zerR�.-+�8sZ�2^�i�����X )~��>n�<���]�=[O�
1?�H�ԍW���L��,DM5M�ǒ�.%���]�%�:�o�_|��۱�ɚ[^nk�W�U~	�G$��^�2���q���(�5Dg��t	s��l��ӎ�&s��1�?����965κw���̨��yY�e)$�=t���_z�
��P&\9J$X)W �K�]Dƅ���`��)���������|�a��=�;�kRwiKi"�om���$F�&z�ݩ�Nic ��Z����'�E
E)l�S��Pr�e�Q����?#�S����2�~�o�9"�G;u��Z�/h��azB%aEe?V�k�m�I�̳ȁ9ú9U�E�K�a�rh?�b Y��F/>����U}����]dH�=ҮU����&��7���	O�6\� 4����^w�1���J-x�fp�4����/3�(2j�o�݊C���4DFh�� TI+����K�]9J*Y�3�qw9���ƫ�2M�B���o5Zu��8�Ց���<7U�Qo�h�Ñ��d[@�r�*�[R�5��*���ȼ�O������E[�r���`!�䋫Cv92�]�YK7a�:��
����~�������{�BJ ŰU0DB�]���t��h��b�����+փ��!�?�?�bR����u,���K�v����0��#˲8J����V��e���@>�����F�^�|����:F�r���~�S������͌㨇�ڧl���V
�mV{H���M�5�,�tpq�:�74�t�s>�|�b�P�Jk��y]/&�?�������9h�J���O����������W?���n�/�~�ܘ��T9�厊w&3�=�n�(;/+k�V��(�<��.G��]%.>Ĕ�
;Sp�mw�/���sV�r�ӗ�(��tM�'��Ya�9�b�#!!�]�o��Wc>���,3�YOJí�����*X��Φ|���sm��͈�}���ы髄��/�
Ķ�b��"�m�������
���n���oӡ�y�=-��F�"�g�����/d���%6�����(�z���hU�Yr���K�\�,]v5I�܅%/�+�~���0Լ�8L�|���}�E���F}C���s������y�-֗���9�$��<͂5�<�/X���+-��t��߱u[��z�ͅ����_6f�����w�5>�m��r�����X^��i7˥qc��r3���81l{w�.B������w����8B���/�qց��\k�d�'�k2����*--��^���bv�Ȗ�KM�F���������p�}PU��m�Zcl8�Ѐ��Hl�d2~e�"��$z���[�J��/��buL�{{�p%Y%(0�O��5-��}�?$����8��u�<M
��_$��T=u�×}�I�@pNؔ�_N�#b[�d�i��3q���4�O�=1�+�f�#��N���x ����~�I����ܟώQ�E�4��u�����?���<j�䘧B�2�!BB\Ы����9�-$�6z"�f1�����g�,�ym�'�t�bVC$M�=��
J5|��5��K8��X8�wm���7���1=�<kv����9G4� 1�W��м�f��ȳx��9P��^�^Q�"qk;�\�{���)�r��E�eԌ�]޸��3#���S.ӱ�(U{��S��-4��)�C|]
k&|S���ˍ}��lo�h�$�^�Nm삘GXx(�E-���.�Г?S�,7Qn+�A��r����ȴ43�#g���a�(%��!SO}�����x+}��xx��&AC���l�PPe��}h(�y��UX����F9+$��a�h���U��`����
7��NT@��)��r����Xж��'���'k�s.�)7��^-����������3�+{���dB�����Q����"���H�h��8m�{����\������ɕ�+mc1��;��mng%�g2�}:��8�'L�[��Sa��B���R'�W*Ů�J���|o�4�PX'�����.|k*,)Qӯ	���)�15���I�jdr&ڌiW�6:u��%.,ݭN�W曨获y��f���ĕ+9R���[���q�C�4�
�'�+�(�7hƆx�n�:'�$����׌�F�m"4��C��;�{�Y�n���-���ϋg�Kn���۪X�fQ��԰������f���f�ӷ�)���{*u��鲰.�h��kk|�5���"]�F�Y�^�y>�-˥mzM�F��� ��_�g{�1�&'1��旾sA��7�N�"ɀ�o��iz/L\���M�y�Go.u��ʻ#%�G���Z��z�*}�vp��&~xe�.�b~��;m�M�C3�x�C-�Pu۝�W�"��'\S\�z��&F/�nՓ�x�TYN�jG64롦s/Bf��iB�����q��Ƕ�� `���Y�x��z�2#�{<��qNzt�2��c�`T��s���g�>m½B�Mf�+�꣊O�h��.۝��v��!I�%־&��7��e,�\���V�������p?�N[��$��\�"���v��h4�~�`�q��=����N�P�Y��/!�v�5٣���z�ez}��M�(��-^��my�]�wc��[!ޚ$�{S��<�o���/	��/���3���1 ��C��[�a$G�#��knw�r&�7��)j*�q������Ť�� '�����}55Cf5̳/7bZ�9��Ě��U/J9 ;��B� ���� ��Cz˳�_��5�N����+)[dYC7-�nnc�:wv�;Dnb�k:i#ШM�Yl��| 3��4/)V��)�5!��|�KV
�Ȳ����������pR��r"����Z��C!�΄�(З�͢���7?��F���z���Ug(71ǜ�&�r0b��i��:rYGC�W�ɻ��O<��?�[[ !��j��D�y"�BS���+]���ZE/�L�DK������|]���O^LO�t�'�q�^�l&S�-��sV�X)X�f���pu���k&U����=�o׃>*"���/W�c��8֖����"��� 1vl��z.w���W��G���pF�T;�t�\+�H*u�������[���l�3rP5 89���bm��� Xp�[���Y;�gKlr��M�r	��d��W]���3ͧ�����[Y�mn^�Uί��`�+/n!~d�'X(�O1�Su����T`fP��x�<�4N����mA/VW�h�x�&�Bb��3�~�N6�jB��ƌno��6[��E��\�!���/ɝe_���h,�ƈI��x��i�߈�b�mHh��DYPP��K������sK��чľ�P������A�P҅��rV!��K�ioNG=5�gs�Qhh���'㬒�ͳb���m_�(����J��i�%*͔F�f	i����"wr����Y���ڎ��ԡL��m���e|hH�񶶾���[�b���0��Uv/�d��ΗW� �����+:��n���=��};�N��YG˧D�����S�b�Uϳ����'��B+�����7��{p�,:W0��7�������9��T��6�y�2ֵ�b4g��G| EG�M\�\G�������/�!U�h&�cMy����#S���;�|Q�҈�iv���&�&_K��{'��d$�}:��}Ǡ_N��8��GS6�c��ʑ4�%�EӠ(iM|��kX}��yM�r�4�qVF����[�Az�}'jy
��4%C��AY�,��O�o����O�v˧+�z�	�J�����u8
Aed���a���1 �+��᥇��M�ށ�c��/��R�m��!-��b��uN�lc;k�7#����8i�e�m�JA�����h\�oӴڦ�P���-?K	5I�d�f���@���-���@�t�qnw�G%�|գד������-ݧ�����
�%0]�+[%1�����εv��n|�ގ��U�^�U �	B;3eR7:*?g>�}�u�<��˺�����	ā_�J�U����k�$�4l��6ն6gԴ���1+�y������ǂ�=y��k�\G �pǆ�f�˼ſZ����n�g��x#ȟcW��x���p�p��ɇz\r�N��K�;�F�y| y���4����TVH�TW�8�؂�,��f�ț�>X�,���������r"��[�S��	���%.m���%/ϧ��K�pj&�#_Xu��u�â�"�R�}-�Y QX(Mݿ�تm�����`CQç����p�"s�9<������Ib�jޓ^��IsIڬ�,J���6�K���M5�c�ω���3�_"���d`s��&��/�ʟx��E'��<�5WZ�s|�>a�ʮt���]���k�,����I+���VP�4B:����1R���XJ��r�.,�b�x�
�5�˖��6ꂌ��.�G��q�<�?5�H�Ev8`d�+-�B�<��H��8`v��|e*�s,Q�p��1�3=��!���}vz(.���`���$;�Lx�hL	I~MbH[����+��^߰==%)(J
H�Q	i�fJ���c����ь��3`�FH��QcCb0���>�{�����~�羯�z���VW7�:rU�+x��:��b�b�Ɖ��5{!vP�'K��Q>.�e����%�Ek�S�A�ÊW%�_�CLT
t�_��E턡M�o����	��F���Uw_�&�|m����6����4��ܠ�us���v��5P8��{X��?L ��&0�uxԚO�U�C�nY�Q~X�����~[�V����/��;o����=wpT� :k;7���6} A� �*4��[����D9)(��La����7i�B�n@q����\��0>�"���Q�j��Tg�_q,���;ͪ)F�r�Eٌ�>��p����m�E�P�kT�E;�v���6tY%�N��N��GǮ����ue�,OZT�%U��x���=!ϧ�x'2���^�?>Q������	�b�(j:J��a���@zلW1�U�SX����N������]��i׽�Zvz.$��rJ�e�i�� �l*�1޻=I�R?Ϋ'ζ���R� EQ�Y���� Y}PS��bd�NNN-zq����-)q?�r�G�?��\A ���!O����)&z�].�z�_?�H�%
*�=r��>�"U��}���u7"ɗ��� ���na=E8����<I3��ǲ"j��0z���N�q�?���-|��/��(UuO�I� ә����C��`��P��$G�ʕ�~^L���?�_��Ljd���S���aa�C}��ʠ f����vv������	�=�?�S��d���,C��O�� ��xaX^zV�R>"��7���efT	��RL����o��?��}��o
Z��u<������L��6�Q������o+2�Sf�cSW��ӎ6�3Sk+�>��a�[�2�͔��v�y�S�!�����c	���p�����`�WCeq[������a^ �j��8Y�9"��#��s�=�(m�C�*��;/V���1�>Y��it����RN+�E溻2a��h�S�5���׳w�D���gZn���ތ���L�i%������'ps�{1�<�� �ء�il�B�8�"ۃ�z�������c��ΐ�Q��|MB&�u�}����r�dm���v="�U]���,C�g�R�����qs�G?�ɒ*�^P'�x	t'S������'д;|��{U��?��z����F����{���$��I��V�Y+�Q�:�������O)%�\�n��[�.�@�v����i���8ό���ƾ	�{���騵u�C1hO�ԋ��c�(����TFZBC�5�'zϭ(�[A�xP����|?�Q ��畟�sr���_�y?#g˗F��L\���V"����y���[z�E��=-��d�!�e����� ��PLo"3�e��>/zǀ�Á-ŗ=V���6�Y�#�נ���!��m�S�S���9@�Am�Y������|W�C�yײ�.������|
�YNx ��s���l1���J����J�Z,n��U
�gG�t��f�O-촕��J�I%g�����
����d�1gnJ�g��ۉR�F�9>�E�����U_NY��%k�2�:�%}�H��43�Q� �}���s��i`�c�W�dP!�-s%�sP�}vbK�ה�(��� R33�a�k��pHz������G�O��M8�-Kɞ:����pD�oK�]->�,��� ¾@�5��y(���/1�����.���K�d�Tغ�6�>`�
�sy����cC�����#|%t_���I��Q���ƾܘ0�W��M�
<G�w]����
�_����i�Hx��G���hQD�62*�ef�\k��{ވ��q %�R;ٛ���H�Nv��1��KQ�� v
W��_Y��;#���+G��+��9M�Y'8�x0�H�@B�[��+舃;c��l�[��(x��޻��NѨ��޷2c�����[���g����H~�rhu���w> ���rM��O�����g[����@�z�x�A{���N���kC�FS2(�0FD����ߚ�ۅm9b��+�����RyQݓ	���ó/�*9�ꐌY;W�`�������ڪ�J�$�Ҏ��pt�2hJgWQNP�"�n3}��?[����=z�����M��%ԁ�x�ֻ��r�����!G�����5��E~�^B�8_���0'������ྪ��>�������I6����Ш��0�������Q	&�?��'bCF�a.I�.����"����>��|>�6�2�{�����4���X�M�*JȂ��0��U���^S��VU�2Oe�cA�u_��i
q;r�����3%��<U\��ܼD�R9?p���2��'��\�����W��4��%b�zG�B�a��Fpgnj�����[�JF~�����H�U[]��������t�	�c��[���G�!��`c��t�pi�Olu.�	�|#��%����P����pL=k�T=��$�(茴=)D��\��;
��S��z��z���3%"��9��,似]-��.��ZP]�}IT�ճ�#��4�/�q��k9s���#�9�B��A]������Y��B��GJ��Y��)�๎�c�smbn�Kx����,j�0(b>�ڼ�x��z-mՠ�_&������n��;����M�DQj�g�5��$��h~5�����U���w�YZ�?��1,;��u�Ik6{��5~�Q����+%�eW�:�y'�6��v3�`O�V�6oz��@W���?������p�ކ�T��1�I}�c�_9�Vg,�=V���K�L��oA��lk{�c��F��e����L���q�Q������;�'$��7 _d��T~�@8>p��\��R��ދ�	YvM��Ə��C���&	�@|v�s7z	rneB��9J��#��>`�z��w㴐tg��c�Vu���$�[t��Ϝz���f��MW9�:�	�R4�涱�Э�"̲چ	w��Ӱ]��y����)��^��zX�(Fg�`7�EN�����әl�)�4qL����k�J�s�I��,oQKM����/��f�y��:h�~�y"��l����쟩�v�Q���%��{c]7�o9We��Gu�	�������#�'�+��O7��$
����T����m��6P�Sn)�e�t\Y���a�R��<�O�}f����u1w�}1��J�%�'ٵP��AqԘ�����A�z���`)`R��$�j=eS�ytm��t��7\#�g����y�YfӬ2���9h�5���I�gU0c��tvb��)���$�T|����wu�ؓ��;��L&�%��乃̢i!�R��!��?�)F��8�6j^���M�Telp����ie"����\�c�y��q����D+P��7�����/Wp������ͣ8	I�=�� ����ke�*�~?������	��쳺:��o�����7H�RJ�)� ���/���8�Ɖ��kg�[$Zl��LI�ȧ�>D �d%ʗ��6��:~ N�=�'�o�<X�R;�N��;־�'-�b�A������O����4)��Y��E�w;w�u������߇��q�N��x2>������(�򟆶O7$<�it+�N��1~���I��2��2o�X����[�%� `�a����(�-1D�W�;�Kɴ/����ƯY���������J�@��2��$�ï�G*�(q��=��ٯ��g��?�׳iK�:'��`L�3d�Gn��v�6e����rmh�� -��i|9嶼͜�Ω�qu�F̺$ꮖ�"o����������hZw��tlV�D���{Ͽ�?��ͻNZR���_��!cq�5B�G�-2'�y: /��r묹���w�>C�W����LW����ˢ_	�e3\*n�����g?
im�/2A©g^����8N��iK�ծ�_��ćU�H 6d��#ݞ�T3NZ�b�C�_c$�X����toMRC�Q��{�����&h�Y~F9m�jw�]���Ͳ_�'_%bR��l:�Ӥ�M�8�.��N��ꮯ>i3up�C�����lӳ��J�}J%�9$c������?�@�Xk�㶓B3\�S<�OU���t
��������4�4l��w��I��X��Ĝ��6�-C<p<�8C��0��C�����P���y������&��#�j���jԼ�����:�QĆ�x�jn����^�]�� }�f���y�(v�N�D�K7t�~GO�����o��ԯ'�WO��e�,+}�53����nc��w�G�.Y8��yk������3���>3���Be����ظ���8A����R�?rH�za�E1����#g!�H#��q��|�D̫۠2�͵�C��oj��S�Y�,Թ��@8�nŜOS9�M!QWJ��(O��i(��7��;�_t�*1��S	�o���\j_���R�3Q`g��VT}�ў=��fޅ��Yp��:ب�7K&�B��!�h��ʯ�)[Q��C�i<��W��_)	1��ߝ�K��|܆��m���H���,��Gk�J�瞢��<Q�{	�L{M�>}VB}C38	��F��]q6'�El�En�3��?�S�a��=!�?%��_��4В�l��ض���Q y͡jK�h��n  Zcq6li۾Pk�K���^>��ᙧ��1kq�;�Z���8��aSwIc��OZ��N�ކg�W4���|������Ž�?@e�VL��'#�1����/��dU���g�)q�-jCOl�Q�nh;Uo�q�F��T"����s��n
����ٴ�晬Fj�$ݎ.P����"g7����6�+^̨2{<����s��I :��f�$A�d�*\>�/�[�T�d���4�^�'��v�����r�_�d�V�R�T!�]��{wO����4����?���-�L*$i�f��4�N�>A�j�*U#�Ȍ�D�@
2]�tv��e�\�ũ��亘P�EJQn��/ճ�K����)2���J�pA�έb��vZ�ɱO�`���fJa�=H��4�/��ָ�7V^4��P�]G�&�M�
U%����#��G����=N\#����N��*`�Č��_$��1Z�@V�R��;!���@lAQ�R�ٵ�tW����z�M�P����C��W�}�eK	�8ɫxW�@`E���2p�4��m�6T�j�f�%���X���䬲2��FɁK�/�G��̖L������?8���[ӰY���hwƺT��Rń��R�[˼z��C��?^�^�R�P��j�O�	����x���*y�,Sz�l�KW����j��"��yE��������rP�kD����Y���z���k��:/!�"�U�Ze�[�w=������:M��Lfm2���`:�3� i�q4ӎ�¹���a�>B��B��g< �(�y5��E��$M�o����/A_�����Ļ�$6��J�����z%^��v����e���\&��Jތ܃3������l�Yy?:}յ��08�w�U�݋�ɫ��f�o�o���w�5]��,�_M�D���5�:7�r�"������4��}��.);&�V���x��"����㴑�| !C�_�>�ո�����?�/��`��~��j�"���y+����9�U>�D���Oe��O�_�/�;kP�2�f��Y1j�R�4��{��*A�"6���A��NST�U�_z��o�60�^��L[7c��ϲ}D���k��s#��R�$���Yg�ꋮL��\�?�xx��᫱�V�}��I鈈������F6�7y�^�J��kM�,�t���O�l�M��~v˒�Y���m�^�a2�砰Vݩ�����V�h�X���o�+�8��@�|c�Cc�O��ý�u
�ǗI�˟V�������XlPJU%6&�NC�SԜ#L`�CM'�䫫�e�^v�o�lE�K�U����7�����������'7���\o�L\��0�xT�X��	Emk=�>o��aF� K�Wf%��0?���@I�Q�Ԏ��ui��K�'[zRV�><Y$�Y-	��y��F�~�+#���C)���z.�UO��ۢG�u�D-��C��y�N9G����'������N�&��"Y˸�
��X3N��������TP�:�E�]�4fa��w.z�'�}7�;|���(���z0j�t�'�����Q�57ۿ�1Q�(��=��ף�Ұ_j��ʿ'#A�#�E�M��(�=�	��X-d[yB��u�̀�.c�Yn�����}����G�'��*�����C)�Ib�	�~�w��,�C'��;99W�%7����� 5� ���vO�o.%�!k�gT��m�iV����-U#�g���fԟ�ݟHZ����=2#[�l��Ì�k���d�����Rw]��R�"z�{�	�ǣ���h����b�kKζt��(����2���p�F^�H�v��=iA[5c�y1�Z\W���J}�ii4$(bSBGU��!MN�`�;�ݘ�(�8�ߤ��Y�G<��T�V��^�(��v��7k�\�s(m�H��횉���}.3�DV��M&'\G��DAA�J�a����#�ߝj��������(����6+�M���Dݧ9`6�Z�G��k'@!������]��Lѕ�������Sb[j��P1zJ��p�Ry�,>;�^����u* ���ҭșJ��Vv��(B�̚�J�����^����mHq�S���I�S�\1�.<������oW�D��T�/`bN^Y_�_�����AFB�뤐�:�N�Ý��l�X*�et�&s���_����NDPDtX�Ҫrze}���V%|d�F�����F�� ���]Ґ��lLvA1��]���h�F8@�
��%g��PX�,Rps���kw��\�M*�f�na|A�9�6Q1��`��������W��H<�/G�ႃvIb��;?�}�!e�vI�B��Hu��[��Y.���r�?L[�)K �W&H�J��5������h)c���n����>�����+���=V�UQ�7x&�n���P;p����ͩD9||��%YL�a�JS�@vLq�Z��<�5nj��EXZ�?3 #�L?̛W�~S�6�Z7y/.;��n9aqe���m�� ��|nF���;q�T@.o�("� Ըy8��R�a.󖯡͍ț+u?���xG�x=�A��f��͞i��ڋ����y`���1{%��&���@־��U�;Ly��z)q(����D��Ŏ=�_=�L�<w��J�ֿ�Y�`{c�=O�T���+�4���g�;u���Z����ʢ3��o%�z���\�ҿ�*5![�t�a�Gx'j��E��C>^E�M:S��/��5+�b�c��>�th.J�?Z8����tǺrUlK��}�U��/Ϧ�҈�\r���(�Y���m�罇_��*�Бsv^B%��~���E��J!p�D��y7H䓝����Rv�B=+!5e��E�~I���=�.w��Pw��RoV���w�XσxYPw0�n��Ҁ�\�=�ǐmێ�]ꐤX@P�͟��1dx�1�;�o���>(^��ޤZM���l��K�?H��L��Ծk�^x������	�����֟�^�	џR
���ҧ]XwO(L�oK=���f@2�|n��8Tx���h���@y*3Ko�����<|5*���qK���!��xpVH������M]3�sB͖:~��4C��.�M<�0�����m�J}-���� ϲ��Ƕ��]V�-&lΚ���J}��jr�6:�Pd#<[,��Nw�$,�ٮt4�������"�'o�?���5N7���_���F�V���ddf�$���#���"XWި��KQM����>ħ�X��<g���å�zo95��䎢�k�����
'L�J�6Տ4#
�ܷ%L�	���aU����}]��"Qe�\���x�$�>����,$A�?�0,B6g���+�v���q6�rVPCK��4OK5̺ە���o�FH�n'���
Ri�.f*��E2�i�߱t�p��}w̳�ޡ��Tǿ�d\��,�s0{��*���Av�w�Sx�=��ڻ�	S�����e}��U5Az��%Cg9�|T+��'�6�!�6�"��n���8�h��sR�G�ɫ=�αa)eԛ/�4�|��!?�m���S��~�J�Z_
���T;�
���Z\�Ѣ]�&ס3	�k�4KS:6��ZZ��n��� w���*�M��E��i�W�_�i��p�+f�eG�x�:�7~��Ս�L��F�_���;�`zE� v-�H�O����Z%6A
�e�N>��x�XPdU�D�W$۞�t$��ţ]B��ol�D��M�!}�R�WD����!�1�>�	@���W�����	��pY�u+�>!@��;�YH���d�s��"�C���c:�	 �Z(��I`~�o�L��p�Y�t���y���<auƚ�LkQ'�$���K�H���q�̝��NNEq��i�7�s�7�y�
罴/[�.<5�~����p{(�ْ3�AEQXm+��h�0t��p�%��&���g�Ɯ�n��z:����A�n��,���ND���s�U1��2%�ë�"��ʱ�縴��xw|���@�#e6�c��Ξ=ݻ�3�ځ�/\[?֧��|�kL�ZZ�t�8�>Z�
mu�?�ǌ����s
�1�ɰk�<$�$��L*o�@㻫J~B8�ε	?�/G��ȟ|`���3�7�9Y͹�{�{H~7�)S��E��H���4��HB�-����o�_4���U%*d��}B#´\��i�FQG�j;�뀹$�͛�f���ze���[���0o��Fw^�ٝ��M���)���ۉm&��2bee��%�Wu�}��O�B+1��>{�z�7#�XŻb�4���&w�B��Dy͜��(�6���ew�u^��<e)%�u"���iK�k嗩�[k�3�k�u��*�������"�W.�=��t�lL��Ƌ�(��%�BQ�'��1��l�2J���x����7�Γ�֝�fv��%��OGm�>��}��m��	OYk�}=��]	�gs�:B:���q^����x��T���:�M���Ç�[��&�����x1��y��7��K' 5�@�!�u'5��u� `S�����r�!Q4�ٮ�z���g��D�G޷],ѷ�����+�h�+W�:��ɩo������Ͻ%99XU�YҖ�x���5`�i���ϩ"���*b���Q�vǤs��t�L��@���'�w.l/�a��C�����MbX���x��g���� }kK�-H����0C��D{Վ9��������5�JtfCp~���vo��'j/K���t00�H�F�=DuR�U��\�*R��R���?��E��N��5o�[e���a�Q-�4�EW�(b�b�fՙF���8b��%��9�k8 �$�������N1���k(4bq#˪��=Z�W�m�1a�)������l�+��tUM�l.7���k/_�#⟽F���'�[�K�6�2"M��P�;۳n���8�~�bM �j�8���)���T�
��w���a��A.���b���������?�vw�{I��g�|��k%-8/#�ni���s�uH�ҁ��XX���Ե_���>2w�A��n2�>p�D��ǜy"A~�vX���w��Ч�d=���m{��w��C;A䵕�߂ǯ�����wx��GA�Q���g�u����s�@F�qy��!����.	���_+�|�	ը�������:
k!���
Lf�Ḝ�޷����`�ə*�ϡu!���@�`�P��ᆻ�p��B���u��"]��\A��0���盉��o���?�|Q{d45e�ǅ�_޿U�*^ӽ�р�W]kc@��pCg:f0W����#�NH��A�\�G����>�h��y��L�� ��<m̌���4�eM��sC�m�%���y,�M�OU	x�M���]��G�ez�`��8W��%��3�G��e�^�+sN&qR�7[�P0?,�.T|�����m��G�mr��v���q�m3�j�~�-��ѿ��P�y#�W�=*��[6�g�}��i`��L�E�kYV����X������<�[bd�.�-�ۼ3ѷӒ���8�������ԊlZp
�$1c�_���4!���Й�6�S߼�j�sR���A�BnA���l�W�dS����`Q$7�"���l�e�qy"�,��C�-���zs��x~���B}z�I��"j�'k[}�.Pp{Mx��I�s�ʫw�'߬v'�\����a"�2,�-:<���=-'��T@=h��%��8�s��l����ŋ�=A�Uv�}u����ەx��:���3����	/�D?[3��&1��Zt��Q�;4��F�i�E���.
v�' ��pR�k�9)/���5�c�,�t�i��∟E
�5�*xZ�f��Ԩ$��E=���$�Gع{ǿ�
�cB�U��u�� ���� ��B�ZC"��%����m���K���<�� ғ���ٝ
6f���W ���ܢ�W��^���>�َe�>�PK_Q��Z^
 4���ʭ7��p����'�j�m�CVb�N(ʼ�Թ��<�c���3,��g�Q{%�T�Ϫ�z٨���Q���h�{�=���[�И�b}�����U�#7^���ѐ��R�����ZCWsXA"ٓ���6������Q2�rO9v��e��l$����Ǚ�ɰYe���{luο��2WP�o]��F��<,�+�mĕ�s^_�Đ_b-(�m�a�����`9��z�-kM���Q��C;�{
{�	v+��VF��VS*'����(L)�60~���q�Ex�B���L+��OXΈ�y�?�+�F��_��
�������,`��y �a���(���Ulj�I��a*u4��eV���-�$t�y��ej|�f��L�n�2�eG?��K�pt+/�'�f&���/i�`
�Ȧ�V�0xr�휭��J��Ð���wFQ/�[��#ɣ�9߈���,�)(��yqE���I���t	���9�[�IVJ�Y[U������*�x���7�fϕ����描���_o��o{)5��h8wԓ�I���*��WF���)ߊ\��٪}�
6t���?�?�?��g�_V�lz��ݲ��--./:�ܯ�\����"�A�c��`-��ֻ��#��k��N�V=0>�6��2d�<w�CH-���b�"-EU�N�*�*n����U�67lSSV����/*~EKYL���e��u�͡�,�Q�|���~����/1�C};��,����M��v�����$���=�������aV����T��BV��S+G�HG�b�z��� TJ���?���[�X�3����76��l������~����o�]�'HC[�G�C���7l���^b�g\Ժ�c���k\7��� �&�á���01�~x��#uхȈ��H��!���t�q�h=����DJ�0����!�� t�p]�E lͿ���l����=�պ��"���@���i��/�H�[ޛ�xa�B�?�F�&U���s�9�a����ƲW9�`݇*9�*�IBʹ�W��O˙ͻ������ވ��t��5��Rq/m^";-]m�|���Xe1>Z}Tp2	�h�;�O+g9r̼1��Z���j�ZfK�� ��t�X��`&ܘ����a�d��?�)&L93)�h���̬�&�X5����#�Dq{'7�Wg��S��6H�ǰ*
;��/��!����[E'ܵ�*�|{0����p�ӥ��a�>�x�{��9�P�0��,L�uA"�|���T��t�=�V_5���� o�({!E9��~sj>jYԚ6�h�J�W�g���D9�"ߵ�������ڙ,�*ǶM��	�g8bܱujL�*9�P�� .�9�fs���R��.d���N�fi��`nl��)}ǟ!Ƕ������i���g�l�!V�,���:#�P����Ȯ�ڱ���Ɣ;!_�կ�p�ɶ��k�CONw���[�.:��œ�EV��]��ب���!����l�@, B������������	s5���"�L�w`,V�i�a�gg_ˣf�RzD���$�Qh.�]�����my��q�g؅����
��H��_Ɋ)��Zvg3��	N)��ο]�=�0a�[�~K��=&\�o{PWɺګ2�d�y��;&�������c����½}��VWxG��U$ެ�)\6'�>��j�6c.���i�n*˷�Yh��J/�٦B5��Ϟ(;|�mǁw�(Q^-t��6�]MdC8��Dx8I�w�[`���?�5G�*�k�'����iq��������$v�2u��I��[�n^��^��?Z\6��v3]:�#ފ���lU7�O��9�>�a\	��3�UK� �{RӔn���������l�N>6؎����.)�R�[��5�G��ni�`��rH��z�i�\`5��g8~�E�u����y�#2�R��5��9��6���8�z�u��u�>Rz7����.hV<����W�M�%�{���B4=Aۺ��ւm�Z(��=�^�>��"D奎׎���1Ҫ�@�P�X�y�g?F�ŨRh��k%����>Sv0#�I�37=�r�������݌��2��նȼ"�4\G]Ϲ���z:C|��W�Vc��U,O������%��N�j"�6�((���r�7X^|������
G��O,�_�<,q3�2iC�c��߀��<���ٲ��ƽ�-Y����mC���G"3r���a��2c��#Zus�h2����|�:��L(�j�'�M��)���Τ{���a�4'�� D��C��l��.Q���a i� 3Gr_�Q����Zd���^b������9�q%ah'��ʙ�B�^.���N��Hf*ԍť���:Cz���G���>ɯB�[cQ��Py���?���P)ѓ���'u��oK:���0~���)E��
�:'�=[��hd��@u4���}������5���g�}����^�a��TA-HX�%t�ƻh���56?�-2J�J����x4���T��_�F
��4��� c�q�_��.��*d�.��b�/L��2t��u˛̱h���D�p�qd�D&ϛ��f�&}b�o�Ą��| $����
�U�K�|��d�v��ٹd������;���׆�'o�:�Q�#��4Rc2H� ��z�%�Iŷ�YY�R����G��Ã�#x�Pk���C�����0{�/>���9�������5]�$�$_W��{;~�Ggqﾸ���hI�j�hD�̿�A���E�I����(�7�L�:}|�L�e�8Ѭ�3g�UY+������-����b�uz�_sb��;����γ� �X� ;Ҳ�/�M�W�_�*\2���ކ���~:n�����]Q�HY6?���O��>�����߉�v��-�7Q�x��¨�Z��Fՠ=�@=0�V
Z'Q%s7Օ��M��y�s�iI��x֭�Ev
+�3%8��ojKٹ6�xc,��K��cä����0����_rE_J처���h����L�Ir�i��z�V��j4k}�D��I��;��wbq��>�"�Ά��٨��4l�lb��M��9\Z�ɠ�l���Fh-�o��N6� �%��O�`Do���~�<�J-\?����(����ʉ��n��$��8�\��uK$�<��!c/�X<7)�/�<"^�y5k��g9�kgph�
����Gu*�8��j�ڶ�͹Y��T�H�5^j�K���*b�w�uf{o>�;��oN�jG�G��T�C\\f0�nxn�}�Ɏw)��o	Ox��M�I��u�r��>��k��6�N݊����&8?
�*8���<�C2J`�
{铰$,����]���H�ӡ�� �2-��o�!�?���H��;�I����ͨ�̴�'�;^��k���V��+��mZ�t3���/����t�� �E�R�K3f�j���_�I����c�7��եo"&�W���dx�A����۝��?���Qjrv�|��V[y�neW$6/�ˡ$5�?q٧rK?l$�����;��g�Vu�x����nd*�Mo��&��50�V`���l�jd�pHֱ��b�l�o��]&�����Lz��EEgPf�e�#/�t4DTAB��x
B��-�o@�7`ֳ'�B�Y!��7A��R��,9r�q�H��!���\�@�|D~���9v�Y]��t�]}.d�®z)/J�7��[�?%�>R�-�x�F87�}�X�k���~�0�����\���b���:A���|��2`X�hRh�N_q�BH"R�؇�0�,<r�wIr�kB���_��0��Z�]��d�6���=���	��|��2��p��rQ�-$��HS�	��� ��o��c�1`А9Q�4YH+�)Jr�ge$t�"��q���Z�y-�HUe�'�%��O�	�À6�1�tG���'u�V����>��\����ڰ���	�+���K��B��������EY����X����ZAQ����cТ%�Y���w֡ ���W�C��7�8%y��%�V�����MU�{��N�	��������$2�7����ޯ�,~�dC�歭��\�St(�Ҽ@umn��7�'t��_���|ˋ<B]���t������D�����&YF;��%����v��t����ш!I;��WNZ�������2E��9"mTkqf��R��2�'�'�����Z߹�����tp�\>��2�=��:��Z=�/��F���u��Q�k�GOQ��0�7�X֮)���F��܆�J��B��Ν-̎�sLY��Ug�W�$����X����c��Q���>�A��a6�����
�@m\�&�P/v*f`$y��"�
����5�_�lay=x�4�����1_o�����mư��9�1 �+m� ���[{Or��t����W2vX�g�jy��%�y�:�:���'-��p?14N[���*�F_�2����o���FZBJvӶ����<�	m����,��E�k=RBi��>Ү�6u�t���Y�1��a�ş~��M3��ID}�Ŝ���I>��U���%A��?�"���+5k�W81q[�����"_����nׁR{�H㻹`:	�@�Ѭ���o���W�j|�"eI>d'c��o}b���J��֨?���y�-���@g��t�3b�	z���ԡ-�/)I��QP������]�����`6�!9�����y�W7MG��r���"lZ��R�R��l�iVwbV�;炥���P�o��U;�&{>��cTtx�8JW��F�Cp_��& ���]����Ux�������Λ�	���b
қ��@����.>�m��y��8HJ_1%��/�k6l�2m�Ѧ�R︵��a�9�|�e�2f�G6�"b��������_�9�=��[�$K�zj��^9�M�T	l߿���K��9�b"��}[����|Y���#�pA"�A��9����|��@�T}�K��#"���Z);J�?JVT7�ػڢv��Ѐ��m��q��-Π'P��}�@K�Fŷ�rt�o�ļ�	��e{6�뷮�z�zշ[�ϳ�s�8��c�w6���q�Q���$��<�G�u��c�ѫ��!�>�.����O�|Ҙ��ә��{V���S,s��::˵�g7q�)`J_��Ħ�uO}�3��iyڜŇ)zde�%5�Y�A��u��M�j]$\ñ�4�����p}�Z/���7�w�x��)r�[����t>R������w2)_����W��� n:h4~��rV��=Aq����P�sz΁�~3����o�vCXu����v؄0�fjoKl׿w[�xm�"��EVJ�o�a`�	t!΅P��D�_Ώ{�*�B�=<s8�W�����7S���]�!S.�����S��f�BO�N���I�,Yaj��0wy���)g-@H���Wb��k��p�ˠ��#|*���ׯ-A�Tq�&�>�9����11C�i�ͨ�����Ϸ�)#Z��)D���v�y ���Z���~�J��K8��R�6��� ��f���s�FW@OB��9�T|P� P�1�Y��&]���e��̡�-?��5��Y�������E�}���<̍6$-��E��C�����<m���_@��t*���vB��qH�%:$���X���%���i�Ʈ��?!��c�~r��c�W!\H�2��#�mu4d^��L�=��wjXRùrJ�b��7I80�����"�]��S0�w��@����پ��>������3�Oг��8w�'b��;�j3�:��Z�9�A��4�Nх<zˈ�x<��)���Ue���p�!�����]I�� �p���x�(��Xo^����	ɴ�?T}w\�KЮ���#�DQDAAz�QzB�R�7�$�(�4B�&��^B	$�ޤ�J萄	I���w���ewg��y���}��䢛��[t�.N�I�Wx�gP�f��n@@�"�z�Ů.�wo�0����$�u+]��򛚣�Y��8Gbz������2������u�����kG��%}��m9w蚓��OЮ�E�w�������EG�-6�a�N�%�1�\)��q&˲ɕ�K��@�����Q�h����+���XǭL�H����`��뭔������cHO����e�%5�,��-}��1�i¢s�͉�;^o��L�Ӣ��׀e���\�#H�7'�z����ނ?�,����FMak�ҺD��~4iG9"M�A0aP�A�4{��]��i�X���Tg���.?����s���
*�X\��%ԎR�$s���U-��B���Ǳ���/���"7'�z�0��+��RL>�׹�s��.�)p��x��9-�h7FȑBZ��k�[�d5�MRG\������ˁ%. /m�0�Ï-�,ΠEN�wZ�oH5<����6͓T:?�:lé�Rc ��4�����7�}=�g��SV+��K^�L�n/��ϵ��{����=+G�������WR,ys��c�TuO�E,�r-e�����������q(";R��w{*�C��׽g���+	UQ&=�eĈ��fŦ��ύ�����_�������V�l���Q�-�p�̀d�pr�4�q͚�k<�N͗�2=h�t�g�~U����-eo���y_����fJ�q��	ǗU�������EM��ɼG5��I��dc����=�R3��Z�Jc��J�����u��%M@O�8��f�U@#γ�>�c6�ok��v�k�������x#�u�Aڨ�>�W\���FR\c:p��ä�W��"�s�ӝ�Q�Qd����HL f��@aw��"�1@��Ua���ʦ��&5�|�)~����"\�7�YC!�w}x������������w��9�v����I�[5C�җ8�|�T��K\tb ��}��cqhK��-\�dbF�Z�2$�&&}�u� 6Qw����'Ԅ�_h�
X#�>�٢��]�O�"ҸLM���O�����<���g��b����_�r��TI�.Ǡw��V�/U��<\�[#��T�Z��(��e����K�������ĵ8'©�g�ա�U*\�\m$�2%��`��0\��9�}��S�!���3F>�ss���sZ�@��Y�|�X@���A�����,@��e��g�������_mt��\5���2��'�ȏRof��fq4����4�������)֯�C������殹�{<�{�<6��N����y���ہML���>˷�cQ��0W���AY��|��O���m���>�!����d�#���x��E��d��|���ާ0e@�V[:�J�Y�P\��)�tg��?�՜�r�$��}p����.�)����L�J��K�!3e�lV�.�17D���:'�LJ������A[�t�r��s�b__��G$YǷ6�R�x�pݩ�<�7��V�Ռ�$%�R.q��*��X�_鴥m�;���#�ss�X�X�W���1u�o����A��r~{f!�Y�0]�����>7�,�#��c��(�o6�J�C�Zh�]��Ɍ~ڽ�~{ y�tR2{a�U��]{$�����[�I����Ľ�2.���:|���<�)7cb덀��ID��o���7߄W=*�B��6����6�jk����@�P�s?b��/��"�]e8���V�@��.�fb���W~%��3K�=��ɥ�I<���'w���l����O9īӆ�D�/��8�A+?��ҽ��h������3�'��-�|Q���q$��CEI�݅���l��&���f�@�O�9�}��_1�\c>_w=p��2�����4a����Uh���ެ�ƁNG Y�k]�^��rm��SA�_5�Q�actfdK53����A@t�6��</PC)�v4�,\`,=P�����hF�(R�3R���,�.|��X�<׽K:(4���)�K,H	��h�w�FB�V=����(��wVW�E��Ǣ ���U�X��L�����U5n�A�}D���俫h �����%���f��4�ݞ�o�M�l�*i�4c���5f ���aYK�iD���`���g�����*3y����KJ ���E�j��crײ��8��� tWA��*��;T�R9�yO�o��[�g��;�n������7T�b(o�{�p�,��n{׍����o	�R2���M�=���2���e M����2��y��Ƞ�7h7ˊMr�JҢwWO��j�vd���>� ]�L�i�N�|�]XYZ����8�J�)	7}�$a۞������\��p5����A��`��ӂ�\��^[ANv��	��0 � ��HM����?�`xz˞�_DB�H��u�
�{�'��+z+�c׵�H�O�4�2�;R{8.�5���~���}oy��kt}���$���uh�:i+��V�(�vxUQ��
���]Pbؿ
����H.M�5���D��4u���̴?u"-�M�C�1��7��OB�\B�a�21,�T��sb���U�y��d�7aҿB���ּ'.;�a����|��%&���\8YqD�/e���Kjl}�@~��^��>�h�p��D]n�;����#NdC�'9ޘ�l�w��J�.K/Z�1W����?����7�%R��Vۙ}]�����fs�sx�lLۣX�X�/-ߩ���֍J�-H��_��` <>D!2�3�v7�M����'�$v^Dn�g��iuA�h�e��8��Q��.8�u��`�~fo�ܿޅ�N�v��VN�;-�&�>pG��|�n�S�ʣ��8��#�遗��������f�֣s��яR��y�X�#-� �"a��@?��I>�?�_�XG��L�5��++/����y�n�����������ݷ��l��`�7����t?�l����J<���*���S:�.˫�=8���TԠ�}g�5��}�E���	^/BUT�N{�3rF�q�j��g����/��K]����Q]K��������歩Ƌ?y�b����ɥi��{VG�#�������P���;x�\��#`q���Ѻ�XLĹ����Ļ)�ӟ�;������}.�����~ ��G�-���$���芳�~�~�PD����2�ݩ/y	��9�Mh\_n���B:�T�f�8�P�]]�Ѭ��j����耕�i�.��7Ic��V����L�4�+}����Z����fR�L�z�Tۚ�q-�S��2w�"=j�`�y���zm`�aZ�ИF{(��`T��W�%�RK.I���9��]��Vóu{2��m>�n��\-ĥ13�R*ҿ�[�
��xY��O���ޭ�Em��If���	���*�i���y�� r��^�[`8�ʣf"�Z�~�}�[�"������w�����{��\x��ܖی����oFSK�����%q dQDAIH4����6�Ney��ӣnQ,"�l�罻z�Zfv�nMh1Y�Y�����E��/5p��>�+-<M BHk�_:�Qf�:��N����c�����7�7e�Fq���-Nƒ���w\��� �.�.�{D�, ���$�����˒�S=U~�#k�T\p+�M�["]��
�����+{��/��e)��R��\8]��J��C�QL�=l���U���#`x5�4�-���ҭ�fs~K�k��7h{�,f��bǡ��W�><ё���n��9,*W�)�7�`�W��X72�p��4�=�.-@`�I�&�J4�l��	9��k(\\5Il�^3�B�[)Z=襗.�����i	+��-�uJ����w%~(08�yq)���Ki����ѿ� �ɉ�����"g6�m,ID2>���7�|�6RYk"8%�Ĩ��X�y��n�oR��}�!����im����ǌ,��:�t��ٜ��3�W�ݒ;����S��s�4J�ٛ�L- ���]�v>��P��H��t*�.z+h�M�NG�Ub; �(Ƌ�xR��vl��rdZ�7RH��/ۏ%N~��($6wjT��@o���	��>�!�1���h!�Y��������A�:o��g���["�/�Kg�nM%v���fڵ�������׭	^�,+-:~�����{�ۃ�݌��	�i߇n0�7�8IN�G��OHG�z�4�aW�����1��i�;�y� �e�s��ۍ5��䠧z������`d���Ë`۵��_���s\얒J�V��2��U�J=0��OT;���ħa�~�Hx�_����7NA-������xN5zQ��+B�Y��OT��t�✵`̈���ߐuuVU��j�1�g�(>n�~�MP�n���]�K�L��aVz��]��%�/�q�޻'�G��5�� �e�6��rc�7��0X�Fmhl�%���I���������b���~������ɑ�9�U��^�v��q�N�O��*���(�]c�l����w��̬��6�,��T��lN��J�LM.���M3�ʕz��a\\]��Ъ?,#��[s<~D/����O��$�P`��6���I��`�?o�N�\��^���5�%m��[���bC�� 	��˫��w�:d�?��k�v�lv������@���J�R�lG_dQɑ����i�,F��%�2Bʏ�K���z������fd?@�'F�v��wB��-Y��q�SeK-E�r.KET��}H+3���'~_�X����!�~�i���yq��.�����I�F�G�V��狟{:ГU\��&�ν
#դ8�*�{��t���L&=�&	y��z<���e#�;���諾�o��8)���Xu�����$�m"t���A�Z�&�-/r5񥩽��S���"�5��tACG��Y������R�.��Bz��/�":μDPp�qH��c��1H��tؕ',��(M��l���}��rv������
�Ss�����^�O�u~�i��	u	���eD�i����r��wL䱰K��+^>s���������m����*�)�|��9��n&{zv���(���;���2���OF�@/��i|>��NP��-��4���C�ov�+&|
������u��ɲa��v���je0�F0������c6�{����5rr�Zv�z���[�.A+�ή��U�o�k������|�i$ {��!��Wջ"�	��b��M1��xl������떙!
�wõ�Kq(�؊>�S���e�A��K{sb]�d�����Wu�j�����B��#5 ���hr���9���v������x:%���{�>��i��Ƅ΄���h!�u��+�5�n�ć�b�;3"(�"z�k�[��6.l�Y�N�ąF67j���֤b�t:�6m;
qܦ����wY�v<.�#j*=�v>a*娣������+z����|��I�����uӏ�sEpћ�xl��وhȫ��CpP���K��fe�ɔ�k{�
�`b~��ܔ���V$��LfU.��*���bs���47�~cH�?�M�$(�-9��"t��W�Q!�ﴍ�-�����#�%,��\��������QTԴ0
	�f8Ua����8�:��R1[���o�&�gk� ��0bN��d�)�:�YvCsCJ�X�ٶ܆��	��.�����7t��A@,��k��d�.�I�&�t����e��/���$K�a0x���J�� �X8�Z�L�}��X�i$&MVb���Yg]�@��|V�TR^�k�[��j�Y��p��z�g�H�*	���_�h���RF�MvVm���%�~R0e7�0B�S�>^��3撧�Fx��i̛v���frw��Cl�&�y�{��N-�'��Ey<�X�G���%��㰺{R���f�`$�v���F�2#6e�|�6< C}�(ױDx����\�)�#�9Z*�E:d��>�o�:�B���P%2�3�%~�}u�o�K�N����3���iV`��U���	7�-��L�t5����04��w١pU����M8�-v�7���?��H��ڷ������D2�3�ҭ	��Z6>�ݼ�"\�N����=�/\�"���Y��@~��������lgsw��&h�7~�(�;���kp�{h�O��Ӎ�RDT����&�i���k1`ʷ����A��(�NNs��/�ٰ��N���e��#0ZS#[׀�6����Zh��my���7\�(��(�M�i�QP[Oq�2��GPs0�-rY(�C�o �5jd43Q��oǌ��";�%G��"��<�L���o��q�pŋ�w������̈'�����u#��iY��G�}�S��91㋱c)G�{qP~�%��T)E�e0�%���y�4pʢk�d��F�.��ڽ����&Y&%��B�2/,���N&çj��a2��h�c�P�ڙ\�a�E�}�X�<^��ۛ�L�a�b_ �8��b�;{�G/��/�i
��%���oE�.k�R�uiTNo9D�\�s2i|�B\kD��v�Df"K�~u��CĊ���Ы��*b=��v�iB�:���iv��kT�쬑��[�6"����Й����%�zٰřn�@��?M<�_��#9%~�*N��}���Bxzit�I��z+kM��h�7l��8���r�\�ȳo>$�J��L|�k9�(�A|[��>�f����VT�#�[��i#�/d�!F�2�b�|s:���מ�[5�Q���x���pt�1�ko�5�����K�O;睜8�5�
^�������U6>{����Q���0���,-��	R�5.�Kw���5��\�뫧'�u8��qq���vJ(_��xK��=�����G�q�t�����<6m"�%� ߟ��ǺT�2��9����w�;q�?�b�2`�!��{��8j���Gp��XsD�7�Guu�}�}7��A�y޲���ZA
2P�6p��1�X�)Z�-�~�޺���0�#H00���YI�V<�*�L75�\�����*W��"L��������v#��c�����@)x����䒟;(d�ڄ���K���S�[�mX7S�W�W��Z�s\Z}G�w������R�\ ԭ'>&ܘ�G�ď��'t䑳+7�Ւ��I�A�2 =g�z�꩚D���{۾~M�h�G�{���+�����Z\61��V�}?!G#��b��oh�gx�����a����UL�yE�R�{��9�\L���%`XW'����lR׎@��E���EQ����sPǌ�MQ�XGb��������L������'��+�4�6��r����uV:V�{;�s�6�в�	���fJe��1�޾�9?l�o�w�\d����e� �ʌI��u5io��8~���~^o���m�� �80�[�S�66�d�{�Q�bV�ublO�z��S`3�6�2gxS�6��0xP�u��V~����(/8'M	2�N2���?��^��g��]t�
� -��9�L�N�6�9��Pw�Y�+�!��~*�3Z�p:���Y��^��Y:��;:�ƴZo^�[)�`0�.�Y�����:(�>���I�������<g����]r�7ݴfF �FZlb
�μm�J��h�5�wt{�V�BQ��ݍ4�v����e����h��>{�q��>���DTPC^��U����n-�ɻ����4\�<gN��u�	ܩ�f�:q� ��c)��7��1/�r�����e�v�h�"W�+}�~�fh��1�Q��b�gt�r�m40'���9���Pw���O"�O��Z���"$���o�$tq掆�j<a���6����ۖ��_�eX�U�J�����p�����3泇Wl�����eڦ1����Y٨����x�M��\�a:��ƨ�:ܐ��;Ca:'�.���l)J�j?rI1.q�F��6�"=z��@�ٯ��	�hٖ16EZ�St��M�_ e�6�'b�4p�-%�,aR/�{�J>R�߲�5"�7\���I��̬w'>��nEJ�c#��8x�(S֊8�c�0B5=\NLl'9N�ת���
	� �\��z��g�ʚ6��.�I�����E �ӟ}����f�w����93������i�W)Z�m���x/�~����Kfʡ�kH�e�|�sjhh������;���h���լŮ	٣�.除�Ĳ����Jg�SRgz+SsR"����\�D��KK���|̄�C��2�ɚ6��3~�տ�t�L7M��_hh�4��֮�Ha&��x]�CQ�#�ޏ,k6S@�����Q�0�S8#�c�*��������vz�g�Gu�D���A�l�|}D���%'ˣ�#6U�����R�	���Q�.��&wܰ��2q|��kb��k�I#��-�;%�](~B.�c���.�����*�<e�����@��d�lxS8R�<9s7�nvp��]�H|B�r�vz�j�� ߟ�����kc_8*�s�$��3�1�E�.�=�ߖ&̵;#���p���0C��gD�����~��dޮH%�#V��)���y+4q�&�r��B�N�y��j���v�*�>�{�s�l��uԮ1���ߟu���I�
�� 9�ۋߚ4�ۣ�:�7�o�?���� ��� ���*�.�%Zɛ����2��V~7]3����>5����a�^�Y_��j���������������{�QOm���3Q���̫���''`^--�1C����C��|;�1A5mgO�(M�7�E-��JF|Я�̳Z���l6�d�	&m�[��we잓A�*�뫋�~'cI���f��Q�p�CɄ+ �Y�S��~��>��ׅ5ؽ��K�X�u��ΧR���"���#C���]�m�����)�%$����
�P)�?YY��	����b�"�m�_�G�GǏ{�s_g��j�{�G����s�2Y��78A0L�Q�5���� ���K-0�M�~*(���&��m)>��߲ �" ��R�%���-�k�`�p{�?/X��)$������T���5�c~�@�8��#R������V���Z���*n�����kÞ��������o+ܞ��	�?���f��hO ���������J��[��ϑ���R��M^
��
�Cu�Cd^���/&Īf1�K�[�y�� 6L_�Q�����R��
��1����VwS+��<1LFV�{8�}<F�����+���j����k�ܪ��M_D3�a���r���
NL-��U�,�؟ܗMa{���fS�5W�uƝ�U���(�<�h�LCd��xˎ�_5��`���D����̍��>p�h�� ��RI@�I�InD|�,?M���)F�wz��GT5�>�{��{��6�[pd�G_�R�G��̊��֟��/2)��6���D���K�M��w�����O�C��T�j��yc��s�diX� ����SYT_�&���X8v#>�6r�*�#oee���q%��f|i:j��$�⭪K_F�$� ���h��n��S����҅�^��ݍ=ٱ́E�A��q����z��Fy��d�UE!n0)*�L�I��D�*	��ŮaU�z�*#��}�zu	5��NG�yJ�(J�D4��S��E�?|��f[�{r�E6�����y�?<�!#P׼�
��=��>��`d/�	~w����VZy� $�2���c �Kӿ\���HH��ϨT���\���B�ڲ��<SƷ�%Ζ
	&/�_م�����KΈ�=���D�ǖ�xo;{ڈ����M��T	�"�7'�?�wz<��"Ɍ��X'6����G�|d��;}�q-Ɯ�a�w��k5y�6ܲ��A���Ûi�	1�)��5��)�IÔ�J��I�N�s=#x*�،���ɝ>�׌}j։��һ듦U�{[#Ԯ�D�)�I;O��R0�o��P(�8��+QH�ڦ*+1���a�޲���6WD�nWO���C�>Qf
�ߓ�3��������/
4'򹀌�Ҫ�h��?$�!�N�꺏.��KxC�n��W�M�R6��D�y>�|��Fj�R+��Sz�4��AH~���B����-t�<�=ۑ�1{��/�C̔t�(�F�ɿ��|{9Nz$����1OtoG�2n8�/���ڞ_�r �y1�|�:�UK�ZXW���Zo�N0c��l�əVg����|�����L8����L�#�k����S����W�G=��r�eJK_&�H�W��B3�F�;1>��o6��śڤ����Ό����'�����������7]�9.=&�r�K0���Q�B'��k��f/��Ӟ�)[*��p�8;S�Գ#�o�p/�x)����C�# :��5��}��|g���)�3m�A��5akp`"`*���i�T���a� �Oh�����n�$�+Ԅ�B�ix;��8���O����'��{،X��D�o���s�n'F�B���Kv�k뢟/��V�E78}�&s􋋓ʓ>H-*P�p�.�锄H��6���E�&�ۦ���AN1���>���Sc���dK�e���x������]�NG� ��^{l�N�!�v5%>�#�>ɍ���S"G0ۈ�^.υ�U�,ߐ��Ti��30Q�E� ��ef.&R�, ��u�ug@]gFN����5������*"�:�^z|5�D�DԿ��S
��|�R�F��{�dV��d����S�ƪ���5a.S�R��=�����d.�5|x�jݳ�=.qݗT����H���a��\#B�E��Z'��q�nM�
�2{�����ƪH������0�=�F���d� ��DD��؝>!;0�1eդ�+b������E^���ˠ���q篴vڤ�$�>������ǟ*ī����`aM�����c7�2������E̒�����x��햰E�X��z7������0;CY�_���rر}~�"]�-3�_����\�,\��~~���גv���Ǒa-#��H��B�a�~����h�m$��3�å��&̷VvhݶZ�,�FnO5�=݁�W���6фP;	�u�O�S!�#��ƎӼ�~��hHٽ8���F��I�����~d���'j�0�$�13�V0Գh�ա�@\ATDMT��ad��uflgn�#��l
ﰹ�,��w�C|��<��N�_����s�0����k.�;F��EOo�$T0��*�=K�����Rm�-�;a���x�F�9��3MΣi#8���\3I&��-�J� �դ��)\'���!7�"��j�k�����yR]d�JI���tf^p1
xw���\�LzhK�צ�=�w��éտ�٬X��	���,���c�J��*��jr����������#�^l�M����ɋ�%b8�-����Y���U�xVo�ho1�����*��HZ�s�F悼��$k�O~���|hg:
�y3�^��:���ώ���K\���g찡f����W��-VT6�\pޝ��gl���{�:F� >^K��o����wV=����E<jy+{2��EMK�ˬ��	�o$9�bF�,�F�>I�oe�,k�Jo���]-����&��+vu9�����6DP7�n]4u����&��*�o���:�5���_�LRpNY7~�ua�W�I��3�O�r���H�ٌ���Lp���?�ƺ�_�����
աBT��\��*dE�"��7@@B�ű�C���Z����7�L����P�,��L��G���M2 ���������[� �n��0����V7a�)$��Z:Uy�>���)��`L�� ����~_wx��R���D M���v�
���s��3O�ht�l�����v���g�3�g�9��e!��g�{y��t�n���Y[�9ҹ���Ժ�% ��>��ybް�w^�9s�X=?����@�~Y�ߟƾh�='D���H��EK\Ƽ��|51ܾ]�L`J���c�S�`�ֈ8�m�(�ac)*V`]^����+��౽.;nV�OcX����Iqx��N	��'��v����A���Ԡ?�~��دsK�u��-hK�k��iR^��5�(k}T4C1,��>0YuV�]����v#E���{��DV�ؿ�IwVf߽�ͅ/R\���ʲ���7�p�d�K1�Y�����#"��%�L���J�柣�#.�~��2�dCl��Q��KD�/�!\�ê;>��f�H��h��P�g�!y�a���]�W�|�!m�](M	����Ϣ�g��1׉�K�&��!��<#��.��&q��݈oB��5o!�x@���v�EU+�;�<X�c�����N��{cj����A�� ��nD`��C������X����<��n鋷�56��4@�ƨR0���;k3?��B1W��M���x�;�q�ݒ�X�A����\��'�R:օ��䆽
��̏�|?��WUK2��]Hl��wN<���<"���eK��K=˝��5mf_"�\����k9�9��}Gq�>�~�:�5�%0��iBjvt�����R�eդ�9�����f|{������lt^�~�_�q��T%��۷/ˎ��۬��{虰���:�B{c��m�SI��
��t�3oA6������-�ϸ��ֻ�=E��G�W�c�︹=W=��Q�>�<��T�����}�-���,���>a���W�����B�*�!I?�s�hU���a^�����+�VyM9��yof��d���^�� �+�����:�]�͏�eGs&����E���np/���.�����:��q�Oc;->5H2e)��N�5�*¸���/S��c#� 4 c�J#lo���A��A�_������������B�ʱ4C����L۝p���:�Ru�&��P����&�@�����Mo��^o�}&�ZhE��^O�R��K�$>�zeHi��ack�07$�̐F�ᕜ**kx�.�/ 1�?� ��=����^��ɡ?�7)���mݵ�C�kџ%|㒯��}���^�`(�z���aU0�̆��:�{���<�c�`��h̡KoOF*ݒ�1�6ڲsh����GM����]UQ����M���j��C?��'A��L�.�m_�$��:��o�$�Mb����ϵ,9���c�]wYX���x���[sU�up]�5J�.��ڲ�G�ᅾ�BGׅ�:N�\��5�������$���'��//d3�td��r����"�Z��Z���[���m3�r���,Qh0��y�ЅӼ:�(ٰwwD���R(���+�_h�C�.��?t��������������-˵��X51�ޤXu{f�>w�q�iC���w��5��U#!w�QW�0M	F�!p��>z�'ة��XmdJnfV�lnB7'���,��Ϗ�f1��hT)`� }-��Y�ٝ�S�jOz�BH܆����m���o��Z?,K�[K��\�Xl��D�S^��6q�U�r�=��7�-����nR��ZS�Ꝋ��1�R����,j�i�x�S:
��%��d��.�zr�S��B��F�1�7���[Gl��8GXk�L��;���/g\y��^%�"+=��A�NF!R9:���|��=���k�X���#�gϑ��=^�	;(P��!zs�8�ߕ���NY�mY��L����z%��d?4�ƻ9���a%N	�/�`(�[����&��V�)άɩ������ŝA��`2Hi�Z�����Q��:ѩ�v�?�x���H�ϡϽ6���*���D'I����v�$]Q�����s��	�]�~mH�D;�78P�F���|�w�6+^Xo�	��5�*^T4�wz�\�p���/��",�@��c��b9,#Ez�lj{N��3�_�!��y���Z��^T魌�0� ��I�U~�ʱT�qcVk���͞� ��z���H8����_g�{#��ٴ^�oQ3e�*�maI�%0J������9�v�����)��ו���̎�Bp����c��; �`��'��M}�y����O���{�
Ń�'�����Gv<W�d��S=7��	6�H��K�/��@w_��L��c��u������[O�X�c�~aC7VC��
'��̥�^������[7�Q�(5ƻ�s��/廱R�����N�{��3���׎��$��B�N�]���F�z����KuI�Vtt)�\I&���6�0x���i,=���GV	�y��ߎFho�Y��(6�N6^�/�{��d�چ1�0����&:�߶XWc��7�{G���%��ko��p9T��O���X{���~�M<e��(u�ȕ\����%:{K��:$� Z���}��/s�{?�ɗ���(�y���� ��wk�gg��ox����N�g�Wӿh���rWjc�k)�<�id>ѩg���^����)W��m���/�B�i^Dۢ�Q�n;g�?�?v�gK�jBwj�3j9w@14p��:�pf5�Xx�]��S ���N�h�9���4\��V���@n0|4�n��up	Xi�Y�o�(Q�Kؐ�5��y�5�*S��)��	��=b�)q��B��� �����F)����M�1��-$��z5vd�\���d,�Wl~�'�7��� �:s�%B����?U�YǸ*#�I�f^�{)�/B0��K}�v9_V���sn<'8�l��%����|{3Pkސp�N������������r��::6L�O
_��?�C5<Rح�X�Ȝi�0 j�G����Ĭ���l�9�VL	�t�Ww��n�����	��5����'�F- �!u�;
��?ah͔��P����CQ,�ؙ׳�;�ѻ*�S��0>��]��ՠ{�T�+�;�}�Un,�LM��2'�K�����
(��L����]B%���Q��E��ٟ/��e+�\� �k=�iE�^��R)�qT�v�1X����8�����.����q�厯�ܝ��1���`�t���h�Adxs��rl�'���׬�Oo�#���]�fQO�u	�]�b,��꒶b�Me�~*��?O�ܜ�s �T�>��]���
��_U��3�Y���|�k���#�/z7�9� E�����R �Q_���@/�fE�"~n��0sR��^zQ��z������4�YR��Hиj����Z�W�����4��V��{)%ѝ�O0/�3y�A9�Jxy�n�״%����J���AS^v�P���w��j6�U�N6����*��/շ��c��_��'dK���퐫2�&�8�y��I�����?���-���mg�U������ң��p�ȝ�)�1N�Gּ�+�j�;��&^�wW/�G�e���o�|��4@�F��[,.��𗸤Oz�/�Os�C�Y����Z��r9j,dY�p8�'�k��;���H��H����$��^�ţ�S��l�:� {'v��<���jK�[1���2/h�}uͷ-��'�/G�oK�Ĥ�-���͒����U#�'�yyG�'�Z����^�q����M�N;G_����\��jCl�K�|�Ri�
�����y|.c�'��8�M{h _^�TZ�݆F���N��<�l��	W��r��	���vk[�u�O��&x��I&���uZ������<�r�H�D�e��qGq��c��J����w��{�b��i�&᫪�E6�Z�����u�K�fa���m��bæ�ł�1���u������Og�2"�~Sa�n�>�#�K�d�QL�@�;j`��[���T�x���<�nӯ���«��}��5�h����+�����l�Vn�0�5m�G�jw+�D��E7�/h�/Q�ʹ������#&g�(����釒�5��H��`2�C�z�_�;�AC�\��9ѬY���Ѡ�y%ɥu�3�7l��냯�������e1�X���`"D����4���1!���S�'/�'z��7Mj��5s�+�z> �y�{��ݹ�;�BB��*�Ȁ�vXΪX�#?3�A���Q�݊w�:~j:Z��;IW��ƫ��{��/�7n���ּMr�#ĂezK�bٱ��\�x��L�A�=�/��©-�H��y�_V�/��kyb�F��2��rj8�5�ve{l8���PK�)�cެ����r��(~�r����b?w+p�S�~�)����Z��O���y���v��7��Iҿu�O��aH��G-�t�#��U�鱈+{���rO�/��;6���5b]Yw����M��<�Q5����p�~��J�$wa��ãD�{��SPg��F�|k�;)����w�V���o�5���8���*ì������ve��3#xw�~I��1U������~��\���dG�}d���?*�<Y���P�W\@,�a�?_J�B*1�lem�%jt��.�3��%��G_�j�����lD��>N8���t�2�W>�_~��w����g9+jtT����{s���;,�u�&�|YJ�����C�k����F>�Tj��|��̍�s(�t����L��i��V�z��=�l��a�=�N���]�Z�"���R�I��k@�=!@�
�H  ��I��^��=�&��������*�f�3s��sϜ�$���ʑ�&N��,��|w.�Z�j����7�w�Y��l�-S��"K<�z�k��ȀPu�*�^?T��h�C�..�&�,�\��sFi�;d���k����a���N�K��"���R	�b������Dު�x]���Մ�_df��s�c�E��cI�{P��i�ּ�~�b�a��^W9X��=L���:d��0�}1�G��+��ۏ��`^�p)����0��9�G�%�'�y�V߅�\U�Ff-��(��/�h���f�5��F/k{k�%w���#�օmV����.��L� �{"|6Ϩ�s��އ�c�ˑu�p�vи�Zxrw�����sj?�6�ƴXy�(j�[�=
-P��z��"�����{N�����߮(��糇�MZR�%k���j�*|^��^�C?Owa�͂���ä����.\2�+[��+(���)V�֨a��HK�5�,��_���զ�h�����jpHl�+U�A"�=7�ۻl��y�_�N�gb?W���&BCW�^�[�0��.������`�K����n�B�q�Q���2��ޫ�_�䥱��
}���>=a�sk(���͂�Y-�i��Q���cSJ�M�Z��DXg�o0�TmN.�:��;qq�3�yi�r�>`W��|s��H���:@�����9�b�]�r��V�ua�E]�'�`��V��t51e+D�{���8�
����I��Ӳk�I��Q�A�zt�s��(愺Ԭ	�@.�nC���p����i���$K�l/��h7Ot���^`�@�^�|/�m+�٥�U�I���C�p��a"j�Յ��ϲ�H����������Qv����u�-�eC?�Rd��tl�ĥ8o7�@Mqeg (ҍ��%��4�������*3��ʮ].?�0��K+'��E�L��?�/�F
w&�Ot�]MX�(}ӻJ$��\��P�:��]d��ڊ�4��p�9T�>�@#�ܸa���!��}h=�Oջ.t)[��9���ձD������[)�P�P4���2B�g�Pg i��v�Ԯ����c���rʶ͓uֆ8q`��Q��uѥ֥^O��iٮ���;�'f�fuU##��s�.���4�S jS��Ō�3x�D��X���4D�.�W����x ��V�{C��*��m`����ԅ8�c, ��y3�u3�LS���&�*��I8V�%6cS%p������ч�BaNl"\��)p��4.L�٬��@��ʗ��O�zor҂��C�~��f#��_��p�j��^�jGQ�-Rh���C�R������U�댑/�J�mC���K�iI�Y���֥`�|���s��V�6C]@\=��T��F�$a�5�A�=FU�-I^����n�υ/'����Jq�9k�4B�^KƵ�a_��Ԉ����dI.�؅ �)���>m�����o_�7\y��F�� �i�_���^��e/V=����a�Ƽ��Гp!�WL
|��l�����p;�0�UՏ/m���bR:͟�ؠ����!ySהnǝ�������o�՝���Y6����7� AR��ʞ)ss���O��d#�˥N\����n�)����|K��
\cW(6�3tx��׈���͹��l|��;�Y����!:$�7#u��gM҇��;��*�ps�D���D:Z~T{���C��$��CW�羪����|H���3������Y��<�X����Ԕ��Uj:��G��{�х�����ø�
��K
���V[hE�b��
�!pE� �}(x��黜��e�D�����Я�&�\��W��)��"J^������d���}��dEY�v��rR�i�4xˏ#ib�<Q�F��0���0!��l	ռ�:�n�C����d�s�&��)R�K�1CE�=�[D�280i�kŦJiv-#����o��i���C���?�w$,{j'�e�M��>���[��������,�W��3X���ğ�e.H�޽��F�ɹn�*��Ș4/1)���8���ܤ�׿hFG�:Gu�W�b�n�ý��[5���
	�F5:S-��-�Mή5s�D�x��8�"�Szkm��..�R�O�P�Ip`����wkƭ�0��y��y�C�Fэ�#��3�MkҿЈ1�X����W6T}R��#5����t17x�@���L�+%x+V�vp��d]~��u�M�U%�]�T�y4ݏ
�a����.� Di?(�g1����z�ق
C���Z!˯(�WK�ϊ6�J:N��'�<�:_O�5�R��^A��3���W��0��-�WIT�s}��_2(�gR�3���
��$ۚ6��K�G�&q����WG����c�=/"Jjj��$]Q<A�L!���҈�������F��?_Dq0Q��C�>���?n7�e�Iȫu�~����2����_�1M����u�
%0��@��o�f�eJgB@�IuY�"�q�����O�]�װ��ݯ1H4i��u��ZKX>EX�˦���.?֥%�%~�h������]���8ȰJ�����:�(Dp߹kE��-���>;X��?G�W���ޱ�41���M�s.��j�zz���ŨM\�� t�F��z�u"�Fyr	��$���oA�9=��b�ԓ`W��2!�eD|T��"�n� 5H�9�,Qͽ�}���>سr�1�#�R�����I�<5cE�4.���"B���.ўL�s��@X��	���̠ζ�J=�k�������axű���Ǒ�R.߰F������4!�B����|�a�N�^�M���#e�Y�	�p���^?La��������h���l�A�Hb�1<��������j0<C�ꠓ8����ˋ�߇�3w��F��~J���<\���ǁ�{�����k���M�����~;nF_{��~Xb��jV)0:���$t�h,�K�"mӱ�����J{��� �z�)	!�͏M���]�y!w#mX@CF�_�A�}���Ϸ`�����+��l��ZJ���C�z���94�~��!�W0r����#�=z��2za
�
�3��?�5$B��t��Y %!^�%o� @�E7"V��r2���r:���;�_0Л.�1���*w'=���l�� ޼�қG5/U��g�/Sjt�s��`Y���E^��/�r>;�pwmC�UH	�z�<;�� }�Z��7�p�|ol�۳W����g�:%�����'}X@�m�o���E�9kE���R����9�/�
�AOE�W��g 1�R<��#v�p��9��1-�9�͖���"�>�r��Y��=�覂i��(�Y��a���L���wFz�r�E ��Ԛ��Hw,G�^j]1̵N��� ������G6Y��.8Q����@�� ��G������5|�1>�kIl*�#Ql�hG�D����qc������}��x�9�K,4�Wp���rG�����F)y��]1���Y�T�Jw�oa��p���̉:�1��S&��R��q{��ļ�����{,�*X�Q�?�������y����@7����$�?C&��Ǌ��(O$~~��� ���[m�)<ˣ���#נ��8��3���
�L��"H��$�P���_�u��������h��IT"M�g��n�y�
���!�Wx�����nu�WMƵ���g-���p����#qi��ǫmK�.XQ�Z�?聜<�`��t���D�и��s��e�<���O𫬈opӑ�:)_�Y�%ʢ�K�h\�d�*� ���z1#��Rqհ��p�ɠ�]@J3�$)�Z���x���=�m+�7����0Xx�t��@k�i��c*!�I}&%���
#Ճ�ˑ/��ת{��k��=�UT~3�}>Y�b��pA�� ��GX/BF䑊;��W(��V�����g��"��vy����/����1�����G�RSa�.�<�Y��z��\S����NA{�+� ������<^���P��JA�Q��)]���D=Fb�)4uy��zx��i�������[���h���M��\��0���I��I^#n2��'�Y�g�=x�_��e�yyG����XJv|���4��Ev�맟y��Kuab|�=�ZP�Vs{�V����lm�����(:���'u�4�/?F���W�r���� �X�C�-+� ɘ>�3ô��U�s�W���az��nܸa>�!�{U,ϩ�9O�
����@Z���J���Sk�z��XdB�lf�4e�+ۃ���Q����Xy\�TP^�V�%:����C��)���0n!k�S$����×�"3�O;����v3�7�Z�0ZۼvG�2�"�(��Z���;�a5�SxВ�s�~��Sr`���-?D�b�u��܉�wdU�/�8,C^�rN�r��G9;g͟Sk���&:\�v�>;˵���]�z�~�CGm�B��j
ԭ�W��ʧ�Y�=��y����k������f}ѪH���Fraي�"N�=HΤ��&��3s ��yW����˕����ot�:�9�-)۴G���b�/<�y��Y�]v�h�<-t�'�:�>���+𩁢:��#W�
x6�i~t�|w�\���Kk��pgke}�Ɨ�=�pZ��q�As#)�d,�d���C
w9_��AQg����ƫ��������O<g�Ѥ�N�]�+�nM�Q\�����r%E��|����Ǩ ��e����U��R����v��zZ*����>m>�G�j��a�(O6���Q�s�}7�0I��'�ݶې�°`�@ųXf�{������Ub!�kS�\Vu�G�8K$�OY
'9���s\�"=���o[�j��S�J��[)�������"��龒`l������K��C�����ڈ���BP���!��8�؋�nuy�Y;�(��2d|�n���$C,#�l	�M�┳i�zI��s�>R�V��֜_3^.=�of�8�P/��)�k� �R��̷��X(*�7�z�E�;i�7c��d���M
�2𜆈k,˫'Z�U& j��Nˋ�U�OPft���R{翑��%R4�*=XӮͷ��@��Dv�􁔢�z1�F�Yjg���&�ݓ���tr²�JG���=��l7�z^��z��y߇�)2�1��;zso���唛Lz���J׮|��9�V~�r�t+v3�1fm>p�$�\���u�qκQA�D�~�MN�qH�k�_g4!��������w������g�ciS�X?���_�fwQ��a���T���Zr��l��-J��7�Bu����|����S�)J����E��9����R�CÒJ�Ep�����T�'!Z>E���6�@[���q������O5E�op��ݪ�Y� ��
�Sy����3�w��d5%��/�5���o�(D��C�W�"�hFèc�f��&RH-60傑mh���)$���Yۗ
��cu5cEk_���
�8�p×^u�.uS�(�qF���nL�����"�wȋ%�Qr1������=��J�)�Ù����h�&��g�]�����{#�(�ې��	�<GM�[�E����z�/��}eb�G �_�h�2<���`؂C�2���$)��!L��lf5�U�]�Pi��	��ޜ^���P��f�r�&VFG�$����kc�T2 n���-�'[�$�F<EhoE3k#�.}�-1?W�({a+��a���\�c��W�!}#n���-_/$f�f��?�G�J$�K�G-ި�Y��6!��Tr�huR�no���kjJN������(���$ �����_e��$��뙱��D/Q��@4��L9��:�sP*zW$�"N`�Ԧ���x�L��u!��)�����#N�STn��aMb_*p$� ���;4�&6��g�V"i��j�bkVD���K��YE������%,߆�a�#�ѱ	#�p_M��t �w3��i��޿�9 }�
��i^�c�&��-l��VJ��I��t����P\���]r"������xe��o�4�P������?㩎:��y���͜mr3�s�̨�U�k%�y2h��i��w�"�����<�6�~Itw� ���GN]K��;^ ��Rm�>�dF���K|�����%����m�F��G*��/8���85xg�It��v�J��)85�{F�"�VR�%p1'OԸ��g����&���`��nO�A�D�
(���Z9�l�1w�{ �H��0�� �ݠ������½��F���}��J����k[��x�j� .)�*!qf����*�x	<W[广G���&�[��'%��+���q��qI�-w��iG�!�dv�o51�/M���h_���3v+՗�D'&�J*�&w��ms[�ǡA��"��]-��P
kz��mj���d���[��z�;i{ݝ⽇(�#ha�CX.1�s�; ��3���/O�V�����E�UNt��k�WR���U*i���b%n{$m�g��K0$�fm���My��,AcJ��IF<�;��0�IvVh�TBuV�4��v/Q��}�[��v���=��E�f@�n{�7�m V��-���0��@�i�C��H]p�у����W�/��.�����D3%�1~)�� �<ڦ�%���@���x��t��T*1�y}����Ow�)��k;7�Y�O�^��za�v���犆���7��??���d �9]E*@E����=b�	��A(Qh��JpJr}m�̞���^$�~��)��^c��<�!���F~5���p���1�$�Te��``e[C`h��ъ=>;�(§�E43�9��^�B'�xq+�x��6%'�����er�y�����[LxߙM7Fם�(�C*,�G����|�j�9|-mϑ¢��HZq3�Y���\@�|�&+
fu�D��>����.���e� �ѧ?����y�� ~�Og�ժV���;b��3�f;G��v9`��)�@�đX�J�DJ/�����(���$,�t����=��31o:�w��yWaQ��l������؜��5V���G������B�m�;��Al��ڋ���P�qP�m�Y�������r��F����^m�n����.v�U��n���g�Tt����K{��qr`��t���AL����2�؅�Z;��d�+6n5��u ��_j��6���h�/�v+e��5��2��7���ǷD���[�a�|�7�G�F�%��[v�'멲�nuo0¡�][��d����^*$xp
m��1*3�
�H9����rOgGl��Q�5���X�_֤v-to�3mJҥ<���<Y�����2�O�a=���Om�a���u�.7��y!C�*v5���v�d��[􈘰/Û>&x$r�D��U��-#���H�*�6`Rq��烈X1��^�\�b6&jBob��F�Ġ�Lg͌��S�j?��_��<	���ZI�!��#Թ/�\�N�4=���.�����!�ة��V�o�:��k5�l2��[{m��&��d
�W�h�=�&طtx�
_���#&??�$���!��P1��^��91?c(?a�{�ymO�b�E%���Q�y�I�N9Q�mf�$�`y�i|-Hc%ϑ���T�S'�G��NU�ZA��f��a]�1z��(�Ԁ�M��=*�l�R4��5ܺEO��_�Q�OK~\�V��5�N���桳����g��O~6X�W����B���	0�f�Eabm��'�� ��w�$�B�Ψޔg��|)��)�~l�@��ų�ݞͦ4��6&}�ͫzDf#A��t��^�A'�iMMaK��B>���lG�;�����v��7���ۗ^�~�-�딦��<=�ᾚ���U�`A�=�@�R�(������IЂ�Q��4t#ì���m��*%߾�����{����m�}�����Q�^��kI�֝���{��d�k�w�܍�)�p���bAF�I�� ����kT�F���΍��QSz�#C��u)��x�}[&���,ҿ_n�c�
�Y���PǤ��nK.���t���j�i�(���YYE$H�ﯮ5��H9�e���ǩ3��X-e�F!{T���Rt0��f��]��e2M����K�g��4��<�d]˽~�O�����7K�C��PDk�"q36������@�_�{7��W`PȟFg@�olM�>_��/�H���f��!�������ޛ��S�aHK���.�ܖ�Q���T��y��?�]�����7��[PN�ò�B����� �"c�;&��B8��bO��k���|�`l����/U��^Eu��}ʄ�8m�	��>"��sR1�_�	óEwf��W��!����5����B{Σ�/^�M�;Jc/���Ҧ݋�CT��$T�8��لZ�[B�ʺ���rt���(���y�!�y��f��z>G��̖E9�;��sX�$�a�;�]0��K0�ޤ��$��p}����]�=����&��9\\�1j�]�����4V�~����l��4C�y-+'��n����]�?�i��jh��Fk^��	��P��B�\��*�<�Lo�������b�{T�.I�%Ϝ�����S:�K}�L9�N�/~�d��	�'xT���[��zj4DD�X�	���ey���u
��(#ۅ�y���S��^�ч���x���z�WM���vh՟��~lt^*3�,�eo�2!~���'��GhZ��_�����6�R�ʉ��i��OZ�%���*��W�a*�c#�@.��_�<�<�כ���nAvL������]���l�d2��h��U��R�������]�g�8�Y�UP�V�����X���%I�����E��S?N%aK�ҠӀ����m/Y�u�<Q4e����tr�@pTX�PY�GT��Z��`�n>ܢ	�����&Cc>A��X۽�_#F�=��
,+��U��>��8#�3�vv��X��Wx�!c�mF=��sD�_+����F
a����	j�^�]��FFaT(QGBe�]3T�ʠC�dNg�B\7���M�s�*�LHu�y�;�e�t�����C�Z�(���9�8q��O���������Kr��:�:	u:C�l�c��mӣC����8
��v�s�$�-(�s�h�����d������ϳ�#��J�殉n�|����S���*|�����*�ࡼ3�]ͮ�rC�EY�P?H2�pu��a�����Js`�c�:�4N��K�Đm�2�[*7f���J�n�����t"+�M�Qb|��ư��)e�ϰ�-`��Mއ��"��^i>"c�1UN#�;^�tZб7d}��/w��h�q�����[fDM�B�0m&C (�mWY_$,��a$xA�ly�m�5xX��t}0|�rY���^m�������⪘��Az��s��h��77?�^��z�i�=�l=���\A
��Z-�|= m�3
���?�I�c�����IC�Ͱ�-4����E���5�Q]�]��R���R�����>T�g���2]����(?G (ֱO��<1��wr_����u�ܚ�����^X�2ʔ�789� ���ɿ�U<(�?13��9���Z�D�5���A;{d\�K��	mÂ��+6��#����s���v�]�-i3��k�V�zH)I�yg����K$w%�w�Z��o�_x~*fg���o��6���u>��v��S�a��y�o�6+�:������~v"9��zG�G��J/[�޹b&��3	S��x�zvjؽ(�2��m)�2�R� kT1Y���c?���ْJg�-�$��^DO��oH%"��꧙�yݲٮJL���}�r言���[ۋ�����[�z6ڛa`hy�)���ɑ9>�h��KE���\��tgi<��d��U�Q(�'���}��*��k�2_ ��\���{=}=�E�`.�2Mi�5���Ct�nq�Gbb��KɋS���y���Y@#����g������Qg��{`�~�����~�\lډQe�$�w�ܣ�(��]ϿTC��>�=A*ܴ�ǹ��fמ�hO���iTb1����WAT?B���gt#1�p��`Q�[��V�B���G(����atW�Yf��aB�\뚪=�����;B���ʁX����B
xҎQ�+Ȼ�,+#1�������M���W��K�MP������p̛�8a7{�G}-��e��7�� �3ן;�R��_sn��iɤ}y_8�$h8��$��Ru��9K�sa�jP�[��*@��iB�*�H��<��
S�CP/tR�a�ń�?�Ө8!�ju��:.e���_��;&�b]i�i[�i�����h�y��z��(1W!P�C�F�n�8])��l�E���������/3�&�$A�	�1)Ɲ�y�VF����WA�I��,��L��يJD�毡!4��큙f�S��?�o�� 8�9��s?�Py�X=���)�8tw��f5d�VO�F�A�~��
Sl"�أ�bx���ys�g�s�o&T<���F���>�����}C������*�.}o���q\_E��u��
Pt��0�[��'����~̘���-g���]6�X���C7�@i@�︆���Y�g�҇��Z���b�G!��kn�����/�Iҥ�\�l�-EN����2ɲL�gy+w�Az���\�2)�gWXza�m��Xۗ�+��M��[2�A�0k�Cs�� C*�/����^E�Xo���n���{����s7\7�~>���Yq�^ ؇":��~�/t�]B}�Gg;7g�k���n5�HtR�����uO���H�\��Q�ٞ?���2�A��W��BW���[d_�Ud:m��A��b�B���&K���.8�t�v�{�b�d2N��O�}*�����	��$����k/���t��^�����I���2�w?ѩi��ZXO���.��*�wԷڂv������ܘ�KM�?M� ��' _y�[ma�+_rTG�)I��?ޯ>������>�el��ͺ�9�P1�K&�J����`\)F/ "j�,ϸ���]�ھ/���W#\NQ��YeJ�P*(.%zn5{VG���<se٫/�+@1��`vf��ᑤ���):���A���s�W28���\q)�_��lڬ���{�����?P]��$~������Z�C���F���53���H=�2|�殴�qa�<�̐D�>ôoNa��V_(��o<6�R�رtwy�g�^����51��J��6l�T�\a�5g�����K�ћ����%j6�A����]�S�;���[�a�r=�e�yk�;Gx������)�/�@<���BT�F=JV޴9)�q�ꂣj�.C���465�N�~��{�}Py��&W%�ԁt�Fi��w5��Ao�*�59�����:ə{�,���Ő���P�K ��U�y��[>�3���39 S���kJ�ڷU��Y�Z����8N��o�����`Iػ�R���Üz���+�B'(^_G�Eo�Q(!��c)'+�8���7x�R��G��JF��<�ps��y�4���]]6��0��Ñ��)��1
�5�?$�g�Z�轭ء�3s����`U���10�W�B��D�O�1�@��H�u��;�R�1�tu���%f��:ҁ:��-^�#lQ�������Ic/�6�e��!���h���uv2+�N�ۋ�ad%�w���y�n��,���{AG������3�3I�/���n�I��Q����)p z籊���_�0ر��ٝ��"�%�vr�ꠚ� C?�^0���U3�)��x˰Fɏ�M#}y��#p��Z(rf���ݑ}#���<{���S�8�yw��u��x
�m�q4���ƛ-n����RՀ2���M�=F�S�lgmVCT���ߛ�9@]�����յ9�7�{˲����f�l���������¡�ퟅݎ�U�'(�w7t�S̠v��������+����*?��h�½;��o�&���=�� ��_ a='��Z�]��2�g�5<<=��p:��(�p
K��_�0�,��헱;�^��k��Y��� je!</�6�%�G����iك�N����{\����A}�����(a���Ə���φ�Q�T��1�ӆk+��Ae�f=�7n(߽��&p����'�x�������7��T����@�H�gkKvmu�ضhj6vIA?k�����_��FVmI�bt#�� GE�vy������6u�(+Ai���FO%���:��F�����#���-�+5�(+A닉o�
w�ID�~���w͊��^�L�K*�g��^����\p��ȶ,{"��^���X��8y�烂k)��й��� _׹z�Wf�3ul����'m�;{x���r+~�ܲ,������d���w�%7��^���G��+����{����/��6����N��h̨�[X�zu�ɑ��D��9>��\�x�Sv~��XV��z���Kdj���u*�IN�0d�3�j��U��|D����V����_��Y��Q򌢴a^�CX����TU6\����A��x��!�̆o@�����~��כ~%^[�o�"__o9k�D`*v�៺2����p u7��́nf�f[U*���D�&�]Zz�{ʪ���HR�j'����F�R�8kD��X���?4y�^QM�W��AE�WZ�)�9�p��R����[����z_ZeS�qE{�ŷN�J}�T^!`��(o�l>u�`ԋoGA�3X�,`�fg�4U5�!�)򒗄>Ӄۭ*|�cT(Ƕ>��@|ƞR�0�ާj?-�������>��W��f���ޮ'��"��nli@U��l8o�S
��"T���n���w(��kҰ�e%$._2X0^��ŗ��/�pIw˩K{@�rWp��30z>�`��w���9�[�������h߯1���ǭ`����2�Ɣ�ڐlS�򶭁ٟQ&V�]��G���n�3r%��tyE�8.��U��� ��yUϺ%���Q�+�⻹��U�� ����7�o�G	Y:��$�b<%7�7/�s ���Є��,%�&�s���)��%9�u�#O��o�ӎ/5�
L�w������{v'_@���*\�J]���6���p�|�4ۅP!"��wn`��=,k��z&ܷ�S�գ=����t���Ģ.��f!�E{�������-U�7�,��+���[X9\bZ��_{󗸝�%Ȧ�.Cc/�:�Y<�o��|	��R|	�z��Lo(?�﫟-L�Q��Q����N~V�x���"^��גr������ʣ{���e�r}3K������*��^�nO�;E��X�3�!#�&�h��̇%o_�	�!0�����X�K\�뺆�	���(K�FY⟣��ˬ�	~� ��N� s?��d]�,��U���jL*g8�1���t�z����<$��u6w�P-+�,�K��\�1V�G{
%�����U���w� �c�º[J����]�Oo�/8�����Cp���l��Ycl�~&�`s�!��xV�}g�/���s#��IC�ߝ�I�B�{x�B���uE��LV'��f��4��j� =���@��承��p�[��ط�溤H�����/�#���-k�I�[q�?!��gۮ��㈮�4��� ����1��{$�-��L	Z{��Tǎ�tH
t�u�E��x������w�0ؾ7�~p��ا�^��N�r+�g�?���$�kQ�\m��{����Q�����k�e
������Ҡ�:�kw�S��-��_i���Y�LĦ����7���e$�ύ���<��ب����J�Xr�WÎ������M��b�래睜����!�ԗ1Ihr���|ex�&�'+Aqf���!wɑTvnu�#�$�j�pg�02U�i�z(��X綩d��<�?���Hk`�U~�cU�uvjx<��0���c��s<�G!�e��S(�?N� ��>�v�fe6y������� /ГR�x��z�$b6�WI��g\�Dſ�h��5�c�g&E+tx��w���,o�Jj3�!1�5�����W�,~d^��-�1�V{��j����뇵3Կ�bY�V���=���̼�>�-�Լ-��R�!.��9�R%KǹNO�-��禼�;�y�Ч�;ū��#�u���}s_�$}�Bg�qj��~m�J�%��J������}�������9�����,��Բ�S�e����h���tq� �
u��.ժwZ�c^�~O�ҁ�G|��[�����õ:��6�;�e�K7
�
�f�?	(��!�l�B�b�����o���ޑ���p���؄ٯUT��Չf�H_)�{����f�,R�Qu�v3训�?յP�>���G��_,��������U�NA�����k<9k>���2����� ��K�˿K��d��:V�P^xX8��87���ء͖{��+����uzsW�����D��q��e�{둕��!�pJ1�d���9i�п4��c.����.q��\�����|ol���A�BgZ4�W�(W�g��XI�\=��@�T)�8���N�'�Й�[�W�w6S��܁�L��ЛЏ�J��s��'�G8��
��)ª�$�5�W.�N��<��sJ1��.�N�J܉�io�B���[�S��i�ſk�S�yq���;���q�+z��ii��~$�������v=;#h��Y��y+ �6}u�ɲ��C�3d�����A�n�����N=-ۭW2���u���f������=���s4��)��_���g��~�-q[��g��v�f|_�\�����JP� ��5���$��M�u�R�r��3?�qGG�y-=�H�0L0�?�p�(z%7| ��N����ܴ<M@>UDB��m�sQ{���'E~��3i��8���=t7A^ʨ8���
�qYm�p9c/�B����ۆX�(��L�8��8�ڷ_�)fĤ�/l�5s�y@�wH��B��$J])�ԛ)�X囵���'i�� �L&��33�K92�I��q���=��fT+���bc��O���W�w��%�4R�%-nW��n����軌����3+��k\n���uj|鸭�wrBi�_ެh�"w���.�oE&���s�]�!��=s6q��A���D�zCAK��`�2 ~s-�Ι9�5�P��)��Q�r�r�N^���� ����~��.��H�Z_2�@���7�4��L
��.y��{8�\3��57�!�3�ϗ���zHg[nn�$�Z/�6ԔG��k�G~^�|�;�l��7�3�� %�؋�-K��|um�v��
���e=����q��Dx��	$k~�����/���ʲ��*BL�����
�
vE�-(>�����|Y��i(��_@:��xv�$���"�C�����Wn�榊�����:s�e�̃�H�e7��^m��$ʿ;���Z����m_'1�@?b����#}8�������X��1���H���F�Ia�+,Sy��^��T��CC��w�o�/�E���-p"8Y�-��@����n|����0�a�w\k�WF��8yVH��m�� Ct^-j	�^Zd>����H<��<��m��WxL^��Q��3?�1"�_��1�_�56.�쉮s���	�@^��"X�*�K�f���N\)Ζ���y�)$NcS����c�	q����H�?n�Ϧo��|V�3X��p�m�]�n�d��́�����*ob���j�?�9U�)������0|cxO�f\t��&��Txq�����T�H�q���8�#>~�m��_)�G̽�����Fp��i�a֩�φY�s(����Ƿ:J	A��9�7A7Ӕ��R�����W`��3	F�@�RqZ�)a�k�:,?�����R*��|��N
1����R�����%��� ��{I�Y���1�[��Z��5]�c�c��kBj��7!�o������Υ���5�v���Oi��Y�� �D]N5<ZA�ʲ	@�R�Exʎ3�I:L˓�9Φ�l���ײ�~��.U����-��CG-<����}��qRһG=ݬE0�J�ν~��H�viI?�ֺ�;!�Ȩ*�
ߌ����(	��{��U���3/�O�0_dx� ��)���H"�!��y��/��VRF��S�Ђ}�����̏�wLwhD���V�H`Q�nsQ��g\�e��a�19l�UD���8� �s ɋ_������>�������_A��4�a�4�yî}�zm|���8}�����+Å�4a�>43���m�ɒ*���u��A���ϥh��.�{�6�	�>/u|N�:PN��0'@�7`�v>C��W���5�s��A�/#�Xm����"��(��gA{;|�kŜ��DeU�P3y���ء��0)�Q�Lt��������վ�4��8L}n�t��;$0#a��4ɨ�>3����>6��'u�'�U_ѣ�P+ŽlY7��s�F9X�y���Hj�]�u�`���ho��yJ�y�1�!�?�Qub4�35�u��($�sL{�"(���2-��&��|��1�u���z��"P�H/�0�� ���/��
ƣZ{���ӯJ��c�[�����IE)tA��D�ߊ\r���*���3�-�TnI����f��.�m�w��n66�����`�=o���yy���շk���S@�œ��_-ގk����W2�N��ҫ�ʘ�q��4�jݘ��S��YV���_$#Ӻ�<���7Jm��N��ʽ���	�ΘbC��M��®�t�<��\�	�+3��S��pl�[!1�0�J�d/��{�&?7(�>j���KߺZ��~��u��8�廇�,����\�������>,
��-����e�v��A�yM{����@��n��6.��8��읔�p�~��*^х5��}z��w��I�PO�vI|�K���2[��6�JN�jDq�����s>��^���"�{����)���57�
�J�>�4��a�Z/�A�pC��?{i��qԾeZ��tm��o��p��|�YLw��a=t#zp�	��\Z�A�-�8�� G=��wc�=&Y\���B/����g�6���*[+�B^�G��RmM�"Z��B�I 7�}�4~�#��>DR.�x�����t" ��`�0%�M�	#'�#��S��{m�M�k{M��mא L��j���K D~��A߲�P}������|>�y^f��_Ȅ����:������_,�
���2w��ʥ�8���F�Ӧ�$�72����
�q+��� s�����=��z�qN��Z��?7p���{d��+�9寍��	8��e��|�=�_uo&km�+qC�
�����H��}د���.iD4,��GZ=���}Sv�Y�mJ����c��)MSJ{�F���	k���ő0�О��o����n�{�V�����z�D�Ck����w�]cqЯ�nȸ"J�2͗4����f^��W���!�ow����M�L��r�E�A���nC�R-���Q���5���Ehl���웲��p8�/�X̞up	��
��DO_�fj��Ɇ�V`w����^�i���B��
�I:�i��|�9܈�nк5zT�G����V�Z�YbV�YT��~�������
ň��o�NWhmWj��z.WF}F�?vx�:q�[��S�t��U�.�@�9�tu|8w�6��� �����Y��QU�+WL5����S[;rj|�i8j#I�K.��%�&�zD��Q8	�[�>�<�K�H��a�2�˃�i�������p΀�t+pe"�c�DC���0=O���	� ��Vо��5���X?��ƪ���6.�d*�6:-�#�&fT���b(Uu��+�s+K����o��hس�nj@���c�K�D&蒬��K�v◕F�`��<U�Ul�)�������}�_Qkw ��3�X�֯�$���kH;�-G�T]���qw������	wx��0<�Nڭ�u��q-[�4�D�
�M���f�wv@�"T����3=!O��т�wid{x�¼��r����y��D[��Mj��6��>�/��0��t\�}��l�B��5a�c$O2��ގ�A4�k���]$�P[������ܯ�y�Y�-4v���<qg��,�g��D�4�=$����,
�}0ݯV��jޝ9��	ZOV#��Ӫ^�0;e=M^��jCk�)۠<>�������>xm�^���v�ab��Zϧ�*J(M-���<*
�^����Z���&pO�/Y'F�f�h�
	���(�ӯ�`�^��UMCg������]��(�6��s��߶��6��{�fU7�o��Õ^���z���@�����nf�`����Ik�E��n�*_��P� ]ŗ+%�dְƇ>O��u�����$���GE�ή� �غ��)�J�i�ܤ,�V�10�]�F�4����-�ѹ��+WM��-i ��H�ش��c�HD3��e�U��0>�0z��1۞����y��hq��S*��˧0#`��3����w��t��2����H�X
�z�<ӧ"�A\���\�����C�8����������vv|��r2<�>�X>D���
/"�q��X	��/�~7b��	�֫�a��ղ���N�����y˵��aF�u-u�z�"&z�Q�B��`����M���F;x��P�	%,���S>���p��JE�>W�}�t��X�T���ɿ	,Ê��Q�}ءj��L"U[�s�e3��Q�o7ܹ'cK��͋_���.�e*)�_��yB@2I� Q�P��<O�)���7#�bw�p���\F�<��3+�g�GR�,,�<�[
e7�薆,��xu�ŭ��y��U阖�>�@۝粉f�����g�˟���Lh
�u�=0�O:h~��Ω�Y��;�R�eK|�*�h�lm�kA�у�����,�&�?���|Y���/2��&k�Q$U%��93Hi
����Nl[Lgܴ�^�)�� �&f�����$�YfrE��M|�!��(�LK�p�t�F�)�JG=���M�'�M���U���p+��V�qݼ9��ç�Q�~�3
��Us��6�t��o������*f�� ��Ӡ;�ڡ����n Ng}�0�H��Zyz����Hw��E=?l�T����Sl,^#�+4��I�����$���y�c)\%L0�k�a͵a�d$�4bIiq�jЖs�0h�������r�u��}3�*�ګp[��8i�a���F�2uRU�m@���&�8��Ec���(��n�j9�E"s��N��q�d�:�-��lx���ψ{�L8�~|�lCمnǸ7+��0ّ�y3�I�}�T����ދ+��?����?����(��Z�"t��vt�+�m\t��#y�����?lR�o�@C`�ݮ:bv�� ��Pd'��~������1���	�yk����r�/̂vɜ��Z>$��lt�u��1c�!�t��eVU��#�t+<��ECXbc����h|%��	l��ô/ ��?�|��-�<u%��u1<�����wc`��[�*�ps�4���SzK"9�E>r�K�Qb���\k���
�㘰w��`.���sY�hֳhi��VM�.���Eq1*<���ƨ�I3>���w� Jv<���u�z�߅}��$55���%�Q�I���	
P�f�w3�����g�l�ߙq͊~J�{5��71p���ZR��4�Jdb<,�0ۦ��r�!t����Sf�� 	����-���;fK�Y�7���n��9Pf5�p~��U��Qowtߏ�����h�ߨ�ƧR+U0���h1I͙3qq�E�=�׫%�A�ּҲ�fS�#�(�~�f�<��h�V\�8�F^�b�:�r�P��f�$N:�y򷞵e6z˦�<C�f�D�h�Yt4�%��`;��&3���Ο܏)�����"m�|�3:�r�w559e
6�Jճb�i����9<�\�����v�j~Fh:?\]d,�.��#Z���ּJ�r�c?�`�¶���ƍn[�����`���G&��	sg%�������V:����s3fuЂ��"��q�F6eBCi�і5̈=�>$E��ne0�]4*�$��t��Z�T�c��yܱ-����J/^&u=�p=��p����!��e�,����Hm��+c�58�J�寤�bA���!J�9�Ѩ�\�M!�Z[���'���>�@b�cu��sZ'��{� H�~���۽�<��V9uR�ɲp���чHJNS�#d�N�b&�p�T�P��l�\��!��\�F�n��8t0lڻ�$i^����]^卌����C���3�2CcMA1������xI_�?2O9']
p?������p5��V|4�W�ݝ�1�n�Iw�:���}9L�����
�-t� ��~�ͅ���ͬ�0+)�ܴb�}9�sV�;��۬O4��&$X�F[ƛ�T��.��1y������Af?��N+"�I��~S�Q6N�M����F��]��R� WKğ�Yi�҈/\n�P�=�D㚊��En<ڭkfL�nE>t � ����3�Ϩ�w�,kY�V�?��̙�.���Gy�p�M�u�t�7JH�!�#���g���'�%����y�ױ��ԫ���>q1̇�B �Abu$�+S'�{�L�N��W	���Z���]��LqC��y�x���*�vw]`�m
u���3�G0�
�$�~���W��}�y�g.�����2ieJ�g[�;�B5k�dk?�������^~����4�Gm�R��p���:e�J�L�+�y����z�ʟ���9'��xA��=�͇g�� T��ڽ&�(B�hàF׀t^-�o(�Q7{M�3!����tw�`׀b>~�����B0�9Кw��i׶��P�掀HzP1?�-��ea�W筮u3M���)�׃�A:�W�g���<^~Jq��I�%�q%�]�� �~TN�F�*�T���vso�E��:�=�@�1U}�EO��N��gR�E�	��&R������Z�ax5��$&ihb����{�	��SCUs���?�ǽy��W��f�u�oh��g�xG f��@����TAc���YpL�GD,�ڮ�B�J ��W�2�+�#���=L�ιY	㪔^S�?�A�x���6xp�M�����
����YoKL戇�-�o`�97i��4��x4�	O��߹Z����v&M��"k -�#�CӨ{KR70o,�)�����es_�N�x"ǼN�/5��֕aXTb���ZN��
���qr��o�d�9���y�e���'d��1v=�]"*�A^R,�~h�Ra麗�!��(޽i���G������k<v�@�Q�t*�uu�L����#����̟/�v�Z��a�pp�8��S��C� �*�c{�����
z�U���u��Qa��]� ��� �v�n	W�1��9 ��h��4RZ�G�9_�9�_ɱG~�IH�.%n�)��qb`j���޻kZF4���<��t��,<��F�$��:8hz&ϚV���N��GvaGlA�m��$���9����̒ݲA��}�fE�����Ē���CS�=�P8w�%o�X �i����/I�Z8���z7T�H�u�	u/U����U&��b$]>��l���Ks�/���K���1�_bmhy�<-O��>2f�����i������A���eʯ�⡢Z�TRx�2��������V��M/$��vCPe���:d�2bO�vu$���z~�<q�W~]�:6���9�&��ӳ��=�22�)�>�ao'=��}W�%���:5�����t��.����^n�z�J�cM�Ug>��5��.<7�n��MW�p�@OP~�+�*ީ6>0���x}�R����/��X��Ya!$p'ҰŊ��ЮI��\�Q���
�K%2.��=-4]p��h�ZyRM������ｖ�A��<�#�ppYc�=�I�S�	�֮Pq1�W9�k�v����U�`v��!L۪҃��4e� �C֖=�15���k��#\��R��dP gt�w�N������͆�Ǘ's�;���e��3`<�jl*@��xd2��Pa�6l���6�>w7����;ƨK�o�R�fp�5��^�%U�̟'q����Ȃ^�����b/(+j�)n=4��V�e���(�����9�Zzz ���:.�#"ݜ����u�̿���U�.K�!��
N�D�������WD$�
d݀��V�>e_�Т˦%a�f�p�a����9���'��y�]fKLn?��|������"8V���|O����T�7CN�U��ݑY��4�.�y&}COM,|MJ��ּ���tG��R=d��D�nʰ�/k����=@�f����M���"��ϰ=nW���_�Y"����W�!h����ݳ���2O��v�ԛ\>Ԩ�kJ��1�����b��egr���w�Ŝ~�f��+i���u�c��5)o��H��U��Ž�$���P�-8�[����+V:OW�]!�/ĻZj)$�_�W����#dH-%�m_
p#/˧����Z�<��T]�\tc&���E �*� ��p���$v�'7Z?|���e�[�n\<� G��T��7Z5%3�Ft+�i%O�?7�[2��;�%�����5�ݻ�ء��K����
��g�*��j�ۖ������Al�%'����BA�ڮ�n��G��1�����_i�+2�nŸ�@s�����I����o�'����J�*�)�o�=&���)�H����Dy�[�.��z�r�v8Li�`QC�FZ-N�2
V��:��mЪ��B���uY�
�NN���HM�D+�]=��ſ��	g�>�|���]/�fѽHW���CevҲҷ~�I5Y5�ý�.�& ZEi�[q�ev�wR����WG�h��b"33���{�t��
��i
������M>��/�Xqfl�\VI~��lm唸���,N�bg��v�,��f��-m�;`A���d��k�9پ7�م�V��Q9P��d\]�9��]���K>=��W��V�ꖷ�Dɠ��1��rB񺠾�U��[>���P�_������<�#	��Y���,�y�;�B��bψ\����c�R��Y��R�Je�LW3�y�1⢭I+�����Ւ97+��)jjE����jo�c1�%�e��gN���޷*=��w�@�'�T�d��Mb(暴�N�}��>��k�]�r�ԋ@~&xD�G�N%O9es.�M�.�ie��Q�jj��nc�0bo5�k�{��V�hgԮg6�{w�FD���WQ69�x��U5����+��T���/���a���30��^^`A$:��aʃ�8��%�����a ��ڗV}�8�-_H��s8�j��!q7�6�"8�-).��ܭ4�q�w��;lH�`�w�Re��������o�!6P��%V [�����-Z\���v�bg�p�+܌&;����xH��A�%�G�E�ŢS;�*��]N�&I^߭	N$�5b�F�>�@�����w�������~������%'��ܐ~�!�徚G�W�soŔ$�G����g#�%2�]�%�Q��D��[����n<�ޘk����
�r�
)��ؑ�jw�y�T�m�|�J��G�J�_ǋ�z� 1u����(��C�mY�t������A����2�䗒_��?�����P��k�֓�i�����eg QC��\gB>,��/�Bi2�~��#�Z����߃��;� �����1+��|�E�!���l��[y�t�Ή���&����U'E\",2�k��)5h�0�]���1��S�K��Z��Bk�z�F�T�y!C��&7���k^@�l�5w�.T�m�Ò��t<qj����_�'�=T%���@�uå"��N��Du##�6p�q�{6Ӕ]�Aف�]V����~P��1g�0!Lk���4�󀒣���:v����YV����q���d��")8�/ ^�w}��U"T�T�$�w��T��[�5r��B _��sQΤMz�:�Z����S�K�P쯇��3K��ۅ����K6��l�fkGA�?lZ�b�r�v s�]2�߁ϔ�����U��c0 /q%�cDu�����`�J��*��"-�������]wG��<�{�� �>�n�ާ&{#������{k�G�Wz��S����U�SS·Z�.���i�:HQ���L^
V�R������7���{j�ΈF=2�Dᙎ#.�Qd��;t�]Yh�p)������=�"_��
`���:����wW]��A%[�bO�^n�"	l4�s�\ٳ�^te{���z~x����"9#I��Y"<��	��jZ�)ů�B\��L�l� ��y���^Ƿ�1&���_b�;���)�^>��(��\D=»M����	6���q�@��c��)�����/�Ctk�b��#b��i����'���'���s�b�d3Y��K��@��37<��������%v�9��xO��{�Y�_3�k7GT!�ǀ��;��kj�J�1�r�G�_/��qy~x���DkL�X$�ù*c�,*����q�����C��yr��/=h��z55��6��%'C�/��)��Y�K��0�ܼU,��P��ʙ�� Q��V!e�ba}1�h-�w�����r��#"�R;/x�����]	�\{9d?BϚwM�0��2���[-�0牨�a��\}����m�0����T^9��}��+�t�꺶=��7y��N�s��e+� T&�د�駸B|�}��I��s����{��ꢠ�ּ�(>�˂�QS���TYh2s�g�nݿHg�#o��l�C�Kr۷Uxc���S<^xj�LT3�T)��*{��y�DZW���/&�mT���N����p��ڞ��>�Ľ3��hȂQ�(3!��c�|�!ǜ��	�1�|����m��,��Ϙ��zL�t�-��ɚ��"+�*D�c�����3�(N�d(�����v�����T3�\=���k5����O������Ԏ���}�F����t���w�*owTݧ�N�jϷ�R�?3k!�T�C�mb)v1�/�Ű�}�zZ�����S��oт�����b�-���C�� �m��>J��O��Hr}��R�R7�,����)8*����F;TMc�B�BUb�TkiA,���Ѷ�7��|�;W(�T�|ܲ5QI����B�����l��4��G~��W,Nq�0�$Ta��Q��%����T����m�+3��G�q�z�>�$$���(���F��A�%ڐz�I������<�5_��ִo=r�޶��,��?���V��_�0���l�h~+�F�Խu����wN6QOk�<��<qN����ep���åMf��*GI�6+-�u��"�k�D�{�$�\����=�ygC��Z�^�����d���<�1������w!��9ݪ� �3��;��ʽ��<� �-�O�?7w�Y:�o���?%�_�<M��S�Q�6�dT��Eo蒮�5WD�\C���455*x&��ZĚ_t��H�x�:,)��,�r{��z��h���oΊng~�Q����*﷪X��T�GP4��Yk�\b����Sʪ�a�7�����t�6��rϛ[�mJԺ��4�)��"723!O�����ˮ��=Z�E��|q�*�������������V��I�cH�嵽x~;!g��#��{7���M��#���R���ǖ�l�nb�� Ή���݅��.X��8f*a`*��
�wC�� ������aI�JK1�{,~��W;�wq:W��w�L���'�k�'oB�ӑO>3�3M!����M隇m�a�Y�l�ݤϋ�58��O�77���U��?Y�9t?3»�8F��
2զ��h�?��F�{�?��(���ޚD�l[j�L�ÉٗO�>�dm~<x�vk�[l�"�+(�"CwG�t<�X�Nh>,L:X���v�C�%�浪ϋ��\�������N_ ��ٜ35�����j�/p�^h�m��{d(�I�L!���L?+P;�Ny�;����RB�(��~{b�3���a�x|�����o�s�ܮE���r��)?���rI��Ka)G�ւEC�5�vZN�������#G&��g�n2n��{e2�g�<k���n�Xxκ�I\��A*8��W)-�"���Ec��*��ؿ�UuѪ�Dm.Zl���Y0�W�S[�"�dq/YS�r�4���J�/{��#QW�w[����@U���Q~?����j�9�}�'�3!�r#�eء������m�ҽ�X+׳��e�m?��Af�SfW���G�c�j�g�qH
��_��Jl�3�Ü{�k�k�R�(P_Ff� �5nټ?�VL��+|!�}"��jbO����]������o�W�u��Y��c��o�
1U���H=�/���}Q�w�zԓXv7��=%�d�Z��k\s&�l�=��vô=�Q���Jq@���;��K���y�/.����J.�'��~n�οiW��<%e���f�X�>�T�(Z~?��L�Cֳ7P��xҳ�x9v��W5��x�8_�#�W����p��Ibk������~ďęb.�dT�v�k�S�Lm�z��f��@`_��l��e�����jTL����;b�rt��cuxke���o�{���c����V��`��~���$ϷU!	��d��q�jdGJه=.@JJz6vܡy�����[-������}���w;;�ب@����WZ"3t�2�]	_�k�	�q���Au�u������(ʤ�ۡU�N���ve������gfS��T����;�4�'ǂ4���^�����r�?Ƹ���4`��c�%{$���EY-:�����9�SS��2鼝����(C�6Ky���>�^��'�u*lRb��$'�ePe|[,r�L���(+*q�X���2�.�Z"��p���T,&�J~;^���H�*�|5�Ǧ�2>Őn�Cͻ�C�HW��R8���԰�y�g*���>���FJ�M��Hjac�(�]f�V�K�dٖ|Gm@h�~��ge��GC�0k�m�PV��u9�rQ<��JA���@�[f�B��'TaN�p'�uԳ�,_��"yE��0�	�x��y:�C��������LWDZ�?I�:,��S�����]�����k+)��:��$����L��儶�82Gfx�A�[OzT{�|Y'a��M",�<�[Sfz� �ij0:��ͫ;H�sAV�G�H�p�!&���J-�z<��M�����xn`bpKqe7���k�ZR?��g����K_{(�������:ɾYM����Թ�v�D�5n��]a��u_�C���ez��g����#���(h������+93Q�q�Π�I�{ʐ5���G���o��p���2n5����O���P���pqC�z��h����~9��t29T�-��a�]��+{���a�����F�_��Ϭ}^�@��'}}�;��Q5�n{eeY��x��2.������E�*Q�}&n��Ģp�����u�<�_���#��w�R��'���n�\���^�N7]��D<�����������g���A��Y����_�W��2Ng����^[�i�<���/t�E��`|3��U����Ծ~e���=�������Ji�M]tJ�Sիq�č?[��\2��?�S���0�F�d���-��j�B�!��Bē����Ja%u���0x$��0����EB����w��K��'_{x�j�<N>ξz<��nW!�ٻLt$w6��)�h���y�#�(^i� SsCJ�EcE��|iJ��Y��9�S��݉��[~�_K����ez��%F�C�\v׿~XB��ڂ�?n��rI�C��[]-{!
W���5A8�,�gN�$��� �S��	�#���JZ��B=:`{�d�f%�(�ʬNac�j[�S�-��M����-�����Ű��ѫl3=��i����KŪ7�.!.������y��}�~6��&�n�ϱ �V%�X�{�����du��#��>�����7���?NG@���/��SK�"�2Cϓt`��޵�u'�C��F��sth�g�p�%>���2S/x{9��o�H�BI��1����h�vW�n5sx���E:��⹺�F�]��G�����ȸ��Kk�V��"���&[�S{DHm�PG�!�#^�bǑo�3詳�
���V�<�~$G�ߖl�o�w=������B���) ����|�m����L?�Kg�M��p��!����N�1���}�����FM�L�X�L�*a5ȇj�C���ԕ����4
�<U	䌂h-�Zo��.�xJ�{�����E�1��k�3��$�r����>��V*pOK��?� ��,�>dg%M�����pO�:�!�\�ӻ�$g3�,B�vӗ����ͺ�4�wV�G}%��[����08����&��zS�-��%
߹"�g-���p5�V�f�$J�~�hc��Ƽ���[�8����oK]�Bpi8��e_��־�?/�	2w>1?��%\$U������㋕����Y��y�]���T/qr�PD{�^�K��#�0�K��$�il(}lZ�v��þ�=3t�?��2���vj:��F�ǽ�D2ޭV�PP@o��6�	]iy�����!�xL,��E�Ae�? O���c��Ik���:��)�	K�hg	�8��e��oM�7�_RP�cp�����OK��D��5���m�W�B��KAU�~�L�K���Sm�&V���%K���]�'����4�u!`���s�Ç�7��0�Ŭ_�k�8o��d�����s�%���Fr+��K2j��
�*=�RD�qLkͬ�.���8e��U�b�%�G��{�;�O9l��EN�9�i�O��*Tc��4W� �V�}�Uތ�2�T���cp)!�(�W�ֆ�m��k-�����}��0Wt'
�#���_��bJ���~���KO�nr����qE!�~���3��e�ɟT�����I?5��8��{�;ߤ�]��s�ed�b��4�r�RZ{�fa��)���N�ZJ��^���ڏ��L�AG��	�x��+~ �y�;�5q�����
�-���m^�qG�7l_%OB�V	C�L�GQe����5VZu���jȑ�U��_��>��'\�al��^�h��<�2��,*3�u%~���N/��U�Gu�͎���˰rDK�>��c-�y�˻�FE�
��p���������L���,K�ݬ�O[%�3i P�ɀ�+�?��2.:Q���T���A\��$�_���-�V��o�p q��%[�|��ԛ�����B��sF[= �X�8S̤��ñ���E����ߝ�4~ᅝ��&�O+��i��ݜc�<��c-�Zh�/�aW^l'��F�nT|���Z􋿩F߾�wP��;%���N��� W&B�Q��A
�dd3�v��Ab�:�6�X>ޓ�$T"�(ì����B0������+�}�\=�%2����N��|��Q�SbкK&vR�s:K�w9�O��c��C����%�$���*등U��ٸAzI�̟����r�D�#_��À�`�aQi37���������al�e�'����>��� �T�ব���l.���3唝�>k����M���ﭭs]�X�w�6m��F���/��f�$M���=�2�&#*T��!�>���)l
Ye�?Gn+��!w��u?{r�luC��uٹ����f�4�譬��f����`�0q*^R��z���M}�lݾk�����m�:j��q|=��)va�&�]ԃ-W�����0v�y3�B�Tw�<�fb�t�M��`WCLZ �~(B�ޖsU���έ�a@s#+��ڢ#m�&2�H�zK#=����~厘2����L����YYK�@Q��:�uuؓ{%?�����Z����/�YJ<���R��n���u#8��'Sf7{�5�\ʵe�~xc�'z���y<x���B�'�m�p�:?]�ws�V�����n�\v����^�k�����l׬�'�?*fi'^�G�xP9�I�Tp�5�"L�G�o�t�s8w�m;��5��1fUy��bu��$��$�~��P�C�|��\`�e���B�g��K`g_��@Cb��c���x�׆��Y��W������.��J�.W-|�njPrL��H:t�2!u�A��#������[�6)�wm���O7�Z�z���ˋ�s؄����PK�@�M]�<,����u�p�z�p�V�>@��B*;'�����ǃ�i-���OEfj�EYF�x�[<�p�Vn-ss/D�L�(	@+Ty9 _K�*�|l��ِē�}�hF$�̥���v�z^��j(�(��qc�r���uU	a�y����o�����JDӆ"n�^���#e�z�Š+����OT>��U����GIu��`H(�Z^=��ВH�,8 $}D���á[w�����4�Z�&&��w&T�aַO�.L��y�#������i���X�sd�~�9<�[g����2mQ��yP+��5Th��߀��s���ӻS)�r��En������
��q��OH�(<��Ow��m���	��H�uSJ�~ݨ8��2OAd�$�/�Z#ok0�n�\g�8|o�����7=����u�M�	`�}ӹZ+%y[��Hlwu�`�,��"�.�&���[����?�ܵ8XWOY��L<W7e
���{8���M)�Y�
���}�XÏ�o�z�0�(�3�ڟ��ѳ��J���oh���~��z�����������}9��z�T�{'|�dPj�0U3�MB?C�6X���l5�H�zrP���] B��6�L�=Q�h�pF�/��b���p7�&8�H�-,��Vu�������4��֫����|�šM�?L�GBE����0�p����K�����P�DT���إcZ��R4���[��F���eTi*���d�5"�:S4����S|S�!�և�[�?�2wy�)ōJ���=δ�Tg��V��g}<۾��յ���SPD�����#��L�z1��m��v�a�|UP�g3ZpOړ(��;{�C�[̪r�â'O���pY��ZtFFG=�?��A@��q�I �.�xX��~ֿ��o�%��44;�*a�>�w ��N#m৿�B��]hk����O_�8�ktB���|ٔs��,�����Z� ^�� m�D��Kho/X����^P�"q��L�L^��;PO��n��tG���7�y-C�-�7W�
ݨ�	r���m�6U�H~a\���ݯ�ه���w#o�Xe�cN��ޥ���<i7�Ӹ�q��t����̣�I_Ğ�{��^�����ˊƖ�.�|C]M�ޓC�	��F�����z��ҡ'�F���UQ�7����ޕ�R��Qj/&WD�9Z��`|�=Ҧ�o�O�h��B��UZ.>x_��}��}�a�y�
Ӈ�<a����O�Lb��%oǐԈ�2��0\
�B�r�g��K�9X��<��l��`Vw�{��`��تm$�E�+%��b��T����T�c��	Y��*؟#��ْ�?ޗz5
��ϛηu��lߵ���p���S�R��h����~��� �5� �΁�O�]����CY�m��x��8�C�8��f��\.��"tJ���g�A�\��F���z�$=�4ie�~�MNN�+jD,��f�s�,�����Ĳ��bj��^ޝQ_$?³ k���IS�N���DE�x��.�6
T^RtuOQ%*Z%G��\�+��Pq�i�"G���d��.^��[^�˖+XQD�uJ7�Gb��lFV���t&���nxi+��۹����0KR��a��J����~��7�m�*d�ѥ��G�~�	��W0B�XoN=��iS���Wn�x�����{�Զzc�d�gI�՝��U����FP O,��һ���F<�c��J|�_"8(���YY����I�`����]�"�1R
Ҧ�P�@�k���<n��S�M�:�fyc�hT�ͪ��y4^+[��,y�ȯ3XgzH8�3Uf+p�z�kR�2L��I�|��M@ȟ,O�gĺ�����Ĉ���j�;��=,eF������XB��rb�h��Ƒ��s�a���ý2�޼���e���t�k���s=i���9T��� M3�n�\Y�^�]d��l ߍ��B�srθag��h.0�n��lwV�_���%�r�vuK���z�`r�����s�ME'�����Z"k��ʂ����Dݖ.�+t8)btiR�C�턗�hUXi�~�3=�j���o=���F!j�����ۇ�u����P��_y� E��H7��f��z�9��-�2�I�:�Fw!�`�3v� �_q#�`?�/��f��X��V�Das�3u�d��J�'M�Z���DJ�����z� s��En��z��1�}���pQ���C@������-f�
�4�}bϿ�X�VYM%������P��7�b�����w�-���i֫��Ul~Cح���kPL0<\��p�'���V�XA��3'q��k$���밚��S�%����������m-�6�~�C����C׺z�+VF�6:����q2TN�y�o˚u���>���u�"���E(�(�;��m�M�-�l-N�욇�;Q�ݶ���N��8חp��P��3��Q�A�ߴ`����݉�ղ�i'�y�]����>�l�T���D�2�VUʊ�:�?+A8������_����l��ʥ��oJ���a��'8O�J6��pwN� �dŃ(��˸�\�������
�Zq�z�.s4��ab42Tփa���c�.�9h�ٝ,�I\'	��^=a�2���~�"-N�P=ӗww�}�[#d��*x�ɅZhSVl6cS�U��*q��(�� ��� ���g�/
�DAG�#�w6IϷ���
c~�{fv�ߏ\"!�=!U{�W��v���jQE}��V�(�#� ؠ�8�l�q�����R\/�.1`Zbt(��D2��[��3O����/�|�e���i�*�����d�ӏ���A*��W���f�>J�Ӣ�	�_n�퐳7@O!3�]eD=� I����#��'q��efQ-�ט���J2�I[F�Ν�����u�c#k��<}|��kx�c&@���;� (�nZq��#����^��Ѻ{�v���=A��ΪX�4z��]��̮�{��Ɋ꫒�S+}�F�t�Fkbϼ�E׈(�t�@*�Z�����>�Q:�[���^���y"~��cJ����=��S_����ݮ$*		�B�˾�l#kBd���-{�${e��d��"{vc����1v�S�������s�u��:�=������X�C��C�U�@�Ild���� �t�D�R��S��Q�\�τЌ�Sl4x��N}���9U������_ڹ%R�!��~�a ��?�믬#�6'�oL��
*!�=��w~���k~ZS&zc�!Y뜗������a�&?$��G�ͭE���a�,���
A5�"�Ж˵~w�h����׬gx0}�J������ݭ)+?o�TA)�q��U��}p����A�4F�������`�=R]�te�4��R�]r䴁��y峥���U$5E95�n1f�[e�El�?֫���д)g}�͖�}g�'b�W`��K�З�b!��43JR5H�۱��
��q5�8t�TC�+q8�`�eQY�[�:&)�9P2]�X��<t 5w��ƿ�s/��f��)��;�5�n�h��t @���mȩ]�Ɲ6
�m��i�>y|�(rJ���u�I�d\:v�r���Yv�x�vYG���«�
��] ^?�Y�u����]F��v_>�(z5�Y��ݲ�-N�y�fh௛����,��e���\k�@�!{@ۓ� ��u��I������]���a7�VE��@�"��Id٧	�s��Va���K�bz H���mߥѨ�?��Y6�{z�;���0[s��� 6Z��Z���21�y��B���iV�e"� Ǩo��������]�Ыs�bu"�ܿ
J�^�� �04g���7v_k�#m�̦��k��ig1(Ԉ��i��NI.n��d�/f]�ܟ� 9g�eCt>�x��!墿��kX��m��&AE�9T�BW�D��HF)����f�x�{�hzNo�k{ a��0o�Z�(ʵͳ��a�8q)�l^�J�3-���[�,AkLf�s�o����Ķ��v�B�i�qg?�����$%*ϑ���%��HF����t��	)��Eco�b��.�K%E�c�|d7#����l;N������\\@�_���惽|?;��f�����0�R��-�|g����\fnxxʠ�2��pJY��1��ƙ�H��P��w�++@��%1���uS~����Z3Ɩ0D_ӓZEy̡�x�޾��(�}4̋�3M%�%#�6�왷6��ҘS�
/� ��,���� ��!�D���U8=W0eNDz
��~��ZG�b���/�р	k�Ը���W���'/_�Ř�y � ��:��*S����d4�+!���,{6�/�:x�-����<R�����Ա{:�p@�3U�c_���/r��O�D�q����#��F��;��x8���q-V?�j�"Y�.l!{7�B׍(.�,O|����ǎ���i55g�J�Ƒi��-
Y`B�+9���#��T{�8��� ��/�^�p�- ܞ<\)u,/�;ݙ�L5����??�y�<�Pɻ�|IC���B4����&WZ�D@_���Hٓ2�B2L-�h������N�u]ij
��)&{y��4���Z?/��y��t*ʸ3�yܗ�k5���v����� 4�h��3��o_d�QgL��n�ݰ2HZ��B{fn���Z5�VE�Hq��3 m��
O��mЗ�W��)Fu�5�����`�� .�/z�Ӂ��Ys譺*F��v6��H���g$"f����RI����(K�OΌݨu�]�����j�
��;��\����F�	�k���J� t��kP�u��ñ�Y);�@�'��J�G���Mo�v�z�~3��-׵g�}9���)��3],��ވ���@F*~C�ʏ���2n��9�n@;z�� ��A6+�۳'j�X�\�&�:x�Zpc!��FOP B�x1Z�ؔ�%S�"�7���wb�ˁ�$��ߏ����/�\����[�{�.�\�,f#�K.���w��B`3�����	s�����W�*�E`�ޜeϪɆK�f�F{�B��/H�w�&�<�n�o�<Y�9�~tT9	�5�)=b|���ߠ��w�H�Id���e}-����|���0[qΕ�֡���t ��J���$ꏕ]U�?��	�Ʉc��)y�ys�T��eo�B� �{�'c��:��Em��^
�M��S�-v��a���v�ǝׂ�}��n�aа���=<���I��npf�Ǒ?t[(���6�Q@��9�XC��-�R3�����g�r;����Vv~��"^�wcfm�S�X?)Nf�]r6�ҞLk��l���hbto:/eYZ�9�r`��זP%WXX�#Ɩ�F'Nh��ٝ��G{�A�j�c��_�͟�&��w�Vo�C���a}���N������"�#�ձgSvZr>À���U]ʽ�ï;�fǗJd��8#��'�ƿ����Ӹc'��8*���a�(����k]0iJD��@F�w˷�ձ݁O��+3�c{P���U0�4��J�B�R�j��A��.��p���E�}5 �Ž-�K�΁���;��&͔��Ə;2]���E%������a	{p"��r�	��-[c�o�o�ىI;e�ٕX�խE�l�>'�����Yr#�fA1�UU���pZ~�3 ��.��-�	��m T����g�P)�݀��i�1�_I-)T*����(�ߐ�f�wj}���	)�0�G��hC��/�C�����vt���C6�F5<�PĞ��?v��3�y;�⼕<
��R���g2̒�<Bn��H�=�X/�2{��TK�98ٔe��W
NN-G9^����ϟ�ZV;���(e-�~��J�+�t0�t�ӛ�Pr��n`&�Yc.�ҽ���QE�3���ˏ2;b�W�1`���&��<?��tx�y70)հ������N�,����lb̻ZK���ՠ\,:�9	9��pPD�i�c3��2��jM��##����ٰ����U�C�n|�ErWS�ٶ�����j���4�+:y R���'��lCK",��\?���mg�'l��3a�ЬXhK��q�5��f4��I�m�����p��7"OzW�Oy��>�-%�uc�{�E�t%ҏU�k�I�=	�sŝ�?>HT{�
�o��\��2���F��[YZ�Y�N�8S�7o���`�~|���8ǸNV?�oXz�WK�� ?�R_Hp��Ċ��3�JԂ+�Q��ڻ��}�������#�9t�X7���<��W7fn8|�3p��f>(t���
��9��?M�O�����6ۡ�FO�$�-w�C��(~5叹r����C�Բ��ٖ��0��V�!c�5Ln9�ь�&~��E�K���9�KP��Wϫ�±�03�:\գ���8l�R*UpUG�0s<��|
��v%�D�;���!D�R���[&���E?h�[\��?�yS��˭�Be��1�n��A���H٫F�4�����a���y�[���%���9����"	S�X���I�)�J��S��K�)��_��g����?u�9,�Qb�s�ǒ�%�*k�x�D��6�ٸ�����z���~2�����w� �9d.mS-�"���{b�Vu�����34a����&,ǂ)Ѐ���?�k57��?	�]1Xs<t�q�rϊݟ���/��x�6��h�;���Mm��(��>+;���r��KNN3C9�)��'�*�
lF�I�!�>����Q2qeUV��#V��+`�F�_���
���]��3w�(��|��������sNנ���l]��{d��i�BI�+w!E<:%=l��h+ROy ��\W�B�2��#��"�m��q����=#y0yEp,2ܽ�+�b�'~�.{&3�w�N�3��D���Ū����,ͣ�r�y�
'<�"����?�$�_b:�_s�q||?�C�+�yGg0�{r�.�_G��Ơk����~E���}��S^��L��i���ɾ_�\}U����p��n,�o�+^x/����ahJ�b3���F��"`������8�q�
���9��xi�PD'J��q�P$�<���FMC����"���S,��)s��Qr&���H�yx8'p�C�\"��g j\���<RH*�������!J/*���4�e���dk�ϙ;+R��H~5Ho��������:ʯ��f'�"cu$͊�w����L�G�n����#�y�5.:�>�@��:�ur94mo�W98#�'hx�M�v��v����N.,�'�7g���,�8�m$��=ợ��^ U�eO�H���z��h?��XG��2ㅘX�01���߻ocC(/�A^�X�\X��=#�?�w���(u�>{�Q̬?fٳ���A�?���>���Q7m�p)�x�!%��G
��B�SZ:������W���������4��Yg��ϫ6��ƛF׈^�p��
[ :��EG�J��\Ad�U8�~��m�ChA��-=�]�@��=zzҒ4C��̕t�M2��0����" ����_:g�,x���3�����9;�i�޳��Sˊ��;� ���q�P�q�g]b�������k��	�L�!vCp��Q���c Y�ghז�i�D8Io��V��ܴF�����j#�g̳>���q'����:9��A㟽�\f$`�>��I���NI���'l�pe<1Eh�^�[�o�x�.����침Z�!ĕbc�S湀�G�=���
臡�1����6Ww�{\�v��>���ʂ�=a�CI_W�ʽi}@�m�l�9��e�ު��W/��~Vu������t�(�.�5n�pj��[w.�}(8�u	�gɓ�r�������TZ�x�)>&H~pc��fV����`/�}Yw�k�w�r����u0�ޡ��\A0��f�.�]��/���6yS����-E�^{I�FƬoO���Ԡ��K=��hT,�~&�ץ��U߅,�+�a�m���a�z�+�eݩ��L<���s�+���j(�HZ�C�@H�Dޜ����oq������C���W�F��� �ާ��V�%][q�Y�"f��;�&F�Qy�ָn?,��� ���E6Й�6uK��)��?��-��aS����!G�D"s�����g;f!5�v�Q/�J���[���M�Y���ȻZ����J��&3R7}�B�	08�>�;m(�o0�I2�!}�{VB����|��LS�@_Űӯ�U��f#`�Ͼ���>�D��{�S��ȃ��}�,Š:�y�q�$��(����I����4���_�Ԋ�$�fӍG��_t])��*h���w�G'�z����� �)��A�R�#�g�	��naiل2t[ܪ�_Zq8�g+�_U���Ea�K�g{Tm����[g�W�;]������Yӯ���ͅ�������3T��R����T��K� BL?�$�V�K�G���FP/7�MFא�#���c��bU���?\�|��H��1_l�'��������lxg0�lӟ��l�2��+Kq,�D�X��w�u1���-Ǿ\�)���������X�5�]�AW~È��ݍ�R?]p��7�S��Zi���,UդD��NX����{"�\�t\pv-6�μ�>��n�����`6K���D��^i�9�F�y_����=j��k���_��m�������7Z/)̨�M>	�C��K��M�0A]m�<b�2|B4�!����ex]Mzn�>>c]���ah�5�0 �t��Gأ �Pa���P�3J =�%�����_-�׵Yy�W�A X+���!ho�T�Npʌ�㝰!�vL �o�+�ĥ�1P��f��� 9Y��ƹ��ȅC�O%�a|7�"�Z��Q��]D���桅��~E�tb;���|�9.k�̿�ч�ņ���~_D=��d}���a[M�L�0�z6����t���̭�������o	�p�sm����7���K��g�&MC�Kt��!+T��	jJc��T3%n~,��k�^��g!ؔ�s�T�;h�Q5w��ÿs���[sս�˾��/��Rz<��2���\�8{�nL�>��_d�U�y}t�GC�B!��k��̭�J�K�}��a�IoʦY�_��=� �������ͫ�2�U����V8
W�N���%p~>m��A���~��?#�^|7�+J�wJ��U��mBU���u.甄Q��h)3�v8ݽ����מ�UM
���}�N�䦔C�Ҝ0?�n	V�	��S�����~��Y�Тf�"�=c��S��V���a$�)��R�gc��|��w����C�k)Y�#γJW_S&�k%Y^�
)1���B��*� ����f
}��r�r���F֚�z�<,�d���oؗ�D�zV3���L��&���k��v���HBYiU�_w�(�aWt~����ҽ����ڋ	���+�FJ2�^	r3:K8f�4{BPջ��[9&���i3l%�Q���?��/���C�2;C<=�Ș�4pD�(��=�����tgW�#�����W-W�t[C�Ĭ���K�}G��F�[��>̢T��K��EĊ��2��AE����g�e�2Ӄ7^4~�_��F%�o��r�/(�q���hU��E�%ǭ� ��Gz�5��O����@�f�'���⥙"Lȯ�
b�qЂ���Sd#>�:d�B'�&�M^"h�=x�5�7�v��9C�D�L�å¦�Z��c��V��m(���|����Ao����^�|�\��(M���s�ǆ�,�����#\�{k��<�IQ��$��q��QQ��9F�}k�N@?�V������댢��Į��|IP��^��IO�u�&Iϐ����z�Vr��B� $�����W���M�^[$��vB�{1\g�?g��9�dp\��q
�3K�Dx%�%2������:4h�^����"9':"̄���k���M�Q�q�Oemv�"�&e�2p����l���We�5t�'(s��~��y�-��H�z��M��,�!'m���u��2ơ�n�R��J3���ԥ+��ʃv>�7+���n�;;LE�\*��ʮ�O����6�Rj~ї���ݗDf�܍�Q�&�4��^p�r�i�æW��'�w�7?>_*J�"O{�1�6��%�� 9AhF>W�QAv;O5�yQ}��ж\��/.gVʕ���"�������}��`$�\W�N[z�K�4Z�L���qHy�#�7A���{��ߎŬ�?Ԟ䉌o���NT�*��Yr��]C��$�ҏ�0NH�S=�#y�~>!��/���3(�Я2q�y0��p
ݶ��pw��^}�����Q0�s%�{	V>j��o���[E9o�Ы:��
��a��� /��4�������]Ik�s7�$����z����CG?Ƀ����v�V,�|X���5no7���D�a�im�ͪZ�����o|�wQ�!Y��dB��Y��~,'��#9���!���O9�#��㖽�$>�^��vП�x��h�8�$�VD���&j�y�������Ҟ[�|��٘Ģ:�Q�Ǖ��f�*������q�v�S��"��m%2�
M�b,%*�9�x�,_�� �G�����܄�xE%�3�Z=��N0��:�vCz��ts��jA0bm_�y.�u�Y]�\���7]����A�����CX��X�J����Џȉ4m��_Q��{iu�ye�;�'�~�v���{�K9�{?y��1?�/�t~S�:4�ƴ�d��q#A�����t�-
gsv/�Y���,�-{�DW��=M��YV ��:W�*䦻g����oP�q��M~��3t��-{�����طA����&����Ԭ�����?w{��]��s��Ikq��-,�o��\�Dw�Ԍ�E|��H���c��~�[�@�G�綢(�T?s�A@(�0�wgX����Aߖ�=��&u{y�2>N��{���ڮx�ǃ=�AV��lE���Zx��!_ӫ�}~�@�٥�N�W��	4�<7��5��d���4«�uo�0�-w�G`e}:��&��]�QM�C��y���㰙y��0�1ɑ�ɽ�ݩ��"�L'�?^�Hg���G����3`�&S���m�ؤ��L>��~U��_Z �n]	:\�i�s�|�HZ&'���[wQ�~^�޼Y��i��������ߎ��؆��VǾ��s<�a���w;I9tm�k�@�siRN��ۻ
�U<Y9����Bp���*���*�y���q��0��z{'��z�����E�T�����H(�Ƿ�u��}��~Z�F�`s�Nٳ/��U��=*�,�Ӓ�҄��~<��WL�G�.X"���l}W�>Ǩ%s�!�7��f���iP�k�?��x��������.[@i��z��6���H�]���<��,�x�y�����u��k��@l�E�&���q�oZ��c�uSW��X�+�Qg�`����\��3�L����j�vS<��7��>0�d��1�y�v>�,�<���v֘�^���;1q~\I����,5z��+t��K��
V�ۙL��XB�s��I�]�4��I}Y�r?���_������%�2�y��?Q�Od�=�v�K��)[�濵���I��g5�֐.X��4)�[(y㻭T(��=(}�%���Ÿ"㯏�ܩ;7�r/���)�V�2��	"�ju�}f`G^/�|��+c{�G:�,��`��G&�_�[QWǯ��}��;:�
s�{�J�S��3��s��Zm�J��mQ��%'�_VX�;���@��'��)��eF��ї<vy��tK��Q+9�xq�E��j#��]9ރ2\�J��뵛]8'�wL� ��F?ux95נue�Ǽ���e����f��/��lX���(g����@�f�J|�(K��q]ۤ���qe��3ZE�����ݰ��]����^\�Z4lW�8�赏�Uf��o���0e���j��E�ޠ��m@Ő�%�ǀ�Ti�:7���_�c��A��!�f�˩ιoSV�K#��{[��UMk�L���"������Ǚ�_����SP߾�Ln���Ȑ�7]���"�Y���s�������\y�f�f�g�]|�����������'�^�N򎷕���-|F)�i6��Zy�����'�^�q__q�T��(�����>�=� L(�^�O���j�(m˕gJ@+��
aӓ)�)q��^4���z�i5�L,����=���AA�$��b�u�#��e+�G�2h⢆���P�I��aW̺��a<�͙3����_E�q���7��Gy'2F%n����?�>��e>���r�N�6�	�E6���TC��
��ۡL����z�ۥ@�\	���?/�д%�-��8�3�o)Q�sB�:��KWFؤ�t�UL v~��H�A�?\�0�+��%W��>�;���Nh��[�`O�Q����..t��9x���]��
^|/Z�K�1�c;?��̙�5{�-�{f)<�V��Fw�t���f�O�e���WW~�\G�D杭���tT��|��v{��1v�3����2<��PØK�	V�!�z9�,�����t��7L:큾���g�K�� �� 4Ӷ�v�.���_r$�b�r���|>�)4�ݕ��;�Zv7���-=������F�vhUĻ��-�Q��>�f
3���TT�%g&��/��R�V�[Km2����%�v��&�l�a}_��n0�H��c�!�y��]M��.�`۴"%h�T��H���a��׵Kqo���A��Ӑe��7r�)������0׽�&�m������m��I��l+�����Փ�LSY�� �<�9�{�h�����y$n��z
�TOv��ݶ;�N�J׺�D�Q4:�U��x5�������P�%���o�vz���q���@����zl��!M�/g>��d��v�BAI�c*@s�����/��E�EBS��#eD�#c�K8����6�w�����*����i��?��������,��7Gԕ�O(%��~:���kx)KS��맼�:6��!�1 N%���ZS�#%P��EY��t��Ƕ0�aOP�kq�͹-r��\>�����5��]TRo̻-->f���~����x�}�U� �L�}�΅W�9� �i��7V:ٓ�Z�8;~�3�������N�@��fNTP���:���AȄ��fI��,�D�i/z�F
u�=b�N���TJ��)���޽���C+�C ��˵���~����3
��#�ߢ���}_f�v��w|A��m�E��7� ~6����o'��L��0i}K羪Îe3 jr(����+�|����N"�1
�F���N�����{~����Y������&F:��r��{�H�=�,&�l4�D�Ɓ!uE9;Lx6I��u��΅��w独?[ցe���
�nǶ��g>��%�;���c�����"**� ��#=��y���AT�sY���-ᕗ4+���z��J4!ԧ9!�u�j
���nwا��Z�U�����_l���'��إ9S�񷲔�R��sρ*e�s��b�k��wтb�k힖�q�kjr�9�4�}�E�E������(7�O��x�?��?Sd���P�4��Цx웴?&�{{�x��c��B(�a�	+<�Jc����.���g�k��
2����ڞ��9�nd]��~*�j�5:���vz-��~m��2�N
����\X���1��k����b���Zmy�ٴ��UX��R�k��iRݍc��JW��Hߡ�9�cK,���o�������r��倯�_�ViY�>Ú��Ѹ�3�;���I�"�/��[KYi�X��4��[��7�*�װ��vh�b}����`��A�2���u���y�����ՑY���;o���_{_5T%]��a��"����Ջ��|��
�	N�W߫	��� 'Xd}?W��r�4����s�� ov�d:�{�Yej�J5?3��cMp�Jݎ��t��B�$�N����b���J�Ӛ��?��2��tR�/kϪD:�����p�).���4՟k(taSһ��)R�ODe�-���9�������}��0M�D�d��؆��i�ah�ff�gGŧ��n���{W	ފ��~j�ެ1�x9��RM�>\���M�z(F'�}X«Xi��E�%P=�?&>SlYw� H�I�j[x��Ȝ�̕ꦱo�q��9���65��QCB*�����T���]2�����i����zG�
��>�
��0�C�]Q�#�r��v!��d(F�w��X�uE�ue�S�j�~	wn�:���FO��epJ�E��q(�b��� ~���#�](V�̟0u����`�?���m����Ԕ��`Q��A>�M��3	�E���Yr#�n-B5̸���)pe|x��h��Ҥ(H��ht�|�;C��Ea����4�P���P��PЭ�洵��K���6T�Q�j��-���J'M's�w%����n�hJ���џ:���j��eu1y��)h�2��M�U�E>��4��B�z|����{��vG����N=;Ct����@͇k?8�I����x/,q��i�9<���L�	/���~��*���TvE�T����U>��2�P��2j�aM�4>"���
w�YÞ��!�M�Z��"��|��[me|�&�[᣻=��/�M��ݣkh8z-.Ӎћ��?��}l�f�}Y��x�}2�B�Y|�T��Y�W�g1�"�89�t�2<;�+�u�^�`��9�1"LP�V�*�gO�����I����𷞎{E�R����v�ˡe�k������s�mY^n`~�V$����bC����ͬ��6��dM��H��������������r��-6z>M#��Qr��F�Qd������J�g�Ҧ��s�K��^�Ұ��J�<s�h�^R�o$�,���ө����4�k��a�*�����[�b��~���b�˟g��*�`X������� 󏒂Ф�^�w�z&���c�Q�LG��$��{Ĵ�S��z@'hf	�[{4,�	C96��3MO��vQ�Bs� l쬿F�0w�lH`�4D�4�㏉F��Q%�G��ٳ$<6�Eq��ХtPmL�����r�V�Pd��N�.�¤'eVhx]�:�oVBC
�l�2�y�+&�g{o��tv_�jsv0֊N�B���$Hl�t��jē��U.rZP-iv٣'2V8f-$�+�����FQ�f�9��jDA�f$����T�w�<�*�X��9��9E~��J\O���J!�����/�2u�Q������Ӳ���}jD)�������|+�+����Y j@B��	���YT�ݸ��6��tI���hB]��s�#N�V�&S+�~��*�!af����q=Hk\R�Յ3�������'�љ�� �/ݮ��;�ׇ�����AK1�f�R�	Ǒ�WO�E
��7OE1�v��&<�{�^����6�'GN+�0��t�^����[~+Eփ��K��~��:�����D[y���j�d~�Q88���i�=6����;i{*�����A����Pm�N����U���IJ�6��*��+S�g�#)ώR���{�(�(�.�@��eڴ�3��hJ4���l��V��du��%|��薱��Db� �������C���_BOm�?�x\�v��"ᶓq��όM������E��u�����cX������[��M�8��l9Oo��Hi���T��D�)��	&�
p�h}E]�j��F���/bld�]̵T���;��%Xú���N��6���`vû6D�Z�ⶵ#�&r�/��V�D���	�5cSg�n�*����+J�J�wQ����q6В��{�]�ö���5]��fl�/�]J���5��p��i3��m���~iMk��s+��C�ƪW���\�>{�i�V{t�U+H���<
p'c�	N�}��0[�;���H��~�"6& �
����0��<e�< Fbu5w)����[w���
����uB�ic@��,�|�!��5��uJo��t�J�fUD�ܮ[�b�Z��MCB�٧�e[͕w_?��l��p�f9��pr�70gi�:�[�<\䏦��s[�	 s�}$�������{������J��^(����~��Z�R���o*}�V:S�H�7}��-�Y����>>���A@���y �r���~)�r�{L�IG����L����K�+9;��AT��CkWw#��f���\�]	]�J�n�c\���}6�{aȩ�`����!��;b�T����@I	�3LW&�ϰ,��w4��٩1����������i�s��e���a����|S3(��Y"��*�n+�틭-���N&��J�ŝ���s�����Jۺ�:�YnK:Y��;+k2Yx#V}�'J*n[��t(���:��^lK�cK���S�9ٮ�f��(�}Sw�
t��k���M��Y8�㧠n�5�������g��[Y�!�뱜���b;e;d�#h�_]�9�mm��4��c�QS�� ��ݕ�����)�r	��6uu�!o5M��ޘ+țӷl�-��"�8?c�3s�:�M�H���ﻣI��c�e��A����~I�����_�Vg�`����]�3뮴���f�r�
%�0;���Ub�{cz�R��3�L���P�\� .n�	e^��& ���������o�ۆ�س�c�y�@1�UY�����������n���Ŵrs2����_���'�����Q#�p������f�[)(�sͩE�S^��&�����Ҡ���l$�B
��/����s!��V_W ���������bk�M��:���6
g�.�`��#���8����n,��x�&�{��/�
  �����#6�m"�*e�"9�m��O�|o�l��P�^�)�k���D�$R���)r�[�I,-��'�מ2xw����j�A^�}N-�Qa�=P�0�t	�d��������g0F��c��c�*�5M|*?����5w!Ř���w��x��{Q�q��K�Na���}����k���V����}�𰬛�zU؜^7Ve����O�ͼ���%�C�$���{}���#��&�;+^y2�xtb"ywW9�v��O��O��!{����	��~ڬ�/���/�����m���9�Ic����Х{���S�=�����Te��V��V�λ:��C[:�b%f#`�7��a%��Z	����ѹ�D<Y�(Y�
��M���; 9w�7C|#�{�-R������[ڴ��0�b;�偬ρ�
eN�h8	M�g��OGj}X���j��L^Ϭ��rK�g,s�p���w$7m��v	���J�_u��coD	5���O�d>��Q�S汹�>;&���I����}͝��*b9sɀ�}��~��$��F��^Z�Z�lE��X�64��)!�%5����+Qڏ����O����~w�L��=0��k��Y�yD܀�;5��-���
��cJ�j3(��o��ɐ���wk�Ȃ|!1��l_g�ϧ����}�T�rgF�4��lVS/qcg���+���X7�J�υ��g�օ>~�-%i�Ҳ�kϾ��~%B��!�	�B�����F�JrQ�'��7ɸ������tB������i)'��}���X�=�L����j��V���: �Q�I�5�q�{�'��������*���X�+k��ɬ��y�)�T�# :݌�� _���I ��Yͦ���>�&:Gw����_�k���6J :rm�����,+zo�S��.h���!�ԛ��
ƚo0�bg�^i�)�� 5�k�0�S���5\������b�������rcQּ����1=i� ��m�����n����-)?�q�4��F��'AuJ/�!�f�|R���o�X��7�m��^�J8��~��7z�_�Q�0i��?���[G%��j��z�Z�r=���z)�f�s������4��q1"$�,�5	o�VEN1dO�����@4}�e|��~�q�4���x�,.�>��J�K~[co�P��b%~1����� _^�u44�?�=ǹ���_��0zb��go�a����/|���Z?�{Y� f�^Ċנ(���s��Eύ�O���E�=EZ󩏗�J�Y��!�	Q)�']e�8�N�!w�^X��i��u��:V�S�F�G��3O�c��C�vJT�����Ll��۝�े�5���j>r���Hw;y�+��/��8�-\��E�CWYi7�#`^��(�8�%��}��{�a�n�q�X�7�����'���ؓ����dU?�ӓ=��y1�.�j~�^��%xu�Çz|{�D[x�P���k��x�nNڶ��[)����1��P�z1���6B_w��!��[N����T<V�ќ���X�G��Ɗؚ6y$�c@�����wm��ɦ�O_����=�.F��N�y�g!�{�L��<!�O�[��)~vn"{�x�{��������'���Z�O/��F���^�1ђbW��1�I��غ�x}��d���~]8�q�ܩ��;�aiz��ZY���urr���-A�-X]���Ig�Oz>�J�e�8�q͛"���d,�!CZ��1��Y����|�S��Ϋ
���YV��~�^�pJ.ӿ��%�����)8�Y�Sa�[<�"y@�c�QC��7b��	�qW;q��i5�س�W��� ���u*P^N`��s�Fs�6�>#\w-v�Tڂ3���z�:!�}���f&<4�s�G�c',<=��f�v�~���J���Z��$�]�����s�����l,�zH��b^\fP��Z�q8l��x"ۖu�ɯ�oU(W�bf�:H�T,��e&c�n�uJ�ɢ�x��
܉�w�K�<�\�D,���Mdٲ�r�� C���� ��s?7ݚ�X,����]�*����
�c��;��;M���!j�u�����)Ǟ������ڶAI�qGp�Or�<4�����e�Q�R��v�e]���WG�=�����琑�o2����mٓ/\��A4��D-��y��w�.�UuuXt��K�Y_��ɇ;I��u|���?Yu�z�X4�i��n�PN-�^iw���!�c���,R�2���،��a+�%���c��^���1e��Ѷ�eGN<}��br��Z����\��;E�{�ъ$ӕG���"�S��E�-������G,����17ç`�NS0wi�W�429g51Qw���϶7�zRf�� ����0��v�P/�ލP��h�"^z�Izd%`�r'i5K��~p(�����PN�9���ޅǓ�m�*����阬�t�%] գhݘX���:�������󫊄 �ؽ��س߿5����D�:�4��Ze*��]���8�c�}]G^���J��x�B�uJP<��/4e�¦S�@!� �Y������G:�
�ou��3hE2�}cj��)j��sd�ֶ;�2YB�Bh��;)�l�qv���{(���VD���q%��oV"hh�!���[P7B����@��UP^[�G>�eJ-��11�#�!PKM^:�?�d��tT�!#`���/�r����7r����e��p�ɾ�� k]��Lj�XN����c�8�d>P��4�Ε��܋{���bc�}�J�u%������{?~<Q�?��$�sq�rs��>6�n�V�~9vJ�y��/MD�Yt���*��nz��R\�*JZ���L��9O����x�ء Ld:����	z$y.,�	\x	K�RB�$\lY�ɪ֊`�:j�L9>b�6�&I��� � fe��U YuV���"7a��܁YJ-�X��6����['kdc��q��_��CW:��7�q>)݂�3,a��m"`A5'QGg ��U����E+�=�^CD��%� B�FF�FM� Q� �D1�(�{�2�����{&����χ�����{��^k����&���̝����D�wJ�*��G=��ƚ�)%y�L����h�&��MKV�I0�acƻ�Ԧ��~P4H�Px�Iww+�(QViM��u�O�[�ަ���;����&�<�ehz�Z���}|�@���J������c
>�b8�Vl�&̜ɚ�5/����a���à���f9�ώ���7E���?�k�*�xF���X|�:J�����ן�*�~ndFt�o�u�<H�}��nNn��U�w��5*F9�=z��z���50W��lJJ�4���C۝�M�m������^�� )�M�~�����\�ۦ1�UZu���N
s4$CgC9�3��M�虼�ɔL�#�o#$�{.�kBwCĠJ��^d�z�h/`x�y��5&�3Z�Ƴ�g��^:�\�y�Si��81�t�����t�h��.�,ވ�dy~��/W���@�Bq�F��E�6��/2>�͏�k����L��ZQ�4���@u���D^-�M�;�M�VՑ9x4S��7���
��t��ϽX��;jRQ���~k�S@~��8����SqIVzc[z��S�p���D���I�wΫ���R2z�e"�N��w���U����9�	U<�u�?�j�չ?� �X�9�3��%�	"U/���E_tQ��,R�U�^�'K��nI�k�����s��7Mk�ctn����`�8%������*0���%G]��;�U?&;+��&H���^�(��!b�{:���)�#�h�G���a�D�(kn�{����<>:����g��`q�4X��� �i�}@��k�
]_�PRK�u2�����s���&�e�u{�)�V�'}�mQa���C�*�(��:��f4`T&�A�7����!���)�s}�)u������p�䵶�';���0Z�a
��tV-S�K@�k�;�_�d���%4�"��[sv,+-k���ԭ��8��W�r��ь��H��v�aޚ^��#�-=�D��§�)&�ˌ�f�I��WQ�I��ɚ��h�~X�Ov����N7%�o��������??�������E�*�Y�ﯦ!�z�V��^���P��cY�@7M�(���j6���H�@|��u��2ì'��\
��Ƶ�o�02��f�$�T��ƶ����}_�[Q�x���~���N�᳓�O�;����i�PT��UZdZ�΀I�|���(ngH�z`� �>�
�M@�%`\�T�Ս�>
�W{��2B����^��7ފ�i�n�ɚ}�}Hm���}�=c�Hm6z�)�>��@���V�!j���)媊�Ŏ%�J��S�V�P� �сTm������i�s�ɭDթ2	�^����IHME����³�%�dH��gD���y+��V��*�&W��kϛ��yT��9�~X�4P����6{��fL�7��t�m�%6�95�@y[�^
�:L��/�C�����#s:�S�HN@�����B��yƪ52(��xh�t��7����Ҧ�|������>�`�{q�4�gX�"*L�|��@�6e��_�aѣ�T�T��'��x�7!��q6�ǡGv]i�XO���K}�c�V�{W�A�%z��[���o�JK��.@����ʱl ��R��=mz.���`}�k�*�nS�W!=f1����7�cv�5�)	r�V��/��<5�M�9R!�9�h���h����5po����8N��#�bZ�o`.�Ǘ���}襱6g���Pj�ց�>���	���;����<����N{{���T&~(ʫ�ѯ,2C�lpF���49�����Q,�X��Q֎	ǩ�4��^�K�=��
�W�h�*p�ϛz�����|i�M#�n�.F0����i��������X�<ӧ�~g,���O�)ƍ�m�iz����H?Gf���ɲR��j�ö�ߢ�?��ϙQ9r�n���:n�Z�;ëN�v�m��}x������_�F�ΰ��E9�䢤�~�l�ʺ]�?�|��ޜ:�c���7������1[�TH�0�7}4w�3ǆm���H���/v�,�V��v
�?��@�5��l>���\
?/��C�q��ö91F���52��3si�m��xS�Ў/0�����L|�V�x��p=�[��-����u_I�J!��\}�<��20��7o��L�;(*���t����r����m�5��9��Tn�)�<��;���17�������Ֆ�N�(�D�
�,�t�;�Y�^T���/Ɗ^�K_ELw�t7��>�����-����>����P��b�/�o����������r�:�A���bҽI�ߡ�}C��d(4�� ��!⽯��zZM�1��)q�����Y�o��v���+9T��D
{������,MJ��t���9�P�Z�,�bU�q�44U�$@0屇�Ԡʂ߇ r���R�r�{	ɍm �W���g]A��F��@8�l�zolE]�z+��C覎�LR��v1땹��FϻLP��;ݧӛ����P��
c%��YE�=J�zK�˛n�g��yZ����*����V�z��n�<ڈ8R��p?P�85V��uɦ��wBo������[O��_�X�4�`_��Kr�:��Ɵ�1����ӭ�ow��P~���in�+cX~���v��\&�͆, MwX�Z���Zy>/��e	$M�����:��N�; 3��)V��A�?N��WGM�b����q1{��#���`x7�Ńtf�a@�:O��mh���^Y}��"U��RV��iL.�_��5�S��������-.*Ldk ��;�b_������Y^ߋ�1N��
��ʳ�� �����e��/������<�bkkk��o�E���\��g�~�?�D�*���F9���s�.ƭ̺,pAO]N�,"�IىC��s0!��p�+��X�2�Z�Q˲h8�3�
�����WII��^���j��D��
�D��\4ZR_<�RR�H$J��p�g5]�)���Yh񼟭%]��%��8rw���:�Y�2����o�)j'��o���<6U��ͫ"��/v� =�~�V/�{�&������^�l5�~b�ؾiȟ���M=�w2�v-Z��*?��$��W�'om��e.H�N�]Ww�J�,ڣ���<�^���#�7E|�mME;����"������/��°o'VW����y��nJ^��̶]�i���X����\� ��e�'�K5��g�=V�5���J����������c	%��Q�e%_Ѐ��[W�P꫚�OR+��F�2�ţ2�j��l����T���K\��E'��)I��Z����T-h���gu[n^=�c�U�G��祺\�����PR�s��E�ξklxPl��鷽j
"�f�>����w5��B;4���"�z��w�v�a���Gd,�\�f*��B�'J[ge����S�^����^=SG�$����������Hw�D��r�
^����*�B�����qz�=�'us30! �ς������v�Jb�N`@�Q9k�9k_pn,�G���~U?�]]eG0(BڥT�a�S*�|?���TI[�X��#��a[��^U*�o�WW]V�������Kb��8c�N_V�B��j\H�Bb4R��c;-zӎ���8��U�Ŝ�,$���O���'oqw�1��z�NI��EM������2�S�F�Ѩ��R�Ţ�ڒ[���s�a�pK��� c�a}f�@@�u��$px�P��Q[�Q�9û����zeff� Ī��1��_���Ω(
d|x�3L���2��O��4I�:q���5���N��6��ym@wOV߽u�	g�1+�C4�:N2#���p�۔�G�aA�C#Vi�F%�����
e3;�9lX����|��`W1rJfPw<� �L�Mbw�3d�:�8w��C1�~ҿ��_cO�\�+��9b@�a�͞�҉��Yв�/��ؖ��td�O��^ת�e��L�0	�I�	�
F��{��C�H�nG����][m'GyݹI����^���ru��}j��_��ѩm�c��w��v�w�^yd�K�f�j�w�sO�Ы����������w>v�\"e�|��7��m�&�����7C+��Ss��~
���� ���������)��$�g���6��GY_p��xr�������퍅���0�b�N����~����3B�K�Sr�D��h+�Y+ �(H�>8�
6I��0E����q��!�!�w�5�σ
W���~��Oд_��?i_�z8<9���!�%�ɏ�s���S��6%A�;ga�zQ���'��NT�ԉ�S�Z�B�E``a����1�Eer�="���7S=8�C�.��ǣ'�t�|��`/֘w�2�3Zi�p�F��"����D�֯.�}Q�X��ۇ���d��f�8�K��򆷐î6��]]Crc�͋���,�pw��K�_S����$�H�J1�qx��С�ņ��I[B��A)�<���#��Ы�Qq�jN�>e���3���Zh�/Bo�֏O.�+V7R��+W���kX���?�:�$��,�u3����Xų����GeS+i�/s�Zc;M[���{��pS�R��"���kSb���eb��|��$:�4o�ݗ���TwTƧn�2ݧ� �3��|�勋�R�,Gv�ܳNJ��5^�Qu����O���˒���ǟ��纎�b���,��%�L��xށR֤��[�iq}���+�U�F�L��Ǟ�z}��١Q��9��x���@�7�ᖋ���R�&��O���+�`���o���{Í�}MlIk7�eo���W���3=�>l��j�R����$���ࠛ.�ݣQ���$=�H��͖qw��$��ҝ�{v��̅O��WYWON��'ҭ(5Ik�;� _�޻ݮ���^��&�N�J94���(�*�֧2����A���g���K�|΋h����R�a�L@ٳF���[꘸�~��!m���e� ��@���_,�@N�g�Y�@ϻJa�	\�<E?\^��Ն��Sٓ��y�H>�{���Kl�g�ύs>�j�h�>4����b��q#L�����!��g}}^=om��G�^�����J���x!��Rx/N�x3薛��?�~�u�q+Κ��&<�p���^2�K�4��`�\��q���;oh����xh��~_��nߏQ�N6x�F]>���d���0TCc!k$1#L���4,n˺��(��7z�i�>�8��_0�x3����o���?ʹ��IՕ*�O
^�5��C^��S�=��Z�g�����,HU��p�%Ds#S��r�i��4e'$J�σ��M=s" ��N���]�����/��n54���Ywj������-~jY�b�G*��k����8&,��7t�Ѱ���U�07m�DH��`ǫW���x����O�c~(�)�)$��#�E=�<�����dny����*��t���W=&�n,��;���m�K��J��]��P�c�FSj��x�Nfq���q�<�PLcԫ.��:T�{���y�阂�}G�f��.ˣ:�uxrb��:�SK��.*����1]�!���Gl�/-�Ɉ����Է���4_=}�x���k��ׇ�������>~ ~ֳ�K�J��pw��|PS�t�7|[%z�%tU���_���Cj��1�۵�Q��*������V��x�"�~�H�^z�T	&b�-�qe�����ۛ�O��︃i8}�>m':lh�Z���Ѫ\��#�7{���_#?6~�i�Y5�|w���?OA�ߍ�ٝ�� �����z�v�Cy#�������d����G�D�hm1*�_'iy���fn%�
����~����RG�����������b��d[pYG�'��"D��̚P��l��r�à5�j�@m
b='�Mњq:�x2�������6N�/Y�d�8�eQL�3m��_J�h�����u�9��1�An�/�"z׆]�ܨdS�b�����+�Y�/'�Z���~�2�3�OFX�%_lÆv�B5j)n��`Q���9��*��C��*����ƹۻ��o��_}�T��w�u����Y =�g1�7&z�k�Y��LԶ�P_�T�\g�cHAګ�����CL����I&. 4�+�-l�	�C����;;]�s[��m�/;\�{LyMV[L�1�х��Ҹ�H@���7*��f���Ύ�^G�-F̠�O�l=��y�CهV<C/�����_@�_��d�M����`�J�F,-`������v���fT,w�k:v�]�z�Yn]}#;�U�A��V���*�罡�R4��`�[]U'����1wLf�y�,�~Sj�d��r�D�	Uv�;�틑�����Ǝ�	���cW�<����!��r;O�v���������ͅ�t_�9�D� ���x:%M`��"�� �鹺13+�LW���VE�I=�R�����tw���M]mގ\��>�g���uI�Pؙo`���.b�� @�F���.(I�C~H9#�����;ث6��k�y��,ZInIu;��F��{w��#O{4��e3�"~�'�6���.;���V���6����C���oGgp����8�v&�y�<sv.��d����h���7��Z�^H�I��i�0�����|�Y��SS��֭��%��D��0go�(�h�mp"n�)C�;��gq��9޲����c`ǵ�3��
��I�Rn����3}��>��>@?TY����a�
�z�v�ŝ�'�� ܲ�r��_�	DY��6A��%ϟ��׹2�3v��qj�}�6����������Y8x
5��D�>0B
	`�����Z��"{��胁B��9�P��󉚜�ҁ�k���MnD��<8���:f���8
.c��^��:߾1�BɡC�H�J{4�=urN������W���4^���:C��3�Ѹ�1音|��,"Me~���ᢛf�?<;�1�LJB�����78��]/�b�\-9���Ͻ=w11/r��ҏBx/[{�_>{�S+ô�=5��VB��=f�g��z�,��ܙ!0P�&���I�
�t�dE�yh� H7��3�WPĄ:�z<�qХY>�'u�I�v1�/. 3���{��r����d�f�%f����n!�Ĵ���y-v���ot�tD%=(^���Q�ݳ����@*K����o�����\(�QjY�Q��V~�t6c3^'��#$Ww�F���7�Mﶴ�Ӭ9Ffgc�Β��$qXD nh�����4v��� �o�b�캊�ץ��L?�)	���Kÿ�|.�߻�h�m}:z�p·�S����}�4C\�q(����w�U�5dV�<�F9kؒ/��il��~Ӈ3J>��m� �E5g?
�K Cw��5d�X%�������2	�����0E��|[-c��Z`�?���1�8�2����u�W�{j/2�[.���ʁIUė�F^�����*�!H�(J���ˮR�>��f���0KO�Ң��D��-��6��=�fKR�0�w�&ˬ�����;M���^sn���Nk���h#F6�o�w��k�rU�鶘F����e5{��Yѿ!�5����>L�Ԍ뵆�s��<J�@)��)���Fe8_�}������������~�f���O�d'�,������Ɲ ����˘�b�˝G?�)�y��_��t�J�nT�s����W�
5��J�7G�:��p\X%ޯʗ�|��v�ˌ\/��="#L@A��������I'B�[j�)�0�x���Mu��(�}fh�dH�����ճ�)���ȝc��b��嗗�2�@r�~�a� nM���8��0w���n����r��9�)GG3�0}��ɏ��.|Q��`Wa�Jm�( ���	7V���h�r���K?�0��侜2���j�HΝ�7��Ư`�h�j��P�0��9AZB���rR�K�䐷*�US�~���|O��/��pU���FT4�9Ŧ�P�BL���5�l�{����ҳ�p]�	��n�ʒ_��N(%j������l�;�?�_>���&��ͽ�nx8.{t���.A��q��m�HdրZ���,9{�yrʐ�"�ɨ��	�L�l�a��-SF	����p��!�㊪o$����7���a�E��NR��,��B~�����;D�> o;N�(�۔� ��k����]�n/�
CkX�.$�]x��U{�Q�_O�y��9���h��0X,�Z5Z������;��U�?����yG�*�,����d���gF�@�VVB���f�ym�g2|�<X"���[�#���D��R�]������&�z�O�z�:��`��Pw�׏�z�?�$�, �����kۓ�ma���0�3��k%�bF�E�(�er�gv[�$u�ۦAy]߫avO	a��m�]ZK�ky����7U�R�1�h�K�UTV��������k�#�C�Gq����5�� lA~��ks@)nsՕb3�p���8����������p�����5��Iw?��0٥#��@洅D�Z��c�����ӈ0�V9���΁�@�ߺZ�\D�=�������1P��MIz��{��'��9�x�tҩa?��ۥa��S�ž+�rʣ����H��S�Tr�f���qP^�3ɏ~qţr��C�\�l��(�3* Ҳ@�Q���t�LXj�;H譟��cc�q`�s��x3�U�m6_o����J>k���RD�Ĭ�|�[m�w�-b2���I�o�-�hg���>�yկ'�TB��%��W�lw[O1{,~��y��\!���� hbݪ�WPJL� ��K�ڀ3Vپ���R�/��6�M���p��<ڀ�g��<�C�����ն�Cnv�%��k& O�khqXY��� <�'{��˓�i��8٧즌2��߼�^�(Ơ����"�o�&���l������Z�\X�BCƸ��3��&VP�-�!���WoU���.3ɅXN�y�M%*ՠ�o<"Aޟ����,]!ȧMQOS5��ȳA5��8q����UUc �����;���e��j���d�	��7�")�Sb��?����֑Z�s?�=P�N�#�2��)5>�������aI���F�Ib�s��t�*Jr��n�!�P���^<���M
N�=����۟�6�4�RBL��Ef�y�Z�x/�o��L��3F*�:5_y�Y�t��A�.�	*�Z�Jo��\Γ�67�'�H;�u�w$@�M)���JP�D�������<Mat�?�_��0^#,�É0mGOC>�n�3�n�W�3��o� T��[Gmjſ�sUʇ�xks7�8/Ԧ�U�����I����������<'%���_�I届ij���}�t(��Փ�)}��e��f}jy33&��l�3����Gܐ _i~���b4Rt��F���Gc샼�[BR�v1���-�O��QcѨ�-��6�u�%x^��w��տʣM�U�����o%���N��;�����Q�ڹA	nzm31I˥�o���fJ�<��y�K{��#uu>�ɦ%_�_���N9wl#a I�Ҥ��H���d�5T0��@쉕��^߬���5����i���6�D��lu��I��hS��A��)� ,;^�~�{3�ЎO|P�ǆ���( 7t�N��� ����T�x�q���Gf���x�(_���%�J@���b�U3���� ���G��9L]!���E��Uo��-����s��J��_�Ï2��+�p/��;Y"���٦�j0%'���`s��xw)���,Q)��֛P��Z/�豯�̢���e�z�@Z/X�bߦb�]6E�t�c�M�j$�=��Xiܓ<�R�M�{�ak7�x����5���d�-����zO���(x��X�o��1�l��O�R`&ݕ|�*�z��+ȝ�]^��*@����{�̧�����e��5��~�H�q#I��a����*�\Ed�SP��f�p#�5*MH���J�h��4u�C*V��|�&�N���$��dd||��ӟx�������g��2;;`���V$jOn6��_�ƾ-X ��11S���[!-9G�\?�#�y����i�Ɣ�wP]!����'zo�]�����An�>d�ߍrT�~%�����`L�c��Ph7���06�I_P��f:h(���M����eP�΋�
895E���"�G�8E��H%�T��'��;>]�.� gv��l]喞�����>y�v�D����vV�#O�'XUՌ���^5a�h��1Q>o�3웯^��q] ��= o�˓�(��7�)(Fnhǂ5L�-��>��:\[������	������"��`GX��F�����C��VM���]�
VV9L�I?�M�u�b����i�����=I�1�ПJ2�d�͚gw�Ԟ��F.�-�x�qK�N��nE�O�К�.��~�o��vɋ<+��_R��rU�����E(tL�l앾~T�����C*�*d 8��Ch������O��]�Xf3��5��W2XO�����_F���.�nTC�|n^==`Ԩe&�#ii�wh���Bܬ�v��Yu߭���O��sN4�����h)�Â ��=�%{��!�O�x]��B�� ��mn����U�wH�!�5��ܔ��$�X�x���Q�fV�5�V0��W��
v0K�=�6?�ٜ-�q�(B��l�B����,�R���7:��v����T�H%Q(��R��0�	�|hk����tk��j�:�d�5M�b�~e9�,���8�8��]�%���4b�ޚ��3xA�;1�t��E�^����e�_ =VgRz6���� �Дi��I�r�w'�8�w���D�d��Rɀӗ��J}�Jp�8���J�=]�X���q]c�x%��uW`T�G�Jv�� �i���q���*fXkƵ������Ų0M}���uc���ٮ��t���*�Y��
/��5�z�������}.�m������)N����/�|:���I�aO��:"ט߮��|Yv\���W�Gw�z5��w�S���+Ot ��d��[u��\��@;Y��tx��Ʒ�sSl�\W�;�����|͖�2G|���B��PR�oo���zlll�9�yN3-j�9Kь'"dh�mh�3���HR��D��<֩�s7��6�#�S��͏��cM'��v?��S���^�AE%W>A,��
a�<�R���6�^��*Ӽ�eO��Y!w��L�x�׫�;ְ;wLк����{��t��8�&;����(�.c���|[`�w(ĽP����EE�HH.
���ny
���xQ'Hc���kf#[xoN���S�1�󱃈���C2ҭO���&�D����6W��3�u�|����_ً��D��m\4�Y�&_��FΜ�u��nb�~��e���DO��W��_�G��k�IzF�7�{I����JM����Z>��F{��C�U�5^�����?*.���hݡ�URR�eo	�-G�*, ;k3��Q��(���j�Q��S�ta�z����D@�m�����"=�b�ѓ�f��S%���\1��1�,�q�.�-����jH|���ꪄ� �j^�W�g[�u�x�Y48��
���[�l5Vj�����ފ}��-M���]�L1ٰ�擡O(��m�w|G�Ff_r�'���o{Y��6b�00Iʫ�NNF] ��#�G1�/ƂU=�,<��$�1
�:{F�n��fyQ����WDd�,��i��}6U��D��΢'Y�X�d�K�|��19V�֕o��VDщ�:=��%
e��9�8_knZ5k6&h*.&nI��H]y�8'���7 ���O����h��ŋ���O�}#|�6�A����ǀnY~t�E�/I{�K t�i@)��L8&������M�߶@���ޛ�9C�Y���x��#W�7�)��\�i�qj���-	��o��Y�7Mֶ6�q��ƲD������0ܡ��cO7�*��1	V˥�w�K��j��Z��0�ޔe,Z ���� {�^��6�FJ��I��ɜYl�
7����ok��)����p��>]��{��syTΓG�k8�^q����Yi���:7�d~��:�����ڟ��R�HI�o�wW�uo)���j+�r���*
� ���EJ�Z�4�+����>��y͖�y��mSB��{���>#
E-�[��8JH�x�U{���m �Can.v���	���)y�n5�);�����zY��Q�	�k+�[p����Ǔ���D@
�����Nem)5ad�LY��	7�*�.%�xa������e�ݠ��E��Ek�[�D���ԻSRN�pS����Ɍ,�qv�)h� �,O9W
��!�s��n����U��/m���m��	Y&m���Ť\0�?�z�'��"!N;8R�Y���s�!?X�[`39070L&]�G9�-H!j�=�n�S$~�n�^���Gg;m�WO�A�}P���z��d�W\p�/��m�Lc��umꌗ��<�!��fX�`�����
OM��(�Ռ��L���V�!�l��+����/�A�0�n�jzu�#�'�"3��<U�OB��U���*:D��ϛ2�c``@#��}U�9�=p����Q��:%=`clN�w�0Hn<�~ qBJ��"��kՎG%w����K�mE`a"��͐�㆛3�E�Ѥ�:���l����R��+{�3�I1��.���)ӑ<��P���Q7g�7_�x�q��[�re\*����c_7��
(���M���q_�B8ߐ�D�a�tĤ���v��f�E��n�KѤ8�m/����+��y�d�$��=��)�@��w~��b�l<�5ZW��v�\8�,�jy�� I�9w���7y�k�j�O-W<x}��;|�!��e%>Ɠ���:ш�,SWl��ݞ��S�ǚ��:5zx��_�

w�|���JWo`Y��p�5�E+@it�k��q#2���9X�U���S���+[�oZ�~� ��Ksp�3C#�-��-�N��]wf��X����R&b�M}0�5ވ�T���w.�\M�����8;�O>P��0Y�1�!�z��xi�B��U��[�{�QO�K�_F7��$L����%��2+��
����T�η���K���<��heԆw���΅����7��/�o�	Ҳu�Lh���ͭDW`O�#��%&P��Re��! ��%pp^0Ĉ3/A��]��p��M�{�!U7���O��1%���BggM��O��JDm?)^JUΨG�"�(�g�J\D���:��#ݦ'������>mt.��yZ��9R�uU�49|���lN�2�!T�������va,y93�r��;<���#�e�� ]�� �����S��lE*�:g
M�u�W�Vvz�jA˽:��(�r�Pm��a��jh"(%C3�m� ��v�ҝM��y���H���z�Ѹ�0����)�+��,Y冊�+?�yB��:z&�+L�؏�a��-+��!�������̑���ᱱw�;�C��<T��H:���۳o�Meu�*�OD=h^?ư��6���~�N4��?>���g���{�E���
�Zϔ�^-Y�|Asa;��K<��,M��8�z_W��Q�Ե]*Y�e2�o�R!��w�#6��ւ9�:�U'&��ŷ��Jؠ�4ژ߿��N}&,L�5����Z�H�y��FI�Bꣾ Co����[�i?.���$�����H�N][[�g�7S����%��
!��`���:�6��N� -�Ȋf�ObZ��8�kG�9VD=?�Wt{�+���9�q}-D�ҒZU��^ɔ_�
��b��U��f�o��ԛ���Hg�YV����ɾ�t���Q�zrOqYb	����^�96��7 �Ặ����K�eLMt�����K�9I^ܗ�W­���~0��Ճ��d#��1R|GG�ڋmXv17�iÚ���v�7�o�%E��������(�%�|V�-$���D�0����wEM3�����O�wtV��i�^�qGY�ɫ�:����:���T��5"Tf��ZVC��R�?r,I��3�qo�y5���۶�^ ޒ�%~I͡q�i�9�ף�ພu2�K/3"�c,�l����m{A�GQgL�R��# nBS�i|�=O��D"������rx!����s]e
r�F�a\
�Zۇ�뚶�H�*�3�y}K��Bf�R�(��s�-�X��Q��J����7f��n���'"���{
�K�ȫe[��`�`�z����P��C�Y�y�f��z_�u�c	��j:C�b-�|4�8V����'U"Zc��7�����0+�6Z�W;��;&;~Ԕ�{��Q���lb.���
\N��`�Ɋ�J�d���"���/z�|sŪ3�SS�yj�L�=�:n��b�����L��IG!0�������a��,Y�q�G���Ø!����g�����_Z��n#M�J��H����K&����z�'M�B��I+����1�����j��2q�妙#<���xݫ��ZW�W�;�&3�v�IE���I`cc�\�uU:L�5�~�86�{�j����`��;�3������a�&~���[��IY��Ϲ��?�T��}���]_f�j����IU<僜Z�*��B��'f���نG�V޻몵6.-o��' *)��j�f�8�Q�������e��aj'^���U��A)� Ą���"X*��{�+��Y�L��@��ܲo�b����	��a�A�^B��/v�:�\tϺ�/�] @u�L�z���6 �]��wZI�55�����a��:\y<�ZL�ۮ4��T�嘐|��Q#��͢�RO���c��gxnܨ����ژKGT��̶��vu,��G�>M<���G>�kó�D^�oH˱v�I%վ��-�o���V�k�q���HA3ǫi�؊��%��O����f3�U-��^g~�l�+3���0�П�+j��\&Eo�9W]v�XƎ���K	�H������H�^�=Ɛ�ۚ���g��Xa���U̯Oy1/��}�D5}����#����B�u]�u��m%�Zx�u��Ο�F鼗�>u��:�s��tx����p�����[�J�!��!�c=<Q�z`���a�.^\W��C����y�a��g'ޯf0PA��D�����v���rd�"�㌮J�k�gY݁(¼�f�X�}<F�ߘ�����L0q�Fw�ثZph+R���a���t�@�(��{܉r�X$̛����޾�F'��_�7�N�ԫ�����0�b�	�Q�����m�cK�Ep�����m|F N����z�������Z[�^�� �ICl��	�^�OC�8�M@��93����ZYWJ�\�M�9�O$�ʗ�OC���\�7�?7��`0�&� 
��,u�l���TE�,M��9��j����f��P�����# 9=6U��5�(=�{���G?0fD n�"?��e��|���p�_�����E�'L�eGY-�v���*z�yE�����.,1Y^ԣ�Ƃ&2<�o	���!^͖dh{�Y4+�L����ђ>��`j��_{����#�~]G�E�ryҜ���,�!|E^'�J�A�}�b%Wl���]�Yϊ��{�ġ|��lQ�\��.Mu5MA� ��?qe���K��mm�ޕ�lwĳ)]~x�W�򔸐D���F���1.dgDF�3�����u�s��
��4�(��~nH�<��{ү7����H�!��'F\w� m��yo0g���|zl�[hT�fO��y�7#s_Sy�D�i�Ϛ��Y�dC�Y��d"J<�+Z	4>��ȇU7A%T(u�8U`�xF�gJ��t��T9r��q.�)�#�@߮{ygҴO1�.u����J�s�b�,���*�^��m�x�L���^�_Q`���ғ>������n��*�P�_d� MB���5��尃$��-�m�\��^��˚1��G$RY"*����m��cR�r5����>�F�����������ms��(��|���YS9��{��BRQ#ToX��w���3ȶu[����T����hrF��C�����yf`���Ԝ�y�ӭ�&?0x/�$ ��,���&�������CI�Գ���FN"s�<==�|�#����~&�抋����v_R},�!U�bob&���䑼\�h@�F��v�xw�������$9�U5�v��-C+�Ku�h_Pu�ؾ��k��^يqBF�Q��tK�P�/��һ��'���|Ax49�ƛ�P;6�/c0M^i\�4��i5/ݢ携V���>����6S~+�9��/����t�2�\PGĊ7��<����F�oh����O��d��VҖ�x��cb�g��H<�p8ܠ���]{�h8S��w�.ҧ����Y����ޣ��wܲ� Ld��4޵3��)��0�O	�h������5&F.Q�Kx���.�Ў��/4nO�ԑ�[���n���v#�y��U�Gh&�Y��[�eN�1㚿������p���V�u
�lzr>;z��^��N�4%5N�����]v�B�	(��%�;<0�`�P\&Ҩ��"��DDD����%��¡�2;�y-��'峺_��<�#�W��w,�����nH20L��.@��D�Ueq�#�,\���dA��������/�?_�u�R$}|�أ��j0ʈ;�E/����j�T�c$48����E�:�ڣ��	�3�\�&���\�
[%9�Ӕ�[r����}��	ͫ8$�����t>��V�")������3�.'D���'ۆ��R����{�e #�w5F�ȏ��,߸E��=_���IQ�X�)i*����3m�I��u�Ѩ��7"!�kbu�X�5��}I*t�Ru�gy��غn��99�&���P����"Z�X�I�,ϻ�,q;bN-�/��zn����e�q?^+��[�o���^�lmA�&Q�7�w�\w�n���Y�X�C�@�� @@�?���ͮi���݊�S\JCqi���S ���V�ŵhq�ܵ8	V��]��y�极�C����ڹK~��3'�.�ee���U�B|����*���������1o7KAU�+��Q�SJ��0�g�.�?X����[	�x	^^���q�^�=�z"�
)s�q^�� j~KU��d��Y(�9/��:ܭTX��0�R�E����{�Uj|�Z�LTr�m����Nʹ�ҧ[6n�Tg6�'I�s��_BL���>`�O�o���")n�J��MMH;,}�`�̋Wk1E��EMN�,�e�J�YV���7;AB�x�V��~��==�_Nru��@#�p 1��O�f:��'}�l��TP�
�[��������$Y�I�ϒ�x�ە��A��D�"���ӗ�$UaE�����}v��O�}g«7���H��_�T��GƶZ��^ �ˤN6~��������@��ab�'q~5��D}�.�A�ĳ⮡�XB�w��@����X>�ήK����!���T������g9p:j�;K���Ӑ����g��������wpd�!�ǌ�	8}\�����_m~��(�H���[	&�;*�~ES���ߜ�ߐ�+�t��,Ѵ1o��ꑀ�d[��z��qWsۦ�6�ZYjeȋĪ�zaT�Nw"��W^{Q�Uۛx�dk�U{�<Fh�����PM��N�`��hU�d�_\Gk��(`�gy��A�R��0v6�կ����Ը�h�{tt)AX�%��ws�4�RB��QHK��JR��Y��o"�!F&5drR�v���i��+5�l��C;��/�=MA�D���q�׬"��U���=+r�P��r���2���O��p�j�W(a��3iz��	ڛ'�i^x�8n������D%J�.���)�rR��Xկ����|^���4�O��
��R��M�Дy��K}�N/A롨�ٙ�y��ll�~u��=���J)nx��A�e��?+�XA�#���v�ŮX1��y�z�������ګ����T��cQ��(u���d#	\�ՆT}�j����l�3�b���P���6��ͫOj`�F'�CP���>=��dX.��o��f,̩��&�䴵���o�W�3�_�%���B��	�s�|K/ ���g�M�y�����	�O;i�g�o��j2�c�]5@�<X׮:�66"_^!��h
j��oA�]�z=b<�92 ��nұ��z*���@,�3�#��E#�(N3�]�')�',��w�_%0�Z�>-�뭇��?T����Al�����y�Wf��4PE��G��,yt��,��H����{�ɅL����6b����udKXH�tߧ�X�=/��LOU�w �Mz���[����7��""ˁ{7��A˿b�}�^��C+��>��~���pd��8�ɫ�#����r��Gx����ڰ���a�ƴ�%.����k�%�-՚]w&<�����Iu5i�r��K���j����-�\�n{B���fӢI�F_$�<�NF��aSv7��d���N3cBK �;O�13�_mv��du���i���Pu���R��Gn�ƪ6�ƮnR#��52t5���f\b�q��9/1�o������#_��Px��s�1��������2�sv�9�2�<9MN)�z�{�M#��A�c#��]����ě�?8�V{��F�V���*_�nB������q(��]���g�6�8I�s[�Х���� �`�V��A��N۸\v2\��qZi%(/g ��Yԯz��#g����r����F����lD���[�Й�Jr-c����FC�(�OD��ԅ �2���Q����#7c>]��mo�.>C���l_vP���Se�ǭ#�O�݅�^?`���z����NQw�\�� ��:���O��Q1UG��@�te�U!Ѕ�B'oG�=O��=�9�����7;S�D;�];����������a�Pd�!K�9���m�N/"�[��ZH�'�-�S�^[�x��9������5�����b����������.+Q�7_�6^jv�
���=�-�We��ۄ�e��BM��O�2����_�`��a�*"�;^�y	�Η�f�&ݖؘ}���}V~/���g^�V���e��+�a���:�����L9�(��g.�|��#�g^,b�E�
B�'3/+ս��p�����g�����DG�5"�F��K��!�	[dՓDS�ry��x`4�J�ޫ�ax� �'mS��p�~V�>>��h"V��{_�d�POe��� ��F�HZ�{}������+����� ���s@݀j�g���U1J%��;���{;�����e�J������c�|�	f���"���9o���%�X.WqԃI}�ڇd��o�i�����b�������L���u�$T���~��q6N���JF#��7#�o�}�ȪAG�uԐPݾ��Řd]���O��#��F��<�A�h�?!�jN^��ۋ��g*o��l��熃ߩ`>Gk݌�u^F����ۃ:�����G߶����8�A���q��{�d�H܁���4����, n��U�*5V�"J�M~k�Z38\���AB���H�3�)k��3R���pe���c�2c��~y^��YVň8&�Lˍ5����H���Y	��=��ŵ�؃�V�H[\���k�����f����u��������||!��{*�{{'X�2e��

8/�i���'�D�3 r3�p�tԟ�KԲR�
Ӵ�Q��$C�&!m���Џ�<�^1����~�~�xL�pQ{�M��
�<G��w����[�ʇ��C	!y�H�Y7��wC���S=?�
)m�1�����u*�~F���b�L��A��nF���d,�M:ƭ����ȞL>jk��}�x�,,,�N|�=xS��y��j{�i��+��虑4}�7�Y�as�����+��?_�i����z�̼g"����*�/jhK�XC��;�)��N�B �^��N�A�ښ	"�vu�F�!X�G\,nՏ��������S<{���>��D��1 �c�U!��-DG���[9МJ+(�sk����s�LKG<r
�p<�����Zg)6�j�-Nt~~���
�6�D�J��h�����`*��d�Yxt�}��II��j��6HS���OĉВX'�z 5"@���IBJ*�M4N�+�=�����r�	lzex��:���r4���ٔ.׮�?W�<i	�k�m\�/�q�4`
`ꬷ����x�ڍ 	�̰�N�󋋍L�jwjK�8�7�Z���䊥�%�_d��U	�B)m���~Y.6�(�{�.�f���3?����?�$l�hjl�R@���B�V�R*�����Ŀ�y��iV���)�/L����ȳ���i${C�䄳��7�P�YgV�l�=��;K(x�>l��mӦ%̽�]��}O��$a"לF[WD��M]��)�ݵ�8�����iG���n7��k�gY�9myy�4I��O�L{�o����9:�"r�v�f�~M&薕^�����
�@A����&����71�2 3�I5��sZ�{ā�9kS��O���xm�K���j�T�u���9�0�F���Dp̄��<mH���C�9`mwiCؕ�6��{fc��k�%�B�\Xc�O��% 
]����魆l��)
�T/K�Zv7���1E�>E���6��9Η��y����ڔ��T����u�ZM��P:�������z�8�^tJ�Ȏz�(2Xj�����Q�0�BP�� �d���ܸ舋�C�����[���efy�1��0�/�8��aO\��V���ʐL�&ǜ'�.)5��n��h�bS�);�ro\������ۘm�� �A��E}pҕ�R�ep�v7~+s+n��E�����Ĕᖮg\�[�>ΩgKp�(�nk��4?L	�aw���RɎ����~�A����[v��o������)��qωe#K>��T#��
u��u$˫��޳IG�&T��_u�����y�A�~ü�k֐�ĸ���Ĕ�s�tZHk����2�����f;���Aۭ�b��\��eX<	l�X��6�e�����S�Hl��W����Z�G��m}6 �X�5���x�h��m�DT��� �>��9����.*N�;V'���b#�p%+kT� %��I�Ml�[gD�&ݜA._���:��O�{~�˥L��<��f���t�~�e�%�6�Jq����zҘ�lW����m��U�Ɨ����jS���S���ҋdۺ�\��)Sᨂ�6L�|
��'�N���}�r�sX���,���E;p�|��F��P�B���[���B �^��M�I`�ː�e%W�i���ճ5�Gx8�A�0�	z�S��L륚�	G���e�zxԓi�~�CV���E#6���ۗ�N&�6�Z.s��s���p�|u�_p"�$nUV��r�w*��Wow��m�%�Y����˴!�k*;	��O�Lټ��5i[�dj���*<��fKQ¾:�ZC\��� %����C�i�| ���"������Y
���t���(2��?.��k 	`���ƿ^��Z+�����R�fk�?��no��ı���]G�F0�D�A�ƴ�~�}|����|���٩�ZY���cԊ�JU1�'�[��13d�U�vY��^��>@K�\L�m�c��h��K�<��I/�3~��4B��'�Z�<��1�;�7;����n��cuC����L�cy;w��]�γuM�~�Dv��Dni�#���W+�o��.�m���oO-˗Q۷"czs���گ�311r���Ai_�c����I�j^c�D����`aqg�0Q)茍�`�ض�(�l�}��Ôp`<�aHP;]Rg�]��lx�����#�k�J�5�4�"2NHU�?�Ѫ�U_��b^Ub�*���S?�N?��v�r��G!�͍LL������D۾����^%t�"�� �'R5R�S�Bf�;��^�s�}>Y�����41����6"����-�dU:�ǝ���@<�'���6M�OY�_k�e�(��
��ǰ�T���@���C> JD9�}�����N���z��gJ�%W�r�~�&A��:�xd���!�i��'���V'F�f��S�/x�O+u���*/�?7��|�T�-�d#���H'��v�ګ��R{�Tm�l�@ʫ<(��8<��9���=�ݞ��8q(�T����M9e�����!W�7��8i�#fǃ�6�{~a�Y��"6�K�ΕW}2y��9B�al�Pp�nΧW�R�4����[�����f��Nl�}�~�eOm-_���6�t�(�R�~��}I!��;vNU���߂\���őD�{�@���uM��i��-e�߳�����1Ѝ���ظ�;S���GJ����Q��K�r����9�ҝ�e.$ѓ�U)qp��4�vN%<��,)�"������h�L%��uz7y�m��`�`�_C�f^b���Fm'�PG�gD�B���9�)��ׂB߻F����P`\N�ާŵ�d��}&�D�/c��פ�dk.O=�8��Q/�|V�WJ=%a���UJ��o���������\�k���B �Ͽ�Z=��"��i��0	Uuu�$E3䆜}���,�S�E��n�\9*Ȯ�ҩ&�$�ʎ0Ɯ�SW�,D�lv/<�����Z0譊���z��LH�q0S͌�?���������f����z����bv����L)1��h˫l�	�V�����\).��3��r�q�W�6ږ)h�?�ʿ���i�l^��T�v���w�m=}�}�i��Bhi��X`l�M(w�Ӎ*y1�4��Ŷ"@���#>Iɸ�#�:�������6_S��c)z��f��/���<��ue���&.bEYY kX�_+3ee�v���P��s��� �{�I�m.)^���f"ޜ�א@e���� r�6���b�ۣ��W�"�c*�k�|D���U�۵�TB��t��+���i����,^��f(�ߥV��6�\>��
��d�?�	[XV.�O`�[GDF�\�� �����71�����{o�٧Fجb����̷�/#�8aevi>r��vN�=��k�B����7DCz�?���pc>�����W��
K?L�����t����O�ǲ�'���/���\�-�0�)���-:X�;ݹT�t�~��,�f�q$�m��B�D���/�R/�������[����%���V��L�i0l�#�@�㰕@��� h�_�������va����YEs��ʁA+�K'�>+[BT��rΏ�/2�eH����2x0xڵ���I���S+�Ab�eDp���1�]š7&�'Ϥ��}��(�Iʱ������fܮ- �Iw�)����'ө=�){=�nD����x���ɼ|ʷᚍv-j����Ck�hu��@�i����F��ْK�O��a�[��['��Z��r�������#~)޹OߛtW��J�+h0�1��Fޠ}�¥��z���K���sK$�*�Xtc5{�o��qew���g�}�HJ�
����(�.ϯ^��,�L��x�5t����,<<��J|gmPN�
8��w����.�@#s*�%b����B?�~�30��Ya[����Ѡ$3�l�E�/;��O�J��F&�Y6F��k9�-НR_X�+6@�b���;y�Yμu)[ŌVP~(��ݣ@I��<�HA�I��'*>n��iH��-Iv�g�!����1=�S����O҃vS]����hy[����DR�R��ˑ�6��c5�ӯ�1�|�H�yFi��F�^�p'	�'��Q�j�.;4��bn9����n2����� E���׍�Q�2��g">:�#H�KKli����/+�hE���B��s\����1	7���Me	���1vx�^��?���X�0}�2�TJO����B�[�f�Q�6_��ч�Ē���Vnn�2Sw`���n�b	'wl\��U6j����6�C���K�tC1b��"�?���f\2���r�9��dL��%�+�l�FQr'��q�OQ�~й��s�z~g�m�v����)Ns���?����<R �m�qCbʧ9�}��#R@W�٬��VQ��*6�[a�<\,��M�V�R���vX�\{V���ɍ��@X"aƟ�A备 �Iaq�t'5��b[���@��P�-���ܠ����7q����	�o9�}^�O+\0=
H���s��qs��|�s�ы�6p]�I����'����V��G�VR[�v�OI�����|52X�b��o���]�U��̄)}�1�'�6���5�W���2�vÛ�a�07�T���ƶD�^��ߋT��yF�5�(�T��m�����͈�v�)���HխA�o�U|`3J�`O4G�˻�~���.%"���]��7��^������X=��;в���oq�f�3��2��}p���(~��	��*�Rּ숈Ӣ.
?P��ԫ�Xf�*�U·�W��Ry$���昕�L�_ ��Bg���t�f���bײ|}�����E�(��aqܳ��+��@�?7�e�dRe�j�zٴ#vJ͎��)30�$X��!?�'��u=cod_C�D8��f8�����O��wlmm�q���lj�e'��K ��v���=�2��b��Y�=�a�p�BG?��0�|�lw��R�g��`CD��}�|v]���-���O�(�"�k>�Cr�
�=gzM���P�NT���<�3�l*ƀ!�R��,�c��t)G�)W�����ץ|�f�C����4���pό(q����8��\�wZ���4��sF����p���gf�R7�M���>�s�AE�a-�q�������D���Ueړ���~zJad ����W"�`�,��+ ����T��l��i7VJ��?��:��Yn�( �S�0�k�K�os�}�\;7&'�=�:��:��6�����
F��3�
��QG�{</=9���'�c!.!֕Os���h��M��p�E������ԥ����!���jS?�LG�@���;���,�a9\��M�Ç�'Zp;�g[�z��I��q8���E�� �qXb�K�/��<$�\<���֖$��¸J����+�:�G�k�N)qS
�秃(���8�͐˭gX�\��GC&`C���8��S�Q��F�1�A���8�;,VW�4�]=4絺^.&�8��X�樏��Wk��{e����΄����=xA|���������QtT�A����ʊ�����Jh�X���kv��{����'�i��c�H�'���9 ��,��3��¶<LNJ��Z����}�O�B��j������F�1��͠n"{V�V��y�?N�j��1ï��UT��>�ꘗ���i���k�л��āI��6��+D]Rn����%X1���%*���qcIa��6i��� #u[�F���$d�g�(.f�$�����@
K��'�O#�	����v2�GO꽯��7UoC�������ߌ���X~7��憨5�Y�2)�&�4P
�VM$~�b�`HB�:%j(c$��k����xbqU�&�q���N�}ԝ|��.�;�e6u�~���`��?[K�x?>:H�*�Z5�M~z�3
�q�u}�f�wn���2�sh�D��D���?c1{�}����D�=H0�]�%���]Z���ᴃ�c��"�	B�=�b�?�'�ž>ݚ>q��IK~�������M�1�B!�������[�]��m��lf<؞<H�N{ZX��x
B��t1�dD2�\�7��7��$2�� ê���E��!dlr�����)G#c�(4-���8=wh��$�B��6�}�b�{�S��oh��x\8��
htd��n�su�W0�b�U<���/�? uk��r�vR"
\�7�u����˝+>6Tk�P�� z)����ӯR��"i�(��V�S�"���f�k1���p%���������]��l���Y9�j/�U�_m��Sa�eqH��ث���d' ?�)/��a�����f�(�N��Ћe�!D�哊4���u� NrYefX�%N����I8�*��k����/�6D�Md�̟��.�n��Mp��8�>���4`����p�r?gY4���Z�V����^��p;���tDb�ͤw�׮ۊ. h�EW��I���7��Bs�:�d��}'�W�Ќ��2k)�����`��Ǻ��x@L��/L����X�"@as.��õNj�6�;͖����t��s��?����眰&��&p��̄:}���,3��Ӡ�<��[��
�T�{�u�ZQ]}�V���J��� T�:� ��]�:�q��%܆Fr��_�����:ϋ�)��4��_�{���(��Š�y}̟@���v�V	��LA��!�H����P�M)0��H*�d�9֩��S'���Ki] � dCV��"AjK�G���ʚ�GZ�s�e8��H~ZDO�P3^�݅�
>�Bs�Q��O�'���ѳ��;w�ąLЪ+�\�P�?��
�����a�)��������ɷH�Q6�ZL���n��T���d/��}���u0��k!Vw{nx�'�$�(ܳf��y\`�(���#sÅ��::C���/}ahHw�9u����!p�ehs��=�_������$��7H�|
�s��ya�W �&}�M!���]�L�qȿE�b:a:i�G�x5X�w����H����Γ���r���p���ǈ�V���0D:�ͻ�jvw	��X�W[�Z4�O�擾����N���U�e�w�cW1�pk�3���4�M4Ņ4�:&��ƛXAl�lHL{IX�[��1 ��Z��µ&}��a�<���^�C��p�#Ϩ��}�Iu�˕J<���)��'���Q�(�+6�4��#<Bx�`�|Dpld�&�i����I�]7}�V��}�@��xA�_ӳ�>�+�m�l�2T#ny�6������f�;௛�"~I�%���� �[���S��aqhh��K�!41�^-���d�ŉ+��>�5�����q�a�0�R ���f�z���ƹ�NW�<���p��	�{i��<�6��s0�3����CG~w��^���N�k�0��K�>��z��#�ں=�A|����d	��@+�����vd経��j$۶��ESd���ZI�g��7��:学>J�_a�zp)�'ڱ�T�T{-J8��X._���UD�]���ʿu�i��Z��Ia~O��E�?�\F�Lr����޶�d�67�^f�y�Z�ܶ2�����}:/�\7�[':::4�� g���p�9ﰁ��o���Jp9'Q��?���Ԧh�'#�ku��j?\�s��^α4�Y�Fv��9�4'�� =/s�9�w�z�Em���}  P�
3�'4�\���r�	19,��/0X�ʁ,g{ReNrV��%6)~ءG$�8G+������rY��$."HJ��E�+����py��ߊzQK�A�6#��@7���,�F�,���R���վǇ����[փ�je,�=���z���87�(�I�T�������A��̍�0�,�J��_5�	��Y�ݧ~"9匘���0�Z[fs������a�$+��[LІF��/(��i�E�ǝ�kymZ�i�Fl���7k~��@�w�+���9��x�utt�õ��w��+E�u���x���<��X���#�|}q"���E ����g��%זTYj�I�wS�?�2X����U�*˺o�6`����[�lIX(�fOl�ÄE�� �,���7h9E96e޳pǜW�M�ө�KOD-b�%y2�MF�
��)��
�����Or�R���J�vu��A��f��)�/�3Լ[Ϯ�W��@W����S�5�ȱ��$F�i��C��&´hG��%�6ȂP�S�z6���D��`��*�-��-�o�c_Ӯ�M˛X����g�cW�R�Y!��`��{\U�2ȁ�c�!=/{`e��_�MŇ����P%�WN�P=��Y!�˅:�Q��
*9���k������#�8ǜ�$B$̝ &g�s6�%jq�i���WBب%u����A�Q�I�Ǜt��f*A��o�E��xy�bM�:o�kx5�;>�* �/�_�|i�ܹ��ZC�X���<þ��[I�C˵��@���.�F�5Q�#ݼ���>`@���EA�g���y�}�solXm����FJ���js"�Ε�P;�E͑\Ϧu�L�]��u�A��L�-�̇7癡_{[���������H1�V�]�k����Rs�g���8���m��GR��A�x���-3��\?��XK4ti{���]o���'�IkI�c&��?f��IL�����^+�8ތ��c~5&�4�Gl�%�ǃX��[9Xzh6�gd���%��j�/(���1��+�A4�թ`E�@�	-W֜S`��� s䄿~�B����+T�]��y��"�c�aR?dQ� ,��)�:Ơ!�Ѵ�� ��,�)6�}�{H��2nje��~o=�W_�Nj��׈ti�e��A3��%s�<��G
!T�{ŏ����hd��Y=0A�P�� 3������%^Odl!J/Ϝ6	���L��Ac%��
�&$Σ� �|4D&���հYZZ�/���@� :3�D���]���޿���I�������=%����G%���Kz?/���E��$�eKE]>*o���OH�A �8�t�IX��e�ʖYe������A��F^ꇻ�_���6��@����E�=v�λU��Yޓ�	�[3�Q�q��$�Q���3����lBA����J��ׄlON/cq�\��@�2�0p�S����y�> y!�Hu��q�������������U�,˅����T?�Z�	�� ��Z�ɡAߓ4
�{N�7��=�q��i<��r=�G�Xi,_u)ι�x�/�6�]~A�ē��!4��F�A1�Ft�r� KFc��Ɣ�Hܵ!+�b���/)��3{��K��6�L�s%��R"%]�GJ�y_��������_�(�sW�q��u�c�� ��3�v��B�E�m�n���`-��
�;+`����d"��fQ���9YcL�ĽF���^-G��U����B_�����h�;�Y����0�*�����b{S_��S�z�3j/���A�,4��ϕ��REƆ�ꤤ��j���w/�����ǩ�Q��
͈��*;T��J�Q�b��]˔����+@��f�par���Pr�Z���f?I�Nϔ��$p`�ދ���F>��⤍���q���2���ϟ/�np�DfŰ�3�M�I��B���/��v���v�Q���R޲�i�`�}�S�	�K	zC����[+#`��y�j�$A�*�ưn+G44�:�@~zzz>�f�Hi~�{Ǚ%�!Tz/v�i�I!�o%���<���ķ�����5F�n~uh*�6S)�]��_Uʂ\ԅA��ĕ�.��V���@*��G���I�w���/Lb����9��9��������y/�:ti�sV	��mQK.4!��A�),�ִx�[�msy�Q�7B��?rz���>>7G���ؑ���xn��B�Ecw.�d�${�*�ڍiW�^V�KU��Ta��r�E&)��p9ʲa��K	���x��-�L��@Xls0,���V�����"�湤�ԁL+�)w���q���t"(���2�ȋ�ܥ�Zy�ݦ.�*PS�Y�{E0�G�@���y�)��4�`����iB�ɜhS����)�������/�捉ؠ�/	7=�huPpJ�+rM�z�[ЛC�j��'��l+"IT���w�'�-�W�-���eT�����[AQ�#+~�u���7w��+oX;��*�2L±�Ɵwu �ް`a�n��`�Q1��j�v���w�����tS���%�����aq��aS[�wv�N��4|����r��%W�7��X�R��,���-��@w��;|��b��ҡ���b�B�E���b�K&��y7AFs�~������77&_��zu�mrqb����;�wi�r�e1N�3a���I���\�5@"�!��QW�"	�=]X7r�9�|�����,|��A� ��p��33������<'�M�t�W�*�t�:X d��E�q������+�n���� 2����^Y0~Ju����?��/l���Y�ƥ�l�G��d��.uTV��*K�.;�}��p�&���[vk��&��ps%����z�?��ٹ%h�ݣywN:<�N��h������ia�/��A��ỳ�Z:UTT�p�"���f�n4�F���e��!_�KC	T�c�N���"��>��1�R.� ���T+^�:y�/H|lKtP��?H9��d{��:2%^�3z��z�%o�#���ZG��W�&����d����/�Sj��bZr�p�S�ؾ�0:)��� ��{ҙt�6x��<�=�]c*ĥTB �n�������t��]�8y �����qe�A��7�LP�	���P��zql$\� @���חY8)|����Ȁ|Q�C{��G��e���� Gr�y;PP���߮]�l"���Z�b��}~'��d/�%k���܂�wj��m,�钸���sޙ�D�2t�;�K8��/���Y���Tze �b0���+� �Ϡ�=����C���KEv�����x�a��Kŉ��0��ǱF��?���F�<3���2R�_Ah�BA;y����+���?ի��F-�2�!�Ï��f��Uܤ��/>� U�{QT�ܡ�qdٝK/9�U�3�
V�N��ɥ�7�y�c=��0"�?����C#9����ӄ��n�	��>?����2��N9Ed��?�X��(���ѐ79��F��IFӋ�ȦN��JU��Þ3��E9O����"�;-)q�}R�x�ʭ���m?�t&�̷êO0��כ>ɿ�<������تb������� ~)wD�2�1&W������9~�{_2�Z�@z.W+��3v̌�U,��[�c�tX�j/��w���.K����ҳ'��b��p	���Hd�F���9���@�z�Y9c	�����V\�$<۠k+�k6�sAFv\����������C��t����q܋-
<$Of� �1�ڴ*�u��V�������߈�r�{%��O��%�7/%	`T��9|����+��G�
ı��SsQoph�T��5>x�Eo��Yԡ� 2Mpf�X^��� e^�А�K-�È��D4�B��_l=Gz�t�����~���ʿ���U<�t	��tԎ�F*���C<�ŵAd�N��S&!1CW��x�G�wF���0������cP?6.��Ǖ�[����p�7��ޚ��&���Nm�)x���
�j\vΖ��ݙ��C.D 7B$�8C�^+�Vi�>EbH�f�[oYZ�V�#�L���s����W�����إfg�xo/ZIi)�T�cݛ�o��cB<YtCZr֣��'7�k@Q�g��Ѫ1� ��Ԃ�h��8L�U?�@�8?Ĭ�)��㆏R��5etB��<��M�^��cfj5�z�N�ww���ju�qR�0LS�P|���A�!�x��n�2��=�(p]�_?���=����4�)�t�l�$�u������{o9i�cU�:uV���Ŧ���.\7� v��ٸ�XP�)���lH��ޜ�����y��Z{_G�X�5�:(�Ғ��S����}@�̶�ٚл�1*p�ճ64A�0���B�"S:�s{+�t؛SkDk�@:�j���4���l)�4c���a8dXޟ��<���سŽ�~��G�vw��M<�I��eiw`w��(31(9s
����s����(������XѾቃ��l{��Rn�\/RG�Yc�[ϐ����n���\澴4�ޓ���LRx˱���F��,�u���U>:���|!H���?�.躽T���EѰ���"f�L�n�C�,-FU��O��n����^r*�pL��7�@T�<2�>3՞u�	�ج�wZwgm�&��]7�v��3�y%����7��X1��rNm*��լ����M�KMD�t�0��}�+���$.�z��P.Wu%� qzɲ>��m�R�c��Н����~��മb�a�i�݌c�.�y6;���-*!�A֦C�g_��p��@����4��8�z3���V+�[n�������h��Rm��`!�Z
���.$�W�[T��Mr��/w�*G �gF�4ۈ��8jJۓ���\nPݥ�rMQ��+>5��wڵ��v��R�>m[�Vf���h��w�'_�����{�y^�<���������$�k�~_��;�mt��>��H��H��e��?��SP����Xw�R8�PЫ�~�Lg��}B�C7#8�M���U�b���V�¬i��D�B�{i�4:uP���Uׂ���R��<�J"���/���E��a6��f��#A��(鱐%MH��Ĭ�E��ó?ۮ�*9�P��կ\:ux+s�C�X���T�W`;��sN��'�R q��hv�1��8�~Dd��q?*���Ӎ5��j�+�4Ҵ�"/-2�F�X�5�)c�X�S0�
/�i�g�=s�*A��V���zNj~��.а�E�[�~���ܦ��޲@^��\=����u�cqS�����x����,c��q�;C|�!�-f�N8QbDy+���h|�I�}e��=#�)?�"Y��v�@�ʓ��'/�E�|�Ghʏ�+v�dM����$���Z�C�m���X߂H�";]��j�����ȝ��.��&�;��O9�W�Lۅ(�vK���l|�0܎#���g]dE(ɕq�&�̶��-�6[��`��3��;��2�g��&U�&qSBg���r��;��m�9��;��8O�aP�C?;�`���+�-�zӬ+[��!qI�8)��s3k+��7T�WWV�)��+������4�[��7�]��6�o�J:-�N���@��,�M��UѱnI��]��P���g�cx���=�K�=��E���E� �m��%����"��8�9��kf�+������֓�;���?�L 
8�ŕ�҅��V�H�����H�����e�܉L3���T R��Gl9;*�@�����ĩ2����"��A8`�eH��0�oE��|� �|�H�E��S�MjK�7��d��P>/ ^��:WN�K���������Iim=�&��Z�(�qt�In�ڕ"F�m6�Ra/9�����͚d�]{{���`��v�}PIB+���[#��4[��A�EZ�U�A��!����>^v�W����lې���!����s���G�ru��N=��>T;�m=����K
U?�J�0��-�HLyG'�,�.�F�5{�]b�o]!�(��%�v(�e7�W�W�����5>�͔WN[�����R�&��:_{����TǍ~�7LUL�, ���������֡���|"H��j5��R��m�:e{-�c���P�%9w�y"�:)M��ra��U&�PO`��\��^4�[g�O���ȼ�����C�ɹ�Y}B�'��ƦI��ձX���õ��q�7����l�����	�? �j8?Ĕ<�{X�q�\:Y8HR������� Y&�i�N�̅��p�8��/@�&)p���V\C&�Cdl�wM� �V���I`:7A�-*��1�����aM~�� �"H"%-- �0P�S@iҍ��(	�����56�cҌn�F����|��ϵ����y����_��<�9g��n۠ϛy���G�M����j�ӇY���R>�����u�z� 7.� �[�z�9�� �L}â^<�}�޷*�g�l=�Cdu_�F�E	��4�]{# ]L��/�
2�D�-�e5��l���x�g�JzN���V.%�T���5�G|9�� �%�#� �fI��yxe��{�����~�����Mءl���������_��|�N�;��^s�WI��(�[��ģ���շ��*� \;�|�v�?9��1J�f�s�?K�8`�ĢMZJ�򬨣���B���f:��w��ּ��o��~��{�ڟ�g�A�ݼKݛ�?:��z�۶VS7�`��sj��8U�邒.^�H��(xq�V�@yyz�m�-�I)�A,ǈ��
vA�>������[;Rj��/��鍫�x���7��'I�Y���1��˂e4�yPږ�v���a�����{���i9-\�J��n'�{�����.��˷��	4�ˠ�HJ�=Xc�%��ɭ��m��ݍ6S�Ԛ(�~�O��������u�(��x��S��}���3LDݳ��p!�*�;+��	�N�u/+t��'��&~-�Kɽ�GZC�p��E��	���	h�)��1c�:�u�:I(#sz�<�M���x���Fz$��2f�>���G���X.��� h�/d�#ZT�l+�;�22y�I�'�Cd�m�g����{E�|��=nq����z��ѫ��mC�HD���;L:/�` _�n�*�9XÂM!ȅq��0�ĐK�t�=8�\)�ޓ���?���J�}�@��˱ǖ����5��h�,:���럒}s����u$�u��}]��摵�`Q#�ȓg*��ۛ�*%�������Z�!G9����� ��D�I�@��NLB������C������z����-�0iǈ�4�g//��Z�?LEz���
9��#��'��a��7��L�5ng�_{uC���ւ�[C��W�i/.O��=���(��J�h��Oz�H;�3,��NE|�Mi�d\�;��~�:/�5��	�E=�.-P[`9qN�W �8=n>prT�ϸ�:�����9��W��o	y��Y�t�qT��߂�V���0R��Xn!���ָR�B���r�.Jw��^�gcI l�N�4#>}=e��r��k���:4���W�0>�^p͡D�3�Ӑ�'!:\�XbkŻzjh��G7����,�E9��ID~�,�=/{�A6U�����7{cz����0 ���¡�,@R)q���\U>Jl|�����I~s�-s'8*�;n�n_�s�}U��ѳnc�w�r�ҵ.�<�$Ty�x[�o�} Sg&b7L\��dXp��.���
�i���]U�?e3���oC
��% a�<+5�j/r�O�=�2���ѥ�yr�}��%����&
����MY:T9��n��T��d��og��Q�5�6�W̌ח5���M�*�OB���]V}m�LE�B�����Q�L^���j⋼9l��Y�Pwe?U���I��f�4|��5����WeJ���l2e��I3�g�z0��r��^K.E�������q
Ċ^DR}�M��܂�Yk�%�_��uKىrQ)����[Q�B�q���Ie����/x�{$�t��z�az^R��E[!9�������y�a	݇�{��E����a�Z\���Ř����k߿��?�v�ͻmd�=�}���n$'��S�T��դz���Z������
���E{&�>%j�g����������o-@�R��j\�HJ	�:�I�qљ�S���QҖ�!/��ǥ�T��S��Ý+�L���1�}�����3��n���kF��[�g��������D/��-DD��)�{F*�e��=�%����7l�8�*�HY(yj�1�$igw�sZq�0_���3 4� ���ο�������8��h��P��6��H	�H�[br��7�����N~G9	�-N+^ H�8�����1D�l��D����X���囈Юo���Ogr*�ˣ�e*i�M��o�sC)ԧb�]��C-�m �%�Y�z�fD�g���3�����K��^���=Vs�"����\��u��1��}9c/�[��N�z��X�?�eF���]�nF��>�UkY4�9�gψ�ˈ�YV�����ڸ݋t�ͷlI���}J���gMM�8���.�|x?��Y�힟���k�憊U�qC���A$��ϰGֳ= �e�+��i��ހJ�2,��ac�ޖ� ��ė������'�=��_{HJ˶߇x�o<���U�|B��y���j,���ݲ�`�T��H(�n8�V�&[qdx�S��\|��s����w�G�-��ϮL�yx�y�d	�%�w���s�)tzo�H��͹?���6���F�[�$$~,�~̴� 
�.��Tj�n�,���`�ѲZ�7��"�CO�:f$�����D�����-���d�����'��⧎���m�i=a*}T���o��'�L�	����w�0c�rRN?)���b�G)�&���3�]�3��,���9yZ$�����KjU�a�w���t22�V��F2����l�9_�{�͠�i�J"d,[(i��YfS_d�N�sui�̬��^κșs�}��SPa5-p ^�I�s�[9�C㭶P�數zvw�����=�l0�{�0�KCbr�l�	�����j��ì��*�(���&��\N��8���� �	��>��L>h��"��RIE�i?�;����6p�gQ2]x�J��N�($�'陙vo�5p��#�
��Q3r�Ch���2�QU��W���vf�:V�����'��/�j;°�e[p�^��P� 7d"���ǲ���sxPis��%�絷���ˍ;ɲTQw���8���^�Ϯ����w�Ҽe�w�-���sw@�?�`̷�ZI��j�i��$���D/4X�FkfW\O̡86�ԬKЄ)
)`�q
�e�B��4�}Ob�e�;|[��G��Յm�aq�g�tPDGb6�05���)U	��.+���!G��5���O�=<B�Y�O�mm�@�Q�ȁ7�����]�z<;	ųLBS�k�$�Ԗ��?x�[�YcF��_Y��o鐜�M��q��څ:Q�J3i��p�~qJ�Y�;���@����K�L�#��S���|�h�����d������F�zA2㊔h�}br &`�������L�����W�x$fL�f��/�ǌ���S���s�%���+ �/�����Xc}k�R��*&���F����z��g����zc?��)��.Dkh��� 8Uj����#^������h���q�-��&���?�,�s�>�o�,xI��e���is��̦""4ݳDz{�H��~te�\rY/#Pݴn�5�>�u[T��+>Y�W�e7'�7REI��H�r�sF�5z�=�ْ��nw�<��<C/�6�Gb��_�e�ܴC�.�[���
4�ɥ�T��]�Y�d����А��0�9PG2	C���̑m���N\̞Ϣ�^���K}��w|�t��U�D�{�M~5��V|$�ɴ���*R�W�Dk�ݚ)�&��<�:n#�����z���B�PS��J��G.��'����x� �=�Pm����x���5.�v�l���l��(�|g1�l���̅�.�.�������L��խ��ݚ2�1,	!��l��!&<³��"_G��k%_�9vN��1��z���.�oc�x)Έ�6ņ����]�}�6,^�8u�~�|���X�e�
cJ}��-_����ߗ�뻗�;�R�[ 2��q��2-���'7[�9	�c3N6e&	�s�i˲��S6�m�!wM�.�aB�Rt�O�R��[T�L�\3��m͇l�����E�n��T�z�2���#�?�3�so��I^��]jFj������¾~�����h9�V˅�n��BHm���F�dn��^!;E1'jkm tR�ߦ�"#�S����zC�@�����ȧ���ֽ���K������m�o�aDYc,�O�؆�G>y�y�L��h�A!�B�0�aFT�eS
F�1GӤ���'U��@/{�<?.��te���8��gJ�Y�s�z���1�l��$�;�QY[��_LN��.� ˖�Z&Gu���:�pR�S��ޅu�犜��'m�ݏ���g�$#���""�b&�/f�$���[�r�f�j<��x) p�d���ϛ�,���S[��"v���9D���χ�,�I�m����R���U��B� P�oF�U�3�}M:[��)2��d�O9Xx掭��� '�t
�����S{� �{L\L)��o�)"`���i?+��z�v���(<6>��ώ��-��B�G�/�^�џV���yTS�Jͷf��T�pU������� ����	o�	�V>x�/�����*#�ڝ5:P'=���]�ݖ�N%߳�#^kA����xT����!��?��-F��r��G���ޖ~��̙�)UX���IV:V����tS��y��\���>L��Z��݋�vgv��H�����9,6FW�U�6�/�v辞�y��ަ��m��/�ʽ�8f��1x)�+f�?쒗i������wy���kJ_��� �3�*��Y���^�z+�]fa�D�\x�?��(�y���������ß���+PϢ��nߞ �̈́�`FJ��ֶ��4*uJR��u��x~踶*�+�~��k�/5��Z�8o���<������k�!�H�N���������E�-��=[c�7t��=�ǝ<���������gW��c�Ԗ���D���Y��G�E�DF���7��Fy"��ワ�%�kL�&�1r"!�f)e��ǋ������co^x�e,��	+�.���sI������s��~��E�-y�\A	mFM�����M��&�vn�}I�w����r൥�]U���{��.�"R�HO���兔���S��r��&��/m�0�e'y���;�<0�<�I��VW���$F�,��!���^��F͙N|�̶�.���o���s��&�ϙ���M PjH���B;�������cpl���U�;�*�����tfͩjn�U��ڗ@F���{D�AW��#$���o�$F*���Pi9r^�.�=�	/��u?���{��qZ�o�s5_޸�}�fh��#�
yߦ}� ��Nt�Zs]���4�,�u_A�:�hR�'�j8����<��.�c�l 

�¶m�ͥ�T7N [0�cE�GU��UV�ќ����d(~APl�l�Oc79�f�rp~27�����m?p�������z,����sة���xʽ5�n�ߴ��	�2�0��砽�(��ʐ-�V�� ����޽`b��;�])�z~drhh(cWW���K[��k�'�p���g��;n[�N�w0� �'UpO�����ĕ��W���d��^f�Iwn���+������ey�����z
��w�n^�bK�r�s�"���W�B��x�'}Rٳ�&��/�(�}��t'���4)���Qg)ה�P�ѷ&��������Y��Qzڨ�ٿ����j�O/xy��Q܈��(�Y0��ݠݚqW�y�j4R��6_��2-���3v �9;{C��|ܯx˙��������{Ny��x��6&��:5�A�;�w��?o�lu�V�Rb����P�����M�Gwg���:�r��u�fy���S5Dh�J��E�m����o 1 %󺙏�h�G/)m�l���#�]f�<4���[�G
�Q�ڑrMe��<FNe���Ĝnx�>��^{�d,wz���W���UĘE{����f�7�߯d2)�4�����Uv�Q��h�1E<�a����W�	�[~Y�=L1�}m:WB�H=�+��%#�ss�S�)w���[����m}�<yl����`��[ie&�0O}Uzq@w�f�SCWdсc1�k��*b3�n�S[
�^��P�Rz�Jfǲ&".�Tȷ�Y�B]��f�f�Q�,�bhRM��o䋙ἤ_��n�o =!�R ����MAb�
$��0r����? 9����<Cwg�+7+�2ԥ�GɵF�׾Yvηb��#�Ut���dk%*?;��k2i���JE��d�=����S�[�\�v�;c��N�%/��V\,<�Ҳ��< �߾�m����2�ڶ�Z���kɐ�^&ܬ8��]~hχMXG�hL���W��ߩ�@xZ������Ϟ�����Px������BKR$�U@�~/�`]��Û�$e9b`����d�25e�&�L
Ƃ�Xh�����3�_(P���u��,_%�d���i'�M�k��RP��:��DS�����툰Pb����ßO�8�iv�䃻��M>_$*��5�_)͍9	NW{W�[iox�G�7KEZ��=ܡCo�
2H�����ޜ 0x/�tϯd��(1:������d+(�A��f�e��
x����L��m�ܳy��D���������0P?wn:<��c�r�Sc�.lr��=]�.b�M���Mϻ3""`%�>"p�&�f�F��nR�<�k����*V��ms���>��\L�ܑ6�n��p�gR��*�G|K�aJ�����;X�}���K��#���M��<gY:h��v�2%Z�T�#vgE��٭��k �t:��;�_䖑g�4�9:�����n��q�C�U�v�;X֬�!:��r��JD�~�l6K����kF��V�^u����T��B��F,Ssh�3�-�YT����/~��ސ��"m�=���w�a�ڣ֬��Yc�Z>�� ��}�r0��L������J^���)C)�s�_�r��Զ��p'1QX%�!��)QR�2�Fޫ�E��Z��$b�1��W�t�E.�"��=�(��[o���@ �%�p�a]E��̫l�m]��I�T��]����O�Sx]d [��x�b�>�JP�"��h��tP?���1Ҧ��lE^��(����o5*�~�&���w�m��m��0)�E\1�}$K��C��#(u����J����gd)��;p~�t
ٹV>|�#�����=g��$0�,��#l�z?�㒝�նb�������(Sz׻�'�����˂r�\/����LH�0�����=9��]�aO�/��tn�J6|O�׳�"`C���KF-��M��|e����5��]��	������1?�]qD��iTu����S���?��@%<���x�m�%~�bB���-��Z*��	��^�s�د�f���m�m7���=Y|���h�׵I�4�7�ѥE�H��aR��f�*$b�������Nv�-��3y�`S�AD���/i#��S�����\��w�3E�pj
����Qæ}y��NN��d���Zz�~��ސ�߼�wې'�j{cV-F�c�O�mX��o6�?iw���k�:P@#��d��1��۴�
�m�x�>$J�-�Z^52S�ߵf�-�P�ճ��D����������cUx�6�k�K�+/�t�d��W�:�^':�{�j6�>���v2�;�x:��
DԪ}.�M�y�@�:�QQ�����Vtmv�w�e���л��}�=�5��R�����9dS�������IEj�d?p��w�=�cQ#���gW�k�4�;���[��ƽ�%E�or�[�k�K[�.&����{��ҵ�H{���������ly2�k�(dv���	JKC�����]j�k,ң��պ���X�,�hH���������̓�mz'�t㹮=�`k�����|:N�|r>�C����7 %3�z����{�QT��T��w�O[W� �ڰ������R=����(9���§�M�DK(a��h�qZ�A�����	@hL����vd���Vћ�ƛ&b�0����>��'zbh�K(���s���Et�m"�ɨ��կ�QJ���XsZ�_w��-j�O��'k�e'�ss��ÜQhC��O�'���}D�A�@-|���K���ڸ^�>����	�o<W�n;�7i�|�5�'_3J�>��.`�9����yL��uL�B�{�RlB�s$�@b+����NNZ�� 2db�qJ쀯���ƃ���	� x�+q�>`4�{��ǡ�%m���C��/;8�_�G�]aE^�t��ж����]ܮ��w���������+���#8��P֣�/O�����{��\D6@u�bꕖPmd��q�%�����S�}��)*@�0#G�4:� OQ�:9��ν�b�Z/
i��<f�����!����m�+��Q����}~�)�ci���ޠ�l�Ԁ��!f/�X���"�A������X==[j�`7&�DW�<�4�ֿ�C`ߚ_�錴vi��k��̱��/4Ɨ��^H0 �ҢR8~��Z���"q9gr?4,?>�Z�E��aF.�L� G�ILKo���y3Ju�f9)o�+T�`̊F{�jJ�<|H���C�~jK寂kT�^��<b��}���h�q�^0MrA��<�)����M�@`2����f#�^����¸�$�����$3���:3xZ.}���ͳ�юvM�ƕ.�M-���w+���� d�C��܎�zp�~9Z�e��dR%�E֙5
�D	@9K�eib��｜����'����{e��]-&�R�X�6j8�RƎ��Q����^=M���s��O����"��m�rE���Y�#^pc�h�h��D=Zo���MQ��4��x�A��'o�_>BN�(�:G���0-��߽-�.�뢚_R_�ܝ���z`��9>�Պ����>&U�n�>��(����;�q��-20Pt���x��w9�Z0qN ~��N���u@�7�����Q��<�>��3�f��yHF\w��%Ә(�,o��R,��b�E��)�e �@�5�TB��:ne�B��j`nC��_�q����5�^4��M����GͶ|җ�֧\��'��j�U�2#��%��3�<�;]'O�BL�ڟ�O@+*h�p��II �$�n]9���{�eU.*�O�^9;漬V?K��=�2~��"�����d�RTf1M�����tJ��G�6o����^2D�;��ⷼ���_;u�B�d�s��%D�e� �G�U����t�F����?�˨�'9����΃�S�t���O41���c�<�ڈ�7N
�R����Q�u@S�}��������y���[�:�~�#V
����N�@�lK)f{M�6',p��,_����+�+�ƚ�'G�h���K]�8����(3��j�9�`�_`��ޢ�0�,,�{�<����h2��K�&[}���m����v�s�)���>��?ε,�\Ze�>U{hV.a�B�c~3�� �I����]kXw�Kw4��Z~.�F�t���[���?��ޒ��bC��:_&c1��������M��J�����4&z���^�Geń�x0���\��@0�y�66i�,i��SQ%�r.�子&�p��/o���ר��{G�����s�i���o\�<����\"�˅{Bj,7<�-����h]�B{���C$R�+`>�¶���{ ��8���^��引�K��ׂЭ�ߊ=;"�w��������#���o�d[nu_Qm�Tw����T�*�Z�Y�
F�b��]�l*,�jx����=N<�ѣl��KLQ��SNNR^��<H?}2�UJ�5Y��?�������5��PO<̐}�dS�@g��6��E%���E�q�@��1踠�uFS�	��DϘg����5�r1c|��/;a��1�e�T�x٨�/c[k.��f���U��7b։�3��̏���G�R=���KM�(1�H̺p�b�w͋�����QCn!�d�@O���3h0�x¤�EǠ��&+>�&�Qlr	���Fe���lWa��Lֲ�P��{�>�B\�M��bBrmUD���_����"d�#g�{�q-?Fy���������	�+|D���,�l<�A3q���<���lz����T��X��2~�����f&e��P8Ru8�z7!q+֝M��,�	跼+��gn�^"Ϋ���?�ژm��Z�?��t:,ifp!����`�4�5��A��~�IpRY�߷��j�"��7���������O��;�Ӻ|(L��ė��%���nTS��,CGe'(Pz��)�YK�k���Td媳�ڏ�Y��N������i��wr���~R�ֵ(d0?��_Zs^��9���Y�/uk�q&梁��ż��nv��b�te:�7/�NH��a-l���sssOn��D�`U�8�/M�
1��S���;��#sqE��m��8$���M��G�B_}'���~�a�u�8�iq����I�nG-�{��qttR��7׉6��Z��a�_ �,���+8j��K}�8H���'/��O���}äs��sW/�l�O��5˱�݊�2T3�^U�o��,9bD^�j1W7�������@=H<#X����f����=�"Os*�K�'צ����� �����Oacn<���ṅ��,A�����jq���O�wd_�����7�觿X��"VE/��lufOl`b?D�����酡ܞ˶�����e?�?7 �͒���w}_�E3Mv�Ǹ���i�!��_��/��جt�Wԏ�*y�|OЩ\8�D�[�6o��o��'��B�b�_�:����p��B�nBL��Y�/R`;}W쇹��#1�I���_ѷ�7� _��s5����u��x�CT��B7����#���o��0���2ҽn�t����M+�|.ݽ>LL����h������r�����F��gF2As�-�
��Ʊ%���=�۶����+7+�s� ��M� nЖ���Y 5Yx���7���}�%�y,�b�l?�{����L��d��Gc5����=L�b���h��v3O��L�`��)���;��a/8_�y�\R뼵��_j��tk))LJ��i�{�	�>=*�\���غ[�%������-��(�>���pm�s�0�����%x4�7M����z�����b�2'kĚi�3����7����z"���I��#���d,ҋ'�|��5��D�ZZ�u5�� �{���q܍��Qw=o]�F��^�h����B� �}F�1s�c��ToUlK��^"����^�ǩ�������o���^$2��T�[�#����,nZC`��ѣU���mOE"*�9���wd1&V{����%���Q~T]c��8�Mª�('��=���]A��7��H�.-���������JQ��I���M��QM�"q
�no�X:F?�Q����/��{0��=?��-	\�Ab$YM�V	���^oN�'E��7�g�d��}I��f�������:��I��3Zil���S��\���[ 6�>�]��?���Ay.~�����[�*.i�)����>E�sM=�=�"Ke���gzi����j4�<3����$u��AD|�����j.z3 �#��Kg���8�:��d��{v�C�v�mcF��v2�/�0��˾�1�d~4�2�N;�����el���G�Q��c���r��Ͳ���y�$l��_�)ז=�i�~8�5�
��/�� ���ȦcJ�9�T��w�';����e�ͷ�$!ϵ#צ�9�1��KM"�iN7�YZ�a�V3>���U�mݽ;?C��?�x,,����M����3@�r+=(��;��-LSJ�L���#���7�ۑ6i��I!/��>�Gi/�j*�ҿ����bk�F�n����W������g׫yq��?mrA��T����y��P���rCb0����}Er����5t�9�	�:RD�R�@FL
�W���tA��]j`�sO,���]�F)�A/��]#��bDq�w�>��<B�.�cI���Wu��ݘ��x��ȗ�5��� Ts���%~�p.��eޚ���!��0��]N����^�c����\H�b���p�q�g#넍3���?z5����\�^=� 8D;g}/�x�mf�=zWAy��N��~���3Z%d��Q8ǃ��
�ZV��
t��
�����>������a8mp���]E���_	$��B�AM�^g���E&�10���jW������`~$��<IH�6�l�ٶA��{��_#O��?�#�E�F�8���8'���7f]��A�:'��Q��][�g�ƕ���?��nv&���{�^�x�X*�=� |ʟ�<\K�����_sAH-j�|���N�ֻt�yc�f+�XǸ�CH�]�Xw ��fK�yx]qR��G��φU�Oq��SRGj�>���wV�,g�y,[����w��*���ZI�U�`�K<����K�P�vV�9�TM�U}HY��6���7b%��Fq<��pSͬ��gxw����̞!����w�Z�O[�4��|Ѵ~p�����������}��$��5ȿ������h������Z��C�d�6�\3��z�>�O���٨8A�F��U��&�����ѡ`�J]�&�� 4�$���\�N�zoR�UU�	�Z���I�L*}�5"�x�}�Ӷz��1Li_�ќ����7�HD��P Q$�jv��~��j�pV�L�|{���c ���W�I??��T�ۚ��P-���M�=�O���!\���S��ʛQ���s��0�9� d���ydF1����,&)R�ϻ_\������}���_n4/
>���̖H�t'a����<*O�M,�R��ڲ�Q��8��9���ɐI�"�"���v�¢Oh��8!d��w7��H�0�����.NK�����9*5�0c�rb|�pO�D�AV���6�Wd�LD�Mt�
�ӏ����M}��Jd�P�=i�v�R��<�lu�sﻬ$hdN�K}����:�B0%�<>��/��E�UD-ɥ���������8�5�/�D��Hش������v�e{��{�
'b����j�m�9�~H�8}����*�*-��qR�x�3�.�;[7�<�a�~Y�T'd#�ԑ3m�s߶6'��3U��s?�Ts����e^Q���~w4v1k,�f{ Q�$�����ɏWMG��	���jO�����*���h
Op� f���J*�����r�_�W�(%����q ߪ�7�=|�2�Ӂ{c�rD��t4�YdcF�u�O�0P���(�8w��n^|��3)���Z#2'�5J~
�0<֭t�����V�m���mމGzlI�M3���j�@����`1,b���v���(J6��P/,�댄�a���;L%o9[Ju�d@��%�Ȁo�uI�&s_}y�] ���9d���aTU��9ϥT��>0��Id��j�3��^���&K+>�����"r��J�����l��U�F�7N�֡Z���f��Q �G/�j��c_��N����������s�|ا^��cT����"?�<I�Y�E`��cO��!Ů��2���{�J����E����@w��W�N�1#�:!��
҆'�d���bB�M�f���pY�e6�9��#
i���@^M���-��*�Έ�K!`N�VE���/b�8�B�kj�����֨2��#-�����c��\P��O�h1"�g�~�֤�qөP����NI <3>�p�^@ʹ�3��gt4�=�B9-6���7ٮ�
]��)��j�z8�\�hK-�7�jp[�+��z�����:C�N�fEA�ٴ�q���X�����ܿ]��|�W��wc���T�'{��z[���IG�H���uOU�Cެ^?~�;H�X�X�z�*�e/̌$����Ÿ�E�Qv\�2"���V�F��2e��cK�\D�$�Օ����Mz�Z��l�TdW�B�\ū�e�v��כ��$��yLU����9���(��������5q�̓�+.#PKj8m �I����.v����jЧ� V�@���G$�D�����҄H\��	�Z6��9yN-��l^���]�bG�F�B &��O&b�'����L»�e�kU�L7hhHc����sW�����,��-^���j�����h�uF�'}���f���Q�k��l�wgO��W,����I�a���m�3�&tQ=11ڛ���?@����w���V53o�\� e��5lǥ悏�K��i�tde*�N���T��,~���$nb��;�n#Mw�R}��'D!��7��{V4;�2t�*z:,��@j>�D�a�YI��C��짬�c�;�Q]�Z��%CE��g۩&}��Ǜ&���I��eC�֊��.�N3���h�$C�>F?K�F&�����*�����XY?�>3n|���S�~�s#~�<3��fk���|�m��z�[z�J���b9�a+?���$��V$o|An�y�.��^�ힲ���3��;p1�wp?����G����{�L��X�x4N�u��q4�o�?����Gj�}�t�Np[�<@�[����f�'Y�]AS�C���/c�v�HH�����a"�,�5z$��p�7$��K/����a{����[�V��$iR]X�e���읋P¿��,7�ԕ���ʧm��W&�|.�V������*~!����o̫��o�������ם��S������KW�I}���'�s���JgR�s�f�$�Ӿ�^p9�#?���DR�p���g�g����,�,[��݌�XI���h@�1���o�L�->K�dBkO�c5��^>i���YU^nU��ͪ��s_]�
���I�jh ��S3����mV��k���$:U_\λ�A��m2 9>����h�"_f�Z���H�'�����R{���8��'Pc���W�Yz#8���~��e�����8>�,\����ʒ���c;��J[�K����B��b�cE�|p�X�'k�p,��� �ε�27b2���S��^i�P�m�|�}��� D{����~D����}�f��7h�[2Ǻ����o<V)q9dW:E����,�1��XRi����{�ֈ��%]�?365�$.q��p�ߤ'܁�rd���!�<֛q��>M;��&��?/D_�IJ�"��g���{��\�� ^���U.R�_3|K*t�<"�>Y֕tH.Rs��P��3��[�?�V�1P�b�̚�q�@���OzT	��rH籱�R�0��[���Afoo���(�	*IĤg�놉MS�D�o���ǹ5��[��0[8���J�&�hF�f��Og'��E��I�2Tpio���S��}B�{���|����\/N��Ib����C� �S�0�38::��/:a�k��3kTf�fs*y��Ze
����m�],a�Rr��HV:��_��� ?]ز�����\wI��<y��r������)(<�h�7��lK������'_b~J\�V�y��L�8h;C�Dl�o+Q�'�	��Z{j���¢U��jDm'SN�Э�����K^�:&8�$�\��q�w��+ �k b.06s��|��_�B��_5A
Pi��/�	�ޟ�4�z���sΓ�S\�l|X`�#��ŭ�}RX�_(@um~'�:\_��d'0�+�`a=����� �z\~ٯw�"V_�7����ٞ�JÙ�?(��O���A1�s��e���|߯Ƶ�R�uS���$�r/��@f�Ag'�Ep�ì�A�$��d�|�b�q��|�o��Ywbh>ֲ�[=9e=lh=>�`����z����nD����N��D�
@'6Dձ2���-��?���z��Dv짟�\��G`��b)��wD�>����Z#���Y��$���#'1�VŤ�rɝrb�6�[�ԼnUͦ��a^��z�mg�iȻ`�z�գIMBWq�p�xc�N��5-�j�����7��uj���C9m�Ҿ`�)�~�����T�4t��Ħ������#��V��a��tӍ'����~�+%�mҔ�&���FK4�6O`7���Q��"���J��A-�	p6�ϨaO�R��{�`uK��V�,����t�w^�D�UN�����^tܼ�S�۹G�b9��b��Ղ���|�+�K��?+xs���yr�}va��u�+�([	�k;���l8 ���O�I�+J�j���w|D�{ǪF�:��hU2���*�1�LF1*\�I*��$&��l�m�A��;���j	s��/�o���m��~\�ZmXT;�����-��~4��S�Ac$̗�Ay�>�Yr��ˌ�.K���ջ���\���/�x^3����_���њĝ��7_,�Y������ ֭������)߉��Z����z-v�Z�3.Iq�+j�J@d��nhzl���m�C!sX��`hz⌅/!�̮"7[m�K��Ȯ��Ei!��E߸���B����̀b\v�D"�,�WE�l�D��B?�(���;A�.�%8�`ae1����rc_:hHm��0Fˡ�ݐ��uY��5�f�NͿ2T��5c�M0F�^�~�M3�׆�
�,v��3Z��T��׳���EC���,� ��`z��
�O4�.O������7U�k���6��]��&�n�J����JM_�ϝ�i����6�wm�t}��^�y���>�,n��ɯy�;7���_�9����ɏ�u[��޽o}��)C�	��(p��|�d��`���34�����`���_N����o�������)�	 PK   ���X��Y9-  �-  /   images/4fde46ef-4620-45fe-a6b4-d27a85e18129.png�wUW�-�.��]�3�ˠ���w�P��ݝ�"�ݵ�S��a��y�9Y+ٹIr�����*��B��� /�M�_�_TM�b��]���AAa�ϡ�Y0H�����%�|�.Q���ӏ�!�W�����XH��d��P�p�|la�!Ss����ۄ���:^ۥf=/��;�?>_�i��FK�CC�EA>��J�Y��$��׷?	>ia#��ix>Q����z����	1q�������Z�� ����Ӷrð�dy��'
Q�j&��	�*�Y�L�ⵤ�E_A�(�٣��ELz�F��h@ڹ>ʻ�\*ʅ��P�5�-�/�j\~i�-�vu�mrq1Qۢɨ#��&��̆Ɠ�G�9����mty�y�x�Ϯ����e:���U��.�2���P��a~-*��X��r�yTi����!�T�#���7C�^Uh�;r�� ������e���n��0&-c�"�5�y�_ /�P����6�j�ڸ,�]}$���)�����" �"p+�%ұ��<���}Uh�a�ĩ���C�t��'����#7Õ�Z�1!O���U�S���z��J�b��~q�:���Y)��;w��y����,�J��h_�m'W{�E�+�Y}�]8>�,p|7�+�"z�õ��#����-�����M�ԫa���Ph{Ji�s	�\ޤE�/V��	��y#F�]O��c���}-�s�.\�{�&k�?]���0A��4�J0!~����C�X	`x8��c��Ĥ�r�"e������G�^2����ێ��+�vʫZ���j��ɀ�	8�������m�L��{C2ء�I�9ɖh�m��е��`RBI�,J�|��4�Uc�jX�jJ*�Jo�LB��o����	?9q��"�X*T��;+*���=}�5��td����ͅPl4��=��sM�b �L�j�~���VT�����~y�F���1U��M�դ<��#ZaHQ�&9☞�f�g&�ܰ��Lx@�]�$_'G=Q��Y
EEe.�h�pΝ�P�业>-]8?��T5:琺l�k�0�{O��X�P�?��'�݈�)�1����������߇/�_bR;I2ӳԭ ���W8�,�,&���B�ܬ�r���̯��H��j��d��n!jIn�������c�g�o�N2<%^��5C�L��l�m�N�OB�ۮ��<j��?��Q�I��f�!��R ٤�,���8ɻ�Z��yHa~����4˿R2��խ�$��!�a�Bevq�_,ʁ�_=o&/�gqK�A-~�����'�D��'�s׃��bR�M�D6ß��t�>���� ��i&����UN�lʺ�[��7���.Ջt��w9s"s���:Q[`�-��xR���M��	��ǘ��U>1�d���8��R
�ާl�4j`�eW���6x�����(qV䩄#|�����q�gu|�ñ�w��[�N2����IWќN5̮>�+~N7-Wm��jr�m��˱���[���mX1�F��S��d�/�{ss�G�k9���ZF��Х)%h������~V�*��L*����~QV�����	V�,�9H�c�x�~üG�Ϗ:=,���;��ٸ�KСs���5�+�4����ԑ=j�2+2=r�ur�VTZx�������Ĩ�_��%����2�X[l���Fto�]��ZE�*O$��X8<h�r��l��G� �w���Y���`�hQ% �u��E�*b�Ճ����F�2�� ���.l�%�]C�4��1�Ha��M��%6��AEE�Hv�!��NS��tz�u�?�s�7-D�2ųYHǥŌW�E���ٶ����E�~��x�� a�Y"�����v~?�Z"Y�%�!h��<0?Ϧ�iJz-��}GD�d5�؁=B��\C0�	���]��-������d	��#=R����>G{kIM�2�A�R9@"�1̠�$�UbA�AZ�H:SF
�q{%�*}��Lx�%S b�㿍S ��II�,��'��h���ٙT��J{�v0{��2$(�7(����4���GJU<w�� ��{#�	�NDH7�9_΋��n�Pr�6/R�> 
+N�t&����s�n`�0Z���^ٕ4D�AWm]8��7=*�>�t������u�Q�^
Q�2[�"F��1Y���#6Y3&���&+����/)���tFU��y�?_��X��La�.���R��^����Z���2�by��"���.�xj�����^�~��f��F��lW�e�2`�3_.�Z*f\��ifn��Xu���R�?�v�P+���]_0E�.:/���Phe)4a��W���þ���ıh�e��=-� �Oha�2Z]Hr*HB����{���OF����[lQ���1����j���|>m�֘��ۢ���_�p8��xnn�A}�/X�&�Z	�CRG�uV%�!/@\.u�d�Z:�Ϙр-gH:g�8N�3��Ÿ_��A���OF��bj[Կ��i��I�[۪(2F�@����`����O{�ķa��/7��p��s����x�����%���'Pg��
&���W���<A��ij���'z'��9���bN@�Z����y#®M��iW[Ţ���7�6T����4��ȁM�g~)1�Wb�W�Y�))b�J ����k�p>Viϵ�όC�~P��ԌW0�����`��V���Q�����!b��L$����Z3������+�}F��Ǫjʃe'a���o�����W�-XtJ��~�``��73	E���ٲ/ϣ�����)pv��K���	����,�H�h!Ҧ>�c!�v�R�b�n������2�Ş��2�~���v-��5�HX;�]�%ΔG������ǃ�!�gB:��r,�`HRI�����Jr��G��� ��Ĝ!
.�b��� �zT�����4[E0���)�<�5�H]xᰏ��,�1bz"�ˇ������T�v�qH���4q-� �V�J4�BS�:GE�\Ƙ�m���0m(
.0g�<�"V�o����;�����Sj%��QZ��?q��?�ȞԁDlU��\��W���X��b��~y��̲�-���&�U�貵�fǅu��g���}�!Z�����TwRn��('0�7�K>�J�R�BRw��k2�:���Yi�B{5�������OI�x��p�h�ſF����$�S�f���a���X嶈0��x8烵�^����;�7�������Y� u��<��9F[�zo�Y!��l*�Z���9t:���%���^~�J��W�1s\B.�6�
���4��\&�K�=+&H��I&B��bu�s�y�g���ݓfi�X%xIۭ�m{n�� w$y�3PH�;�UnD CJr��:g�C�IS3�L�@�ʃN����)����t�<��Θ�����A����
)�sʖ�=�KӭU���k��u��w�o�q�`�N�Έ�:�`!�<U^�1�˨�����+�2��`�QE-�>��$�z<��}�7{�
V����e��xsz�!':@� �������Q��!�믔�3�5����U�ӥ<���Z6�aۥ�!�/M��[]�	-W@U�2�Y��>����U�rЉB�4��5J����uq5�n�_�Xn�ܝ���[��Oa:��7n*S�>`��:���2�����x.��u�񹠠n�1��m�-1�b,t`5Y*3H�i�O�wҐ��y_Wf���[<�\�$�������;�����Q�C!E�58JC��|3�PL�E�F�ٳ�.��R��h��ħ+<W�A�i�<��FyH*���%�j�'�r��Oib��=S��\���_T �w�'��dP-H�(IhO�ݼu��С��.�Ө[��k��x6؟���vK��?���axebu�/�{`;@r��5n3���8�ea�p�.�4�N+n��P���E�ܩ���́�4%�2�&��0q؛�\z��u#GČ��`FW6��G�>�a�W/�ga�)oq�e9��Ѩ�*��Psm�s��~��@V^۱.��q�� �IYa�?�\���v��A{ؤ0�������L�c���[��ٕ~9xm>�g؉n�$�&�&������- ��ʟ�uć���8�t�\����Ǧ؋`&v [��'ۛ�Tk��dJ}��P�Pd�zi�R��+e@CIZ�wmN�J�5��NFꍚ3v�}]��r8=W����5#�b&~�`�oM�Oh�G�G%br@�B+z~��Mp�� }! 甖G*Y�wh5�JĘ�X��Z��E�9J͏Ө6�x�d?�RÒ�7f�xv��"i�1dTW�Ƙ�6� � 2k�:zi��u��@�)r�gT������Pp8.V�׽0:N˯B��N1��-��W�ߕ�&�Ò%�@A�KB+	H�~�_WX�S*�ػ��l��t�M�X�*c���N���{�u���Ky����^�f���T�e�R1u�#Q�呬�YŤEo��Mg���W���5��3*��2>�s�R\'y��FW��Ra-�Smf�������	�����g`E��E��o�m:.<K�Nz|su� q��꘱�MXy�^_�B��G��)��z��g9��m�z��������T���5�&a��3J�E��3�V�d灪�x��{?���o@|w��G�{0j_�����☍Bfb�_�2�@������)��Oo�'�Ik�oR�5�@$]�i��,�K�l��L��r�E�Dp8��UQ��(��Y�,e��'`ן���׺�^?�e0ต:�TZ��(���]�iK���N-��¿I8������z�S��'��H�y��&\8�"N���ft#�2H$ Э�({�Om�OY�Ciξ3q�Ӥ��	C�(����}�M/�v���G�8�p�"X���׶�������=�Ҧ���m�R��p+�|���qu�}{(�(S[��m��J��Ɠ9�~9�н��3>�{e��CkQx��t�n��F��n�'�h��
 ��l�W��.��|jE�I�8��"��d}F��K�K�ʗ:L�K#>`��{'����n�j�Y,��2~��.fL��[K�|q�m�&a�����!�7�ؿYzq��w���u�XFfFw�-��	�����<l�z�#=Ô)W�#*�.F�M�5��ؽ�.R��������{���1H�]�t��m�d�
| O�����*�s�tWp�	b�����9D��f�a[�M��[����wg�|D	�9L��\�ՙO���xRqGFF��0DC|� �|ۭ�Ծ��s�j�QI֖��o�Ԫ�ѥ�".J��7��J��76������Hǂ��/E��֎���O-2��C��EH�\��[gҿ�cB���Չ�����5gn��8{B��������kFn���ių�0�<;�y�HBT!n���7i�����f�����g�b��3���s�԰������{��6�짵��A����w^6]�v�MD���w�W��h/u��ϝ�0���I����yblrL�!-���f?�}H�w�M
ѿ\�yt�1[|w��}�C��c(,��%p�꼣h�ԕ�׈��a���!�?E�Ijmʗ+�}��+V^�kiC�����Xϟ95(�O�\���񏉎Y_}l��,,��9; �̇�Z��Q�&(-��{ ��
H`J׿��:˧-~�>gׁ�ǯV4�Vy�e�k�����F�SN������5(���yS��v9�x9Y�\#�y��!��OU ,а����8����-�W�Hm�<�t�k��.'+�m��ZM䫯F+�W���E)'P�%�t�*��1�
E�m��͍���a�:T�������O�Нd�-����V�\j<�u�{�˦	�G�b���ZǷ���zI������4�ط����K3�����.��]���P�?g��'��O O�l~<��_6���;"�~S�*��礷� �-8[j��.��j���L�ǘ'4Q��x&A(���|�W*ɰH�K(r�!-��"'�qghTO=sݜ����D��J��jȮMR@�Fc�!h
�<5wKyI�i�\���>�QoQ���RB㥠7��[��k��iX
O��iʪ�G57E��ת{W��c�G�C�����L��\nUX"�k���0U%��sS(�2�
*!̌%nz��O�b²�>x,��!F�$f����İM�sl��qH��C��3,ˌW��I��w���ÔoW�L�ȓ�~�t��/	b���)�&��Xe�P��.y�l-��W3��Ldb�R��#g���`3i�Qh��<�o� )���+1&�
���F��V�&�='�S�c����j��g���h��1��-E���=��D�7ʍHDG� c3�)���OL���$�G%�C/)�v�4nK�9U�j�kL��Sp�9|�P��Ԭ�t�qB=n.����=�s��q�T,?�;�Q�F֘��,�Ց���.Ocvn�4[I^�K�u��>���vev�<H� ;���z�DuUu��-;���F�Cgu�����йlr�J�o`0�6ט�=�-�+�:+7���1.�����A��i��^����:m�ݏ;S�5���,+S2�ደ��;���ݛ�0?Ȕ�|�r�I�:�ϩ��~�jɼ�Sai!z���auקY�Ff��p
yq��R,��=�^� U�tNb� i���N��p�bs��r�"�	��5�b����V��|�T]l��No.���LIEOf/b(����ZVظ,.�9�4ξ�_ 7=I���1{��l�j�޿���z�E��ՄE�eO-t�OaP�u���7|�ǚ皚Kؖ)��n���	Ǽ���t���?�̓D�������dg�:�ꪓE���t,��B�&���^�U��n��\��9
Ѝ2(�-��S�2Xښ��y���'���⢵~�y��[�����lb�Lo�5��;�~4�����N�(�ŝ�`i��+��J#��K/<�VZ�@�vV���GG$�</E�����x����ZY���M= rъ�E��y5"s9��?=�T�P`̥�
�� i�1�$�,�َ��$ ���ӐG�ɪr���)8
��=k���rM�O�����Ϗ�s�=��a��6���g�LS���b|����]�$|��a��l��O�58�Vf���4�A���B�[X�`5����f3٠_ZU!�P���ETo���&�'y��a�a���o+=�qb��zd��*N�񥊕%�MP��޴Vf��V�n	-�'�Q�N���g���9�s��[F�{��C9p�{�s�����cZ��8�H�ֈ)�*>HTx����EXԺ]s�i�����i�27�~�����[���O�c�c����[��X���� ����W�8��b6Ig��������W<+j�A&ZY�8Ã)��^�`�ּ8aD4��[���c�c������ՏX7s�O<����9�K��=[��3p�ǺJ���^[*aT���[���-���-U�.�f�1��A��`(�G�o �%�@t���J�H�A�+���5>��G/��]l R���ɖ ��<-��[��%���Q�͢Mi�h�����~��D\�
� Ϫl�	�1�K���yA��ɋu�Yg�:�~6ө 4�tY�" �C���"8,/�|)���q6��PJ������F�����K#���f��>g��C1�-�W�y���۷��*2[o�~��z��t���t��,��;�kc%5]�xI�E�,��9��e��!r�$��|������r�G'Y���}�� 4��a�J�Gȹ�(5�zK/�Ƿ�v�G:f{�K(�Y1��O�F���U����yp�`�;^��K�j�mn��P8��-����r0��Vc�E"���K������{�U �
�|��[8  ���+l
:�&�
?KU�����֭�,C�9���,��tH�4Yf���T�gYụ�ݳ�8^�68�O+�Q�����ѳ��D�D��*�`�k�Bl�X����G'�&�|�R�Z��ʧ7 �!Ȧ4"
��D�+ͺH`�����l��(��W�?�yAB�)^���)DJ�����h��놌�T��d<B�%���OhL������w�ɞ%� �g��c��[>:��je��՚���(�[�<�b3�`��ʆ���G'��pJO�o>f�u�E�h���Pu��������ʏ6z[<�#��mh��c��� =rd�F��ڌ��<�"�!�_�n��Wl��Lt���4F����]�W�&�q��̉��}���n�����^<�3��S��2��-�~{�mENƻ�^_�����t\-<]l/�k��
"4�}���J�=��Q9i���fw���X<��ivpe��m�Og�a ����@�<}�#]F����������ʼ�觕��N�W{� ݆~���7oǅޅ�8[L��`�Ȼ���L
�+��P)$�����a�e��٬���R���[��8�|i)�SȒ�I]�<r0�=�K]�aM��{�N��v{l"�N��T���9T�ZG�l8z
jZL�\�}��" 1�.=O�]+�r��/)-����Pvm����\y!rc�?�>�w��$1�vx�yxq��t��u4ǚc�U�l->5�1�(U�o6�ah���rn���]d�|�}KǱ8o���*TN���&�G�_�k�{��vhkQEQ��*ThRA�/�@�dx0��RR��=�[.�Om��G�.<��.������C5�ݛ�hJ�Я�vl���x@��b�D���,�5٤�Y��,�� ������tR�Z#\�:2��=e���W�:�+�kצ 3hS3557*#���� "t�k���"Ȣ~=����Y"�\��xdV4�7� �o���|�#f�𞎢묂�c*�r��DUN�,���eI��l�P6�s@oҨ�?� +F�	�`�n븓����P���Iq�PwQ]DP�����U.��Ұ)9/�q���y��ׅ{35��00#�N(x��aM��"1pKk�/��w��m7~��HY�/v��#����T3��9�1���>�K+��V7ü�g%
K
��Kob���ve6Y�61��!��h�ĉ�ￂ�a7�(�/Ev�5�XfP�d��^�_��>R�Yt����y�&v|,�_V
+�?D��(o.����3;}�J^4�1P�7Z�\̄��46�J9i�Q8K�D9�E�%�qBܰ���x�m���RY%���'j��W�`%�$OƝj�}	7��:_�v��L�*���]3�Ơ�
)˾�	jz���*#(VT(�\�GQ�!�n�G�d�p�5�vMH����L�Óh�1�V�K�HWd>�V�'���Y��c��q�Wdj��D�
���jD7�p�>J�?�#���P�i��f��ވѢ��g²kꑺL�%4v=ѵ�)@���O�]2��,i�OJ�����nkSCL�������H.7�?�����G坯�u�_�O<���9���G�럋
O})��k8�Ş��^w�����Թ�\*޶��-S����V��*���mČ��ʲ+���qIy-S�����9z׍���	�󯔴���4}�]�╶����R	R�4T
�rf\7�7��U]TU�����w=���"��T�~�t��lQX��0j���Df�$�q�4�re��j����Jx�U��a�*t��b:����Ȩ�ݑ|�>w��3<٭�Z^+#�Sp,�!4��H��[�
�q����n}�X�`��z�n����m/;'g���~ٴ�+2_�u��M�X(�0��6泷>�_����k-��+[:������Y�n@���ʓf,QY<��7SS�t�^����2�<k��wmh<�	T4&2�v!�7��#�&\�f�"��\4�FM�������g�h�Ŀ_|�|�u��5B�9�Zz�_Ἲ���D��m����� ���_Wt��Kw;JF "��]���/�-�ÐE{Y��~
�}�-PV=�W{@ЮA쮸�a�Eas���*R���T�0?!m�HK�_�A�x@�L�uKdFA��˼ �Y[i����ׅ��Ӭ8ɽ�)|���M��P&�'�����7+p,s�m�[���[�h)�˿�����합{߹�z� 90�A%�wQ+*���b����K8�y���~@�O,=�9�`9@$�	����
f[�[��H�-3G����,bof+E��}�E;m"!�G�/���##�J)���N�U�Y�E	�m�ZǓi/�q�B�?U���Q6��rї�#�sd�����@G������S�Lx2����U����f	��_ń���z�����T�.P3i
�R|g�^�n���휦iJ�AN6�*5����� : +��j-)]uݜ4=C�c�� �l�*��Z8�`0t|ų�C�A��=&z�� ���}�O4�3�{����ׅQf_�'�������e��u����r�Ң(1�2��F���\&~H����O�E��5~���8Z���%�~���~��ǒ�zBV\��Gj��~��ڛ4���V���*Tv��Ҽ˒��(��ڬcC^�"���r���O��"���;�l�&Us���$��uV�0��WVe�ف��^ܟ4&���H�~)H+���\�ׅ���`��H���{:��\�
����^�)kC:M�Va�I2/�X�+/�.6�#����z8����]sj����|�����6D�cZ��Ǹ�T�i�a:�+E5����d^����a�|�a�bVzI�����*�o�}��_DA0n�j[�`�\&�4ę��|Kn�q�ș��I� ]X{&�7��a����/�?����s=�M>g	,����#������T��*���cRV�Yn�$eQי��(�C��RS��i���C��~m¸.�r@�s��-z?�g���v�A���sܾe{|�Y�����-���wV���!��^a�T�K��������+��Ɍݔ>lP0�.��%z��M���B3��|B��@��r��A�������Z��b}��=��#�����1����5������_�R����/�ߍG���41���Q����Ѐ��h�}.���t	Mޱ"_.�����Wg�Am|�-,F��_��]�|,gg����/��ecÍw��D���J��3U�78����s��P� f�p�̴U�T�EY�va����U����s�r�;�fR�M@2��:}�d��/:�4�DM�T�����gz��
�t�e����#�I}U�}b�<������bV���cdf��$u��j��Z.���/�7��|/l&�-k���d�gwm�:�6Lv��5s8+G#&qm�4�*+�K�;^�2EKB���������,Am <�[���	���	����=�����Ox�;�J�[�42c$��ݱ��~3��{�qѠBia��b��)ȨJ7H���PK   �<�X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ���X�j*�o5  �5  /   images/5ca6391a-909f-49c6-8bb0-8f0a302a1c0d.png͚�S\M��qw]��!�,����X\�����w'X����l�Źy��'��0gNW�3�S�===5_�U�1�1����e4�������P�����\�^�^�rRp��pp4p
2�ڟM��SL��!o����0S7��fAk�����&5�!�Bj�p?�r�e�2���nm��5OJ�D�u:-�4O>�����$ܚߌ��Nt�^�{��o����H�9����2��Wݺ`=�狷�Y��d�@k�q�s*���і��4-p|��4-m���>����U�"�aZC'F���-ð�זwgJ�������\��2����Z����w����G滟�_k���&��E�C��K�bg��o��8c��������v�W�?X�5��J4��3�.
r�O�t�����m����=_�"J3vV(���~�E�q"��6��%`�Vd�P����d�-L. �ju:���a�଺������~^���O�E�s�rN��Hξ@�"ܧ��G,`��������L�{娎�Z�@���z���'XclLL��7BiZ,*$�;CG� Q�k0^U�/ku�y�e�Ke�]{y�˃�m%k<��>9�%���ai�Q=鶁���a�IY��m9S\���4#QAl�ǜ�.䢄~R��*�x��z�W��4��7�T8�!�gk�W��퀡ϣ�Pt�H�t���}�3u	���a�`����@�+!9P�I
� �#o��E�qf/WS���V��C)>�A̖i7��0�&!�?��|7P���u$��G�&�<[`h4��*�qp�|���a����m��>�f����b 5�7L��&KPJ��a<ܥ�>�����k��o�������jv���Qs�ba�����!����ߧ�.c��6b����)���p̏fRo�.h(�����u�&� 7���_bYYf2�-���%G���F�U�8G}`��1&������0Q�z;�x���G�&�8����o/�HيH�r���Ch�����8[�G����� �״��iH�ȣGo$t6������B�3��5>���Oo�T��z%孯�W�}��|��-���_g�=�4Q���M��>�Y�?��o���4q2���d U3����rS��� r�����!�)�z��/�K�m�J�c�j*7C�y�S"��V�n�x��dH��2>�M�9_����'r�����<~���/�c��T���C&��R�,���H#�1F�}�Z�O ��^�&���6�HT�d���g�v!Q2�޺SnE�!�g5��վ��m��䃠q�˞]��Q���W|]\���ye;�E�#ީR:bv���P�6F�T8TZ�XR����/Z�ON�!�6h�+�CR�LI�юb�'��,	r����z'Y�^��WI��O��a��g����`g���zo��-Gⲻ����>�ĳ������T˽Om����@:��ob�Ƃ�����\����<��T�G]o|(���'ݤh�:��CYJ�t���2��mH�Jk�<���I	M�|8�G#�t���k�:.��m(X��r�?�z*��C�/[\M�q�x���W��Tt�q�"����>zCY���5��9v�5B��j����>�%eS#5"�f�\����:1<��QG}w&m�k�s�7�FƢ"_p���D�9��>(p��७�W'��,x"���Bo�I:/_(��փ�t�UUo{��N�'�?�����x���U lz��Fڛ�r'��`lqjTz�?�%��A�CG�5��T���B���_���Qf�"Pw7��*fL����]�V�� ���WM����y^���,���o��=m&7_n_㚸\��Y�љ�_��1ݰ�P����ƤF���o���$�Z��J;��X�4���R�V?� 6'�����]R��a���m�݂R?PtPH�N�����Y����g�D6�/| �++͍��=��5k��=�/�����m./�n0�YM�6`ؘ��F����x��kk�|��{PN��B�����ָ9'����Z��
IL��h7}����~�� -�(|���sθ���4+�B5�/ͳ�I4v%,\��d�m��6�ш���7���)�(�&b�4����_*��H��e�������4"�uz�4��0��M��85a2���Q$�����|!�)���ǯ����w�ȏ�qy�Oy��� WF���]ii�2�ϱ�r�r��[7��k��!�i�s�/jmؔb7.�e�6(P�dE�����Kj�P}��$��`I,������,��:g�B�d�ꕾ?�,X�W�F��P��,��f�pNf�V���(��%f��=z-�MJ�8|r�j%a"A�i�z%˾�P��>�Md�ͭ.��7�=��r`��f~��c!��P��ג����k�\òԕ[�����O-�S���;u�2_ .�1��!W��]~Wf����:�J��}8"Ӱ��O��y7�<Ab�b(9�7�G-�H�ͬ9����!~B(˿1BP�M�iL�E���ЦjA����a9{e��up�ޯ���#g�z�^Gj9���}���I���5s�����Eݥb��?�y�����4nʈ�q0���חs�>!NV�_���Q��&�DXJ����O�g�Y��m��ѡX�*�o��At��u�������s�:���a���J��AVN��^S��m|�fu>��I~#ɂ�����-Z���B�$K�jZ�QC�ֺj��H�G8Ͷl
 ���4�d%	�g�Zb���~�B��������ƍ'�̱*�BzɴY[(�?����%�z�}OKK�B~QQ�ÊE2����n~�B������g��V9X�,�i��8��:Fx �k1Ti(�7@=���͵�_��;���xo��/}M��{���_�n���=9w�YwV��� �|�]�yh�}Y�����7,P�c)���!���13�w�--���o^̲)X�ܽ�6:#,G9W��$���`��@����U�{S"�]i�}�aݿry���?V�L[��>������aV�n3��8��ޕx��i*�@8ܿ�g�������lE�8#=C.�DRX�F ��K�C�_KK��.L�ڛ����ҥ`N�f_	z���S�����˸�>��!�y���	%-5x�);�O�6H����m�O�!���6�c�ZdR��Tߝi�.�;{	ȓ���4��i��}��pr�ۓvgm�KN�4�2�E~��'��`��W���|��L,Z���}GD�dV;{�)7��j��`�ȭ3�ώ�T�K$�Ɣ$>��ӷ�RFo�*	�\��)���=�j�O��L�b��˻f�3��{�\SP���}!(WH�d���Za��Q�- j��i�c"K��R)�x�TׁP���?;�J�|	؈�x'��]�X�B+�"'-w�ǄSU:-���"dڋCy��m2���U֢��R���;���|b�Q����ǘ�Q��W~I�һ^0'F$ˏR�H�D�����O�j�R�q�64��STe`T��%Ak�WM���{��$�η=�����nM�eX�@mc��X����w��c�����+MI�A���G���pv�4OL�B��DM�.oH��&���B)�f��i"�`�ؿ��+d_��?�ϒz�z���=̨�YB�=7c���~��_����$F"K�KbԷ����닔��y"$�P��3>�����e�"w��:Ӗ���'�Q4ƽQ������1�
��	���g�W��u#0�� :�{0+>�"-	4�_ns)��f����߸V�fsq_�D�|�����;��(R�"�w�5���&��;,]�$�i��	3"�9�ɛrEn��}[Ah���m'��C��,uSL��$a�Q<7>p��IQZ*wOn���/(Ō�av�[�9��Q�kl��o�����\�����|�gq���Pm3��<�o(�sΡk?̗��cD�����2�.H;��B.ЉB���N�`3C�e�Uة=� lw�IS��O0��D�CV�
�V7��Di�p���	��"�ئ}A�{��B~̱��)`��&W5ڷ��L��l2�_Jhӥ�UĿ�ϐ����[�%L��:$1���`�r!�VU�eP���=}R���D�T���9��$s,�m��Uأ�<Һ�b�;���Qfw��%k|� ��.��	/!~�I��;m��8d���k{�$;��p{�sӧ�W�E��$F�)��ֵ�;��\83�;#��q�
!b�'P
�Tw���۵�˦�`Wxb�����n�D���,d��0E>hN�[�V4�A'Z�￙t��~y�*�L]`Xef�X���؉�K�oq�,(v�d6�\D`)ژ<� =�y@w�����f�{LD��z�l��摊�$��+��.H�p����C3?�U�[��a
[�+�f�uVs�b����o��9�ʄ�N�+�-�~���%�ǻ��7-�^���)�Ι神���<�! #��"�`��J�=��A�:����p與�Ɉ�����5s��B�W���Iϭw��;,��L�C��2�e��s��[P`<6ɓ�A���'�cKQN���c͞	eAx;�s�{,��$wpJtr�q/uz���7f�i�}��0����@#I���d��n��~���G�|˖��z3+�*��o)4���`c�[ky�ȸ�F���G��s!nyu5��-�P+�2� dM���)��ڮ����G�i�����~�x�7�(�'y����2Z0�����Ob��c/t�ُ΢�et�e�ruZo�m{!��94�L��:�ᾊ��d�@�C;K�ux�t�m=�[-*������&l ���cc�o8B�9er,҅6����_�c##	o�2�Mg���zዩ�!o�a��j�ʘ@�G~�AO��bLr����a�i����N���ߞ�OBB�8�O��Z�*�S�Ux�m.�Th�-�� �A����OmT��!;߆�M^-�T��ɘ��R�Ϫ�3��B2�־�{[�-��@,hw\\�3C-Mr� �%�"��W�x�gR�32�_d�ya2?�1)����B��3�dd�B	��Hjd���TpWL+�:*�Tk\���#�&�-��7F��	�< �+�8y��b��m�A�Ζ@��y�������g&��R��� ����8 �WtC�ઊB$�$[@)�"�";�{Q��$-w.�
�w������վy�Ot-�r�S<1BK�� �1(�e�q���ⴆ�J��Y�?i������9&Z�A�k�+��KZM��Q��c��ݺ�u{����5�X �_;ܽ{��s=����hB� �uWa^�d�Q�[���w��1`�����dl)�w[�\�";��W�jQj,��2�2����灎<��ͩ���%{�x3����]&(���<ԒZ$�e�, �gz�u�L���@p_��T#�D���+ݞn�/���g^�Sl�}iDs���x魟٦m���o�k=����@�`��!�Y�:���ʋ�s�J��@|��\a�zɺ�y��	V����W�Cz��r䬰@��S�o)�y`���x��q�D8Hb F���H�.�����q�||�Ng��e�^.�ˑz�-_�J��o�ݫR�[%!������x/�w.ڡ\(�W��t��d낚b��&���d��t�b�S_�DX��Q����qJ��Y^�M`��f�����@�!�'ܷcLS�݈z�w�c�)���[b:���I�P�P�*�i�mG<��܌��B� � 8� PRt�v�h0�蘧�(M�[�t������B�ً5��2p7H�i�7�у��g3�H�{S���]|�c�S6d��9�
��W,�X�j�-N�f^SY�Z���`!��0�x�K��Ï��t�kMa���l�b, )�U��7��-Cvm����Fژ-_I �>C�/tV]:�Z�2��w�4o�g_	㌭`����� g�,M�LCn��]�UY
z*�&|Wd�J���'���}�λx�%u8	h2<��s��� E�%�\4k���Ld4Kֱh�$zϋ`��Q�>$� \"�g�O7U�����枟�ɱlpLOq�ق�X�x�9�ҡ-h�!�d�5c���;E�hC��̶�|I'�X�W�����BB-����bN�MkLY��)ge�E��e�Z]A�/�a��j���-����V�BZnV�t8�ҋ14Fѕ��wS�}`)�Ǩ��x��xx���v�͆��d���0k-��I~�9�;��C���\}zKl�
p߷��"��c�ʒ�#!�QI� ~D�	�{ݦV�d����|��c���qsy��T�j���c�K����M�]^��c���T����C>E"q*�s�{Dm�R�:ؔ����
Joxx�V��M�]���� n/.�zo��{a ��(�?�8�h�u&����k���\=�;պ��{�dNO,��@P��mu�?&cn}R��-Umo��WEiI����ң�I��Z��<�|���dƍd^0g�i��b#tʷ�zB�$�Z�0�"x��}8
'8��Iم�J��R�̘���r4������lԵm�*��CG��(:(���>zp���]��V�?J|����]?8_��y U:��N�~����2d�Qh��tP�k�8Sy�}�~������O=Q������o��؈�|�nO���:L[�[���ܽߪ�#��;3k�TBs'E������s>�����9�P�㠆��VY��[�G�<��&1��C�}�U����ͥA���%;�J"���������5A�j^���ĉ��P��3%�2t�
'�Д�ZW��%����D�/b=K"R]<V s8�|[q����&W���d�ٛ�6r�>�3���^�2ڝ�����QrUP���;����sa�S��p�ǯͷ4�F���C�(9I����L��X���v����3M4��ZR7��b�r�gG�6	����W�4���KЅ���s��qࢿx���� �� ���Nd��/��x������~Uڥ�%�Q�Ļ����:|��Z���/�݉v�^��[��u��V�m��1{�r~�fYw��X=���dm�D)nʳ6�D��H3�x����~���X��:��mW�h�< ���!�չ�Rn.&��r�jV�?��[���#3f���Lы�	~�ﵤ����DƱ���� ,���$�ِiHz@`
�6F��u�6N��e-	ͪ�,��d�3{&��J�	���\�!��[Viu�ʇ>->1Y������'�⺴��F�{Chn�Ca�����F~T��\}g�x�����}k�JRC�ח���� �;�VmUY�@�R��17R��/㍌P��D4M���ǩF�O���1�*s�ּŘZs���B�_=�у*h)�RA�i�׉k�������@T��~��RI~O�a�S���;".O��u+S�{��=w�: 'w�B>�1>�q��Y���9+�Ӥ�Q�E� B�,��UO���B<�D�D��:�G��;,&Xo�3��Q�r1޷�}PD�^��7P�D���/
�sC�l]BL�6vt�c�u��'��5jM 5�נ��@K��/YwX@�aW�� ͮ����f�XǏ����Z����Wg��!S�b�@��LprA�#<d,��,����ok����K�wX�)�]�@1d���^���;7i�.�R�X(3`{R���@+��}m=���Q�j���Ne��K�QF͌�L��V����qZ��b��8���'edؔ�P��0�\��O3�f�̖�V+|0����������j�i��d@�'�G7~Q����?�_��\�������
�R�\��yC�{���h�DN��_��v��Ĵ��W��C_���	1U�=+@[�E5�� �&U�4�s���ټb��r6�(�^�ɳN�=އk��i<��U��_����0��U��7�O��4l0'�6@b����Z���ƝUa�bE5&9IZ�8��_�![ p���X�yP�|�7�����~)�� d'�:ؘՆw�Ҷ�:�2aqO�~�n4G�Ԫ���:��1�ڐ��l:D�g!0�q��y�Fɟ�*�;�*-���>�V�>
�]�N�HW���jf{����5Q��V�9{j�$�X88����0��b�OeT3�΢��2~x�-�v����o������.l���2������<�-�������F�i�6���v�*b�q�@�}ҧ8�>��^��o��g��?�k��-�2��6��7�%5듁�&�L������+k�ǒ(�nW���5Ċ>�.�6
�Q�ݿ�8J6���(��!`S��)�����=����Y:����V��D��w��Ox���oJ��H佨)�Q�!eK]g�\��5�c�O�(�{��g�&�o��ޟ��w���~��JC��`KQ�X@��;m�9ب��
<WE�)I�P���>��;5ϻ`�b,��-�'=�ϙ��
����������V.��̌+�Up���~��y�[�5tܒ��Hg)�K0����HdK�����|z���K�8�r�$w�Hg���B� �L0��f�>�R��9F�3�2���J��<}>��Pܾ!;sZ������I�*��ٍ������;����@�~$A�S=?H�.Ƽ�4����$��|W�xT^�X�r>�a�7��U�X��b߿Q�c����L�t��mh��jI��-��X2g�c`�^B763��V��D?x�c�"6C�����^vI~�;�8\����IƗ�E�T��D)���n��`]$GC��q�W63\�*N��C��V�/̺�fuK.�QO���Nԇ���U^4���<���x�Xd��S�A�ZZ� ~S�&KbfCv���n��=z�^3#�A\Ɔ�е�{=N��A�f�?�~�����ɝ�IdV�̲�>4���T��0�O���7ɔ �ю�����H�eC�J��`"�)��f�n����ڈ\�y�O�
�a&&�9��s��玕kN�	|N&���ϛZ�|��Μ��\c�,;-��Kg
j���n,����▼�{#2P�bt#��+u<b0`�P�ZҶt����}����n�q(���������c���i:o1P�zt�]�Tփ���˪ �5����HO�d|Q�کlUO^�v�ۮ��{;�AI��#�Y�|�����bcP ��^o�R����;�b#�eyo���Ѻr��z��0!|�ܣ0�{���%���l��5J��`��q3�;���?�깓u�4{�A<e'�����5w������!����YV��U�p/�8�N���O��K����Ŏ�Y��ˇ��2e1��F	��NV�'8<1���p��e����;�B�-9i$:����pv��cp9���6h�:?BS�T��xZ� �3k���w���=m�\������9�d�Ǫ�/V�l~����̔�l�|�c�.T�=4Q�+1���e�L�@�^V�b"�s;M`�b��'�J^��֫��
e�@7[����/��'p)���m�{J���U�q[x޷.�����X�����`�d�(EHs�\<�=[��B�֑�VLL���P"E����8���=��Й%\-AK1�ϛB^�[��09�q�/5�1�4ҒK��I��{���
9n.:�qY�񌇫��e�}��Eү����(�WC(o���;���I�?�Y��w|�;(�3���g���$`�pA:��D�p���Q���Q.NB���H��:j�R����I�7��v��V�A�̹�{��j��2��c2��Y�D�6��T�
D�W4w<�2�t��|3���_Mލ��-d��ϡE�R�����3������Ƙ ��x�m�:Wc�)�e���D�I���GFJd�����DI�Q�O�j������*0&}�1-t�T4i7�9�)ϭ����&�`��odq~u^����$6�*,1��;��x?\D2Sm�H�诮��	�UPJxc��l�sB��)���������n�?]�}T��$��M���;�QS]�u4Yl��@Z����14	�V.QR9zDH0"!�5��9�L�n!�$g��>}��14Tm�8NfZ��O��d����� ���'�(�l�/�fL#���P��B�QWR�<�id���)<,n?��X&��Ox,�xv�
��L
�]�J*}�g�/���
"g�MKS���~n�NSoB�=9�`iҳ��Ӿ��+˞+��T�F=�x,:�@����m���/����hq,j�аsQ<j��4������Rlޚ�Y+E��$@��(�o3�zR�$�	���gѝW���Ӝ��ِ�(x��(����`��.��X1q)]y��
�2� $M�46�KAb��G:���L�[��d�&ʡ1���k�����c�zv	�����_�"n������ċ��b�fu�Zں�K�Bc�%��θ6tC��S��\HD������x��v: �wf�����p������5'[�-G��d/$]�P��0�� �ڊZ�\��L,I3���dU�'E��m$�&9��Y�X�a�>�ރړd~���DJD�*7u럀ܐg3�abJ������l�����{wt�)�5Y�[^ߺ-��o^�{��^�)��3�����"1�x��4��G,t�+��_c�F�hX
v��~LQ���V�Y�����.ӈ�#��=|�����[�&�/7���~>�~C�INl�4�\�xƫ$V6���E*�%Sh��3^e?���?O��
57@hO������SoG]�9�Ƨ���:�����Z��Іj#S��o�cm�>��/����}��ȶ��Qʭ&ӣ������2W%0�� q� ���x��V����f���_UNN��Ж��D_/#��c�MP���99GYV(��Q�XI5AH�A-�����L��[�QƦX�;It�V񫝒�K��#��6h�p>R`��?���������zgc���7q���@E�k�[&���K����e	�6��M|�81,u?xQ��1�����V�����jAf��Gdo���b�'�(7Et���-�q)ԭ.t.j���F�UF���wɺ37�h1ׇ���K�ܫ��$k��yf;����	G���	�����p��/���2E���즊�����E�aH����	�x��)�\?9)���+�HSZ{�ǧ�����'�o-d$�F�[�ϱ�
��������qe+=v��2�	�(�lw���ɯ5��oe�o횚��d旸ڳ��)	�����vm 5&I���:%�|�P�tS%�bJ]A9�����}WU��f|F��H�����	�_�g�q3�d�s�"R�D�9���������6P�1�B}�������\�.��g�9�0�0Ѹ�h�c�R��X[=+<*�o���x� J��[	�Yyֆe?�@�H<��l��H���&
x����������#�_ɚ�2ّ�"%�7,;j����%i:�5w����E�}+��O��KY�Z�̏Z��V>��4ݭ����Y�/�G#�{���Q�����g��9R�Qd�e�T�I��a�Q����G���1e��.tr�ǀ��p������)�l��Y���t$2>�
�m���o,��H�F�RoC�}7gn���$�����=�����^M�ˤM⧻w.m�yl@���+��"���OK5T/R�VOq~��\��+0��e�tW:y�]_]-����S�����-ǌ�X� 4n��` l�1���vA�~�)��,R���5���Y�ӪY!;�v%����1q��fr���W��uDeE���DU,��.OR^<߻n��$OyQ��H�Z��q������� ��n����0�^յ���=�FҶ�ms��a�5(�:T�U�/@���^iU�u�� ���G�0�ƭF2��Ѯr�,�WF���L�h ��-wt�����lO�ƔԾe=� *��\�+O
>���M]�9ܬ��دb��>Kh-`��
�=j<�[��]g������,�j�I�)S)��p'J��:H�ڻѫ����b�� z�plJ�ڪE&�w��u��� r�������XcB�u�����e���2�C�b�O��� ���3/L��쌃���o"��@����g?w�|�A.�\.����o�TR�WD}���f�Q�"�O�����;e�w� ���1�b�5QG	++��zy��O��ϰ ��]��(�ʭ;��ý�-�=/"w�7B0���kK��CQ��jP�����������KX��7+����f�n�䉁?��Ʒ�N|���� �-F�),�|Ѳ��.��I���t����5�_x��P=r꘽y+x)��fS��X�8a�a�ߞT��e��Q�č-Q(R�#FA� �qW+1�ö�Y��ō�it��c����[	��Gjd��ʃ����MS3�P���=@��v�ɋ���qa�iI�E�A�{vv$޴�X��B�4���-�>a^��e��<<����
���=�_��3Q+�?8�v?@��i��E���Z�,v��|9��t9\˂A�X8�%�D�Ǝ���Č�^�;�'�Ufy(�i�J�����O]��6�)#�'M+	U^�2Rß1�=MW���V�X�H�ϥ/=}ǯs�u�Y MBЩ�Y�Lے[W\_Bs�PZ]y���|�%8�e.�R��(�����n���^���b���G4n�	B/9�����8���������$�=p^>����������yͤ'�����ӳz蘘&9[�Z"���?P�)�����Ȝï�}���ߚ/O�|,:�@g�_�CUF��c�;�J�����{��Ԡ�!�_�u/7�v�k'=o��e��c�Yߩ�]����t\!ҭ���N�
���.�$�`3f����T},Ƿ�����lA��Jd�lD��`�i��0i���;f�b��D���zZ�&:;��,�����_�Zח�t_[vj��}�K�@����--���I�#���B�����F��:�^���A��d���&� ��K�_%�?��E�T?�	h�ީE{<C�._���!�c���P�K��������u������^��1=b7� (��6�%���k-����
�*��j�T''J�c���ʶ=��������/_?��]�RO]5�[<��|UUs��?�n�e���ۛ�e����9)řJ��?��7�^y��0�|M���a-j��f.ae*d~��߯�e��CgטK�x��:}��J㥣���b��\�]��7a_��/)�lꚂ2�:��H �Qg'c"�ԡ$�#��շ���U�;�N�߰#��}�|+���"��견Q�Dv�M9$�L�U��!�+�nz�;����������A�f, �u��\����M�\Y���-�~�8���Q�W;��'2�=ǣRA��mX�C���!o�jfH��op�YU�)���PK   Ŧ�X��~��K  yK  /   images/7ac84256-6e9c-40ba-9a9b-c812e48c1c94.png 8@ǿ�PNG

   IHDR   J   �   q�   	pHYs  �  ��+  K+IDATx���dוvߚk�U�V������I��9�)��5�%�!+�X�
E؊����H1�P8�3�0G�Br@ ��. �n4���k鮽r�|����w2���*k&�_ċNd�[�=����s\�6R��Fl�Ԉ�W���
P#�_j��7�'�|�E�ق���/�v\��b\.[�0��(j{��ݮ��~�'��a��'D�8���L�X,������F�X(Xnōb��@��>+��Z`Y���o�ߧ_�$CG�������;<ϋq=}�8^.��t��j��gϞ���P���7^����JG�������lGD��8AD��-
m|�:������0�H\7���4d;j��n�Vw�^/8}b�Y��6V��g>�~�Z,��ٹ����v�^w	�v�N�D6���n	�q��§O����88n{	MN�t^Xbbb*�T*�f�V���w�y��^|��W	���Qo������Ӌ�67�.	+�H���-:�]�,���+�����ZM�z=A�)�Nt	�k��K�繞399e�54��	��	�b[� ��H�c�V,ױ
���Yx_��4o��c�Fkkk�����|����C=t���2v@� ��������?|�l%O޿w��๾Ł:�F��")y���3lT`��W����q�0G~p��@���1�C��V�����-7�����s��1�[�:33[��:Ͻ��W���㍱�^�������	 �'��nz�D��s�P3`���&Q�u �9\ 2�@8ƀ���}yK�lv����!ە��ͺ�y�x�ɋ����bcsm��?x�?�ͯ`���Fc�D����O��?y��h,Z'OJ����b�d��1|� `�)�J�����ku�a 2@������̀�c��h��=���c(�*oz�hܚ��!�H��ck����Go޸񟀜677�_�]���e'W~�B�����m�s!�����@���D��6�.*���ꀑ3�R�E$'l~~V��m��a����+ݼ{u1I.�X��� ��ݻ���~�[]�����[���?�C �sӁ)ÇIPo<@�E����0�>�f �տ/�����*@��KR�,.Y/��[(��7�_?�&O]#��s����<��/^��������w:	�V���xB�Q�����|)V$C���.��d��C��k���p���q�p��
b�uR&��.\����o~�_?���,��H�4�N�\	���zl[wH'�: _jY+��x��a��%��]&f�uyM���L�����'O% ���$�c�*Ւ�h4'����!ځ����>�i�T*.�{�J�x��k�6I�';�D�������>p�ɀ��2���ߺ^�N(���y&&��C�'�J�����uq6��S@�3��۬?N/j��Hk�(�E	u$�(��>h,�pÚNF]��a�����x���xO�X�~�������X�Ei	P��եwm��������c �-��t����*�ɀ�&�ӱ��Iəb6�t,�$o�>��Fԣ=�_�Z�FcO"2/�+�juR��!�N]d�����W����˓��w���Ki�6�v�t�굯8��.�,Fl#ꩧ����O^+|�;��f��\��l*���5�9�	�+��fj�\�@��]
VM�X^�;y���/��L�E��d���0p[����o�֍ۏ�KU�%;��v����ot��C�Y�Ӌt��ӟ\��
y>���S!���v��t7����1*�FTڼ�O,]��҃H�t�֓VV��Ԅ�Z��p��:�M�Dc����[�uO�<�%��dfj�3�! ���@�RGI8��h�+���y�� �f�纮���J���3s~����^Z�$����7;��8�|-��ցi��I�y6��t=}Vڒ�m�و7������N�'!ѻ#i�����h�dJ1s�N6���_���=y-���$C귷��Q��t���#�����������<�	�.���}r�0��� ��3������&��{�o�%`?�`�>�����/<лN���{�����8q���g�ݤو,;qڝ�2܁���u��Àh2�<�1������y	 |0��ϟ�?���?x��W-����b��~�����������m[	�S*D�\Q��������wl��̦�$�Ml��3�R�jU*��a����텅ʺ8D�gn߼�q�0)M��I�
�S��<���%�os�y�K���1/Ͽ��Ǥ�0_�t�+:��a$�Fe���D5���-�t ;���n]y,�!}&�7�ә�0�ӥLr�X�X�k ��FJ�M��,,,�^'�}��v;��&�:[�̱^o�v^o��2�9�0K������~��}��*'�V프�8�R�h�N�G��X�-0�^��8}]�� ���n�q3=��[&6Je�u2�t�>��G�w���G�wH6���z��&����ba[��#���^^m)���ޕk}[.�<�[�]gz����c��ԑt��9$*����G-�aB��N-��+��͂~ml4lzy/١3�Qʕ��Ey��,S9�3viP��G�	H�c�O�(����0�K�����Q
����ٴ,;�{��R���?�@�ac����"�����!�h`�a. 433#*�
t)�/�V$#T�;ׯ�7o�|Ĳ]F�-[D9�f2���%|C"��^�0�.9�=�49���-$4�
�q�L޸q��	��+++�:u�5
F���M�O������œ'OK�y�R%�W�s�~��δ����;5b��tJa`;{�::�Cc�����~�{�����{K��;����/��=w�{��'	i����M}*O��?�� �Բ�)�U�rИ���"n.�D�fV��O�\����K�:q�d�������0h4�ӧϴ�}��Du����〇d��t���#�G�ُe�hy��t����9�@��j����I�"��Л�c��tmx�^ ���BePa9��JC|��s4�n��o���6��B������8��K�X�Z�b�������&���X�f�%&_�t||���v{Mn��ð�z�N�
S��b_'/�Xcf@���H�l�L>�sx�0��b\�>Dn�:Jq�)¦/�������I��]�G�q����fj�:)��&�nj00L�2�r��w��V�%U|��;;[���J�������U�dml�z���{K��mnn�qZ[[2��Ѩ��t^��u3�ԑXid����Z֙�T��I<���9¨f�T^�K�:�]1b	P���烵�ť�����w���[[;����p�q3�!���7 ��0f0 t���\�KI4�����l|��ZX�����^�W}���g��ݱ
}���	��Oָ;55!�5�X}�c���7�4� (vH���I��3	2��$gF���~����|T���i1��h#��l���8������R?fsX�����r���¤�:���q'�1�����f&
^� LH���t�QE���xI�ѽ�W��d�`Hש���H%>�g�J�G${�'?כaA:��w���I�{���GbS'��E�	1��Q����W�XR�b�_�v���z�b�p�(�S�s��:_��{]3�\�H�?�B���� =�Z�$ ��Ǔ�S¬�T�Ȁ�N���l��6փ��P�&̰�S������c�E�� HG�Q	1�)l=zí���d޼W=��4�����n�sy&����A�Ea,�l��Lz��|P�R��v�(JTH2�^h����b��%�0>��v�>NNNJ^H-ƥa�zk˨7�ͨ��������-8����5��sހM������k�40s�Z���O�<�������G�V��dЊ�ayQv�)�06:�J�9༖�u�fm^o*��3��ҩv��j��o����v�N�$��[@>�ŋ×_�]���{_!E���ӟ!S KK˙��1J39L(���M��%oJ�;!� �;wn�޽{���N�u����=��������t�lt2���m������&�9h���s�����Mf��z0
Rܙ���������w=���c�>zoei͚���[*N�\�Z:;�L'�N~y|Jh�)�+�y6�����}a��J�k���<3���G��$W@���f�����0�ӱ�\1�����2|5Dv�ϊ766�^�Qr�#-�*4�0�15c��b4o@��a��x����L���l��`�8s���i�v����#�{��%���>z�񥥻zihY�`�G5Z�=<d�b�y�{�b8u@�q��k��xm�w���O�گ�.ѩ�\-#����o\y�ը���ڝVk�4[A���.P13����a=&9�)�:����YBڗ�ٳ���>Z�sFl#���٪�j�������w��Ƿ6j3�JI�O`�b/��M��!���`� �6�!���=���k_��W�ţ�^|��iMmd�jmM���T�ި�c��0Rk��%O��2�:���<eJN�?��,���o`X�b�ߑ�a+����s��i�M���{�A���yX��<,�7���S��H�ǔ�KE4��Z]�����,��An��<{��$Z�y�x���y�&0,K�~I��v��!`��v�cĈmdg�P�I�����]D^��d��ޏ?�u 󞵟.���-�+����F��ɡ���#^g��M/ú^���`ny��a�<�S�.U�{�k�X� I���#�8��t4<
�>�7b
��F�$	2X���p��d�<W�������H�{8qG�zvb���^��K�r�5]lb_��an�s�߆�<&>�9�x:�;sG��v,�dwIQ>�r:�Ȯ�nt�6}���)`�}7Y~8�5q�S����wnr��I����	��A���ڪ�Ͻ�]C��n�K�.>���ȠL$C�;�A��0 ����m|-#�����Dv����㯼������u�܏���a�
_y���׮���)� �ǧI�ΡA}��E�ʐ��p���$�$ɒ���^�V�����?���g�z��x��g����Οۺ����z�8i{3������=:���1]�6�qƙN@Vc`�����z�Dt��)�T?�@2�<p�܊��[���XY�/����`�eJ�|�g؎v݃9�k�|7�������x���i��	�Ľ{+دgC����-^��;������<����6,v})��Ò'�����6i��I�۶ƹK��t{x��&&�byy)�z�b���*�T
��a�0�B���������iy< #��k�zawww�.)9�H��u�V�ڵOol�̀`aA_���2,�H��ӲM�jb���l�p4+Y]]�_~����ַ�~G�P��_�?���s����$=�tl]+�CRy$���c�;��\4y�])�H1;;+��@v�{�?����?�����sպ������]���{_�җ���?��g67�]��\��3 �y��mSL[0��Zy^35u�KPM�ﹹ��/|���<��3����zn߾NO_,��t:r� T6�bsy�$����l�<�օŠ:�*�)�l>� ��k�Q�0/��R���b_*b�κ����f��NR�}�3���Y�|�AX�� I�ޣ:�p�2�3 0��X�'���G�$n#�z�-�ZH�P��<�3d�o��QZ����kE��Xj߳�L�`�J%�x����4d#�R��a[��d�,�<�$��A��Þ�[fS��T�S,. �G�M�k�(���Vx���XG*ڄl&kss[����ɽc?F=L�&����f.���d�I
&~��
�Rq�6"�&�b���
n�]�0X;�Im?>��<er�'�#��y&�ar�����W�
��F��/�W��qWO���^�+.A�j5�ر�������=��i��ڰ]���+>�����|�u:=�&�X���H��O�w����\*M��vj�Օ����L$����(�����<��d�H�ӑ{��ML��V�:�y��sp܍P0/_����_����KW���y-i�G�^[���V���$���/hqf�Ș@�}$��}�}�����Օ����������qw�♻���nDw�.ە�T�Qux$��5ȋK��8-�)�x͐-�Ph�y��P��v�q��tEƻ~�����;,��̸�~�[.<z�G?z+���:R5H3Rn��mJ%���:���Q������ԟ���/�����#i�LOO�w�v7�s���OH�!5?I����>A���+���T�o�Y�)� �7B�Oڻ���C��	'� !-=J+1#��PD�^S��
�3�C�i�餧�1�R���[ٴ��	��-�ψ����tNH��)n:��G��������9P�4�� �󀕧3���dL1�?�PG^�o��8��3[�����	a`�ۡ����ݻ�4I�34��Eܽ��[�������w�ίO(v8!��[[���<`�Q�I��q}ˬ	p3_��/��*U�Z��$^�zv��t�����7���Ԕso�ve�̢�T�{n��.S)u��m&`�a�����Xϻ��k��QȢ�z��-�mZ)�ӳ ,ο~���3�=��c�=�����xw/���ܗ��|�v�O�._�Z͎���N/_g3�S:���<�bF�X�U?�\�OR�~��[�%}��r���fK�*��3O=����m��1qd@�B;��i��"q=b����BWZL�����z3vN��������k�^b�rj�^�c�s=O�|�6�
�vH�+�Z��-����z����Zr�89ǝl>F�$���%�e*�L��&o�%�Z4\��j�P}q��ǬH���2��I� ��y�q�8}O��"o�Q�C���B'�����+�qWԹ �ɺ,V�U(������d=���Y:3fI �$��l�������k��PqG#
H�8I���!����,��zo�ԁ��[��@q�k�pg]�b��$ȃ��D��2%����vF��r,G���~nA�S��<p֣nT�˓��3|���wvS���T/;��b�k�*�ϗ�� B���x��/}\��ml�L�����u@�yH��d�A
2�] ;!� ���Uy�\�^ej�|�%!�7�����6�5,Y�
|4J�\L��D��+���>K$��n���,W�0���J&c7U5�@[�Q�X��p�b��C�n�[��*��$!��lj1�^7����C1��s�5{��ً�۝ ��Ct�Ocj���ɜ́�'Aϰ��Y���Lu���B֗�r�GLdӈ�YH�t�zm�x4�ň�`(�ލ�W�x��+o��]<#��م�h��i J��miz�{X����K�%%^c��L��u�i�p}RO�E?�R���J�n�j���Uo�D�������f������D������.<�rz�����m��Ïɥ�N��� ��D7bY�KH��ax���̝^v�0�8��%|��ہ��!�T��T�6ӗO������Sb�3�ʥ9g�'�!���76&ӓ�}����/�eQ�
bm{W��QAH�Q�K�nf�< � kT��@�Ii�J�@���T@S F���N�5��T��w�9$�����v���&��S,���p{����f�M�Z�'s�	�D�8Ba/҈�&&E���])ѽ��9�8��n�,�T(.[�W�T ��e��)1�	AŶ��E��&bO˫woj�zy�ر��pN�o��JA�)�d��4 �-y������1�Gj��}K8�~� �q�wl��i���I�oW�x�)t}<�R��!!H�R�6+�#�Č��Q,ׯ]y(���`�XG,g�^�������������1���'��Q}!ak��
���$�ecz\��,�>���_�T��G�l�Pׯ_������/����'N��Sǉ��6k�4��`F΃g�b i��3��s�4� �ș�+�"T��0���RYj�:�m��9���aF�Ν�SO���2�������3���Ok�.z��w�SPEd)�J��!���\�c��e�\��@R�f[�\%tdɜ�@���J�����\m�����4��|���
E�i"`�,�)1�~�B}��	 _������?���/>v�'N�	�F�g?�ٰ^_mLLTw�?�=dK�m�&)d���҃��T	6��mm%�4��Q�f�P���fٕ^Wt�*A��%�bYL����A��+�Ixt�[�^暪ek��$����It؂ޕ�vW$����r�!t� �Lo����=����V�'���-2����	B��XQ��X�G�e0`�R�"V3����Mjp�D =�$��\*@wIO�s*���ltD�$k��jy?�1��2P����^�"?YN���L_�I���r�H��ɜ����h��C���,��[?L��$A�A]L�̊p�H�=D�n��e�&q�U���Vؓ *����	� J'�l�^�+��e�����@��Œ(TKҟ����J�*J�"�Q�&w��[�D�Uo�R���T@�����-��.΂���Pyd@3w���N��![�mwP��$
�jeB��u��bUZ����P#���V�M��U�̀��0�'e��ب�N�0��M\��[PYj#�%�D�,�K�@�
Q)W����\O4�Q�҄)��u�=Qo���
'�@>V��ͅ�b�&��\7�}�^J���dw�S�gٱ�RUc;aW8�X�|�ƈ( Yt V9{;4�6x\H�	M�45B��a�Qb���F[��z	ن��%�;*!�`��������D.8@�a�#	p�4Q��.������w�!�H��lm�M�솑Et�6h^��2t5[4kMi� �f���HD�^��Z�`�����30S�B )��@�'0�c��nؖ� f�#�� Q�Q)�yiv �
�Yr!"��C���O�t�.�]���F��tcb�8��fs6�'��(Dn�ْ^E�:��u�!�י �H=p��k�ds�o؍��&R�U��Va&P@Q"����9!�&�;5SbO9��b�~�Qip1!�E��2JKG�;C&LXhy�S�=��:@JU�D�M
#R�c ^�e����&�L�o(\*�mA��]�\�+��旄B�ÈX�=���}�]�q�ir�.� Ɋr&^Q����v���4 �a#�P"����߳�Np���5�֭���Ϗτ���b��?n������X��,
Df%�8���p��p���(,a��i��L�����[(�4�l� �C+@:F`�tO���(�J/�����dǸ �@w#l�+����KOt�OLb �L^I���.M^R�������Z��ɓ߻|��'�88}��n����������_+�;� q�L�����y�TIo�d���g���<N��"�'��B9�jt>��,j�r�IjC�0��M�#,��ZԊv�=M`L�(5��B6 M_bb"'ع03#��n���~�����U���Ϯ�[Xk�6Rh��]���|�ؼ��C�O�MN$�`��N�\:���h�Eʠ��B�W�J�
 &��@I�� 
��.�b,/�����8��`
 �I%��Ä 8�Q��@%jp�2Y��!=�\t�c���O>������+�F�(<p��Mϵ�������([��RC��!�sZr�&���qJE��1@��RXҒ�N$]��_�:�N:�0����˞ �T9DO��8i�t��%=/!��u�2��S��-y�M�mF�z��;�J�A����;��* J�s'��+M�+����0L�<V�8R�>
�sKŎC $��ɕ����`ҖZ<(X\�Ws\��Z�ءr$`�Q���jםN��:���h����)" R�S�\*hA��(� ���X^J��]Pb;� �K$,5p������^�cΕ[8:�~�hRn!ف\����MLT��풀� p��-W�WW�*_]��^{���÷���G��6	�X ���C���R	�cɭ.�$P�	�[Y.%���X�A>;�,%��D6�$M��(;Ib&��P+�N�h����qm	�V�K�M���jh6����=^y⹛c�����/ޚo6[�'OO�JƧεЋ�ő�n�{9�D�n�uÔ��r�����$� p�EK�cK/��NK��Ldi���}(�8�f�aSAX�'����k��b�9ލ�.\+���<s���~����^!����_�ӵ�P�
�٦�Y	M��IƖ� )�5	�M�:��Z��$�|L��^Rl�K�}�'�*$��P�X�I�y7��]����o|�k�痿��[��x#��n~J_V;����$��^&\RI�x:��_���%�Yl�5���L?�J�Ʉ�+���a���%M�mp��)l�m�������CBh�\��}��{�6z��Z�`caL-��/�pB����Q3������z$��{�x�%1�U<[�I�D�~����T�Y�B�đ���
��Z.1SK�r��җ���t�~���%��j�^ˁ���U�r2K�}�h}�cBՋS�$ͽ�!�*�J����¦Cʗ!+�ĝ�2���1��
��R�0��Q\���"�G/��C���x5���4�p����Bė\��Җ�?R+�W=�d�kkKx0�D)�"3��l�@��hB�?�\q�c� N�����h�m�Vj�`�+�]V-��h��Z}a{�x$a?��UV��9��	sC�=p����|Eg�jЃc�R��͘�?CZ)C�LT�]*�e�i`$�')�~{f�
:#���ݻ��G�0�8�B�ب�M
�e��cEE?�c߰L?\tG��;0�f��&�A!=��۽8SWn\�B�T�^����j�D0�WNw_��e0 Р'q�,m��=����|x%�I1M��?ϡ�(�UE���B�E*H/D���j<;;{���Z��p��7�������̜X��я}�cK7H4st����[F�
ց�KY���iڒ}�d�z �k���_����3��M׼n�{���|xu�z�嗽��~v�ʲ�2;t�g�u)����B�a
1��y*c 阢��c�Z�"�Բ������_���GydA�Й���'�x��v���K�reh 4fؽ^����rp���PD}W��Գ����.zcc\�����c�[)W��[�N��j�v:������D���&DQ6BW�lR�b�����e�XL�y�f"u����[�%x�U�W��=1��=Ǳ��rgzr�&�h��juf�<,%E<I&��@ژ���.�`3�&�j����AY��>��k� ZG�d�� e�c/-���C�ccG�����cT�^�XYYy�#xQЙ�E��d�U[3ԀY��σ�p3�Li냮�:!u#�ң���DV��*�A��V3&�y����M�?��#$	P?��ϼ������}�ϟ�?=D���������c�V�E7�m���}���T�$��셑�jYֵ�	���+ѵ��?�%�b�6���bw�����ƵO��W��Ul[y5�V0�hQ��r��kpX�������lK�^E҅����Tm�Wƶ�!̇˛��X�R���b!\��n����������Ϝ�m�P_��W�Vks�~���_z/mnlˁK>�/���������";h�j�����<��@���4��䔈�1�h@,H^��K��8}����}�̙�e=<�:;;�N��>�j�
�)h؎[�c��T���o��ٙ�
K1��x��DK���M���,dGL�x4�;�p$&i@��
�k4,�&{|Lz�t}�Qw�� h���	�0H]H�?V��:a5R:a��Ҁ�ey��K��H��+����U}��FQ��d��^L]��5g�&N�<�G��n��d�| �(��qm�=��� G�����&��G�
��MR�w0{:#f�N�(fU��L�+g@���67A�i�y=��7����<B��d�� �<�a��qɌx�Λ��䦓c	7]u��1��%�n���J?��m��	��n�P�ٷ���$o}�kR
%�]��w����S�0�b@��9����3��VT���Yڗ�Vv<�O���S�?
����[Q��m
~ĳ�o"ԱKw��>&����p�-���@�r�z�y��	U����>�	�����A���FY��*NQ�����%�כbr��Ǚ�Y*��F߷ǘ�$Ƣ�I̴�Z똄!����4��_dEzIRiP�-�_�j6��?��?闿�2���(:R��~6��2�2i2��Y�����<�}LJW�p]�Օi�Ӻ0N��=�������ݭ0I���e����v��ӛ���+?��O�s���RQ �lv3e6S\�c�X|=o��In��u7������ufr�
�*��WWV�-aVB�<�wy��/���B�����4o�X�=���R's!����ճ ��yM�U2��
�t�Ɠ��(�Z�Tz�O/���S�Tc{{��D>�h�Z�����ׁ�@�d:�M��tL�=r_����@Pl>�q0�{F�B��;Ns�? P�V}V1F�(7]/��c1��k2~]E�c�l����2�*`?1�'�m-�f�
������� 5��i�F�����d�ĝnKbB���P�@Z�=nI'KS�ߺ�ƿ�8*�>V[J�qHfIK���\|�8)�#���S�z�Ɠ����F
������?��^��D=����3�\!ݧeH�TuFku(�b�8t"����ڠ/�2��Vc��	"C��³SS�+�����v��^�ݷ�y�μI���Ν;8Η>�p���������g��7"Zw�/Y���(`y�τ妣��|������B1�v�� L�R;'X�	?v|���ֿ|�_�#1nfN���V�c��m��t�رc��i��N5����z�KQ"+��3r]ߒdLMT�(+M����[[[��(�m$�W�dv�e��+6�9�E�<:͵��JD~�����ޗw�N�y~u]������ʝ0��x���II���0md@��fw۽Iz���j5U�[RE>y��u�$8��*������L�M�Z$I�ib���y؝�uHl}���G�B�0��ѸYJ���nJ�37� ��6u�,��z�c�����	�<�q�5v6��G��g�,ͻi+�!?�$8������*�𣩹�q�$
ܨ��F��������S����u-u]~U#ـ])���?��z b�kY~�H|��� �����b�u��~W˒�	��7��HoL�rIS׻�0�o;�Q�;kis`�]I��Ť~�.��B{�E]
���!0
��Q�V� 9��=f�@�L�|Ӣ�LǠ��!� �l!2�v�w!�[��R�"���JVWt���ʤ4d>���^�A��zўg�@kÊ�C�`�����q��֖u��B���@ش}4�d���V�
�n��Q�W��^�^ߓ;:�5�ײ�k1�Κ<�+26��lkp�R	pX����p����ʅ��$���e���W,��n�3�������juZb��!ڤ�aP�u��ߧ_�_oӿc�cY"��rx]�%�!<��_���v������wŸ�bRܚ�O}���T���جV'�Y�O/g���t"��Ub�p����k$&i<y��
�O9.b9aY�>�НӧO�w/L�"�C�I������&���;h���T򎛀e�Ϳ�Hy��a��� S7r���G���Id�9��;���&�W���10.4�70���7���ғyG�6c��b�x}�T�,�Ն�U��ъ��tt�����nw�:�J����b�L���)}��T�Z޳���yӃ��	N� a�0����N������)Fh#�����;?{�%۵J�U������D�����/�1gT�g�$�������g�����y2�a^urB��j�Nm���{�p������xF�*��?�����w_@A�f�.c�ʕ��7{7��կc�t?�?J�C��	;���J�/�����$]*�ն��m�@�������o~�㏯����ns��L�֏�j��<3P�~��Ǐ��y������'��7���d��9 ��8�îK�A��Y3���|��y���د�gf���j�|
�ȁ���������(��&�e�٭�;kJ�< ���F�����b88 �3�EA�G�լ8LP��6� \ �8�=g`�N��!���_���Y5ga�񣈶s��Tl�=�q�o|��B˙��zGu2��~� f~��N|�)��^	1����V��xP;�+ز[�V�-�"0r}�H�Am��Ӽ�{V��� VjIԏ����|8�:����M�L"�=���|�F��L��K�r�0��8�HU��>#��m'��!b0BN��#����v�ym�"��vZ '[|��4��dj�x=�E�~p�A��Ȩ0s� �BK���T�Q��~}�j�f0j?���{?2͓��]�m\oB��㦜���|Z��x��(/�h�8���np��K^y�U���.�;�q��L��P� h��)�|.k��7&]^��ݭW��7����ݻw�}�̙���!�^��{���X�`��=���0��< �i����sk����4�ÿt�ұO��~������ų�ӋZ�Y�㒧�s��0og�uh�r>�}��|N�c�ȏ��������s��G6S�:rd�i �1�Qm��x�A�k�M��l�v'q,�4�U�|� ������rgg/��ydb��3����B�͐"nI����}1IK�0Ţ�O��[Y1����;~�]��>s�����x���e琈��igƃ��3�g����u�"_fc���{��L��u�Xղ̚H�BBJ����9��Yz�y���nr_}��G^��~��S�5@Q,b���Yw��B��:�t,ӱU��D��YI�D��FS�r�C�Kw���˯O���:y2F ف^�Q�t;�^���3�X��=غ|���Pc}o���כ�q����o]z�>�=�����x:@�ǫ����������x�e=<�JCH�Vr��g�y��Տ?���+Wd�����ă0�����<����{�=��k^T��#)�~��'��/>�C�Z궍�۽v+�Z�f(�q�����Z���a$�̃��<��sl��<k𼔌���JT����b��MZ�8v�bҵ��� �LP�n)>���w�{e��+O��'�O�V~~�:W���&''G��v�����y�}�PJ{���@�ߴ��u�)����	�*����F�����>s7h�{whfԁ�n��
����3Q�5S)�c���l�����}�<ԯ��4P�3.��^A������:2�A��ng�I4�ҷ����`�:�5��w��N:@tC���I��#�pj�-H'#�躮ϗ�G6_(�N��Q�`�U��G� i?џwL�n&`র�����|,�
kZB�v/�^B�h��EI�TiV��Z.w�S��v�)�=gπ��S�"S�0���و=�FF~�I�C�=)JĮc���0nu����jJ~In闝͑\�yL`�qݛiJP���e��Μ���`��Ǻs���C=t��}h�{tq����N��������Ͼ wV�dj�$3�� ��M���`��o�e��s��f�xi�$���7��o�������o���4�:t�E�����c�NH$����H6��I;n�+�^<�4�M��7>�}�5�m���R
t�1??$��Ђ��n�$I��b89�E�MSY4Ig��l��Ϗ�ɛıQ�`&�����Hv����R Ӎ��M�^:7G
�/��c浲(�P���g�g'����RU��1�'4�#'DPسG_���f��CY� �[�I\�Q'#U�|`��qM��;��<r�Y2���+�C�<:�w�� N:�^���@�&t��Q{=	9+c�yN&���:E���Cj䍍�u���KU۶�jh���~�c��k91Tb���)��sz]Ļ؅�%��*K6Ń4GvN�����TݥB�aQB��KKK;6s���Z�
$k������x�A���;�*���Y�����c�gb�lfi�Ѝ��:a:p��\֡,<����c%YzN��^�t��./�}faa��ٳF2FGT���p���3g�<.x凯���=�H��̓�m(��K�駟f�뻉m;�H��ʥ'�p�K��7V^����:u�{��^{��'���珡��X���LMMޱ�Z�݉�\JeB�|u@'�N1��Ů'l�}��=�u.��	�RD�y�'@��p�L?�ܫ�Q09Y�YX8�%Du������w>��Z�t�F��챯YUJ['�y}fY<�1�B�`��]�&����WJ�0fҔ�-)F
��i�
P��Y�� 4ҩ7w]�j;�51~�����e.[��T�yS�=�̳���%:���,Μ^��Tg���k��F�m�Qr1$`��|5�P��P%Sع�s�nGŞ�#�%
P��k�{��S]���x��x�J1��qP�ܲ* ����3g���6'd�c ֺ���Q����@�#�ƥL��<Hpw]��ݣq����A�7��¶�#��
��:�8�4�h�tj�fj0�s$�Q��l;N_�1�I�@�I?��-����T�n��c� a/��0�-�>��z4�Va�����j]��U
�Z���-O�����y+{���Z�\|Nb���#KGN
���vY1�1���E���Y\@��)$R%/i6[joZvq�,���^K�Y�J�oX����XR����{�7��q(��>�^¾���q���VYd������$�.
z��w'�L�r�#z��t��iD�BG�M��A�d�ߋ2��5P
��
j��֊���ё������x�'�-�]�|"]u�	����)�yהy��~d<
�E,���T�=ϛ�A%�Gݼ~���O=�t�����s��u7k�����O�n��>��EY���0�ُw��O3�{Oۻ�F/����C��v��.�q���ƯG�K�_��'O�ڽ~�:����":�� ��	2�Iz�l[v�>i�{I��8LS)ymρB��+B��%��鏺_BF�r�*+�v�0��oV
��q�5�ϻ�J�9��%+�f6W+���J与���rQ�v^���
��Eӓ��v�h�[$Q<�:M�FEk��b!J�4u�ʿ���k��@|��Me$D�S���ĠCH0W�ش/���++_;�4w®�vPz�2�N�� ���;;;{n���+3��"<�wS/���=��'�g�%?]*�Ma��md�a��(�#���w��M���G�X�Ѐf�I.�8�Q���Y+�ۻߺu�i��AE�G�'�|R�w��W^��~wii���̜'5s2�Q�_v�
g�H�
��B�D�����mGf���ڷ##��+��;������V&L,�X^�[۶�����W��׶�^���|��xw�ӑ�n4O�|����>��뻮�޴m|�Ća��=z3�V>z������(��גpY"-N�긣>2i����T�����b��*N���H���qzǏ/,=�����oݺ���S���SE%D{;+�xp�0_}�� 7��J,� VR3��,��S����~�J99�x����疗��\�x�j̨wэ7jԧ���f��nD�!̨)������MW-Ll�=m[K/)��OXS0��,2_�^v=KI٧���I�� |�C$�8P��\t~r�	���|�TZ�N½�ׂ+ V�U���ldľ�2{f] 1�JB�U����Q���V��-u-'K���������@��̱�s�����(����p}m�Hr�6sm���
��A��a��Wy2t�)/[��8�y{�ʸ/���M��;�h��~׶kK���RJ@�v�ў�E�ȍ��M�*�����z�i���y\z�c�X����+C�u����l��<ȮX�Jc�PLH2&�o��I�t�;w������/������RC*�2�p�jf�l�q��~y�헊�.J}K2٠�L-o{�����g�</Qv^j��8�v�kݼy���?;�{��r�ĉ�fҸx�b��ۛ޷���"����#��h���j�vhR:���k����j�ł/�v�A� GV��UmaY�0�%CF����	�A���Lv��㹝vϾ���3Ss_|�?u��5�/M�̶��B0֞��k��OJ���ĳ\�T�������'�a�a����:�
B,L��a}�L�nF"�J%��I&���OO�	�����'f���% ;D�4vk}]'�2H�n��ի\!��^��^�T�e	 ,.p9�4�K;�6N�B%�KE��'�����^'݊��x��8��x��#?%#|`�ȻC�:����߿w�M�巚m>)h���&{_�1J(�[��i���ͪB�E�S�t�ǁ��ky�;J���uX�����S�dss�So4�[��?��z҃������3b�_B�����M�N�#R�K=����N
��]��N��J��hؤ-�}�$r�� �pM�"ǂ�:^��u]�}�)ѡX��w&P����.��HaY�-5���Df��xxknv���<��Nݴ,�h�Љw~�Λw?]~d~~�4M��_t��;2�I�[vB��%�$ͦX*Z�v7�Vʽ��3[�f�&� �ְV�T�t�q7A��f���n}ww"��r��vw���-��-'!��-��"�j�z��H��cǽN�"L
|��|䑇�J�O���ϼ93��s����΋_~��Ǟ~��th��F����մ[-�y�L��t��6�Hќ�4�hrrRf��_��}	��X�ܰEV�Ϙ�K���8I�xg�1�Uo�T����?�vh@���~�ۯ 5b��Fl��An��ȧ�    IEND�B`�PK   %�X5�3$ �$ /   images/8251b1b7-c97c-4929-9682-a545aa133660.png<�cp%\�5|b۶&vrbL�dbs��mcb۶m�Ěض�=�~u�]]�?��w�սzG()H"���  $i)q  l�?ゅ�/���#�?g/��  ���%�#  ����"j�Y�҉6:��MO�ݑOGݩ�*Zf�pf��pb�Q/BH�Q��Ef�8�q��8�9:�̶9�����Gk;�^f*�Wx����y�=Ow'��W�������\N��������/�������rb,P}�_�O8�B�wG�#�6�����e8K�Ż2)4������] ���( S� �\�ޯ�s������?�����o*w]�z����s�Mv:񛮼�B�Xn�Fe_����B[�	f�W����f�I�����Z��2w�is���9��F;��Z>!��xS\ْ�s�ݏ�M����3����7)�U'O4˽Ħ>�Ka1��ҕ�G�"����P����QK��?_g��n5_�x���I{ڡ�﷣G=g��?)�]Kۑ��� P�����E#����f( �r{�j֯e�wjY�QȘ�:���`�]��RFԊ��&&�y�M�8��<��s�z�9R��[O�ȡ���*�	^OP�oR7�H~�Zo�ڌ�.�L��1���&c�2�4�C�8�����[9iӔ��rܝ3'
G:��~����|~�Ef�H� x����F�gs?&����Y�yhK?��Y�x����s�v�m]ߕz�Y�>i$��oX�:k���^���\__������}B�����'��_��T<�ɽ���`�u�J,���֪�Q9;�W���Pp?�v&#���t�b��)����=�����y��p�v��BSȵ���Y��|�V8'����UE�����U!�%/�X�#��*?�6X�\ͶnԴ�G"s�����Z�Oj2����g�j��Ƈ%�vmk�犹av��0'� 䘙V�
�s�|�=:�gK6�rB!�z���{�#eؘ�z��#�ǐ?"�uJA�(#�t��+���!�]��7\�W��g���_Ћ��)1�V��ʭ{����@��H���S�����Ͽ%�ǰtP�����1��w��c�w�X��i�B gvy�e���e�u?؞�宪P(�i�.wK1rK�՗G)��3�	J�	%S*3��th��C�5\��or�L:G_@��/m+�Mh�Ry[V�0|��������|<�4�ZZ�q�`��!8s��H����W"��m�Z�SD���4�Q�/?�a����t�OiVS��[� �_�걝-�� ������`<�[#���������Fe��F��6���Q��6uc��ޒc��L���ς��& ����_J��;5��8����^��5~�7�\U���+>5��O"B�k͔���[I�������q~�Q��s�����=/{��(��3���rfT�@A�W�%�Va��N�v�h�_<54l w�����kQ��.Z�h5U/5iB|�jV���b��'���y�*B$��dGf���us�R�HE��2����B*��,�����O���X��Y%�!.����b��S�kw=H�O�n��-�h�Vw�8�����_	�t��Xm`�]�!\��R�q,1���^�h���<6 s�o�E;��7�`�ٲ����0���W�ݚ����=�p7�m�CZ���BNk��~+ܢ1��TY�쀦�[u|4�W�76Ma��إ�i���Ke�bԝn��MH��	��֨���:��'��Y�о\��X]�L^�#s=���v���>�U� "�����&�K�@����G��i��C�j[[�V����}�U.M]BN+�b=�޿C ��g�t���`�y�^U�+�jG����X�e��j�2�f9�%���XJ˛��v�~����l�`*2K��t�S�]��L~-^;%����7�����v����%��}���.�U��5���ԣ�y�n\���z�=�?�ǡ��W�$����O�9���a8�^Y:ð:T�2��n�?o>���@�����v�=fϦ�'LF\|,(������G��S�}�-0�Vytk6v���W$�O��r44�|���1;����L�����j`j��_|�G�<kN9��{�{�` ȓ�����0����ua�/"�aە1Q"��U���ld�dI�Z���q�&�Ja�:�$y'l�N�DݿS��QF�XGڧF�o�si�H=�D�d��$��!��{|f���7�knWK5��%��(Z�?w��b�mq��$��t{��&9�m9f�;�]��%�BbF��V��m�6�=-t\�dk�������(�[���o�=L��h��-sb7hg�~e?�W>�h��g�_6�`U(�_�~l��(,�fo$�6юv��j��\�X���r\$����$��\U�:N����P��$��Pڕ��'f�T�dN�希;��fb������mj��4��KI�?��W�K��WB��e�(�OA��O٣��ϫ��:�p�^�՞�]�>���`���	E�&bpeb�x�1&���&aA�}�mX�E!=�J^B���?�׬��ݣ�\0/J*�c�q�?^%��{B����J�x�
�ď6+��U)���I���П�5jO��PҊY]С:���%,�ϣ���?�����V^{�GY#۷^z^>o;�P�vbw������#ο���0�`B�tFT�R�+�p�93�8�K%G��B�x�}k��Usp�l�C�\�o1�o�˃t�z0�!��H�jf�];�2�Q����B�<w���X� �
%��MI=���CAo&��PRg���*{Oҧh�	����� �ϗ:�J�ϝ5������rDE�<UT�%<f7��� )N�s���&k��s���H!���-����S��n�C*�Հk�{�8��\���:7���_S%�5z��C�D��1l:磹��KKM�w�~����tI���c�n�Ol�f���`�e�
���=?��9�+6U��Mj�z������q����xY���<� :�0$>M�i�����MO*z3{�e�W������_ϝ�]:��i'DxX�PW�%V�"}�C�^b�3\�ۗ����߶���uoWU��~[ز#H��/�ϲ�D͌�+�ëhC9($U�A�o$Q���"�ʻrr�+O#�ҩ� V����֤A]�@D쉥�9��]NN}
�~��Ax���@q�@�!Q�kc�csÀ������P���tQ��)d2_�di��mZ���cr	ljlC7�4�t�p�Ѥ��^7�����9��H�Dds��ƱC�	Q:ǿ�AS��1����Q$n�����y�|�X
��LK��w�!Q�hbmhY8��*f��H�D�d��2���I��s:z؟Y<"�y����~ͷ�Q��K`��@����_��x�S�7>N��Q��UG�ֹ_je��y'�F��l� �0X�L�p��sv�9�?�r;�ED��#�!?��E2�Ne�~������J}G�}�2�N|�;	�c������ϙjaι�[��>�X"����.89�m�z/��9}G���3�ْsf���$�@%��2]�'SZ��
D=ݨ�~NZO�2��~� �3���.�ٗ.�o\��w�=������W}l�Һt�ڜF�����U�m���0@F��	ߝ���d%k�P};�J�<-A���
�x_Mn��j�d*V�Gd�Mr���[��+�_-�/z�^�A{̔7K����fR5�UX�J�H�W�%Ջ���R��h�F�b`?�����(�8��z��J���e�'޹��;;"
8��ቢs����=7����;r-c�OЃE	�����iA.������x4 \�:����p��v]�~�I���]=������b̭>H�T^��x|�`=�1�#{m�ód�+X�	CO{�eE���
�dgR�'{!�+���!r�'<�����l ��HJ�p���6�X´z�t�!V�CD�������� ��hm��햑-�:�=�U�0Y|�t���I4�v�v���;!��+}&7�ݖ��^�.��Oc�3 �uĻ�r)���]1�,0p��I�P[`e����G���bU�/����|`w'ڳr�8�-k��5Dihe0^����9��V;Y6�����p����]�+LX��E�:�ܞ��U*�;��֘Y&��±�!=����.F�w�T�Lcc1����>�����,�[��y��(n�R�^��M�������k�UG|k�)�s��}�����C�ag���|�j���4��ۨ�ѿݭ͊�<
ѹ-g����'v��v�.�r���|9Eގ�a�����iW�7��Y\���㛞�L�_�?��$�t�mҴ��!U��P� @����Y�����o[�DO8Ԝ}����*�|�U�:r���G� Y��>E�*�&�4lxլh�_�wy�I�se��['n���Jw�:W�ޥ1-9����Ks��X8`�D=dܑ�ڋ�b�U\����9�POʍؓ�d\,��o�ʦ춸`M�7��ۉ�֟�Ce���ry��V�x��X��-�aa/� 4 0?I� ,��R�k�6��?�q�?q.���]%8e]��@�@���O��c����֝�tBjT���,�_��IN,�� >  w�ÂY�qb��=r�j_�^�vn9��:{+*�`y��=�вgc��7��@@�`���ᄘ�c��
�ƌ\t��v<�k2y����hpd�ѫ�l|�|]�M7Q@��\R�u�1;
��K��YW������;&e����֦6Z�����`N�r&�Ŭ�ǭ�|��Z�<F�ʣzV +�ܰ�D��[~��y�ə��ũ�J��׻~�M�*hnc���8�ARN����L)�~�h����һ�sD��^?c6�������8��z�Գ!E*���gv}�z��A+��D��G-��ϣR	z=:w��|q�h��ú0P<�͇-����?쓁2j(�� (��	%O�7���tX�r,V5�,��߾)����:
nU��R:�r���͍�p[T��kE5�}��'�� ��z V�A���#YJPB�Ya���n�ow��!RS�T0a�������q���?���3�b��M��b�><=w�a9;P��O�Ff�0��l�.���4+w���h�39#紶Pg�cSB��Q��я����a�v�Gܹ�g�u�]�� 2Z�/j鳓��"ݐQ.&����*?+������A���-vf�[ߞ\$��Yr�GGe"Tio�6�E�3�x�J������{�܉@j2��cj
�3�{��lu��VlіT�F��{�L�,��Y��]6�q3���Ύe�'��櫑�%�UFa��q���[�B���x���6�g�b8ϕ�y��"� �i�EJ�s�˷���q��F��q{���B�
(�;#���$���p�I��'\��W֑B4�^rV�=���+��U���tn,G9 <�TT�o�D� =JB��3v���(��������$$��B�!��\��2܌l��)`���`k&�j��H�X�Y��z4Og݁\iDe�#�d�^m�0f�PNn�!�^���[�l0���Ć��h��nFٶ������1�D��2��G*��/�e6(4�"�����?f�]�K=��=��=�� �<+�(`��Tg��B:~Oڇ��?˧�M!�e��e�۫]�_怋�ԡ�g��Zk�+�8�4�'T��8�������}}LG����U�R�/�)X%`z S?̓��$��J�v.�Z�{.����� ��j�M{��g4"��y��l_j��������"�>�v�@�������7���[]ί�Y�vT�zo09�9P��^1+�[Qf���?��+�7��|�y�o}�������>�2B,Mw�-���Ay͏n�=U��^B��wo�(_�7�� o��+!n^������'�%����#����q��*�K؁�>����k.a�1L���O��~.��F ƞ\?v�ÔF.5buí?!AN�^� n�����F�j��y��ʾ�Ͽ���=�sjT0����<Q����B��_kW��'n�o�D�8{c�b�p&��\��d9�&���pǾ��ظ6���;����9�]�ӫ�4�,����ԑ�f�p�)���(�D���-WD�եD�C];���ܵp�s�s93�-ˤ]�2�ii&��,O�����r���c�GU2���ՅD:���e�r��P@�Q����<���՛tm�� L~�@3\MU��������eW���6_.3�  
�B0Ze�ʙ�튝��о<"^F7ٱW��V���%�V��m�,����׾��=%bA���f�֪�幔��74ha_�̰�&H ���vEb��ս����chjV��z�xp�Y�w%B�ޱsuO�E��<��}����[���X(u}�����`",���Z�J��Cs��qR���q`Lt��ؚH�������+���~�B`��3f��?֎�m��x:K�_��z}K��!�����T>Wnx[q�nݩD����g<���h�j"�c��i/��h~ �8*$�Ku�b;���x���	��X-�k��g��"P���ɕFrϹ�u/L#Upn�q:���M����F1�C?�wZ�!Q�(^�g/��K �M�8

qb�.�{�5� {C��e��f���̈́M�2��zp�o�Q+�Y�5 ����<�a�P��7 W[���A���0�jn�YJl6�bԃv��4*%e8cVGVg���4�OO͎�a��*7o�	m/�}[���B53�b6p�L��\�@؈[�n�O#Zd��C�;��0J�o�����!�T�П��W�}Іuh-�,ďۋu" {���P��='f$<��}c��a�9��߉��Ym���2ϒ���ɨ�~�>wcX�/��W!v�]m�]�E)|��}N��n_�(o����2_.�	��t���5�KkO�|6�˰\~.�ǻ�/^2K�7��_�31r}�Ю�ړL,n���jhA�}���C�럟��<&�x�ŷ�2$�Adⱐ6��U(sR�<��|"�~ަ�݉
��������'(�`�*<�D����n{T��D��8u���v,6l(.lY��Q.R�xs�-�~w~���=��ǡ=���1'2�\Ҁ���]�ts�+$��T*� ���=v���Ddܽ�g/M�\Lb�Uŷ������JB&�nvIi�`�}�2�yr�/�Դq%6��%��q�v�>^r��ڹ�/fy�{R����O�Od�.�˗�+���zWbz�h�8֞�{3=��'�v�yh�|^��[�G��-�.!,4/Q���/V��ٵP�]��\��_Hܽ�P��?S���>���>��ri?���#k�N��J�j3]�t���^:�~� 4���ٶ��9�U�Bĺ���y,9�D����,��N�i�0(K�>8�"
��\�Wg\L�H�F��MD�[LK~7�%�o��3�� I���Y�r�z,f��?ڰ�/ϿQ���A��@k:�&�:�D_v����?�3��Tc�t�@��g5��62�������#�ĩBXIפF���K@4����3"�D�pg�a��P�H���<�Pd d���ª�Kf;c��P8�օ����]I&r-�e�ů�7�Q/�Ԑq�2�t��Xl'N�]� ��G�/�9�kN�����S��H|�:�/ܣ�^�����Dg���_�Y��N\cD�D����NJ�)z�|�a���d�Z��X��'0��Z��NoZ�@"έu�k�F͉�Cc���I�I��_�>$:a��mtWA`X�kވ����ʘ�L�S�f�D�=���N�"*�P
a�vt&��(HR�|���+����o��M�4m��-���m���N�r!�$`��$�t�I��-2[�{9�����S�A_�v��̠�~��1��(4G�S�v�k��t��+�fN���gObK%7'���X�{h9L�&����c@`.�T�6Y-�zP���g��r�'_%���y�c2��k�v�ҵ3
P]('���Z,͹����4��lQ���uľ���C�٬z?�Z�AM2s�1I�����dQ_��Q��(>�*f��C�J�:�$�\��JP��<���J)k�y���H���1*dE�:����,�sDmGW5b�����)��'�r��,m��&�vM���moy�%�VeI9I����$���X䤣�&����Zgm���k�������@Rw�Z'g0�R����� ���Cz�#%�*��ÿ�|�5%cl��	<n��=׷�"/���ߧ�&���$�~VB[Ew����&�u��B��k��G�Q������*;z@��.+
��A~��	����(���2P���6 ���9Y������Y�?O���9ߞ��6�X��z.�D���T�k��t �x �Is���2tf�R�Uf�wâ,$��!^�7��js��s�\j�	'S7$�n�Hj
m��Ϥ���a�H�d���n�)g�X��]���S��Bʜ�q�
Ѹ'Gq?�f+��Ʃ	f#ax6vbS?���*Z��Fm���w�xVhO����7�8v���l�E6�Pg�w���-���h+�����!73/5:�0D+�m�5��s�k#�֟��4Ģ�#eR
7�II���~�-�]�(bNffg�������!$��,�R�0�a�%�R���À��g	Hyf�,��� _|��\�!������-F�݁�@���c�-$M2��M�۹I�M����gn��f�x*��!�v��&,&0-l)ѻ�sҠ�o̊L�zL���I^|��Rv�6fҍ/Α=v+�j�	�]A���{��?Q��C��]�俴`�|p�y��7�0 !ΩYڨ6�m�f�� Å)%�s���U�"�W/�O*����LU
��{N^H���ϼ�C��L���Hx쩈@��4P�v�g�1�3!��J\όut󒅁o�����v�}&�w\�\�7<�RcʑN7�V��z����!��y�w��� M�%��5Å�Z�E q��Ἒ�rd���0;�O{ _�̙X�+<�h�N+W���)��4]�e��_��gz`�(h��6[V�Q;�/�g�+wroo�#�Z4�ύ�媺-`�a�����F�K͚Z��+��ңvl���4���: 5�A*?��x
� y�#qTN�'�����p#���k"{@��F�Lꔑ��+��ϙr`�����dϔG��zd������B7�J���,�7)r���Fl�f��^�sC\~6�h:�K��߶w�t���E���m�Ϥr�r�g�I�l1_kH�1;y&��zZ�ë�����޲˽�'����Y�������{��,���.��7�޺F2�<�7����qǧ�F�dɁ�k���1�ą�%ޒT<�M@�ҋd%�p����5�O����Oo�����w����F�JQ�=�JH?dK#�������lY�� ����Qu�"k�Fi���>P/x�l�h�1�;LG7�������Ҩ�8q��@��dU?�� >�	<���P5��1bh�5�N;Y��=���ԣ��t���`v�������4��% ��x�5n�x;���B2lٴ�x, ��z"պ�Zi=D�E����D�{�ʡ�<�a ��:�[!��Fp��	�aX.�:�|1��NB�U�,�K�)=c��Y�4�	�]�,��ß�S�L~�����t�P��z��ϻA[�GbćfO�l��2�D�(�ׇGG\���d���kv1�}^��NĦ���7��Ƌ�+�OѦ�U����7.?���!�]�]����Nn�W#Gچg�5z�7�>O:��r�$�硼����i��&��R�D6������1U�K-�N@Ln�{�6p/B�*m9!9�>ìx9
���c�� :A��C�k�08x=�r�=�����kS��>P���^A��>��B�k���޴�N�T,iP���8�ә3��8+lK�rه�,���㮨�������QA�ZO�k���dt�^r��:�}�h*b�����]��j�f�\)>D<t|�E(�z��k��80�gS]s�
��J�.�FD�&����1p�����j�v5�)������f�g%P�:@b�I����|��Ղ,��z�,%>�\1�H���NvV���iz
���A�iс�� �@�d����EF����13vE������圇=��A� �}q��B��_�����Z�m�p.�v�JS��a�Nc�\_P���E��Y�iz�	�!�\V�"�9+�~��Թ�Y���*������?p���@
Q�0�LB(]�+s�1���1��%G���Ȅ�R�(ui�X��G>��/��'�*��S
J��f"Y�P�b��O�p�x�Rjo�1���%�t-+{��8��T%�0s�I[��Ǜ�3&�ǩ~�˨��Y��>��a�7�|��q̅i]����Ғ���@�y���W��3<{[><����79��]��+zdSPp�MG֖`fl@#���-�ْ5%���I]�X'��u1"���W=f�VٜQ�k���GØi�����솶��,�cQ	aᳱ��}aBdщ����Q�����9.d~|5�p#]�����¸�%�=�}DY�:&�.�Hn��6���&�@l����x����Ǡt��c����6������0<�A��r����������B+�!	����U�o	1�oPҗ��߻/[�U�-����)�_^�8?3]���W�R�c�m��iqƓ�(KŻ�q��#Q�-�!h�f�#
���L���ʆ��գ������@��ŃnhW�܉���2�Uy�G�W[�,m��K��Ir,�8fJA�@N�ӽ`����ɤH��g�C,��X:�&P�v�<Q�=��� =B�JH���1��&��N\��'\Ҭ�5ȳ
�ñԊ����쉗7�Yix��	]�M���XC�f+D
�Q�6���	�d�r)
D��F1�޻�I{�d6�q�!���_��G���N{��l��nY8F����&��'��B�-�jxv�� ��ص�t3�`�2*���B�x���9F�߫�V>3����),z,�y�P�i�����Iq�7�5O���Ÿ��d����s�iR·��J���귪��ү�&�@h*���qa��.�c�� ���ݷ�u�5�A�	�!!����d��\�|�Ecx�W+��Ӯ�1Q��Z?���+L��i�����.J����c���G�6-�`sj2��7c�4�ʒc-V8�x>C}�pN�ߠ|�[��-֞8C-���M�e͍�c�"9��V��}t��U|�?i;H���V[ѫtu��U��]�cծ�侻i�WA�9��J���I~�3"��צ:&_r��	,jr6�)�:�(��m��� G�}�%l����0Е�nb��y݊^��5w�ڻ%	�$��DW��Oœ/��L�U�k�O;�T�s#�qZ�G���\e���*��*��A"eE�-h*#��ⴰF�e���}w��bA�h�Je���F��"v;�/<r�r1�!<������I��S��y�B��6�t�cĵ1��z�yQ��0�Ay��	V��v����n�8���?X�ʮe:[�����E�ɮ����d$ھ�Di���������[$������!n�~*�@���ˬi�n���h&�]b[cI�� �^0��hץo���T#7����ovN����k0��y�ݟ��bL�!Gx v��������7�-����1%�R�c��?6@ \����k��e�u4�wC��A`/q׉�S��dȈ�URѵ��"�A��y�ّ��ߤj�5��Yb	T^\�!KXׯ�X|RF4�9��n�{�Ɓ�V�ʁ�(W<���[/��:
�++�x��x�0oB��t\�(212�����X�_&��ղ@*�Yټ*)����^��sJ�m9�
��v��G��N���aC:آLMBY��Y j6O|�-tke����(y��60�����r����Y~saRX�׋�!�h�j���y�Z�<��lQ��.�
0�s�է���6
]Z4Edu6�MzsZ����☪H��d��7� �m������k�Pg����.�I�@Íez-a���e�h�9���k�����&���O��uz��Yt����'�@���\��u�H�r��P9Ù���=ƮҪ:��"}!�4�!�Ta�(�������1��P_�>�ˊ����h��9b�����>�WR�2!�M!��ϔd7BaőV�/���7q3�mc�L��I����)F	!p�%��s�KBx'��d�iv0>�s�"���������f��_N�A���e=�����蝬ӷ,.�?�\�h\�t
Cw ��q�hj�&|�놪׷���S����[�����_C�i���i�r�[#���"TȋR������T�Q3H����P�!V��u3H6���cD0�SBa��Cp��n�:N�2�7]W��z���R�pA���c�����\��r���x�G�Ʞ��nI>L4u�YY���ތyd����0r�x�0�R�a���S%�Na)̒W���7ȝu���+㉁7(܈z-��W�_��"���E��U��ZE���ú�mLp��j���츍Ȱ�3k:/�$2%Ư��0k� _����D����!��s`�#G2k[cl^��V�g�Gύ 8�F$�8��l���a%Y0I�4Ȱ!��!�I��nJ'�&���ķ �5=��y��x��Ӆ4#��L�<kK��9m�rީ�uK�ҮŔϣ�Ӭ�B�����-[`l�-����q\�h��`"�6�1	�Z���E]�DŎ<-�����W}ܜ�Y�[�z�4���E��5�Ph�� ��_��^YD�g ���8���y��~��n �$f���R6��UֹV���y��:t,��!{M�`>��\q��q�6�:��z���ڲӭ��s�;X.���%j�:�&�0�����BC��� 97#�.��r��0�E�cN�\~��{��	�&#G�� b�z�%�Lb�ے�v6,z�^BQ)f��HN27��H.1N:
-~l���mu��+Y��|'�/:\'"������&��V����WƸ��`)b���H��]�3���D�Ǎ�6ч�F\����˹�<�2NrVT	iB���8.�$Ƚ��nKa[�'���b�!�W<�r������hr����~��$
7�Wmi����W1vn�a]&6��3����H�d,V2k�^���&7�X������XzG/._C`V,wm-�;��i�F`�`�PEo]V�!fB�'��Y��߼	x���n
���@�h��X�Q����r~�m*�����&tr�a��)!�/j�9YTR(��(� Ơ�FEw��LK��*���֯邨�S�"cC���β&�>�U�
��MԒ�C���.d�R�٢�&���c+gc,$�g;�����H]�.�Vt-:��*V�XczFǆ�̽ʸ��]���0�&d8���֧��`(<M+�6�yx���HnH8��������R䩐��H�,%eM!�����k+����B��ޫz���;V��6��5�C��l�$��PM�gB�����'�w5<.u2��%��5������	�M�	��`Jҫ����`����j ��;fȢ0�:Nry3����)� �EȨ^�Dn&�sV�h�#�3���`�E���W$�] ��,���`XiRl��Q����s���p?}<!�)*�����}�3�G�%H�D��[�0q�?@�.��Z�Ktڜ&5D��6f�='O#4pβ��Jf����z�IKF���u 9�=��Iv+H�D'Z};�4��;�%�bL1퐷�b�,枹�M��|�9��2���Uգ��W�'�Q�%������/��0j�^k�9����?+���:��b$�\�^�썶!$/��s�_�ޯ�4�J@R��������k%��2�����RP�>VCi#+s�5UU���A���y�Eü�٨x~���t���N[�hT����_�}x:~HD_�E�᮫G Be"�� ̇�GϝNOx*����-�5`���QY��?!�歐8C��K�%����<K���I��tg�CkQU�wI���o���('����#��|@��[��qu�|U�����r�XFgS�MO��3D���JS��v7@?rؑQ}�Rz[��yY{>?��f곀��՛e`!���h�D4m��Γ?�~ы�����~��@1�{�0�r��X�_w����B���!�$�o�k��m+�Ǯ"W@�!��KU�#t��0�2,m�e�nRZN���>,�Lo�D���C>9Zv1�=0֣Izj��k$V ����S�ԃʢ�.����tX����`�i�����^�RZ=bMbD�$�L��W�7v��b�</�7W�0�kp�HDќ%m�]��e;:Y��e����uM�����v���u�U�}��k���wDH���~;�I=���WլKcEm<�s�*���P�S��hԃx��?�懋�D��5 �C�Tmc�kI���1A	4��]����^,;oު)&)�H����T�u���G�m���AEs��nd�M������-�����ɧM��e'�^���.��"7���؋,�߁9ٳtA�p�mY�[�;_�(��p��%Rb�)'�7�GF�������DĮH��κuOF2P0< �$��͠iZ�K�P��lG^�z�m�ռU<B�R.rW�����VOC����v��bI5�iW;0�p���G6fs��t�]s�$5�/�[8�h�v�!N�4���&Qh$�(�����`с�8�%=�b�!����!�ʬ��pa(��i�?<Dc�3Ex��O�M��'�ɍi�ӱt���|D��E�p�=�֠{��b��ܓ��ll7�g��ʕ$B�r5����0�M��©ߞ�Z�Υ���ΐ��MZŸ�/")ȧ��F�j�ֆ�t�\W�	����~r
��ڑ+{lx<Jh7��y�;0@S��Cc�6Lx2��@�7{5�J1���:��ݓ�ն��W>@����G|�W�d�;�{�	��	�M R���k�8����c��-~�qG�=%?�\���[J��{�Q�y踲X�G[i|����r/U��z�U~��ލ��}��@�Eg�GRĘ@G�5��ɕ�"���]���[���^�KF>�e%+�䣰��"�q�p`���9�R��ʟ�'}��`�`�G*�3�|U�;�\�P<o�$z@"x�5ͱ�|���X��z���;�Xދ7��nw�eʫ�m}���^�~����UD`S�{��Sz�E�[�.ß�%r�p:�A=�F
bp�v�+@Mj�E�F��X6�����ZTO�k	;����y5�$�h�A5`�s7j��%��]����3�}���ȡ+#�nƤ6�_t?�Ё��W�_�H:�AjaU�z}���Ϥ})�!)��C2�?b���^N��bƑ�h�c�L�����n���+���I����J̸Z�}Xx��Rݘ���OL���2Vb	�Ui��)�c�V�&��*;���΁ư/JD�e�W�?�6P�v�O2R��(��G:�z�h�7�{g�,�O������G��~Y世ʒ��a�>�;0-<��k�'��m�] �T�>�U�Ёs�w�Kd��e���-oG�E_�3�ȫ?�OCͥ�����v�(��NG}�������!��y��ٵ���X�G�:.����u=��HK�����1Kޔ�s���Tk��姁�}_�{"�Cq�@
�E
�`��'�#�&1J�����n{�n�L		�c#nYn�V��cﹱ��4����:����<p!A!(Y�O�j���L)h�nAK_H����4��r�f&�Yg�B��£xI��N%fu�k`�'��i(��V0él�V��>JL3 h�����D�U89%��T���U�a�|F�򅯲˙��1t�ƺ���$�Ά�|$��g�ܭ'�Ǽ��lo&���/�!@th�盙�a���A�s��W�d���^{pu��Yb����l�5�^
ŀ
X���~W�%�����1-�U��O$3��� �I|ozjVHBO��Y��"�0<E�g��46�	����uV��}l�+�j�cOp�һ6{ݚ�7�{z��~D�:�.2�����K��yq�@vV����p�k���@�@��taLm>u4r��xSvj�=cAbqA��P���W'cc[Uȧ�AZ(H��~n6-�(�yS3(�ձD��X��H���D"����#
����L�]��n��H趞������n>J��������4��n�Q�;�va�Ka�D`� L|�n���b!O�hdd�5������J,J�����A混�^�P��"-ʌ@��G�G"-���v��Ʋ,�u^_���_��E��@F�	��� p;U����J.�����t��������A����G�i�9�hɈ{T�6�)B���T^_��WW�4ܸ�`RY �>4�p=0�_}�<:�W�[��l0/��+�cܶ+�I���-�;��۶�`�I%6�@�/�/�\�pgUD�pÙ�9��joOSNӲ�a8���y�U�R�]8�(��>mEV�˧5��[ ��� ���:抝��OG;#j��@�@�p���:�\�A��Z�~��j@���{]ОO�5Wj3'Xg���������@�1�Pv�B��µ��i�e�:��5���$����v��>�7�����P-~`aX���;��@�:��q�a?yS�ȉ2ۓٙzϕ�r��tƨ�u���[�r�F�+e��N�Є��WЛUkF�A�5�wȉ�WֱY0���cTU�|5��U����3�\3Z�1V6����^JV����<�ab=D\L�������,�gc8)�L�s���{�j��w�˗_�Z���� �jX���M����syyq"g�؜�1� �瀒�F����� A�n[�%�g���R��,f�,g��8l���f	C�����!9P+O�{�kg�Őo|��f,�YW����>ԛ�
j3)Ǐ�0������u�4rw{#��/�\���e���p��y��c��y9;?a�!Y�2h�s̦�{�׾}�V�zۗ/�b��'�gs���A�1w�q?ڄl�-1wM��8^�����# ��w��#��g_��,kC�h���>z�u+��K��>�󾾸T�l��;gB�����!8��,�oC�ʊa��(���0'� q�BՂ���6\�"�`�ZJ���vw���b:�S�� �R�h����ŵ\_��]��9�w��ӹ���Gk+���x!?��Od�v��G�³�
�
^��rŭ���7���c��$v��iF
eS纆>{�R~���x�	���|9Pkր{�Pۅ�G�}��Ƒ��
,��X��l�PF�(���(s�>	l�Y$�MKR�R��n��g�E@�Emc���&�2(Xj;�Z�������w��֤��X-"���w���9r���j���8.y���O���G�	m�|�!b��B�]��Lc���A����tg���#Y#����hZ��K5���v��5dJ�ܺ���M/.���;2��8��<2��@�����s}��.n����D��7��g�}��)C��C)�2��u�5 T�}3u�tani���ۡ[�zK&�dz�V
�
����@p��EΪ޴w�_���[=���$0�>��£V�3X5dg��}^"2<���Cޏ=K+e>
�\���&Nu!��߯^��@~����b��/����%�u
����|؎��uD��7���n%��G�AeI�$����ޮf���7�˟�\A�b�K3L8->[�{�0���؎8�aS� ơV��E�0<y�P���Z���0T53�$�ٲT��C��0t�${!�����+z��i��!�dSJ
��c��^�m�V�C�V�lfrhA�\.���F�LJ���̬����A�0�&T�%(+�Ѕ���q:���r5ГQ)�'����zs9�,׋>��>����K�p�f��Yx�m];��a�B�&�[l�����V��:�u�l�c�����.S9���	����Y��Grrz"ejM�c�p�RrGfvD1qo(#�C�����Pk��*S<`0��S2}~�-�^k����;J#�=X���+����� |���H����b�_���m}c�Xat̐:��4���@��iԈf��\&�)#Poաe	R����ghB��Td�'�<֟sn�"�=e�9���x-�f��,�
�-�zEq[��
*�Q��z��=��40z�N�3��FJ,C���P��p?�#�{7���;u�d��9Z]����.��.x�b-p�%�M�OK��ɧ�>$��9�"S>C"ւ�����!�E����ñ��x��^��~-痧trp��d��vA����c���[*��������z��ѧd��@Gq!t��Et�*��Aj�A 0zy����E�����γ=C���L)i�'�u���r���P���X���Bk1�D�,W;٬?r�(����9��Ȅw
�s��Qf4�Q�D:�
tB�2��D��#H(e�X��v[�a�:<�M`�J>>=��~.ˇ��kn7{x��$�A��1�g����F����&̠�X��M��{�J�Ņ��IJ����-�+���,��:��f���J^( _�\ȏ��^��(�AM	4���5���cNF��ݦfȿs�H�qؗ%�ZS�u:�żv����}hb�"������&/�
A�
�J�-��Z���Ҍ0�;��5��S2eJ�]y��z&�;X  �������)�M���K��l�y�B~�/�\_�P*�S�L�跺жd1Xlӑ-�qn�E����Y�5ƣ)���b%�w�:�7tP���gz:����p`?(����=k� B�A�b���K�0���5�������#̖�5C� 52�����W�����KS����_���5�p��Q.F����s��md��NY�
n�=h0�ʀ��F#�T��p_>�+��S��L�L=��21��7��ulw�+��-��J���@�!���[��X�^�˺ޱ�ߜ!�,���:յs��� ׯ^�� 8l6�DUHG�-��2�[��BDӞWo�`c��A��0��l����Ϩ���͋�@�=hk�ґc��ةDX4	��
y�� �CGB�r���Ш�!�V�~�������g���IH�Bҁ����ղۿ���q�S���?4L:f�" ��j:��u bi(D8{SkYK]�����ěp:���/�Ky��;��Ws:ܸ������C��c�{,l�49�q=��d�,�[H(��B�֩$ϙm^b�y/u�1'Ԇ�]V"?���L�*�Vt0�n)M�����p����u�l�X'I9!�d8Ԯ�@�z�޾�(��'Y?����)|����Cn��<���p��9�4tX2�%�Vm��栤��u<W쀄��6� /��N2_�~����Jp]�5*?~�9+���!*��Ll�iq�:����P�Nf(��Dd쐕��ˊ�,$����Pg��?�����?�3�:*��e�,��̉[�56X`^%t�)ʰM"r)ȵ����i�?_�3����^W�K��� �Hj9.����zܐ���v/iC����gS�DIy`G�vI�Zq6u��,���J]g�3�W'
�������ׯ�͛W� ʁ���|�L�Q#��/_�O�5`" rp:5ȩ��;� <�}��&��@�����V��[ș���YfWr�)C���
�9Ǵ���~P@}R�s+�e D�Uj��!���`�^�:լ�Np�-��GP��9mu������G���  h]!�^7X�":��zo3������K��
!�[�H�
���L�!΄C�%>D��&{cƘ?<](���x7�Tכ}Dɓ�����:�*�M��.n��x/�����K��qM�� �X6���{KpE�![Ȑ�������LǬ�0N�v��#���F�!��T{Կ`� ��>�E����uM�������Z�@�������F��S����ø'H-���ي׹ �6)@t@�M: 0B#WV��M�^5j_|�#qo~B��_��_�J	�m��Oe�cB�����8ο&I�	�����㽅�$�f���M����F��=�xE"��F��[W�o�́mEt��Z�˿��/��/^��}��W`T� *�:pc��2{����%+V�K��޿c�sߥMP�[�ǣ�X�b�:�c�c\��]�@�+?���u��GF;�c� y��y���4:�F�z��n�"��8���>����!>�s�H�Ij���X�e��gS�v�>(����6<`�Ibpj>�I`Z�O��4�hϒJfj���B�*�AI/J��Js4�ʫןq������7�N�ʓ5��T��P��ȅ�����r�(xSc[8�o�=Y�!O��F&��m�:�%M��^�1?��}�}��E��b�Õ:��0�a(
�'�m�:�ء�6�p���$�X�*���ϡ�#� 5�%�5�uWB*7[�}ǲ��8_$D�����"�[���oC	G`�u�J�����X� Ǚ�%�f�s.���齝�seR��"5É��!
j0ȑ���?Q�$�̆N���lt��m{��F]%a����5���}n6=��L�~E�N�7?��,u0��@�:?A��!Z*����{���>����4kۺ�i���
1��ķ"-���>��T�`�gj�`����M:�<���\{밻��i�\x/c�n���ӑb?a��ͮU�K�0�.�r��3��O�탽Ŧ&�����Eqj_n���5%�0�N`=�`Ajl���[��|ʶ�'�l��:T��1V<����%��W��D�6r���� (t�vv�V,K!$�\>Do�h�:�g�
�:Ok�u���w�N��v�������ڙÉ���&�a��̕��k6 ��{kF�0�32�F�c���_����������ޟ7m �_���+�|
6���#�F�_��Sd�a����G��w^񳏙u�덟��=��yІf��?jH|��
s
���Ib�8FP��D��`}���:b�
������ l|T����/e��H'�7��3~J�!�=�f-I�|����0��ݷ�5�ɚ��L��+}�N��/)k�1������V&�5lwKy��r�����H~r�O��ҷ4j���Z���z04tz���P���\A���M���������t�C5I�h�Y��	IBR�3�zst�Ø@��il���t�.h����eO;�	C�R ���ۏ�R�7��;s�+T��e~{����D��PY�A�YZ� �%�Sc����!���g�Z�z�1�&0���K�SC����پ���?>Ƚ^��C)|����D�~w,��l�-�� �Y�0UEP�(eڱm^b�����[�n56�zɼ�X�W���6�:^�mބ�X��CKϞ�-q����;)�����<�-�X��e�[��[�:j��w�����`�7��.��B=D��F�O[���B�leZ�^��s�ٶh��?(K4ʜ��B*WQ�0���dzv)Y9����|x� WWjfgJ�mW�]�N��I^�w�A��݋���%)E���|��8U���0$�*����D��_^�ۛ��_�U��c���o����	�)��iݱc�6��Kq���s��/��8�1E�eヘ�"#��|:�Ym1v�2�齮�wO�$���T�^���I���y2Q6�5f��w��F�a�!sk�b������m�����7�H�@��_��D�B��lu�>�#�� ��ܺ���Wz�P��9DW,SbG��B(�m^�w,�v����}�qΟ]������z͊
�*��ȶ������k�m`����������������6,�ĺ�|@9!�T�����\ǆը�:ĦK�!"'Q�������j �m=�����q���P�x\��cp=�S��@�-#w�ׁ�l0��db�G�&%	�T��}!��1����V�vB6[����S���d�?����X?�#w�V�~����7߾��x��P\(��k3Y�k�+��c�~_��:�Y6lG�������C�<�����A�O���0W�3�p���(�7oe��e�&l�v<+��}-�e-�>��˫+���`w��ţz%j4�������ԡ'��EM�J���j@0�I���3�d�>��T�;���/h@�`���Ã��[q%kX����X�v�{�'/&(�����@���1|ۆ:h��Z����c�{%�&ƀ�SA�MFF''l��;�/�B��1E�0�6"�AmC?l��֥)a.9	N]��%4�Ol����6�G9��cr7����`?��
�������/T�!SdZlc�$�������S�~��ދ5q�5�7(l�j�X���
���C����{K�A���iDv(g��;�
������t<GaЙa7���&,·��\8_9(��ЇeGp�Ɉ��N��[]�\ț7o��յ,�-Î�OM��� {,�����5�en�0�P 7/�J8���c��߼�����^�Z(�v6w��L�;@!��t<G���9��611Kl�	��^Z����+3U-�jXl�Z*��s�[��F�:��T�*s{�z���`/�hT����R qG�F��Qf!b�;���b�t�w�r�`m3}�s�i�	Zd�DN�	8'κT�z#ద;da
(h��iBG�����D�w9�%W#���~��v�T���ק&|��w����?<�V�p���q@�%�韞�������ku�f��&t&p��q�e��~bTV������g��齚LӰa��+�)pJ,R��oǹ۸n�z��v�����1�m��������c�G���Ci�
��ވJ��)�\]�����;�w�&�+�٢�7�)�u�������쪸j
`�� ���s�����NN�c\���d*#�78�DyN�3J�w_�t~�y�cr��� �zS��*��oe��7 ����-�Xw�p.Z᥶~�(]�q����E��yb@t��7h`�ۭe=)�{�� �*a� \2����B���~���Y���w\8X0�d��P%�:
����'t��Vz�.��7/�SN�>�z��S��.g�RP���~���X�F�^lr��Ęx�P޼Etm:n��zGg��b��'��, 
0?���\l�^��8�ӱ�}��ono����6���
��Pl�t���e@�!'Ǟ�YP�b�����a&&�kp���i0:2���J�4�n���/��a8�-�߷��&�r�mgM٭�ZLBۆj���`��D�!�N��<bg�|eq�X$�j����1�w�[Rh�H� ��)��(���.<Y٭P����W�z�=�s����O��g>�W~��׬7������ٿ+��S#�����z�l���% 4At �i8P��:w!�C���ým����
�6�5�����ؼ"��tSSK�aE.��؃2��1�N3��l0�6r�XCȧa�ݰ-�5p4a!C���$�M(j�z>O+��QO�p~g�`�<��ש:��&��E&��:su�D���o���r�(�Co�f�3�.&�,B��6�v�����Ou(0\�H��#�~&�}14�B��a����z"��l,\�Vm���YA���_q����O���}��'��|�ϗ�p�$��L6��n��h[��R�%�~�߸��-KmͶ!�L�M�=�M�OEW>�5�|�͡s���{�6���>~fz�ݱ��uM����wAc���Hk~�y>>3G���ɔyv����d�����,Wҿ�F����/t��B?ь��$�U;	!%��F���/���BN..��ťEu��g'����9�>��L��Ax�\9e9){sK��̴VC�R�pq�Z&I���Qf
z_��3�ԉ͜M�Cc���Xą�\nh�N����I������m+w�(�f�K�5@*K����9�<[o�Q�'(Sf{�
J��H���%<U�ZV߾�T�*���vz!Ԝ���d-6����k�;��]!j0�F� �b3:g�T�2c�}�X�wQ��J������}~���|�d�������� �]��6%��x{��F��Z�#3p�r8SU�Rս}�z���/ү���?�ͤn��ΐ#��I�CD���v�Yj3�2���<$<����Z�F��f�������{˾���9| ����f���r3S�כ�����?ې�k,��NB��� �u�`��[�&	��{�=k{���@I:��{$\zSɍ8�8�j_"wM���S�aD�~٢;=!(����1^�wRyM`��Ӌ*�{�Z��10�F�)�Twx��g���J#K�F�O�TI��g�������R�e���1@S�zg!���u��9��Y��n-� o3�1-�M��ݛaO
�O8�{ws+$U# H�Iz��Q�h-� �{�����>�
N?Ju:������B��ܞ���u�z��*ߙ tUV4�Fm��?� \x3�M��i����>'�n��L#%��r�瑐A�3�$�f���	ƨ�#�U#���T(���{����P�|��u�P	�B���	��pѠ����*���mO���A�����cX�kj<{���R�OP�zF�<n�gh*�v�>��y˯�tg����v�ono��ew��.+�lW6h��$�UQ�f�`(��F� �������lV�Z��[j�N����Ktt�ٗ=�����<���Z�X�N#t��D��M;/-���?�[x��g���T�h��>ƅM$ SE��q���S���}X�||�`� �}���>�9��]��٢�W%A���ڽ���U?<��O�:��o�}�b�����X�����>�T����� EIR5��]or7\�c]%�8�z>Z�h�dzo���c*K�A
�L��$��W��w�,5�5Z���e;��R���96s:Lʉ G'�� �0��;�=�m���/l#/](ڲ墳_U����K@�h�8�sT!A�}�Dc�*T����Psb�I�XQ)*�dRв����:���xSi����J�4y�~
�|7vЯ��C	Č@r{�g�"a��>qB�E��٥S�I2�0eQ�DҔ��N��(��ë�~ @q������� ����JNb�?�y���B@0F9X�TrD���e�v���3z�<0J|&�=׈���4��~����T_>����|��ѤU�i��d+T5��J�q�QHdA|���m=��P���9��'�A:���	j��
В�i�3g��ə�:����c3P0�-]&T��"�=�I	�D���dͩ|N�+�;�;�r�dʦ;��2>M,��;�}t=\G��^��lG�44;�����\\�m�h�fj�����[�SӲ��d�cɞ� )�	�s$��[�3����$�K��;�nhjK� ��W�R�:U��(	#�{U���9W����"8)H�t�"T/���D�41�)�X1�02�ݞ�h��
����u&������{
�3#f2�P�2�b��®��������X8���Gsʣ03ak0@�
U�u-6/��ݣe QV���A�f�=p�pqo�<��U^�����۠*w���S~�N����K2�����������p���⩢X@�������/j�|"�,���u��>���\ڮ������L؄�W��^�c�m�2ݎ������5�����AB�z:fci����鮇�9�/;�掆vW�cf��Z��
�=P���!|���p�����6����	�ꉣ��S��f��<؇$2���~%�^�)���d <���,� �a�V���X��R^;���\3�z�jn��(
�V�r4����O-��~�PYc��'"�R��Γ��GRwQ�K�خD"1�=]�����o�žb-#_���,���  �h$⨐9�Y�<��0�|xt;��/,Ki;_�ЮՋ"�t�1χѧ�ѝ�
@���� �dv��M�P�58�,3�5��Z���y��@��F$���ݣę, I���I�!��E:���+8�����Xe���e8��A>8I@o2Ɩ#�AB��A8yy���N�(������~0�Ms^��V�W��\�a��̳���d�j�1��o�����T�d%���{��Ə����t$Os9�>fD���'�,5�Wqaey�q��ӣ0/��"��}��x��i�0�A��	p�BqKj��x�w��ï��>����"m"��_L���d֔~d�3��5�jY@c�7��=���$��*Vx�k���������9�ޮ�,��Y�x�}Q}�%�$��PP�`�?ص=N"4�x쎪�#OA)��R��7����^'dA��gHt�E��Ŷ�=<dX�Ah��g��[�������� ��_�. L�
�!����^�z�vŏL e�i/h�!\�߇��G{�;�AM�q7�tb:���h�v��}��{�j΂k�ظ��Ƭ�e�kmیV8�����Xʄ��'Sf�%g�v��]�~�C��Ke��H�X���~�4h�q�����	I�	�����p��M�;S]�9>���lcܧo��h��������f��)���k	�>m�}*X�
U�h��(�[��w»��u+/�e=��#�z���S����"Lw����}m�Ug%�(�8�U�p(g88F̡�+�`)�eљ�9zq�$�+�0�^���7��.	�κ�����vA���	*Ȧ��);TM _�ٙ��"����Ύ,���tS�p�����l������{���m�ٌ��W��á���Z��9�UR��J��|�FhX��AKE��x�����_}�m��=����=�fj�'m�:e'��'��4��XQ��������2�f�u��H�Ԯ�!�X�m�6kN�C�R=�x�xQ�����s��q:����'Zz�J݃�9s=���+J��ζ%k{�u�,���A�n�X=�w7�ֲ���[�w��/��"�V���>��q6 �[�*��+�G
��Հ*�e&��� �Eל�J��|mYv5���H�^�և2w��W��uZ&��KA'jID��ؓ��t�K�.	�� �!�/�!�ȅ�],������o�������GH�(�5��,�h�����Z+���Xr����\���uP������2:s���Z�7��-%�q�ӵz	��F3 �L��t���텽ݣ����2�=�|�'���Q��e�2`C��XT�҂��`G��*Z2��I�4�^d����f�?P@#]���LSr<��R�0��8aJ�cF��A0N�*7YvR_�з�{���G���ʲVJ�RV[�d���9�������peA����-�y��TN��q���z�sU6�Ւ� ��@��+�)b>��4b�G"�y��������~��};�V�s�9M=l�(��|���G�Nt��F��vBc'�j�Oo�(6iL�)Di�����5uqm�SCX�,�1+�Y�Em
�7�VCx��˥+mUT~��څm�9P��^�T�D秬꿃�u��<�&�$������l2�������o�03C��p}x^�2/�A�TC9GG�>�� �0'�g{�e!# �bib���ޓ���b���f��;XZ�׻�£�<��
5��E�͝q��^�Mxt4�P�A$/�_���S� ���K�N$CTy=�QE�@yZ$�G	��b�)���eh��D��~����� y���0����cs�{B�Hٴ�P�|s�04��Zx���76 7@l�N���ZI.t̀[���Vd�G��?��n�o��Vs���e�yܦ:��,��gI��vD�f�kEݕ�X2_E�9C�Z�V>�ۙ���{� {Q����\�����<�̱Y�a{n`�W���(��+�F�ío�- k*�ڽo��g�ܢ]^SABQ��J��J��.�eSFqa�&�e�r��Hvx!�(@�[��{vvN�4����nB�}��ޅ�Ҳ�L>CM�'��0mu�sQ�t��'ar��hiF9)@w�h�9�ؾ�}�������Č�BU��������`�;D ���(�����ɞ�Q�|����DԖu�U ��`��,�ݨ�vs���)ޗ:ɑ���X����IX���6�~T�	���pg�2ɵ�A�G��k��k���u�Q���s�.�
g[��@0��{��ٿe�c��0�I�|�3��`-H[*]KB�p�d͍A!���6{��޽�2U���qE4�pG������>����ewbp�~vaj{�ͩ>��@�rgӊ�+�6C)Q%�j3NԌ��^!�6�g���B��o;�/��I_�����_:�m��I<���	�V�8��,��ڙ6��|�GI0*Q	�����b�Ι �W&B�D�HN�
k����R V�X�o�Q�"��D[���V��>��N��������9iŚ~I#qZօÉL���-%�cƣm%=��Mv`wzmV���O�J�/���pR	���%�t�Q�Hʟ{o�B���7��e6�)�Ǌ�����[�fhj�������٫�9W�c���ڮ-�̝�dv�C�;f9�^S�����L"v3�U��@���]vaj�����T�L�Μs^e���Q���l��*J��g �j�����*Ef� f"�g�����q۱�ke�����
�P�l'9bJ���E|4G�
Nͧ������� ���@��@7V�N�H{i�Ɓ`CS^":�\ѐԫx(��#��	g-�Z��A��:��j�o+�A�"�4	��Xٸe�׌�������lF�<�,t��C��0ǘ�k3^����D8��"��u!0��=�L��&z����TaT�ʪg0孬���	Mŋz�2���R�	%��h�_�����A�>��]�!�� hn�*��q͛�e왱�`�-�[6��T�,{���W���E�m!֓i���H��Y��U`�߷��Iۡ��?�Q����U����~3������`k�5E���-'�OT������!+g�y�)�8E؀0��;;=8s��,h��}\[�����,�{C��3�E�fE)A����qo޾G{�a�3�;;a���'�&;'�Z��!^g����V��|VeöO���}���zaA/�Q�O�>�gx���/U]��u?��=�X�7���vMd[T!Ԯ�HU��l��}.�y���Ѝ�J�IMil��ɇ�vSh���a,h͖�<'2��� 
��2��9�L>1����m#M&����2��DI�F�ܰ��1�U���8(�m�c��\�N�ї���6�%4���z^������١o��U������n@�*~����	�	(�آ���A:��.b8"�o�G^��������݁|C���R���L8�BYt��=�������e������,����W��9\b�	�P�ǈ�	��>�仯�SI�r3��˪��/V,��W�ی�t:���x�M��*�$}�G �68�w�g$��1�ą���3��x�����#̓�7��_P���_��ӓ�]]���@C��Ő"�ilY�(T�)�bdCIo��������~�駰��#��	-[9A�h3WJ�PE�:#����=I��c����w�i��YɄ톢���T��d�C��ss@�rPEX�0��2C�k��Dq�0����f���f�1�:4�gj�
N۞�>.ë�_`��{��������<���]�^�ZЌ!�����bD�(��A��C�rvS�s�@��vm�������[f4��KG��F㐙C�!���d"�Z�D���XG#��t
�0�]7Ų6�.D A	�n��R�K˘f8��l�u�%����vw�����ك8�K�Oߩ�bc�xJɎY�8��mա����˰��G��.ȸFc1U&���p�ƾ�� �]/���C)�/�=������ؕ9�c�=%	�F2�%�0��!=OHl�P8K�Ϭ.�<ٙ�����|vo���ݍ�D{ʪk�������dg2�^�/O_�- 	.
���������ugd��3j�#�}���W�#�߿W�Ү��_���/¾}ֵ(	����æ�Y��n.���%#|�Hf��Q��φ1*w^u�N{gӫǦ��q�tU���L|�#�	!�$�'�]F|�x�	�vjo-�ߺ��.��oKv�Y.}�S��������A�2U/S?;F}����ʄ7Է��f�C��5�Y��ؒ���	f�(��F]k��gQծp<K#�{k�H��a�U��&դ��{����ᖲ3,I�针U�W���d��C"e׻n�_4����yXv2�8��0u�z5hִPfG������>��ڽ�������P��ե9���A��*j����5�`4�P���^9�nfH�d���e�"F[8a}_JF|�m�qb<uY9�YK�NK�@�G�LpAײ��9:4U,�X����m��Y����^��W��pa7�,s��8BGY���ʲq�UD�
Ӝ��oxe�eY��EX�܆�FG,2�ol�f�K�d@EO��.�|\��o���!I���2���g�.o�G;�fNGz-���yJ���7����|7��!�̰؃�V���=�Ge��*�g���5��uP#��f�#�ej��Z�u{B��(I3o;��z��裙s�0�� 	�8<�A���-��C˼>bh�E�\p��Eaf�����#ڳv�&��D���Է\Ę3�!�.��N3�7Ͼ�e�r�:�^Vt��.�9�4wlǾaD�Svcz�\��*3�Yp[��P���#�`��0������2P�����QԻ��͸���c�K�������j:���|�k`T� ���>��j~߲J�:�)'O9dj�Nd�c;�Sw>~�D�89x�BP;�Ӗ4hU��8�-����*x��}��	����'��{{���똙�pB��[;.�L�L�*�������Y�֮g�]a|i����A�4{���l���w�D9KB��+������)�ڱ_&r�h��U�9 ��q��|���џ�1Fq��shK�� h��.PjJ�Z��"�[��2:g�h^~�m~��Ϝ�v���i�,[�rfX6}�9�g3�_:�d��!{֚Gށu$W���x��OVh<M��g�Y�κ'1Ӧ�q-�_gA$�cP�
���ch�ۢ���k��
'T�YU��/G��yfIG��<B�b*O|#B�%� �_(��2��m.�S�&�=g/�UU�ޏ�(���Ko�c�;g�������3�y.5>S��������~{t���b�ΰ=e5И�2>B�W����؎<���um5F�Ъ"�pg�X�����:������ݻ7af��]CRvv���e1�0�8-nv10��46�	�G�lx`�3D2�Q�8Bt֎%�¥���G�R �QE F:(�qfI6��K�cFqjH�C<O�#���7jG-/�kjـ}�N��@	���Ht��8������̛T&�͐o�������T�[:;Z:�i[�9�DT=�+4��0_t�lf�ԛ������24�k�q�-� q7� �Yx��Isx�:�2�jy,�=o�҅l��Z(���9�����5^/#������Q	!�-��Ubt�
�;v i���C~u��o��R�3SX��&QQ��p���f,�һF�-	����&!���0�<��#`�K~�q������ٵFӰ�§�H���=<��E�ĐQ��=�s������z�S��po?�-hI�EB��p_V��q�݅9�Oח������w��f���Rk�,(SS+΢�s 
g�DA+����֫%���^�
���&�f��W�fR�"��a���#��ڳ&)^�Jt�ij`�oԵ(w*��0[]T�O�")�P�r��<~�y��K٪�NE��U��;];��{{[�2:���I/r��Ά�~��e�[��%F�Ϝ붓��#O�eC����~_>��%���icW���pf+��ת������%a���-�s U�@�B
�Q3���&Z��*~$m��x�R��Z�d���%�m�G������Q��>N8����b�tQ�!�<!���
`���B]z��v)}�](�Ț*�fu�P�ax��2�԰�1XO��n �B��%&�\V1j�n^싨��YTi	����u��� @�� >�_B0y�%�&n+EF/1��'9J����I�ֵÌT"%,�2 �{��e�w��J��sQ�S1� �=���s�6��$z�Ͱ��6���g*�8W�?���1׋qiwʍ@?#��k9���u0ՌMgC�����(/¿�1gm���9N�/ކi�*%2: sSy*D>�h����N�?�#�kQ���k�eN���PH��\�uR�NՏL�;i�`�-�!0�sx���8J�)[Ks5���5
p�l���^Y��j�Y��p ]<�I0�LE�Ӎ�E�+�+0z;��e�tw ����Q�پv �f�A����c��8d���M��,�-���o���Ψ��./8�U�`�N�O��;�]9�YIYӂ�o�Y\��A�ZW�Y���g������y8>��9��QF�o��3��r~�9�)�T,�v ]`���I?=���װsK�xV�(�[/#N�%x6hp�����T�F�o��4-�3d�I���]�+=qMY�y�رτ�`S)i�Q#�v��y�����A�Ƕ�{�3��<cj %�jF����}��y����M=���H�J���h��:b{�5�|��I����5�3\ǲ7�άAB]z ��h@G���y� �7E�R�V�x���7�ή��y6��=��PcUMt�1�L�+�"J��8��;QH]?WlՊ��h¦��&B�Q�(�q]��� �[N�	�̒��;�2��A�E3��<{�`?�O��T��7�3����ރ �v�~������,�����}ݽr��u�9��/|�"'\���j�g�(Z���h�X$�g&=�t3|3���Jo�)���V-��Y�@f��� �_{?$�j2��fi��e�4���8�v�_����=҆֯R/�^��E B�N��!�;}JҖ��{��A�����cv�!��O[:X��=�4�YD(۷k���`��*�PR��Y_!�BjQ?�l���cw����k~�6i��AE�Qd�%�*���9��s��W:1��ǜ �A�����J�d��A{�,'�UZG�ʼ���zD��b3����K��s�"�h 7� 8�Z |Ԉ�Q�U��:�ّ�e��r�v���N��	���,��,�wo��Օ��P>ho_�֭��4��Gfp���`��}�ғG�d�r$�;:9�G�B�Bw�gQ4R��Ž���]!��'���e����\�^�ǖ��L���z��]��-��no����F�iw?tv��	u���iq��=cg~]E��"���%�vtpN��.
�j����`�^��g3&K�՗�̹�l_�m����?��}nz���|�z�G�0����n�A]��k ��N0�5��<G�Si0W����U�6�E2����[R�����ꨣַ}n@g��[@fs����jG�b0�S����	��$���}F@�'L�ǿV�؉:�򹢳��ׄ3���I�YԻ�к�:��w"�����2�lVE2�����]F�]F~�:|�p��lSV��-�ѕ���nn��SF���&'��~[�a��#��}9S����>�J�� ��e�5�}�i4K�:�̞��w����ԊT�O`�BD/�T��b�;O�	�`:Z�}� w�f8/�dZ��T�-W�Z�h�ש����2�(m!+π�ﰮ}��Ч��>���X��T��s��P�����К(�r�WA���/͊1~�� ��y,C+M4�I���y�[�#Q�nu7�z)��>�
��E���#�A�j�n�hRsʉ��^Rό�=ϲ�tvv��O��\˞�	�/އ����oB��)���~o��YIn*%8a��4�g��$��T" ��ȑ`$�Æ$��	#B�+@�ܐSG?��z����xnx2O7���f|(�u4��P���y�?�/^)+:3%�>sR����0���HS� L���0�׊�a��밙�X�w���@�5�|#��!HQrxV��S^W�<��(1w�,���eص�udAV�E��̣x�1�����!<~��!�@��G\����kehdnD�
*�k�\��U��NSH������a8{���ʮ@d���v� �Qҳp���!���!$��Ss��l'�%��J�Q��v��r��p�o�U?֞b�5hRa9�����Y8xq��V�[ ��d�,Cl(�r#D��ϙ����������V��J��'rΡ�%3����ZE���W��l'�o V�~�~|�N篿R  ��1��g�����yؿ��`�k���7߄����C�����pfg��=v��O?� ��>*�l���B�Y���D7�>"H�x�&^��չ���;ـ6����=���������6����Q֨@��ډ9�O�(	���
�d�|�ϳT�A�v$�'xtN�Q����}�L>�(-���	�t��Me��b'��#����������6e������ʖZm�<��3�Cq�G�������u�۽���Y��45�0{�il��z�G�^G�ù*v��Q�8�{�x�PLs�k�ԭZ$1��CQ��so�dè*��۰OÚ9m�9*v������������''�vڣb�^[�2�+�T�l��^�!�'�G�1g2s*�3�wu%�J���r����E"nF�Xl�g.Q��,n���8P���(�H�1E��4���γs���Kg�0��Nx�a�9�*4,���{��W�e6�.l�d<�QZ�>�7��#�g�*1fyU����:��#q&x�J���TŲ���k�{r�(�g �N"�﫼(������)=��'���d2�r�̈����zz1'l�Lh5�F�@�R��]>@�*�?@$�>���q8D�Mx�#1F���[�v��52�"٧2L|��'+����ұ������b�g.F"J|koFK� ��i�)<�A�-�==��w8pI=h	��d�.�'�tw��_hi��Ã�p0ܕA��Md�r��<����(\3�h,K���g�k��	��R�K!����@ڧ�{� 2흝�m ��f0��'B������e�Ex�ؐ�d�3��J��l�ý&[�w��/[]�d���C��	'��8pJ ���^���8�>>�}rz"���Թ��`�'�VQ���H�&�kWt�ʮ1�h$���o�Kx�fl����+`�OBd�K2�4B��D\���"�x�Z��v���<��bVF�  �Ү�������U^���`x@��9�o�IJg"��|�,����N�0�;�<��%��	>7�������k^�Sv�`k�1ld��`^��F�Ҁ�˃���6+}��1{f+�с��zUB/���5��S�#�]Y�F�J�&a��~s���S�������� C����(<��R8�f����V�����ml8JT��m�8�a9� ���O�Q��5vڋi��q�e�IO��ES1�M6\��jC�Mq��a�Q��
?_�߄��Q��;L1*i��#���YXH�X��E ����U�Ā��H�)I�L
CO0�o�K�����XT3���6���e�u!�n�B�2Ľ\�TB��_~�_���w���C��J�4��P9��|���)#2y+a�*�p*�㨋��uT�Q�P�Po���hƍ��w�w�Zr��AK�$�8F����wO�\i�H��"FO��҅'r�e�����y�i��Z\\]jV� FT��'�]�̵y��P�B��&/�<���3ͳ�Z@�0SfK�(*�5e�rg�P)/�|@�Ӱ��[���*����FtZN;`;�P��96����Y�z�X)[���s$f�׶����B�v���J���@(gu(b�*D�SG��14�'! W�AOӭ���?q�y�T�/k�"(��+X��B(��98����99p�a�+*@��+��|!ǀ��cCL����e�)1�¾�5�� �lJ�]<�$�=���I� ���S���̿~�]����ێ����cx{�>��s�WfЖ���p�0<yT@z��ܮ������g��������ʾ��>1�S-sr��Q���	��0htÕe�3{���~߂%�뛷?�D��9n1v�e+#iG�7e�%����)d�L�&���>���1y�
`3�Zz{��mfm��0��/��b6�
F%�j�~����~��Φ�[�@���G��Z��]�Rf��猯��v�=9h����@�rh� #�$!E����P��i |e�؋��Q>b��pg�����H�+[ѡn�<��ڮ�y�<9ֈ��������@�QTU���?Dv��۶�������fo�Uu�/�q��eEu�H����#�	��o��y�U#P��N�l�$�cK�3�oA6�q�����E4��["	��١E�h������EN�i�:pG��gm٦���x&\I4���6�۟�~~�s.+�΃� �N�rL�Qd8>&���xQ�M�D&Ls��ߘ/]�9N�q��p���iwv����o^�C3��?��ǁ��y�se�V��Z� ,ﯮ�[�4�,Rz�6��=܉���������T�֫�R����K����T�&��Ne���Ml�p:�dp�g�d\�?���P٘��G���2�����:gjRVI8A�U�'0�p��N�+�c�uh1q�V�eZ{Z"������ ��/�ۑ��g��^w>�|f�C�t�����Tk9r�0W=5׊�k����Ux����� a�������Fdh
۾�ۤ:s��,}NY���ف�dl���j-cH���j�?P�� YD��m h'�G�G�ҲE�C'��,bo�Q�9E�Ct�����ks ��a�Z2���>\�*�#����վa����u[XVԨ<��$����ah�kU���zk�����!�;�?^������G��gZC��c�Tdw�d�w��!�/3g*�|sw����v��Ë��4�Էk��t��2�A/�-� Cм�}I����T����V�3����D��49㚝f�)c~��/a�8�x���p���狏����UY��XXۂ�Y�Ld4�F�q&؝��k'ʱ�p߼�ßµ}6���ٙWdZ]U�R�^A�����8�a�b⢕�Tҏ|��܂�����8����m�[�
��I;g�O��<|��^���Ǐ.=9�v���Y�I����q��3=�5�)�f�dS^��$��
x��r���X���2�8���a_"����d�$Nm�m0�&��T?�+y�﹢�S$�'���*&��ul�����M��?�6t���{��w��o�������`�~��)4iA�h�P����E�:�8u-�ױJ�p,"{AP����7����eNx-���2�$��:�vĹ�T�,]�`�,��T~��D����=m�"�p<,���}er [� $8n�`d+7��l�qRO`�r���՚�4����S;������W!�aS#�n;�ȴ��Ņ�덒�^"awZNsvy�)��x.�׫�d�fd��h6�>^BE<L��ܬ�j�S�c��uYľ/��vG(�>�����ڝ�Gp��UNK��q�Dh�橳�b㠼ǃ�f����K�8a��gu=ZG:ɤ5+I�TƊ��d		]���R�c�4�5��� �pe9���L�_��,c���������Y(ON4k���F�b�;�j����Q�d�D�iNk�1�]���|{.���,C�z�-���!*�[��߿{'��#y���z��8�����Y�qn]�S��ڋ�ً�|-��KIKvNN����ʜ0��R�Y�5�K� ZQ����r����PA��j��l�u9�?�T ����]�Y07m���i� }j`=���ޛ�F#��S��;�l�/?��_����/�� �>����P�����>��H���������%���S�1�3�۳!��aR�P|ek�o�G��[�g��	����ޞ8�����;f\u��e_�&OR%�d:��YF?����mt"Ǻ}aR��HO�Fu$�X���g��H���^�s[?o�9(�L.��K�X��s�d��c�h`����=>�`?Ae��8��M�@V#sT#�ʫ�\��#�#
#�-�2$���<L��4�J�L�����$(Sf��'�/d�V9�3'm �%,�~��*�25�pUbs�3�-��P�mBO�p�S)�����q�(�ގJ�6���T΄�M��޿�J��[@��z���鐩��Z_�ȼB��.i��f�N�pn1IU��=04e�W��
z���ĞJsD*�f(ʛ/"(k-��+����E������O���P��3�Y�n�D�11�0z|
�_�6���2���m��-꩎�H�	n�"�H�	i	ٺm�1�v�Asɢc�aHB��Y���͛��凰lfg�� e�:����PYtg]�z���KkY�7NR}����"�EwGΖ95]C��^�&~c��-����@K�A�|�7K��"߬�6 b{����o,�ˬ G���	�lR�Ɣ�I��ې���#&C�9Q�84��gA�=���T�a���� s"��F����y]?N�����ѣ^��a����޼{�����)�129�~S���_����s'���:�y�r��݃Pͧ�\���C�f�ub{�1���M���������s8�33�"\	����2��ͽOZ2�X�6��x҂�g���XZ"U�pd4e伎=[�"��|�5�[T��ĕ];,eIf�8���n�w�a�0'�(TPo��M��.z�+˴LN���������xmY�P}�`IZ�Fɜ��n�h(mm�w{C�s�	e,�r�JOB��^�9��GX�9O��{���q��t�z�ڗ
j��+]�>W�%�_�maz�6^F�6횣#Ϝ��s���^9��BYi%&1z��� �v�?�^/��c �Mҋ:k���h�)D�4{v
a�'�)�'����\���JN� ��JM��-��)s��9!���p~�������d��-�6�ѩ7���<S�����@�3B����Ly�k���w�j��+�8Δ�:m�$����NG>GX;Q�97$��"�&#�h�bhu����s�ģ�Z������yh���ٶ���"��Z�bљ!�脿��p���u�r��a�HE=�ύ��!(��De/��K�h�Ɉ���Oë�W�l_���\���{������/᫯���B�(����EĽ�����V�ф�� fh^���OvA��d6�9۝~�ن��7�{
��2��2��B��`n1Xf�7��)O>���Q8؄�� �B
��~]��f�nԞi9� y�ͩh0T��{A3_X�L�����k�S�3e򷟮�xY���0���ܨ�$�5�����2";��U���ی,2d��F;@-�Z1�~J�\F����vnV���2�C3l��������^�އ��.�ǫO�T]$rv��F��w����>�#\s_{@bR��{?����۷�?�{���P�D0yǠ݉��B�V�\���x�e���{wsn-#�����?�=_��R�4�}uo����'3�v_�oO0׉�]]���������K2��]?N���+��޶C���]���D*l4{���X�v�{a%�,�ؤr�2A�~+��h"��r�
s Z*[�4�_m���7��F��糥擵'bh����XS���0���?��C�?����"xd��to�fE�K��R����]��� ���\����αʱO�3�,FvɄpFi�FB�ƈ�J�R�@��c"��j��3z�n:W����uߏT�������L���2b֖�������q� T	��-�{���t?�x���zf�ml�$�뻯�Qٝsy��c(��� ^<��=�î���#���g;S+��.����FB����ٖjn3f��p'�}�զ{���9��q$���g{�����Ib�,����w��\��9j� �<�+�*K��>�3��`
	^x�r��݇�㻟��ƌ����;_A�l�Ek�}�@e/�6�p�cV�r���f�R�����e�8!\��}3{e�a�%�-�O�9���S���PjlE�>F3(��ܒ�.�Q��g~#N�4:�{�[�ZFE�J���u|ʷ	
�Km"n��՜��յ]�DB�D����Ww�!w@f]JӅO���#�Φ,�S�(���ӱ���xd�k#�:H&�-���~gIwmf�zj�o�	�i��SG og݄pUo��̝�D�lؔohBJ��`���G��ġhl2\����s۠z���9�^��z�x[����W_}��o~�y�"#�g�{�p~��
��-\ܵ�T(ڃ(�ĺ����T(Z���h���p�p�K� x�y<��h@�|��y`]�8(�Y�LS���Ҝ�	���~3�%<s>�%2<H`D�NƂ O�	R�F3�v�����T�U`�� ��Z�/`py�/t��)@SLG@˞�������S����)����('AKf����t"�
��W�c��f�5�r�|eG;�R!T-��s���3��M�@U���ԍ�����P�Ȉ��, >��=���}�S��0� D�..��o����򵸔E�R%����KK#K���d@���Jǿ){�G��v.
�+^�(��VU���j.%�����:E�Lŋ����R�2n�/P��� �}�="SfĈ���i쟭Z*C��Fu���Ȟ�-�8�ut��Y�Di�A�'�N!٣2����q���(�m֪�HCx�}z�m{���E���忿DYo��dY�̐�߯�vP��+��N��z��ᦂӳ3�HH��ғ)�Zr�ә�녝����{������&0���ަB������I�������`�͑�M�F+OLWE��D[٪3��iф�˽�_ƨ��63�R��e�,��,%���s������a���~7�^v��ή"{ĳ)ǰ�v��	��/�`�w�`�� �1���F2i�����A��4�Da������f �ro�ݴ+;8�0�P�;?�({6L^58#� �j� iF��Q�������F� � �4�7z�R��@�D|�MG3��e�7?`Z��s�T��*�Sy̤͠Վ ��ZQ��0}/��j�?��%����՞ظ���@��K⡞t��\Yy)�|v��ٵ�h�ʜ���v/|wt������A8�u��}��C*0Wf;��3�s�Nk��=�ʫ��ʴK���o��*Ý�����o;�)bfm���P̙k��́?h�6�����b�s$+O�3X�F���Ƙ�� �Qo�=#�څ.%G:mn�pRT��rv�(�>�Z�*@�W҅�n�{�*�),��}���S�ͣ�}��G���|,��#;#G��$6bS�R���axqz&�:�n�%eV27Fr4�����Y��X��0
]���8�^q���h����a|gN��%�`��0!ȃ�j���HR8E�r�恾{cZm��ڹ��~�JPhk�u�vOZ�؞|F�͵�궅�e� ����Vr�-F�������κُ�5���!(1�$%$��ImCը��;����'��Y�e��F�l�a ��0�}��q��?���l�өg{�0:v=��f"������
����S�
�3��U��rz��B�Z�<�#�!�H\_8�"J���A���z�\��v�:Ù���F�<zNL�eX{P���,RS:���奝	;���,gZ'��
��̶ߡv�ID
PQZcLn.~���Sg��1#p/�}v�I�vJ�}(i-a�M\#�3����X�׫q��pȋ֪h��;Ԃeޛ�܆�P�V�C��m���@�h�y���Cx�>�~������I8�?пYh�+><�lǍs������[6�w� !_|�P��h������k���xb��&r�3,�#it~��zg�ԌƽE�h���-8�]	1�qjx��o�<�}Ec�;��b� ���vb��J��骨�3�r����gI�F����i���W�:D��?�����J��2�@����8��C���m��3����p�z�g��1�]���]z���{�5��	�,�����f8l��.4���2zk�Z;��[��^ڽG�G�D2w2|��d��e�����lcY�6�'��R�j���`���u�(uM���/���B�Z	1�C���]����_�?�$����d�����B�4�L��7`*F�P��1�r0�� G�����Rf. f 5�	/Y��#E*B��*�",�b	�B�a��G Ek�.=3��D����d��D�>@N���B���������*�g��ue;Qo��f[\�+0B��o�~G���V��b��Д*h�d��ik��z�d��E�Fѷ{���w��M�'k�V|��Wv�%l ��S@5d��V�}�d�K�nn�AD��ZA\���_kl�-`4c���+���OOe����(A8�4r���u���ݯU�ӛ��{�㈥��ʾ�+�*������:7G<~xT[�}���� �̨��S��ͩ@:�%�Ja0��`_d ?�ưtMЧ��)���&��ck�ȋ�@���.�G����Y��G��*K���lS�H<63±2���✨��̅�[��V	������������71��a�*V��lM�H�j1&�h���i�W��-5nvc�So�\j�NJsPݎ���/�����}��y���	�ڽ"ೠf]������	[Ըj5�sEI�tcɅL��mրC�ʜ�29 q�ԎzQ���%k�.��	�NO3���l�a�,V:<�ww!�����)�%r���}�t���o}�)��p��j'���=YT$��-� |��8CF祈(�,JW�$f�[q�B ��r�+~X�8$;$8i�nz#�XkW�H �<f��sM�ţӥ��p�=��r�(ɛ��1��t,�5c0�t���A�[?��Xף$������?��L���\���H;�8C\�i�:b��;\�2���l3��-��̉@�ݎg��{}9��� �>��N�L�Y���2jc��ok��{�4D	�o��<�kEA�H�"�<�Md�*��[�@�,���=N�Ƚ��rr||�C�,҅�s�������?�7�7���bn������1#�(�dP��� �Y�&�{��P��x?��J��ӛ��$��	Ls3ƔѦ���QMl �f��ͫ�0��� 1�ߟ�ވ8l�Y`��u���֎�l�$ǃ�d�Gˇ����XT����1A�Y���Ἕ��{�(Q�<��>31ӥ�����1V�+%);{���G�V��Ͼd}���Co���LU#�k�蛲�OO�	-�1G�R��7`>�{����U)G�X@�p��<|��o��W��.�ۘ�NT�go_�Gadgl�muxV7�m����{��}����0��WO{e���ec��' �h��������Hs�ث��]�,*��Z�,�v�ߋ��²�Q���B�-0�uE��U�<VG�X�����*��N��ǗNvS:��9��T��7���jd�kʄ�3�Y�#� K3N�)�	�ǩ
拳|Ü�Le��&T�~���йj�����V36�
�pb_p}P���'(xkg��_�h�V�f�Àb�i���G�Y;����"��c�|�}��/����7?~YO�,�,�K-|p�g؏�b�ֹNd$�Gt��7��؛��m�2��� ��hrl�(X��XF�r�9<� ����
����Ĕf��~$��{�ȗj�8��4R�"�vˁ;��)ݸz	���L̹����J&��^���S:k���B%��_�ǔjw|	�E�7H帆)��]y�v�zS�f!��r�'��:<�?��=�MVI���H��������C�.]�>ɨi$�ֳ#U�M���aia~ya � \ǡkWIowmι���P
�2�526��}@|�Fxa�ksX��V�#^>��)rS
�w�E��)k|41����MrU M,�}|�o߽?��1���]x0#ɜ��.�46%�H�rq��`�c�Q�w�Fe<�!�3��c'����2�����D�|����>f"��B��@=�<>�������s������1�u�v�!�	��/-�IF�s��\$e��2�>$pW�w�?cTd��?�g�4
��Щ������^�m�~��B ��會����̃]Tl�0∢�cϒ�gQNe��}��|&�V�N�y�+$La4�xL}.^|�0F��[Π�d�\��,+���S�#j��9g����x�s�)&뤗;6�Ț�s	 �')T�г�z�	�7w�#�0(�
`x/�W�Ӫ���ES]�Ŝ�)�|.,8E�܉�hwd��!9 �:�e�D�����Kض��ۏ�hӾ��S�{�W��mLz�6�:ԟ��#5�2�M��4-����KU��������R}��2�>ˮ��T%��w�eNŁ�7�����n�k�'��N#Q�3���ݮa�J��L���-$�c�����4����iN&���<"��T�E���D[�����&�D���X�)���͋��9S�����N�2Yr�`�UD��w����W��)*� $�=���W�'�gv��D�Yȑ�� ̡���E�+��Pu3X���#���EV������5����E�ń���Hp$e(��a�X�I��>,7S;`׷w�i�mj�J3=);3�X0���1��2x����LpyI�`�n�|W"Q6m������C��s"���j{_�}�}�����_��e&o�h�B+��������̂�^M�xN,C�VO����:Bf)�&�a]�447Z����A�<2�-*BkGL6��A�Fe�w��>}��l]�Ңo�7�Y���yƑ;�S'3jM[bw�p@�����++���K�6F��m>Y��
/��)C���!s��a�������� ˙�������yr�jLmo�wʂCD�GGiY��L�s`K�QKT��Z�FvC�/ }=��%I5
�$�m	�m!�v��UYP 1@��޳�
�
^	$�*�倛"쏆�����#��{/)Ͻ�<իN'�b�G�H�*��yx��&$�'Y'�v��i�7�X��A���,�a�ݏ��r�T!X-&���X��+����	t�ٍ��ImnN��2VH7P��s1�ts�I�kdNw��Й>��^z����A_�M���(�
f��eN��2z�6"�w����o�.j������:r9d�Tc�U\�t��:	')~�����L�01�H�6��Qv��%\Q�7L@�,�V����ݞ/ָ_!��X�Ȉ!��W򁒳0;��Sȃ>Y�;.	yٖ�6�)��~/f�~�-�,Bڣ�[p '`�nS@Jt����U�|���	�u��,jʒ#��(�R?Q7Zs�>a��A��˶�eN��/�gYP�(d��X,=RR��
�k�OO�C~߲�}=�v�������20ܖU?<���;������$08�A7����@+��\*���末v{[=��K&�͵�W�J�����w�Q������2R����_^��z
[T�U�H��2ʷW���l"&��U	����8w���	�#�z+�H����H���mEƉ�*��8������I�ݷ߆�e�d��a��KvyzpV'UF�+��8�����{!g�n���JZ�+sX �V�q���IPHJM���ƫ����Ȏ�����~��P����Cx0�8^LT,m_���XVMs��?��i��它��p��^���S0	��
��=��1ԙ ��Ge��[�Z��Q�7k���΃e�D�d�����ؖ4��Z��ul����F�{ܛ�l�8t��\�oAeI~����Ո����%oA3�� L?~� �U�~nS����;��/@p��b4�$�<'5�C�zt^����e�$M�-{�?�S^�
X^2�-�ׂ�.�лFw�i��,���������u�ԋ0������B���۹w�؎#��i'�eS�;�m]F%o�5�>S���J�
g��v���g��V��Sצn��M��N,���BR�+-�gZ]� xu ßUmٴ
��ƱN��%1h66�x6��@�	A�ܧ�"k��SDL\[����Β�^nl���6�����:�6A�#^E�Q�H�'�,�{נ��L��@�F��O[��8O���3WD��n�n��_n�_0#�)sJ01 ��.#K��ҽ]s��Ph�\e���<~wtX6��j%�M%�Xnu۰�I��f7��J=(��|b1��l�E��%_�:�][�ٰ7-��o�mb�(1�c�M�&އ��hy����9+^�ޢQ��>%�񻼹��ͽ�~<�<�M��,ʆ)��)ў��=��]oIt=� ���%یqU.C6�y���<o��깤�S! d4��*��Ĵ��R�%B#��v�� "��*
dp�����j�}����48�z���T��._�Y�^��Jd��c�m�z�P~��e����&��peN��>� T@
�L9� ��6�1���:=ǖIA�����ûO�4��4�-V�.�zR&B��ʑ���u�S	��Sͦ[�yEVy?����o ��zꩽ�uC�T��������u�yײ/xɿ������ �#G�V�8���И��ӓ�������ɹӆ�nlYW2����ж�f��H��ݡ�Qp
�]���ƒ!�RQj��> $U����W5�RtD#�pa�J%��iB�(&��C��(x��	s[�;s2:�z�{N�(�9�.�}	#E����~ �y�3����M,H�M�*V#F��B�`�����A�S��}Q�#Y��v0�+�)��8r�p�;'�	
�E^��6�@e�,�#2����Jck9[{@�J�
����g��s�ߺR;��J�ɠ7��@�����ګ3TX$t�Od29	e���W���]*7R���DFP�R1r�67ם��y�%e�ۀ�M�x�ʷ���3[��DR��j���1�B���ͣ�~�*S��aS��kJ�!�l\D7�2\����)�mBHR���v�F\T�j�R��t��m���;�^�[>�V(��}5�O���`Z�^'�5�=_YX��f�����RI��U�'��Z�D���x'�3Bm�?��c�~��2s�A��˗����.�f?\̜S� {#���no��� �_2a���b�A	�Y}�r	|`�d�?���8�)K\^�Y�5g''�����vV���+8��F�3�=k2]l�+�CXG��g��th3�hζ��{5��ن:�ˡ��n<�"�����¹֬JB��|�Ol���R��� (�(I7=���m�JPQ�,�;��b��K<���hȉ< ���rS�K�x�������{sH�z�:\��6,�hN�*�A!�8��e�1O�_���F*���;ݝ�:.�jY��Ճ9�g̚��`��G�v�BdW���	
����}����6��W��p'�x
�֮9���=���|�A��..ã���R׈R�L�ʽ����+�n�}���0�������)���-�q�3�q�Q/���ю+75�����%����������;����p��� ��n�G���
G��unn(e�\�|�4��_Z�9�8z5�u�Ɍ���^�o*�cbB����{��|y'rU�$C�������/�'���U�G���;����G����9��f����	�֢��Ϋ�����3-H��9 �A���l�N+I�y[�%�T<Su���y{�rd+�A��^4��ð7�52���Q�a<Kc��U5ڎ�������K��^O	D�.���R+!��#��� ���l����,]LA���2���
�X���핁���ܵ~ɐ��N����ec��3aMhl%_��$����V9O}�d���\������3۶�zcP��k�3�y�AGl���(����BV�U�S���@u��b� ���n3���c�|���*-�.T����J�"�
I�U�:���i��ʆgE��[,���������a�H���m^���8� ��lVo���D�40��'˂�`ᄶ(pg���0�9�hDs��+�?X��T6�������f�;��*��
[�%s�+P��гC���{:
W�WbM2��9>J�;s����~+�=�e͉f. "@ݿeG!n�*)�M��*�W٦�Q�nKrn<��=Ē�X�I��*� "Yh
I�{p��n�?�S9�ü C����jD*�z��Le��Q=c�b����ؿ�6�'	��G3�����]Ϸ/_�����d� ���E��(��� �f�U�Bs�d5)0�-;j��4ON�E���G!�ga %���%i�`�_.u���_�|^��2gy0I��K} [�U�>o>������Q���N���%D����,�(#*'H���B�r�:=����@80�N�\ʊ��ܵ��s�(��� �8�oB�_��8fÖE=����M���+����1(y#���[aسH�2���}/�]�γ�Vt�!�Mp��ƛ��z��L�����j������{������7cf�3�Й��'(w`�"�����_"ۇ�u�� K��en ��@ �i���_#ή훏o>��ŵF�i����F$��|�/�Gh?��|f�n����_m�]�����c��=:��r))��L���r��k�%b)�5\���,�A:cfyrN�&'
�[6�s���>J��5s\iܲ ϥڠ��K��Ƴ�L��w��[��&!����*y���������3Χ�,kN�w�L#���.��L��_K�2j����;�䀫�ޥa>|f��+}R��#�5�vB>	��{\V1��9�V�9��ng�Q�$�t5;x����q/8��T8��kk3;t�YGe�> �����F��R-.�J�48::����;�oQ9s�s"�ŕ�� �Z�؁C�Cw؜�
Ҁ�X��拷��էOr1��tP)�P��P;�6��{14����:b05����|�!g���2�ŵ�`*��ic�x=SX�8W��Kt�6˯'xT��l8	����&���G����&kĤ�f�{���������ɩ�{����{���RF�I�����R�_��/��𑾋�*��6�[�utΠ�Wq�G9�ed���CE:Z�S�Ǜ+e�ޡ�:��۵�U�4Ԧ��2��U���YG��mƤi��?I��9`��^R�&H�b����1�����㴦���<J�I�Ȯkh{�����<���%Ty+��h�Įe����Q�)�����O��cCօ �@����@9����p��7�2��N�$&눌�Ϻ�7�?��ѽd�\J�񐅤�G{a��$ώC{��kᖔF�b�R����z5'��|�
=/� �����=�N��ݖ��y�d�WWW�ݻw�~��޿��>|��xG3a!�<�l��7|���G�'6�	wt�|��֎-�p��~Cקk��S��O�8=�;R��}��r�gN��y�@s;g�B�đ�P��?�z�&�wfԝ���no�3k^
��[,l��`�#���.�Y�8�Μ�o�.l5Vl�Z
Y[��3ٖȼ�4�^�O��γ8~�z���Jh�M�t�	�ϙ�h�/���0�[���f��#����3 ��*?''�D?�xΥ� Na�qǂ�~�EkS�˲�x��4�
,��&��L �,�\k'Q�]��W��]�=0`��*�{�?&цX��^�B���kU7�\���^mU������/#�4^��Z�I�M���_0�T >̱��R�4;|gF���N��G'���\s���}(;�q����?���,�L����<d1�^���5���f�R�>[�Q��
����H��	����E�Wz����$���e,�83 m{�6�a0�HX��]����z2d��
�G��s֧4��H��V��&���3q������e�w2��Ly��O4^���q��<���_�Ɠ0@��m�_9`HJe~�6�[(!J�V!@W)F��2;������F\�6 }0_G��&��/FSe�߿z�����2��Ry�b�
�9Y��&"�B��W��x��w���Q��ޮ���4t./B{�U�Qb�N��4+ae�ײi�:[+0&b٢��t�͝� ��Fۅ��A}e�²8)���1ː���C�2��M�ȵR=�j������H��˂;��S9�����Cx�u���cW��UGs���x��8��о}FvR��N��3�,�Q���L��,闊�۵^�kz���^LS ��R�]*�*$f�d����γ�V�/��q��W{�����J����qy$h��s��~mg'���!���Ƣަ߷��]���CI��af�y޾���K�x��v�{���\*[|*�&��Ⱦ�W��=��a����7��u8�����0k�n�ٛ�$���>��щe�����<�I�Ƃ�ڂ������t������
K��&1NӪ+ ��Z��4�-�]��l%��F��vv�����L��8X29fRlb������]WY����Tʠ�r�^pMY��r �38*��$G�'�3Ͻ�1 �yK-�R7덣L�������#ɲ+����Rg��.���3�;C3�ښ���1�p�-�U]*5�v��w�{��-4��J"ܟ�w��D��Ν	Z��'�4�C�N���c�ߏ�c�K~U�t[�̂ ��s,�e
���YP���N͎P-�Z.�5F$�	*]��eǖT��fcS�~��[gً�q�ʖ��ӻ[�����퇍�/쿋�?���ݲ5.Ƭ^���{�vޒf&_�"��i�_��A��yG΀����A�����u#���ڻ�h�B'��:�C+
�E��2� ���k��=q���ҝ�4�>�m���<e���=���.f��9G�#{��7k��d�o*drx[!eF�"�2�}�r��5WB�����!����c�a<"�[:��F&r!�ɒ��D�1��۶i����f� H������pl�/m�,�Ew�і�|D�I���a�~�.Ա̚g=��Db_�'җ��H��E�s�Y,
t$���=�<�,ۄNo�7�+i㚳�XWν9:����Pd>�ô �ʲ��=7V����Ee,�XP�l�=�z�LAE���_T>u���W��@urs-��0?ϯ�(`��y���;T�0���l�*���;׿���*v-��l`B��d4?��	dXf\qXK�f:�Bo����p�ټF��,bi�0��
/��7aX��t��5�3c�6���
�5v��><<ۇ�a`�oNٍ����-��Q��,��SQo��c��3`eY�/<�����[,(�:��-��r|�!�ɥ�K�k�����'���F%m��%yI�aF���*m���?�liG� S�zFo�v����n�y������Q��}�%&��*NK���m������n��ޱLx�c����~	n�-fO�ӳ�3��'Ol/��K�ް�F5��jTך�R���Z�=�$3���5��Y%�h$0��Uo�$�l�hWN�3��U@[s�i�f?�+��&&!�d���!�9���2�(u���{��ٌ��$Sּz��K���'Qi����g�E�׋-?o
Ft��_�U-*T�4G�m�B�8�
I��vصgu�s GI�&: r"�
9���l;U,Ͻ��Z'j�̃��'W�.on-� �<~O}����9�n�7��vFx\���L}���n�j��Cep
 ��7�
{�j��4P��c������Z$ۃ���Qs[�[�F��[E���ZyQF���r �r
�����B�6>'G����
�l1�9]��RUߓRd^҂��c!��L��z�-��Ĉ��o��}�4pB�㼛�i�b���[��R3E�%!|Ŗ	PVő}��?�Ȝ&�ʓ�$t��BN��.�D����gDE�W��A3�m��;@�TP�*�*J-����P @  蘻R�4N�X�3xrt=R�DlYf�jS`��iC��J!fD�q���_xl��|z�������kEI�uO��ت��o{��o���%`^�{Q=#�b�"��>�it]�U���d�����^Y�nU�j�CjGb�:9/��F�+�F�Ԝ#Җ3˒�_;ا��r���]����a�#�j:�#%#�mw�P���^�Vs��o�%j^}aٜ���FLIbs��]qvom	,"|����v�!u�j�LF&̆�J���<�������Sźo'�Qe:����`]���Rl�E߷}3|8��eW#h��\Mb�ՒA'�MJ\�(R9��� gg��eY��!�n�;b���U� Ԍ틧�Z�L�>,sd��.� �Z�HQ��KUg`v������M4����B�pڔ�A��3B�b�����8�?{n��C��s��y�'��zk��e�]�&Wu+f����VJ^6�#����!4J,���@���*0ɴ��G��ѵ��i	 B��'-?R��L��U<�'J��v�DO%h��"%�^	����eW���O�2[�|4�Ը�G��w��_��J�O�Y'����K��Ad.񚅍��{x��$�Mbڭ�y&�٩����6%_q|��R� .	�CjC�{���1`��8��X�Y��� �LK",o�'\d�E�SeO<o{ S�� S�(fD+U�l5Drn�S�s���/?�"S�/��>�/�l}�\ڔ{q	}����!��o�-j���}�2���_��}ѥU��s���1�"���YF��y�� ���ō��K�tz.���2�!�ly �U�*�M[��E���ce��?�!/p[@�:�71`��l\�<�}d\\���^�,��2ܱ�?���8��w66B57a�I�V�I�� �4�ɂ�h�C��R��_rX�����l��p�����hcS����gmk{su��p��Q���~�Q!����E����0Ǯ���|r�2&�����l=?)����L}�n�Z�8D�F�9`������P��r�2#J�#�X6���措ǹ����g�����iͰ <:y�6�l�t۟�/>{��a�~� �����-8y��}xl��}��:����5�X����T��m�;�:?���^�y7�A�v,�ꘑ������M���Ie�L�%T':�?��cgǢ�Py����GX	�ⲓ�r��pr�*���3s��R/���^rm"����-�[У1�θ�7���-e"��\�#��+1a:�=r?�M@i���r��[T<>V`�z|�~���0�Ϟ�g�B���e?-s��~z�?�jTs�fp�K�){G�٫Wvv�a����F��d6�R�?��<�{~�8<�g����_�,����U�����gD�.*w�n_�˻[6�b�=����9�����v��p�k�3���LG����vO��\�rj���M���Y������ӢX�a�ww���ߏ�6}>�A ��^�A'>l]�����K����y
�X�kd6v� 69�[P$'���z�	��t��>پ���Ʉ���s*��*g�i������[}�`��Ix|�(���� Iߖ����)4�/i����G� g.��R0FT%��g�H��/f���S�n����nՔ�HZ@���jp��GdN:S�@c$�Qۤ�{�aی3�	=�*�=VN܁�e ���b���\Q?����f�W�dx�Y(/.*�l�s+�sf)v��v��0?�m�M�^s� �"
�Y~re��n�X"�a0ʤͣW���yrq�Y�Ү�ekWXBƯn������X�*�-0f!Z63�g��Y��O���~�J��(��݅8����Jq��ٽ���	�5+��e�DPǽ\�:rV��E$=nD��x��s����C��Y��y��G�-0nV�4�4M���s�2�vu��Q��?��t�m1a9á�Lc5Q�}��	������ E騿7O?G{�>Z�o[��g�l���gI�^T�]��FZ�4+��(�4-��	�b������ot�B	[G�GfEo���F� �Z��^ח���ݑ;�V&2�溜O���?�l{��蒠sل���e`@硜.�Q`Ш\Y�ʜ	=`*��P�P�V�\��d3Xgd�L�O���j=��a/
��Ȍ���~;���ƙ�s!U�LL���ef|s|�u߽��限����[Y#�ݲ�YI���q,����F-�����uڿOf�f��Tfe�bhv�7ꇻ��'��s.�n��`�û{�������-U������f�tlg�O�F�������8p�.�P�8(���£�Ga��U�Zc~�ք�N�1˸�f�3'o�DF�XN�5��;���L���,��DU%?+�,ff��m)�J#B�걊�m�p����?4�\�0�,��>�z�=�W�L`T��:=��q��`�?mm�PP!�+Є{�g�Ng�ɪ�Nc���/>�<�����#�&��������mo��\�e:O�sә�t��}��T3�^'qlyaC�@�-�/ ����a��Y�`�Z��7�j���6��Ff��S�.�80Fc�g����f��V�q�C˘����j��/F<0�<���Z���6:Ɯ��2Z.����� D8��K�f�{1jw�me��.O���~H:�;8p'*U%�@Ap�n[�v`���ᑐrU���e$�>K'�|�O����pD��v�J�����At>~r�rݧ��U�A�P �a���0f��ZO��=q �P=.c&���q�=$!my@2��?�'3�������z�Q�����q�2���POunF��T�"� ��[cs7�Ѓ�e�%Yʂ�^q��^w��!�.&3֭�t���b�d b�����1cI?Q�ϟ�y{���޲���E�p����#�ڴ}���IJ��f�5�Fӓ&��7���%Ƚ��вlil6�����ɫ�9�.�9�ϴN?��>��JX���`02��y�ʶq�.l�3;Cx�m�������gfh��ڇr`z�RZi|�KS��C�]��9��#� 4>BEk=��t�r������tV)��[��	��3s�p���	N�Vc�f+�3��)�����8B�� 	�';[˻i���m�G�gV.��]z����F��,yik}gϕ�������Ȍw_wA%�������^�S�86	£�ii�26�7"�Az��eA��g`?{||�ZչOP@)�C����a�s���W�_�/^~f���j��pɪtQB���ڂB�]/,h��-#�*	�9l�܌I!��������׿|���I��%��
�����n��O���~�+q|2���@wU�'B������v�	%�m$�C�H^�x!���n�V�̼��h��a��\Y)�#���o+��?~/�46������}MelmnH~��?{�=[�s��/��)�HI"���p5Q�L��j5�,�������ww��~��/,G�I̭D���>:��KЋD��~�<��/�����f*y�$��[���4z��a`8��9�m���`��<�"f��9��`�	�J\�+�}�7��M�Big!��eby��}�;�����i�8���)mon�/^���,P��������k�,||�d��@3NYˁM�3̼�����m3�G�N��h��Ӈ �^�5��2$tm���H44�nG��G(��xNd���xt�"�Y�:�TXKU=`2g>�@BP��� ��J���C͞��w�,nG����\삞���..�6��ʫ1�MLK��t����VI��c:T�U���y��O�[cG�R@=���%1��3�?�m���o7���[�{����o����L�I��h���i�7?�� d>qJB���*�ީ\�a���k	?�>bU��}&�M�'0�-���k3�=o Y �ږIQ[�h��q�u�2���=y"�]{.�مR���ef0�*�y���N�p$���8�3)Q���(w@�hT	 �o1�����F�6���8f��G��k���T7�8���c]Iǁ/ʾ��u�YC���+�<�7׷꣒�n�:Q2�T��7��f�����3��vË�G�pw�Y������w�W�X���<�nn	D��5��	���H;,�adN䳗��S[���1�In�RP*�l>}�<�����O���|1�����]/|��!\|��o.�|�B� �}�����ٛ�\�q���&%>�����O̹U�̢��P}4J#Hƛ�X�|H��ճ�>��6�jT��*��v��UN�6D�Ud����gZw���oD�;�ZgMY)�C��q���0"�C�\���Mя�����c�_���o�t*R����-�X�S���E$��5�ٱ ��}�˫{9MyS%��+V!rD�|�N�~��~�2'�Ȃn����b���o���m;0e�m��;�!HY��0�E�%�N�J[e�6�ٚmȞ2Q��7�dV�	k�b؅T����|+(�Ւ��+΂#�xndIk���[�6��˕�M����?��G�@�甎*��@�hD��r�R����/��ac�>W�2�i��,DfDp�߿�)���~|�&\M��)4rHl2_o�C��Ç���d�YIy
�L�[U�U*���!"�8D��9�� �#�P�@�D(=�FY/����L��9F��@����mIB��0G�P�-E�l�m��`���?~"�ʲ8+��|��5=[�]�v�&��]_��O�'h3��*�ޓ�-8���ǟk~�Pf���{����[�qr��ՀI�y�Ҵ��2�Q�����B�L-#s����u�]_��M��5�F��~��{�����[77�2�
T, �<#ϴ��̘ �	Ҙ`���.Aj>d��v_s�:Gf�_�QC2����f+�$��R~a_�!p~�m�Za�>w�H�i^N�j�am�������ֳ���0��?�:�c���eB�1��ږz�qse�-� C6o��H~M;@;�B!ci����q�o���N.���������P
�@pQ�Q[��?���d�d��;{a����:v���X}��}�uX �AV݅p�V�$����o����Ҝ�W³0O_����&�ƪ�q�M��v����pEp�\�µ��/w8?��}��"C���O�7�`tGǫ�!`Dz�0������7>��U���^�����ϪG)k��s�?Sk��4[�Z�3�XQ��G�	���� �~��lkG&*�wp��p&��D��ʉ��� 9k	�P�`V.����t���T�j�++��ؤ���������TN��rn�<}"g�=LH�B S*~����s�Āԃ�u2a��̴n�lwv7-�<���~�,c̀����C`1�z̬I�W���}QJr��j�YbDq���٩�"�p(�$��à,���,%�.B"��\Ƕ�T*������/xR/$o�h-� �l�6k�U�L��%a����P(�?;<�}������sJ���NTq^�#��9;�~�I�/Gy����3�ia�b�cyZ���0� ��9٦��;�y�.��Ԑ����	m��s`���9O��l-��Q>F%`��$d�E��!�XZF�q%���5l�Z�kAV��5oݎ��c��?ن~���4�!��=77(�SN>99���I����FJ'5���1�s�g�Y�z!a�Vâ$�f+
�C+Dj�r�0�M$��Q��6|6�Nx�Hk����3�x�)�%��T��|�u��GhO���<)��}^�t�}p$�����lؚ��_`��TzT���N��K����v������W5�k �O)��5������9/��ʬQ�b�%�d����Ap ʙ}ތ��I�ǜz���=�Ȑ;��m=/���������Wt��2l�؏@��@��U͂OV����[Q���M`;ן-^�~0�'9�L�gk�� �g�=Иd�lVДb;z�n⨋Or�1�������0�ӄ;�$��<��H��@�!M���h����c��q~6����,>� ��dr���N�D�j������c��߼{k��:�;y�+�����g��w���ek���}J���<3�l�)�l�h��Q���6�R�ZpC�$pV�Ԏ\��IP�ȷ��k	��EE��g�\�L��v�@ >�`����!%b��YM�
.��|[�-$9��?�j*����HR�f�U����a����*�~�V��w�>��x����pf�58z�H��f��{��eXڳ�M��v�;���/s�u٫�-�e�kC����f+�Wu�\+�R�-�9��.M�c�P�G�bT���s����-t�a'j���`��z��n�^W�w!�ԥ���(�H��?��ۃ/�g!��y*�9�O�Rd��u_�Ј�O]��R&�b�-']B��,Lm���T�ڴ��Z׵�;$ٹ�
 m�Y��]FD� �`i���YF�LwP� ���a�=��(�!sF��x�-ZN�8$��:RH�ZA�c����8w����m���6�mP�:��1s���У���p8��GT����m߂�c�7@]���a hA����w4�/TA@9�l6	w7.GX!�E-���4��Eӎ`�{����=�fɰ0�	e�w�k��-�O���p�8L�]��@��g�b2����ƥ�����4cO��^���E�[��w��I{��y��_��:����{t��H���mK/k{����ր�PS����@�<9p��]ŽG�I�������q�OJ��Nг�3�2-<ݒ�Ђ��R��=ǅ��܂�!�����w��BT�!+<VG�h���Z{66��:��|ӱ�]N�SK��Q���0��3���&X��tV����<�����၂̀�
�a����&x���( g�\�i�R/8P4�n��J�ќٿQ������w�k� AUR�L��\t�t;����B�*Gт� B"��ʧ	��g�^]�Û�{Q�(�{�!�ތ%���9�%�#�)g_c��-u\�K��9 ��
_��Ԃ���`���9[q%�n�R��u�I��Gz�}��T�كru�-&Tt)��*[.��;�5U��G�
�AU�pO㫹���G�l*;����>o�"�h�,���ӭOˀ� -�F�A���Ŏ�Z0�m�Y����&�T��pr{��ϼ�m�v�� R�{t�v�93Ϡ�-
l%j����9�(��jS&;�4'�w�� vq��garw��tJp��d(�,jGD����u^�z]�����!3tn�d�H��:�XQRT���	P��DX_����|n��*];V����*	x!��Ȥ�,��5V8RŤU�{$�~�7�T�0$�C�azK�X��:1?�C`�Lx@��/=�"�[z	�^�|fN��PP����f5�`[;�1[�:J�%t��!"�������u�3C�p���C圾S'�Eߊ^��G^GP��������R��Vw('��d�)3S'%+�>�-}.U���݂F���hUI@��4����2G>J���E��h	`�sx��+����O��a��16%a�v�I��e=FPa��m@B��1����_���?���7_�}8�t���A%��³���~(�"b�2<�{��������5<�0J��&oF���e$�'B?0���P�è��:?�ÿY�~�(+� e�>H�М�6Z���e�����8c%��*��1�����X4��h~�
����;�P �D�#k���4�.�a���h�I���5���������T�) �l98x���M��h-浐�To@�/�W���3w��'e�,sU��J9����L
?�^�y��M�1ڞL��|�+g�"�P��L]�����" A��������&�F�(+��!L3�K����}���$8%XA���*���
�����,*�H�v��^���)Aa- ܩ�<1���2 d(�L߿�y��sa{��9�=��*����\�4io�3Kr����U�l��&�K֡��'�V��U��MIC>9a�����'�7��J8��l\
��idqq/�C�oHn�h��j� wv���:� �P'�Xro�7�ˁ�+1���)[O�Y�-�������߆���p���M�u_4a<7��q�b�
o�݊�ns{W�u�gWr�,�ٯ䄕}����"#�((�n��￱������r��v�VՊCC�����[��9ڒX�Nu֚Y$�ZDf�M�MA��ͨ��m{d�9ec�	4��,sXΖQ�a����LR�ԅ"
0��ԛ�s�W�a��H�5�jܠؠD �N���MG�%{�������F��e��k�z��lor|x�i��H�ҢcJЖe�!�`- '���Yt��p3e����)t@�̐?9:�U[e�U�{��1�oCW�������w����f������d��� �7kwy7�ى��}��{��*ϧ�ۀ�+A�^\c�d&=a+p�s�V�b�|=�*0H��^�1�J���;d-��9;ֆ���%��E�8��˱��f��E5���V�V+�]���Q� v􍘁�:�`4��@��3=��3��	������NT&
BVK�׾ߢ f��V��j��:]�V�$��n�~:<86'��,(l��	s/�|iM�h�*K�XC�����Ջ�� Ns���hEJ�ё�/�N� ����e/�ᾃ��V'"����N�P�{�����\ k쳷F�7_|)gμ+��
{��o
{��N�h�μ��hT�H�}e$r.�gܪ��Gș�Tޯ}�"g�ȶ��MyB�r!h]��5�z3���w������Y *�2��{�nz�Lڱ��!�et����l$�ì�P���ً�@�znb&�zo�\|�y��;s U*}�`#�Q
��}>X ��tZ�{����
qj T��V��d҈QZ�ĸ<�p*O�٬n֙��,8}n���bt�
�:�cQ8K���ňp�8�*��S~&!)ʎ��Oo^���lS�j@&��(!@Bb������E蟼�����w��6J��*�� g�1�A�]w7�#S-w3KΜЈg����]��_iD)�PڜQM��|%�_��뫫��7߄��ONpO�FHG�4�(0�0���=��pWH?2����2���Dk4�D��Đ���^�;J�<JT�k�N,�:��)q,��5g4�yXu\��Q�JY�/�RFP"j�6Y��s��d؝|�q%'��e�&�m1����"<9~d��Fxn�mU�X#�X[:N�1p����<�3e�j��C�Cm��F{�Ik��b�ك����A�h�U4y8yd��;��h(�"��� 4C�o�Վ����m�sv�I)�\�mQ$�y�_�I��6��:�W����=��"��0��iY`���<C���ϙ�µ����pv�|��&@)mW��Q�P���ЩD�z �����c{�4�xwu���k��Ζf@�.u8��V�L*H��PQI�=W�X��,�Y"f�W�9@��Ϩ���+3ʗ��/��
�6�g[��߅7?���`�&'R	B4OkO|8h��|t�X�*����9�A�~�q����\�^�Ha���\��vm�U��{AC�؇�,XT����c5Qƒ��|Pʸ3�F5�o��h�ݸ2SUy ܊%`!Y���9H�����o��bf��8�gEi���uc��2�C��B���Dכҁ9+�����J�� W��S5�2ۗF�(��E*Y�(��΄2�p'��y��{ﶄg��� k���w��b�м��� �Oi����%�lZ7Ty.��7�P����pP�^Z���}��؟�N�l�%e�l,�;�8$/؏����}L�{�t���7x����D~"'Z��;�IO99aٹ,��&I��g��4��j�Kة͗J�1+N���).�7_�X�J��髬S����q�Q��󮩎�3%h�G�j�i�Ǿ��S-���
��]GR/-�����٣��]u,#����n��ys�=�k;���@Hxc��Zs��<r�6^��~��.@�oz7Q�W ��|�΢���gO��?|����W��Ɍ�J�|P�K�W�M�Ulc^_���Ƅ�r=`������J˝q�w	V;�p�Y�}p�0_AG�R1FjE��O,�8E�/�Ω/��ݗ"�Br��5��*��W�od�N`
1�ֆ�ٸr66���v���ak{W�f����\�x��jW�a�kw �|dMەm
��u���MuM]�Qz�E'�$�f�>�?|��q�*��v1BdB�#����ml����4�@�Y�Җ�1ݝ_��3�0��a�.)�]K��l��/�f��X�
�x*6�|�{���BP��`�"(���vM^Nk�E,�E��g���+	���?{&cĳ��2Ck��Y���=��k�	����JR��'*@��V!�k72��~:��á=˾�iy�s�@?���9(9�8�̣Ofw"���CBo �������0fw��c�� �۠�a���tl�ON70"����1
R|bܬ���:'R���N��dU(|NY%��eL���4d�Ih�^с�������̃�%��ʃ;pF Xt�o��hQ߼~N�N�M��xq��*�޴�8�������p\M�h�Js��]�mjq~Ȃ��i���_��p��7ډv��uJ8�1��~�v�ˢk���Z^�i�>oK[袶@�Z(�&����>�k�����oOO��ݲ{��;~��K��'��*��˱.�'�&H�2���!��[�G�t�)^�W�,���_����zzʷ��}?'1;e���R~��^;aNr��~غDơ�`�o)�-�����#��
���&�l&�K]m���_�Ĺ�Ut��x&�j.[�(^I��	��aZ�=����Bt��:��e�j n*�hY>���N���8����ӕ�3{���X~E��vؔVϲn���U�WQ�I Ⱥq�e`�2aP�����"�����l��:� �0�;vÿ��U���Ke"#�� "XP.*�����(�H��p�\o[��g���2Rao:5��	�y����X�1d��M�#���%�W���R��qʔ�Ч��7^���
N��l�r1c��FUk���/ʃ8g@�%�IBd��ix���E�R�_iOrg-�h*%�"ғ�Ws��X�e��6�h�&:]w��(՗��
�x�)B����-�lEŦ�yb"��z�>��!���2���.��7/�V�Xâwz�.��\+����HsJ����f嵕Cln�(��S��@��e7x��qx{y���u�^���؉/����n4��N8ʻ;�5�Ƞ�Q�y)���_�s3��m
���	��H|��gN�����qas�������@ws�8[�L��Vш��6څ�5���
Ǟo��.(.�1G���`g[�6�H$A�ۀ�L�"}e���F��bEk��������4��ԋ�J�x�q����d����z����;�̸��V�����d�N�f0��kGߑ�E-9��m*?ϟG��:܌�"��q�Z�zO�y����m'�~���K-�����s�	!��J�7�����4-a��w\*8�}�:�ť�N�1be�<k{�O�OP������$�����V�Wbf�[x/������n����#cvt�3 /1�Q{m��G�D
\�e�I8�`���_pL��p�����Y�ź�&�B�I��{�Nc���?PFzȈ�v�@��	Х�eQ�5���Y*���k�5�ߎz�I"I���4�$#X�,�NU�Z�s\a��W#p����ni'Q�A�-%C�v�G���Boo+d�o���KXP�-ll���G}��l�
�w��7abY���,�-������p��>y�;>��34�T�M�а<�Z_~�Exn�ik�)�+F(�=z���Ȝ.� ��Yj�F)��VS��g�/ڳǏդ �1�:�6\Ӄ������ח�=��MD�lTлW]��%qo�H�qЩ�7�C��R���e���p�5Yd���N����_��F�+�<U�B���簽|�E��o�.|��KGc��h	⮎;RO:>�L	O��+��;��x�3
A�P�"D(��I�X���c�8�&DRMGҋax���r9�U��T���b��h�{e����$#�� ��|�3��-Zo��ڃnµ9��}��0�3�@6��ށ��
��E($+zƛ�{��<�o  ��IDAT�(v#`�ӧ�f������CY����Ks�R�M��Ђ�����l�m��U��S���婮���s�6��Ȝ"�S��߼7��� @����������'�~��=�x�/T4u�ц�F=�<64�a�#`�v��ɽ�����FɈ,�)�<��{��H� 8dl���2�s���`;1�o������ܿ�0���i��eg��`k(v���J�<�9eƆ��-U��@Z[�OT]�M5��R#e���Щ/�K�-_�@�����ǪUǞ}%���ǌt���E�=�Ri�Fn
WJ��p�+Q���j
�Ӱ�	DS;jZㆪ�^�b�rE2�� _!�2Z7�N?	��T��r�,܎�Q.�P]��5�1K�� �ru��$5���Iʪ�*?��}��^�W��v��!��#��g��������}8����b��a�f-y�L7����^t�a�,�v��F�E�mX�`H(s��e�8���s	@��U��]AM��s���a����N-�gcw��Q��h���̸��m��z�tE��e�������+������ך�f�2��҈J��^jU4�B��"��S;4���|�g�{�-�]ޘ�=��W�!�[��b]���" 77�q�X���5���1Gy`��\�Y?J��W/^�ϗ�{q�>��|�,��a�)|��1{�ӏa����=˾�'�.!@ m��w��z��P�����`M�]��=8�<�p�T�<3����[�|g�q�5��v���:ux�m���Sӏkҡ+�T�q�n�@(�g����cը�[��o�(�(�!3��}/��bP��6,�Y:S*&�M���X$>U��`5荆�^�|�?�-���@I��^Hh�Y��2h`W�y�Ne�H�'�-[?`i�m[�AK}��Ζ=�+E����Q���کo8/][��M)��@�ೊ�YXdS�$�t�<{�@��ZV���o���[�֒uxb����WrT3��E�J�B�������ߩ_ة�DfB�B���4����q�7 �,j'�`_V������d��aW}�C��F;a�����e��/G�� U�}VM�����%;g⹚s���0_�����
�p	�8_���n����Sg��Y�c��s_�YA0��7c��0��Cm��^�4u��k�DI<7NP�.о;���?��)|��f�K�GgEG����N���7��ܱl�e�+X�86	p��I��x��k��`J|�gR}k�I�r����C 4�l�s姖�+�K�	8�Rkm�I9�%����Z��l��#�B�;]�	%�PP��ߑ�c@8��2�{*��NUv�S�
�b�n���?}:���5�mϒ]�C\�,�j&���=�۪4ҙ���,��׌Y��]��>I���6�[�r�Vo�=Uq��6ռ<�CG'�f�����%�_�����x	V�N�2:o�����ɀ�UݸvF)wF����;j!��5���;���(� �x�F������/���m3������F����*3�������1�����2_*�&k�gQ�8s�-��M�5)�Lٌ���`5!�K�D���OO��>�o���2I�aw��B���Ň����[r��f����۷za�P}�Ϟ���N��\�q'����F��ϔE����o�����5�*~�#�4�CL��y��A�5�L*�z�=�|�D� �o�D���� ��.3x�c�lrg]�c��ch�^o-���E�D�P���N6�9.,Ym6��ү�8�kd�l�(�D�(�7@&�wmc���D���û01g@agW-�k�.fk�A���sAo�c��8>�];%B�j��Ԙ\���^]]�Z@�`@""��n�-�Vk��Zyd�rcw�.�@í���-�[!Թ�
"�F��d���W����6{[}��G�j˒0� x�`$����ţ'�l�=q�w�}/o�$DrԦ]'�'׶ޢC�<��͉`�g��ak�7�9�=�5@�#��r-^����\kL�9h�W�������:�l��)����]��a����%c�`O��Z� �#�7��B�ӻJ���]߾��]\�[Jh�)�hĳćg]gWҨ
���D9ҽ���ٵ��Gf?7���
UI�|�,Ļ.�����K���i��TfΣcDJd~�XC��Ț�!Of���8���m1/_�k�e��8C�]ab@��Z�rx�o깦��,w�]G�S~����T������PW�ZF (��i�g~F�r�9���\텏���X��ɒFN�--����pY���Vp��i���,��@�d\�3^%Nк��q��V���#~�S�~����N��ƥ��[_�"9���ƞ�g6���4ʊq��s�yU� ��χ���ܰ�����J$-�ZZ�� �o9@�%\	���d*���~�����i��0�Y3�DE�������g����efn�Pg���a���f�CӦ̚�����<���䏽ai�����Xv��B{���� �<��ž%�E3C������	�=Ԃh�]\<����2�?�����R+y�,��?)#����}{������+�i�Ҧ�}��I
*8zM�36N&�e)2?��8O�������o������9	����d�,���1.���� �,���U�N���,j�E�z�ZC֝L/���(�Q��{V�����i	d� �w������+!��=W6��eޔ*{Q.��u�{��jp��k����#Rvmo��q}}kF?
�gIZ�A)��M�/� ����W"z����������"��Y���d���1�8�3��k�ﮮ���NƓ�$%��R$Hz���R�{V� ��8=ۇ�.����|��q}�����?���@���}쨺��ڞ���-{o�ڷ�"Z�C_T>w�����{ug�`?��I������.�;�.�(�ۿ�s4���J��>��d�H�wI�]D��}���b�<܀����3+u,��{l����Z���Y���y��斪�HP�	�؂@���.d/�D�S���ʇ��d�����"������b1�H���ek���s:_��ܥ�V+x������!�`�k�ݖ+�)���6���y�Mp�{Ԛ����˯�9�3�B�[q��}ć=\�S]%�Ѧ^W�Tyućh�{F�_8j��L�ĽL �R�拳Xr���> `i3��\F	安?�]ơ.�np�W�g!�pe��0��'�LrҺϪZ�~r�8�N#��+��,]���m09z���S��Jrİ�Q��$�s�~o��~vley���x�H�}WD�Mˢ���D�����Xݤ�hM�U4\$!��D������'�\��*2Y�}vyN�iA����'5��^;1���2�T��![F�]fao�c�1��ŕ�נ��R���"׹#�7\������y��C�>�[����c�J�]�k@y6$+3H3���=T5�Xl���"n�1���>�^K��>3G5�������W)��|�#w�f�w��������,*�M�l��6�<�������=��s�*��xV�U�>+M�L)�qȘ��-��v�s��(/��\ň��cc�9~�@-3�gr�zh����GSpP��ڣim�{�J�	��/T��hٖ�v�r��%�XҞN��P�0e��hE�|����2R�J�PF�����s���+��d�2]k8u�K� ՠ��tu!'�9����2����ެ�����eؤ$
�a �D��\������	���}���;ͅ����27gy�l����G�a߲TD
z�2{��A�Df{6���a�Jں����E��� h�Ar���;{>�����l��;�)��;g}��������G�]��Ϛ"����p�D�9d*-es;;�=�鵽��LB��hm/q�=r6�.͉�B/��X�g��}8���~]�������7�!�c/3�YD�&�����3������4"����ѡ�H!p�8)���I��2������S	Jb`�r�r�f�(	�OY\��"�ɬ�����+�U(FU�dm�� �Mgpn�%�A�"$/�1ֆgAK����e���o �w	�{L%�&f��ݤvV��*�'����l[r�����Չ��i�W��j= ��u�:9�����=H��2��>�^<3�Q�,���Fwij��E���Zڋy�WubQ|0�@��d�Ί,~u�\RU%�5����_�-R�ʲ��'<���iv�ʇ�A�Kt��[���jS�!�\NE@~c�NO�%��+Fð��\�|ah�f��X�p�v{r����mZĽM�����!j����[��<hi��u\�1��7:t���h������(;I>��i��aN�"�)\��15�`>ܸ�ÞS�\QT���o*��
0i�O,�8⻛�:��E��J�A�+���.}����/2�[Gz���8@:��lpy�0��s��^��hP9rX�nx(j����;�œ��o�p�]w<|���^ht��GS���ۄv��=��D�+ߕ���}91wv�&�0	A�[��Ï�������d0!Lɛ���2z��(.�~���Xn	E�^B!�2k9�ח"I�f���v�G�lJ��;�1�Dd���I��_-�����j=RG@PZ�U�۳x}�Q�=�'L���0��?m��n�?�-f�]'����3�$�8��~����W��2��m/�,�c�*@yc��=שj��@$)R�"[%#n��gYW�ۄ�hC�2{f[�Q���f�W7���q/m��@�k�۾8:ۨ�l,����
l��_EL�g�zۮ�Ft w5����x�m&/Ȋ�+�O�E��0�2C��Ι�?D�Fs��m��do�����W���'^��b��d;[y�S�^?N��#&5zq6�c�g�\��0*�[L�_��QO��pߗ>>����,`	�5� ��{��Ը�	��˿���O0O%,���j#Vj��+�둡��'"�`R#�1;���ԉM�N��y_~o���W� (?%��	I�����H}�(?�4��h�|����<VS���@��r����P.]K�g�#�*R�ӒZ���	�{�B���W>���v���l5��:�,�+�C��v��T*n�·�T����؁�N��c�p��
���|6��^F��1��aq����WB9X��e'z��p�{=��Q�2��T4�Id�7��q�|ߎ'�?)�s$}���?���f�{�WJ���p*��|Du%j��Ћ��;c9g��pbƭ���O+F�lT��HB�6b\;�A�hӲ[�(Ďtx���m'�z��gt���µe܊��ZՑ>.�C���\�f�&
���§�'�M~�� Hw&���E�@<ϥk��8v2nT��>zr_z�Mzqs.m��捸��oc����y	���wd��gq�87KKd�P^�' �����FI�Q�R��T����u�
����C��˿(S��G�o�kسg�G�dk��CT{n����d>�P������`{���k�\^2$߹���!{��>6'
��� 1Fn�m����5Ϙ��c{��6�����d�)3�#V�e̡�IS�L�d@B���c��^�2�L�f���pz.�9ա��=v]s�p��FE	2�ʜ+m����������csTm�/-���΅N�1�Ǚ�Ʃ%o�+af7�a>*آw��S}�o�F�RE`d{�xg�iL����w~bk6[�r��'"�zΜk���~�b�QAb�=��X�7����w�Yg���>�ci<U�(��b��B�x7q�@=^7�����+��ÿ������S�h��rX$縡U��<h�"��%�G9a�N,���qw:	I3"�yU���n�$[J)���@�!�U�����6�.���Ri��'�����V�GAw1I�,%T��J��JY�c%�K���˭ց��5>!V:��<�5
4���x/	Vx�S/|l�%���BK���a��V*K��-,*��7���2'�~y�`��>\I�5��-b�����g����e��ή�����'�
�K_dFU`o:z�D��<"�Xt�sfN�l��/���Y���j ^D��/q,�Y���J=(�L��vS�A�/�˗����]��GGf��Yr���)_ W6�O9|���ui��}v�������u4.�����2R�qH��u�	6�ٶ�#����P���(9��,E�I�(����ۚ�ؚ��|6��,]c'3H�l���AH��v�d�ȁ��{R���������|R0����ǆ��|��w���e�P�����&�����!`�"��*�j)!�TQ�U��c�h�_�^Je�ׯ߆���{�G�D�pO���_��gn����]���T�� %���)h��)�*�!�)-΀O!@���ii�]gt"2�	
N(��Uz?��q:UovgAX�.�-\��H�MƗ,jo/��o#e�ʁXS:Z����c�5�a)1η9a�c��$��L�%\��۔�ww$ Y����UTr���	#j=��oޅ����Gǚo��}���v|&Nxn�E���jO2M=\���� �8�������|�%�1��H���� ���=�3�-����z�E,������0��ɆHy�y��3�]kGT�G���/��G[�a@�B��#�s+�U����8&�D:1s��X�4�*����>@��ףp��0]������6�$�dG:IA�а���Ŷ��Ź��~��Aꗦ>,U9��V�׮{�1�m's�l��X�̦o��=k�8Q:o��	�l]"�{G�u~&���cŖ+��|-�?����1 HR���4ݐy���O�TD[ ���uӛ�g�>8wgӱD� �(tR^�Ҕ��s.H]�=�ħ��+��f���z�v��ob�� ��z���|%��]�0G�؀��yx6���V*�,�z}�����a4'W���	���܅זq�f���O�E�������w���BC�0�W0VI1�l��[d�0*�O§<���W�^*�x�|���G22����o0\Q��O� ��)�3͖ڐ����|���p�d�E�I��+�����^��P��x�J���mS&���,��̽?���	8x�="¯ȟ^R�,��`����}���%�ƷB,S"��f�®���L<��)�u2r� ]�(����#�����kE���m���اi|d��� @�!���p�d#\�0�u���C��Y��֒�QfP-e�0Z�v_7Z��YA�� p(Ia@)��3v��Z��m�thA%D��dm��aRc���-����N��NeW�@�ܞ��"��ߴk�2#haƁ1x�۬�T� �)1J��	4�F�0�+���9����s�XP�Ѿ���/>�<"�T�$�����c�Z@�т����V�-͹V��-�����p||�j���5�4�o�{�ioAk��JU����)e�U��	Fn�%�z ��C�,�C��L��!�R�H�0�!���4J8�:P9v�av#N9s#�� 1��lA�L}�I���D%�T�b?`�^WA�Z��y0�VM�c�.�w쁖U�D.�aW�@D	P
��{,b�r���4�G?�N2_����^
�@�lbEV��lz�q�{M�`�a�q��;8I�(u_�-	����u����2�_���ys��o��*2�i|��ɒ8{|-9�hk�)	p ��S�g��&���3�4�Zڽ������K͚�e��t�^���������mV���h��4������9�&d"��EbBvƟ�Q�.F8�户�����w�z==H�>WeWd
�OCnNU|�D{���@��20��r�wʩ'N���o��h��1��k�vɩ��|]3���L�V� 9e$�0N�|�o�1�/�l�7"�6�!	�7�^�sg�b|)2�ןޅ�(��[��lmi��*g֓ٺ�A�	����<�4)�7����O-p�_aM��,����O��O���b���k��z�s�*pN�q�,c��5x��Y8<z���^J��gO�
�va����T��ܣn=㾓�t �hwEG�zNlsCF�(=T�B�hM��v�du���F��\1eQ٥v�k��ӈ��������X�y��Č�`M�G�6�-#M��{��9A����������-�ߌU7i#��9�J�JzKw�U�[��PQ7}�[x�7������X��������:4��Js��H�}����S�0-xB7�[2,�j1�z��H�;s��JD���f��I^bq���2d(���uDE��gbh{��i8~���F��7��}89��������u�n�5�K;���BT��}��2\$���ե��Ee�!Է�}̬kњ������}���T�鳳�v��F�#G#\�ev,����K	+�pz&�oH
����MT@�+e��$�L���{�Y`Gb)s��ﻊ3Lh�����tmW��5N'�yc����v�������.4�a� v�}��~��䄖���S�UҔMKA͜63̙g��d�-�V�] A �XE1����C��O�h�9[�5�N��N����	(VĲ8�;v���զ����_�ѻ�eӧq�#�Z���X��^�z�FB�@!.�I�-��QA!X��iU%'L���hpR^�}�ڱ�y-��4��
��M�A�C@���;y���	W���x�^\kT��#�R}_�N���'S���m�_���z2�塓v�RE"�vd�L=�q>#�1��\n0��|�c�lBnn��d��X��QcO3B�!>1ci�D��ƳjT{(�}�����D"?ڰ<��g�����L��h���9��2��|6����>�"'�>��������Q%+I����Y�<"43�<%8a~a󎲶eg7��һ�gf���Q@�|��`�u�ahYwF��v8�I%Z"���Q��+��gq�ϕ}{oӳJ�W_}����޳L��؁9��Z�=��L?H��؂/��*sԥ4�#�/i1������I�E� �kVx����س�D���[�z����P��������Of���eF��"
����`����e��_~��0,�/�h�55}��cV��h~�t�R�H�ٛWEZFy5�wƌ�3F��p��{/3BEO��]>�6��(m'�߷��I#���|aʂeiᆞLd9�(0�Y�E�:����WfA�j�=�z����ty��6���p� P"��Ui̽��	n��U��	a�������	������Jͫ3G̗(`�s�;���7uC�c��y��@u/����BGv�ע�pe����6U�!ڳu� 2���qbO6Ӟ�r�!Y��g���R�E�
M�\W���X��>e�71��������l�<�1UM@1�3�(Gx%�����(b�N��y, ���c� �U����	X]��f��]}W;�8�'/�[�i�����@$m�4�(�	�b�_��B�!μ�ىҧаOFQ�[v,�`��\��;�3|>�����W0q|<7�;���u$A��>8V��({%`n�/�b���l�c���l�;T�����TD�I���%'���C3�߱}�;�, ��hB�'N��uG$b��oM����Ty+����K��/SQ��z�b�(D7N�}��aA/��txa_����)���N61���qH�At�)"�O�]z�6��� ��3���?>V�}�t��2�`�,��q�)ѳ�&Y89;-�}��T�e�T�I��=�#���e�C˔(����)/]��nA�����$�f����e������k�>YH�M�8c\lA��&DpV�F5���r�S"g���e����R��%�N;t8d֗�R�m;H���� В�KKu���0W�T�[k�c�7�b�]��dA�^ڣ62�ڎ���^����8�=��p��$�u�s�?�v��<�(�Hi*�l�f�	dw���.�Sn��^�zA�C,�����'��B D�9��՚h����.�����g�g�E��ǛI��q���:W�Js��p�"��tڵ;�5q�q� ���T�aӲC��-��N�hW<��H�EjPq�R}�����d�I�����#�[����ۧ{��xe�_Z��k�P_�����O��\���Cx#j�I��D�kYi�{'�-"�H���e�m��.�L���=U�^>{!^wph�~��p��c�j.�z� �S��N6���ke� ��],5�v����l�f��kZL8�i�|��^붉e�7X	�T�9�az��%�g��7�u
ԕ�8�߆�Yʀ��$��7��0�ߧ=CŌ��B��>_]d�1�|ȯ�����E$�q��ή]Ȁ�J/֖��M�XCZ �"������3'����a3՞!(Ej��a-	e�#U0=pF�6̆i#�)�'��H �3�ݐ=��0Δw��U���D5��C���Py  �,ͣ=�k��-k��;�ɩD����`{�k!�`Y�9�#�u�T&	@���TᔵSζD��n1�?�y��X5He�4-FB�������o��EN�6�틼�JI\��"�H;	���E!@4t��7��k����;�PyP�prS6�ť� �ې��D5oߪG�� ��=�"Hx��Ge��j}��[fz�L����6#�A�^�h؝�
�<s��oz�֌�R%�3J'v�..,�U����J8�� u������Q���
'���6-C +<�@�Bߚ��%�VQ#pnS��-{%~��I�%l?���=��޳���~.0����8�B=8�ڗ���v��"F?X�,�"0�L_WN���>��A y���e���<����2�b�S��r��D�4f�3/�(-)�BP_���u;��ּ�Yt̅��V��<��̪W�	#�����Ǫ�F�(�Y屽nv}���޶"x�T�gsd�u�@ᘐl�Чϋ�|��ɢMY����:{����t�*�1�����@m)�ˀ��U�D�- V��3Ҋ���,�[���zGu:�sJg��^j�d��G����#��Q�܂�gǇR;B���& ~|�����p�R���	�z{>��NFf�a�+Š�)�nC�`k܁���L�.�����=<��l���X�0�r�B��������Sę�B����#H]�b�v�1��7��2��G��y��E��W2��wc����y�f��8�|٨�R����Ftd`Sۥ�҄�(�+������|�8����O�䛰����H�Y�Ey�>�
cP�*b�R$ۭ�Ȅ������s�9Ӆ3��v�7��QME��S��)?�~-��|�J�q^����Y��S����#ܥ��5�f�]�-�`N΂eL�W��Ӊ&q�|,��c��m��%���=�PVk6�"�%��G�ԥ�d�hONX����$]>��h�4qaP�5�gS�N @�Nx�������s�i:E|A�,kx�A����H_?g=Tp�jw;��/rnV����5�Ԙ�&���՘z��6�n�������G�'D�d�|r��II��f�ᮜ$��!��G�*3��0�p�8D+�\������U8=9xB�;��'Ї���uZ2�.{�墅e�C��_���&����4��8�d�ݖʳ���f(Q���
�4����0(��.J�W�=�fDp�t1����,܊�v�(����I+ �3z�[�m��'�ݏ�K�L���BA��n8��g~l��p d48�2���d9`�N/n����X��\ƞ?	�v�7���E�
κ��g����]�(w,����J�^�mW������=���3����L�9? ���5D��(���f}��� �$h'm�z2˫��PZ����G��Dv���������B��v/S��+�gNl�ߚ�����O͘��jdIP��;�j!鷳q��2�jC݊Z���5R[�ke�EY�l�>�dDY�1��!2u�aL���5CslQ��Ã���Ga����٩9{�g����Yt�r~�64&4�Ϸs".b�*Ę���|�@����]�f߲�.���(�]�s��gM&��."! �
 `���!��O�{P��O��I@h�Hx#�H���?��]kK���[�f�@k�[ 8��1����u1i��t|����w�2�Q��vrr�*JV]f��ʚ�_��=U��\�åo���ھ�攣��KVD=�L�z>Q�8	Q�{�k/mZ�l6�����|��1�����٩kض��@Sۃ��ۻ��ע��*�������-�B@BɃ��3��@4$��Nt�4�Q�k��`w ��Of�?�K,~1;UI�{��":R��o֣�Ǉ���P���D䈘Ded��%3ǎ �j�Y�H9I鹎�W`+[�+UrN|�+�u�th���̾�ٳ����s9O��h�^3]�2ظN���U>.j�p(8X��.�G���g�����?9a&��g&od�q��A)y���@��c��G��D4�����3y� ��޾'��R��< Y5{��N�)-����'2�VX�0-{�����*�
ܘ�_�3�x	/��o��r^�K�YZ�>S�z��ќ5v�&D����T:q8�E�K��7��~g��2!�*h�B�R�W��GG�*�K>M �J�ȇ�>u��ٸx5� ��-:�/
Y�V����V)�k��^���,x`f��T%@�͜������o�a��e�zۮ��ّ9s��g���q����9��֞�9k��h���>��H��-��Vk���E����p2�L�O�I� 6/�Q�4~��cwe�l,}v@��L����0�X������\){��$Ș�ؠ�af�*�*R��n���C�ߞ+AϹ_g'����.t����7ڋhmH`��h{�`b�����;\��3��Ým>�0c<�hI�T%��|�B�h�2#)���&\TN��(E.��F}0�3�oS�m�ed{���vxn��сD��E8��^cFg�eZp�,�,F�1�M���l��ǘt���}�v�E-�������qdY��	�	�Ul3=v�ht��,���HWwz��,@�����a��w�H�Z�R�����,�@fd�9g��@�F�swЕ�9��ڂ��򳸫�k�Iik��0`��l� }>��i)��󫧚��`��pձ5���x�C9}��1�d:��|5�k%����G�K_ctB����f�[�I��nHڰe=h�V�\�>ھ�&)��i����3K�!�������*�~W�6.A��3����.���F2�{�+���鹒u,a5��W�s���hʘy�<J�j�]��r��]G;�pS�*�?{�J�^� D<R�R	�tܐ�^��g<�g����j�b$&�:J_�����T�MUܴ�Y+t��J2����ak��X���R	SH��Y.7��Tܜݬ0w���#�$y��\�v�q� ���:p�m��1�OϲD(�ݭ~�J8+�&��+l<I6C��$�t��O_jf�')�M%Bł�-�yb̥-^���;ٱ�sѐ���շ����UyW�K�h��n�>�hf'S��G尬��pLqίZ�p;2�E|$�c����UH�Q5<9��Y2�i����-�g�re9�7/^iij�3j3�Lc6,��R�>�d�S����Ra?�=�v~�)�z�"l�m[�x�-e��;��N-�No.]h�)��_J���&����v�<89�����(�����L�`Ѷ=C@1����v��:<y*Tǂ���"�C���&��B�giS�Z%��)
��g�N�j�C���њ/�0~�M�vm.,� @��#1��7����Z�Y�ԙ}�:-�i��qߵ�Kd!頚�$�҂��a�t�R�e����!�]��:��Tge>�\E�v�x�,h�	lcmi�1-DC�b��N�>��jl;�:)���_m�� �����,D��`x�{�o����IxytN��Z)zs}>:��>��KkKDF'����	s`���#�ޒ���`�=���2��\�u�鐩"���aT: �8�쾦K��,pn\��{�p3���R��QR�"�X�Z7zMKXd�A�vx>�=isX�^�e�u� �����P�bS�&�|]��Do�B{$������/~�!��=��)�d%�|�$���nvu'g8��f��n�1�-Kۋ������"0�d��w�S��	�<g{��gΌ�$O�)Y��9ziυ.�2�~����Q8�8S�.��i�.(�[�F3�Et�����|���f�3���.�5[��o~�����K�mI��~��pCw�BQ���߄��咊��o��޽�H��t�L���ϵ̢R�/p��z̴�Y��v��|��7��Yu���u�A�5����J��|.iL���C_ų5Im�{];%Ɂ�u#a����"(M���Wd�Rx������L�-+�#�jEU��%���y�R��U3�T���&(�U��b�E�`A�KJ{7�B��S����?�cx5y�Jl���r�(���BH�bz�V�ܙа�t����?I�U{�+�cשG���*Y5mT����ښ����c��*c��Zdv��ޱ�"��V�z��v O���j�M6��/͐�їΔ�����t*|V�s�<�"�J��=[P�i��������ݍ��PGp�!3f���4�W;@f��z*��vx��O߄޿s=�N.>�t�tOU|S�Z�n�́,��o�O+դZ��4���lA��5��R���c*Na�3�ڻ�j�Z�Q2���+�u(7�9�@�
��[� QѤ�B������7�nײt8�HK|�'�{=dKi��V��$�B�g���+%�!�M�jQ��y�ud0�'��m�+�kQș�
�#K@�,`�ߑ��GD�g���|����V����(����8�E{M eOv����3` Cp�m� ~:�jhh�ꎭGa�{�����*i�f�=+�qŒ���܈�K�9�b���e��H$W��|4]�Ʀ2��d��δe� \(�=����Pω�Ln5-���@n�j�D����P��Z�G.�9D.�\O+{o��j��՝֘�Fd`��%���a�Tk�'ڸ�¡�ȹ )�%�YXs;�.-х�ݷ��J�ΡUr<�н��$��E�P"\!�[��(F��pt�v*A��:
�����$R�<�,�� ��G���9��1YzN��/�L��*�\yi{2t��0�-DCpv[C$F�'y"ϦJX	�N�`Y�x@��z�uZ`��3�����%J^h�S!��N����.`� Rȉ�JPYh���B�}~�9a7���׃'n��b�� ������g�㌘�C�D�,��3���up�D�u���޳T�l����/��U�Y�P'���m~�B�.6�"Ze��!�g��������o��g7t�C�l��I�QvԴa߼|-2=B+�����վ^� �_��1nKRAZ�4��#y{9[ʖ��d0�&`�ԏ��D�1�+�4J0И��<u1ˬ@a��$'(�j��sߞ� ����v�fRe�1ACb���@6A������.?_� ;��\Th�Q��I���e��a&��\� \oV�Sj�iT�qA�mz�������A�W��T�vK�j�A��A�A��	5`;h���`�yx���N�F(qX��PpZ�Nsӎϔ���4L|���
�f��	����B�
-�Un�qc��;:;�	��k����v���EogkWq���Q��;Zpľr>+ë���۷*�{�l�g#y$@��|�w�<}f��k�ja�P��,Y� M8�H�  ���S��u�G�j5]�k�=&�y6�@Y�2�c�~��:{���|d�o`�e�Өcf�����Zv��%��'ak��(��P�+`f�#�k�����|;$�Yf	`�(ZrWb����_)hj[��-+'���3��琟������UHW���������u�'�fF���	gA��>Cgw�GHp>˶Z� ��{�	s�J��ԑ˛��qb�x�&
E��Pр��Sw3c�W�!2*�:F"#K�n�������^��ucg4l���6L� 	@���l���O�v��J� t�HR���t��Q<	I�ۇ��;{��C̕s�v6�:��*`O���*��N�u��:�֠+� ��>vsKN���.3{�璑�z�����M+ըp`kV�9�Y�)(�g�pq�i#LW	:%,��ܻ}K��-Pc'�\�r2=;��G�����p����4{j���H���c=�(����Nض=8���j�� �+�}^�|�={�}�k���oép.󈼖 �,ko(��=��;�q_��ES�/�ކ�$%u��:'u����_?��b��3���p<��=W��3�R-��^�ϭ�dI��?��_Y�m�
�Ge�� I��l����ɓprr$> �~�B�+r)�W�錚�L<�\�*"���MWR�rK��sH�SQ�-k�;v=���ҌvZm[�`�-Z�<%HY��1C
nV�K���d���/��Y�[�TX������k�r&R�TbR�mA�ὼ�"���`g�)ITF<�p������O4�H��A�y�:=
��^�#����Gt�\��p���<<����%�e�0�M�2�����<357��D
D�
n��-B�|A��uo����_+��`U;G��r��.Њ,J�������������	�� �<"0$@$w�"{&h
�t��,¡�
_�x�u�������q�m.���pH�bv8��R�@�`ږaԙ��*
�̍�d>-J��tY�Z(�~ߪ��*&8��~[�^8�Ϸ'�H*xP�Q��vpr�wl�m�ڀ�B�*L)-Z�.�s��Xձ��Y���*��~��65ݪ�M[�[o���0�X3׵˝��w���D޵����]�g�&aN�ˮ�vl�"���vm��U�HRI�r��2��CO����g3�\ �@����c����R*��]������,���O�P#�؋��i��4(X�<O�>���N8y�TU৳S�ک�F/J;/B� Ep��ٰ ��to]33fWFq\�9/��`|�4�JR�}��²�V.�	.k��EjZ9�,�e{a!��2
�=	�B��73]�+�21��5��`��	>�db[��v�mu� �Rus.��k�ٳ�e��/.d�އ5�cgסT�v6����I����������뿩��,C�}J`p�~���
�K��oW�K[W���z���0�k��^w�g��6�ON�y�^֒:��6�l'�M'Dݐ4*��^������jҽj�e�����H���U�Z±�� �*[�9ٔ^_�|e7�f#������������`�I�\־i؜d��
jU�~���Uq8�핫ah�am��wqۮ��©=X�}�9x0�e��i�m>�0������J��%�_Z�����o��v0���*�hep1�*���Y˃���&.|N;|i���߉z���,|����y�hJ�&;?;��C�k�M��r� ��������)�.�D�Q�)"jQ�B�\n8��f��]�k<��=�B%f��^Ӟ�I�\+-WZB\�{-���l'�d�^!y9�;U�?(:����2͡ܖ.Q��,���9�y�Tk#$��"U�Qs�P�A-�'Ǉ�7�^)4kR�%����6jA �Ё�������.�beۨ���͵��5��.W t&�}L3� �}�_�5 ؞eE��t.d.�0ޛ�d\���E.)�xI=�
�қ�`ڪ��o��s��w�$�@-Î�é���LHcR�#
��%m^$j�2&aN��b�E"l����9M�*ղ�׳�s`��J�E�/�x��F��֧�m��eAjU��>\Ye9^;n�	�,>��&�:F%G�#���Wm��t��gZ`�쫐�|T3��G�Tr��nB^ՠ��V�} ��F����["�F>��c���wVY����N1�:[�]��V�6�,D7����Ȥ��n� ���Q�F���\'����k���|fφjN]8���4���V�0K_���������L�+�����ވ\h��J�EK�q�$�(�7����N����#�c���?�	� ֤O�4!�l�Y��ٍ
[��T�B\�Տ�����V��`'`��3����|�]���p۝�Ot^�1��=��>�^��~�s��I,O���g@ߔ�3��zM��~Q0lh��#�����}ˮ�R̲�o�?�)����ZM{����͍T�lʹ@_��������H�n�u���o���s���>˴JK��t� )IB�š�Ni`�B%<Y�E�`�qUS[8�%����e���m��2����-��=ǱeB��%��!0��wgCz�R���bBk�9��NB	���a;�p˿�{e��	:����â���	�g��e���V�BmYf��8WD�/m+@4����ZY�E݀
�Vl�|�W��a��#߇2E�DB��պ��X�Z�D�[1Z&��+�2I�%��Z����2�Ϥ�q�ϒ	��&��6�$�3}>���Uv|�|�cױT�[ʠ]n5j�%�������2�t�Kˠ���6�M=��X��)��f�r_�T*I�l@����:4�0^;M^���z�KlPc�:.�m��x�t'[2:��f1�X��ծdL1I�yG�����9W�Lr�Z��BK�'
Av0oZB�0�RgZI	��'H{�,��ꬎ��e��=�c���}O-c�ݬ�����M(l����]���]�S��"�Ҷ8��0kW�
ہXfbU�*�%�����A���GH"R=ʾ�]�s;�l����0���Xj���-J�^�� H�d�@�'�I��`(��y��fV5�Tc�A3v����/���
E�����0�ɇϏ�,�~O�Q:Si�H'z`a�2���{J�~h{p��M4����Z-f)��xj�N���X�1��vVT{}��4!uŵ���v�G��v�]!����Ϙ_��ѐ�HJ�HU�d�6�źV� �[�3�=L�>���	��{�w�z��T3�/s�{���t4��u�k)�\H-x�эS@\7�ItV��:$>SU�
��Sv¶ �-[���g{N`..?+Ѧ# �e��A�I��w}�e�B��2MbG3D�/<��R�9Ͳ�:���O�D~Ư�]	7��'-�M�J����.�nڵU|5�04�kGV"�O����e>�L�Ü�!ܸ''G�hz�ٯ�z����)IfC�(���/ʥ�HY�9+	��z�U]�����V�B���\(�l�Û��¿����ɳ�.I'�w�����Y�p�)�����7m�2fRh��__�{���o�t��v����A��F�
 �
����D �R����X(�R�E�.TY1C�WtP����m�݉�p�Ro1�~IJ��
��.�,r)�P�=T �j�no�Vr��-¿2��b�X�|v�"�4���;:���{��2U�z�	�b�p��%���i�h��U���ԩa��'0D)Jb�:R֒�Or�&��Q]� �w\���kw�UK�X�0�)�pT�&����
}����+��sn&�K���q-��]Ჩ���g����в$e��5�\L(QK�@9K�����C0��D4\��D!fS���7D�O �,�ܝ�*F��[j���X�ހ;�ɪ��{��[��:\�A��{���Ī���%\v�aׂ-3��3$�T�HF�J'G�2��嶺a�pg�/�R�e� Bb���Y4:���@t�K�"��+I`0ؙу�	����Hc�>q $��@L�/)����y׸k�}$���6�c�i-6�I��Ʊ(��|�ϸ�|����GJUvn�v����w5ݪ�5܊Z��C$��Ԥ*�\��G�O��Cw�X��T|��w�I�!�e4��=��r��'m���:�tq ˲J�$&�ݮ�r�$���Aa��O�4q[C�ڍ$8O���W_Y���d���!tÙP�SL�������l�{�-�N?]���g�c@_��|x�V�Bk;�^�h�ʖ�ל}3B+я�8|��>}<M��?n��x�G#���l�Εբ5�g`���a[ϩw��,�+�9�_/��s�Ҳ��Û�+W�ܹ�<���{TB��������'G{a���M/���i�4�+�A��B�{
0"���eIT���͟��\���E�P⒝�^�%�s�R���*������uOL\k�*�í�x�@ �(d�����\����/�B-t��b���n�9-��ӕ&���K�pD'�R�)�&:�@���i'�d�g�o~�k�<�j͊�"�@��"9hY�+5ӈ�ڟ���Z�qa��sv�Ҍ�D�Z�DN��,���,FZ��O�t@�w�ނK�`�77W���:,�<wr��9/>�Pܖ2P-`Dd����ծ���������KP	���W%y�4+�@�-T����2��l�T�M��h��3J�6���FN�C����L*1�9�>���+Y�*�_3y��)3����m��Y5���\��D�h��7R�JK�Y7	f��Ү�+mM��h�-Y�ߊ��^��Z�tX���dR~�z�}�����;{ngP>�A7��uiIO:	�5(���k���X���ڲ�y��ŠM;�
��Q���V�"���gn��s,���:��Z��D`I�Z�
>�!�|  �N��̡�;���_������?C�Q2L�&�.1�slTIz�����b-�6,
��U.���FҪ�%*c���V�@�p;�&���/:JT�7w#u�&h�[0�6߻�M;� PC�iT�d�h��>�`�svt@��ψ�1
�om�;�X{G��*<{mL��qC�὘�f�FP���Z�k��@�A��,�g��J�_���P(�*��y��߷s��2}���U@�ىz�ͬ���<�+�F�p��s���3]�or:pT��_2�!�Z�~f�Z��fI�Q�T����V��ʎ�	�g���F��T�4��q\����zP̈́Y��EɂW�F�Is!:��#���n=�dZP+��������Ӆ~����pa#��\ }��Ү*M�2N rF�ޗ�/��~�
��qS�*d�J��۩�d��fɴ~o��͋��ѓ0�)e[>�<0h��S/�Ga�U�{�;NXeݱ�����2�c�9����̖����eJA�	��2� �R�j)���U��~@�xY؝V���Ơ�|I|�hZ/^	#�Њϣ� �Y�p�oF��� ��OE7x?�u�.?[0����v/�PD��ZA�q�ʥH��3JrOl���4؁�؄��oe��Xղ�ӡR��Q�ǌ�%<��q���CEϪ�7h9j��1P�~M\�����(� ����T� U(Jkt_ �(�Ϻ��3�B���L�(�+����`���v��IH���P��4z���
�&s�xݨ�U�f�q碌��E��+&�H R]r���k���ځ] Y)��4\���ե�ѳ5�ϩ��Nͯ�����`Uh���8���Ԫ�"&"��ŵ�OՂ�6���X(*����|��z)f#�N��m����{r��Cow[.Jl�uE��Ee�똤��;�����m_��J4���sYD����!��$5h�#��rz�\���3;���D���:����7v�#{���$�����,�s��U�5mp�%��ۚ��~_b�H�5^wt�$
kW�#��-�@vO��f�w*����e��o�c�9Z�e^;�@V�Y^�q˞���X�$��k�c"��r6S����ý�ؒ8����ؤq8���e�$]i��&)�=b	l���	�x�a�d�S�]fq�Hf�Ɗ��������;(���3�ռh��v���dÌ�#O��~T!��	֍?���ˣ&yZe�_H��=-�b���P�m�.���Ȇlok�~�ۿQ%�	�������͑t���%&	�����n��o0�([X��J���	���|fE���#�Ptd������]��pG@��	�s�`�{��F%-eg�fa�r1
34��-��E��5Tf^d�H���^X�v���[Y�t[.�A�E������b`�U'� �Q�S����a�8X�i��ZVЉ��M�&�/�_��Q��)W�%u����}��/j��j�����Yx�x.��7wd�5����Wz�.8���V�h5(혊N��ع�Ӊx�M^E�t0���,*�r�)����y2�r(�Y����M�?���&�q�
?s��r�1��4Q�WT��[�� �k�j'�i�M><�U�k\'z� 	1��-�l5���k/�NB�=����K�Jm�9(���8��g�뇳խ 6����
v A�B��n�4��p �l_Z�v�<�P`��v��--�k�[p�[�9�.Z�h�T��,q�Y��ͽr�G�v�����.t��f.L�+���Ba�~�m��( ��ݳD]x�6��8�!�����Ց�z���������(���ݝ����<�����g�l3U�E�N��*kq�[ҭ�m�o�%��h,]�/��R�QZ ��`��p�S=�m��.���w�S��m��#ǝ��\��Y���I�dw���fwg7�X ��.�~t��p=��� �x`�!�m�.*�&��"˾�����4��s)�V���JgF�!�G#98�D��?�d��l[�$&�����m�N������l��8F-�;�"����� �M{ V먡Ѝ�H�F����
�T8`9KF:Y���5�~��4�����s$ɼ;�s�|!䒆����"� -<G��{�����\ER֏.����c��)3]Y����VORm��Ƃ�|���zM(�|6H��V{�Q����ě�������=q��r���p����8�	Uxz�l�����"���;�l�� ����8�f�ɑC6�?��.|�(�G8@����^wv�nض�{�u�����'Yձ���J�tt?��x��;Ӊ��2ix��yc{.hǽ<�Z�Z '!��aLe��w�Hc�T_̿�S���63���\#$e%��!��שF��QHms//�, �v �<�d9s�<y:W�vz@c���v�2�Z�lPF�B�	�i8^�7� ��K���#� fg�Ӊx��E����=���mL6�R׶r��nOA�d�k��t� /��ݍ�&�v\�U;�P�<mh��Yn� ���Ul �d��X����o��W~��3���~*2�6�%��>"`�T��+�$p��Ė�_�{N �]|�։� :.HK:��$�=���H�䑴��l�$�0 0�O*���~�8[���yD�O�| Z�0[�D��5����h����?�c:��=� �U��U���W����Q�1*�d�.� T�e<3�q�jvW�t�$�<����ݽ�b�bt�&��E��P��Yy+�� ^��$�=	-[t��1�[�ugk���s�?�5:�}6I��kd��QV�_n:T:��/$���3&�+�u��E��Q��#1G ��m�Ҧf}��.�=ܩz����h��?R����0�}P�vtOd"A۸\�z^&-G�3걯{�7_}��Ei��e��0kE�F"�eߛƾ!{� ���:�ڽ�O�%ؖ nn%Jұ}O�EiK�=]�2���2x��%�{n�9���<��>�J ɱw - [�%0\�d�($s�nAi�?�5�7Y�$1H��ȭ���]Z�h������72솿����	�y�={���q���w��- �@ ��Bd���HJ0d�F����)E���{OᚲX�-< Ӧ& �(��(��H��l��V���_O)i�QJY�W����3̭����_��͛p����ٺ��
��X$��iю���Wj׬w��k���a8����%�:�ZF�/5��C0_�B~���ւ�fvR�F����>if��)/c�Ʉ���^"ص�Dϼ��KI��Փ����������
�H���;���E>���m��q�a�
?���(вۘ� ��ɛw1U�H.#�S���t�+}��bk���g��3U���%^�H7:��BtW� �/T\k[sX9�u!��o��o¯��a�n�pS+K�j�IëՁ"I�m�`
��T�y�I��taz�j�A)��9e���	/��e�[o,:��HoH3��"��
���8��QjQ'{��w<��k��K�s�2Q���C��BO�QQ�h��������Sun����  ���H��ɡ��S�-��P�p�˕���3�[�����:�=��
nc��.$R�k�g][�p�z�{��O����Q��>D����$I#:=�z+�k�1� �.��C��L�V�O.�V;��a�3P��L���7��$ni�_-Ƿ� �����Z{ z�̆9(6dC7 �?�Z�$���̤u3��޴�zҕ�>&Y?�8��1v�[��:�w��{)�U��-�B.S�R��,����DzI�+u]��^z'�5��lB��+�݀�tD�./��M��]��oFu���2��
<�P���F��>�D��$�6��y������p��'V�$�hX7nl|n�XWH��.��/H+/��	�}�%��7�F�C������j�ˍ&t�n䎿DE�k3/&������XR�?^L���"�9������7\Mڐ���jv�*���������$*���<3���T���r P흜H��iV(g�I-U*�?��&Ӆ`�۱��id�}m������즚��_# Ӂ'�Tcpn�=�������b)���}�'��������$<�9�����ܓ��?^ڡ���"���>ugs�j��������Vao-cA���d�l�`V�gcv� B�r�O�eI�R�݁�ʫdC�w�����B!�LCmLة:��q���iGц����F-�+�= M7zr~��VS�U��E�|,��4qj�Z��#�jЬ�6�x�"���֏\�F�5��R&���\m8i��Zvx�����wk�'Y>���Й���}���5c��c��2lF�w�i��vv�?���K�����ۈ�	$����
ĦUqp�q�:�<��%o�7�]��to{���GZG�� G�hfν.�'���ԓ�v��n��:޶ 2mw�cg��x՚9ZU�N5�f�[���R&����m�0����A�σ��"�.�|�M�t���S@p���[CKF�����H�X�P�"@2���  @e�E��}^��c�N��q�}�<������i�͜.������g���XF�S�)X'v��R����е��-۷�8�~v��v�*r0'�:1�z����m\�V�Y���g�a�ˍ&��1{���@Փ󁳸�9~��ݐ�Q%M��S��Vf���o�lr�X;w�[K轛UiĆ�B�;�vt�b�u&ҧ�G�G��4Di���:�N�v�v{�з�-�0Ѻ�Ol?]�H�R<f�o0��w���c>�����8���C8��vk禨RY�erOi���k4�Q[�(�x�#C�~�ٙp7���}��<b�� z*.�-��\wm-��&'¨x2sG{��9p�?�OK��N�_~��J�V����p�guc��\��@�����L���Y���_i�thA	� ��ZB�k��CHΙ��xza7�n�rV}m���,�8-�_}������]�T��h�����AS�\\^�?����_���pwu�Co��5�& 5�8��Ç���7����n(�����M(Kͱ{�*��ZB2���Q���߄��'��w-�TvP��� - �ɤ���#K"�'y�����������������o��+A�*h�� � N�� ����u��ҭ��r**���&�����j��,���t[��Z�� 'Jk��8�2b�PON��7�E�pc�� u���: Xs܄��w�5;S�jj�
A�%������*4z�Y�i�D�}�R��X ]�J��#thI���\B@=�}�����ݭ=;�ÛɁ(�=!)��GG����\�Q��s�+ſ���L�=�,ZoC�*���+�|��\��/�F/�K�?3_H��p�1OU��'��4�*�&��Ƈv@�(f͑m����?8�[�s$�TK������XI)3�F���j]yDy��7�^�g#K |~^F�f��ݠ�ݩL�-ͬ����]5�Ċ���9�|k��D����栴���7�'�a��Ӱ��$�,a�`D�	g[T�O+W�kp!�;�Y+��EN��|&����Ju8�t>���c˘��N��?��bh�R�r���ħ��\��K)߭�61m�)}�� ף��k�o�3T���"@���7�W��1#v��kfommӖ�
%i\LJ����?�^�[�F�J�� ��� �#�8�`�w�62�>#��R�����V�3���D�DnF��	�}�����4|����yd���5������fT,��R���J�{v7����7��sh�PRa�{;��]��Ϟ*U1H6�x��L��>�I}��F����:�k�E�)ی�����Z�>[k�r���tߟGQ�W󥂈���H�j�lc����W��=۽���ѹ6�Z���|��h�0���B"�����.pu+��g/����oÿ���ݨ��Q7�p(Y�w���Ls�O��=�m�S�D�%��g'����E���L>�'O�Ë�t��r4�<�Gޢ��Yf�1[5}��m��p���4���Ѻ�_�H��������'����m�c%�J߮���}��w�M6�jڬd�d�t��1oYq��Ix~�4���]Q^��m|9�� LR���n<��o����Lq������ح����w��ZG������gw��d�������	���F�D�S��<!�F�%��t�Sr<��E���j�S+��;���F:=�/W�;��'��֒���1)4�H��IKZ�;���˵z�eej���a(���QEI��[���b����hE g�25�pt܃������p�G�Β����ٳJ���!��}r��WE=�k�����|Zj^�C5!H$��¤$��I��R|'KS�J�
UK�2����ZPI�Ö
8�f8���R.�V�X�'Q��]-ML(;��][Ç{�w�Ϟ( �-�U@���޺'�r�5G�
4m8㾞X#���)M�3�������{�M�U��Fr�����_i�S�Rz��k�Q���nFk�a���9Tڳ���皟�n@�����|�$u�6�SzaC�O�̺��+��J�O�hO�uGG�s�X�0 ����eQ%���c��M�FY~^0��3�"��|G�b��Ii�X�㜓W�YX��S��m��TN_�]�3?P��s0�t�X�̈:�A�>p��@��S�2��;�Ԩ݁'���JgUd���|�"�?"���u}����������֏�y�[���:��$��\2�?�,s��-+a�0ȿ�|��jv>��۶�	a{ڞ�$Y�\]��t��n��kjײ�ON4���	"�h?[d�:�|L��,U�Wu�B7F� 15GD�*����V%_k�7��U�x(j�܊vBe�Hڛ�ji�p*�m7�V-�.~}7�v�?L��=`�FU�h��!��B�s'ٶ���{�֚[���=��~��߄�����e	K��+*M����婪Ƿ�3v� d�����o���C5#�_�K{�,��YВ.���9����Xﭲ�]XE�<��\K�����\d�9v�ȯ+�9����И���jS��ti�A��>O�6Yn5	>[S/��}��]Ue�ϮUѳ�X7�G��`-(��������h!�� ��e�܆�K��(��0��-��=o�)r�t;��r�����Bԋ�s.Ւf��Z���\���m@�d��|j|�bz^V�
���U/sgw7��Y@��˻�|�*|�mU=��>V{>^��A���D!�{ۃ�i�t�����+U����*ߥ�T��W����s;�Z�;!�å�
���>���eߞ��>ײ��M(����L��Ē���V����A�[%�o�p��7{"�����j����Ҁ5,=Y !s��J[-�,�Z��^���_�������<J�֏szZ��G��|/�Zt��[�ݯ4}�l	��� ��6��y����Y@1C��\M���_��fe����LZ�X !24��I���e:��|!S N��N۴�z����f�$�lYm���:D�N��SW����"CYFi̲~��7:̲�����tB�V�=�U��VU�Do_�>�yE���7��4�ȢkEL��F?Of���c[���_Rm�i\��%���([�(~7J�`�DQQ�Y�Z�2�p�Elm�����!e�!9�P��!��N���ت_w��])��o[�I��v��<P���r�*��M�^���e��+Ѫ����U]+�.Ve�{���"q?RK�V�h�۹X{���+k|�����$�u�dIx���Y��j����܂�]w��C���aw+�8\�[��F��P���q%&Z��[[��T�U��c���5[�̃��D����+����}8{�ђ�;u��2<����|3K���k(KMK�<]���v�$(qFS2����F�����>˷������Nv���K���ʒ�����e,��~��&܀�S!�� ��	{6NEYWխ'���<*.�5M+�.Q���giv=�l%e5Z��0Y����و�Q�P����^F�@�r��.���u����A@�����X��V�%G��%�����fO|F�՚x�k���i���hm�Q_<Υբ&���R���p���G_9�[_X�ٮ�i��Pӟl���o�
�R{�2_��mک���u�qkI�U�=�l&0�q�]Mҷ�QŊ�t��Qj���z�g������k[K��'���Z�>� �}|��lo��-U���/8�����-�-v �Z�>��ܪ��A��q�@&%-O��^����,��+)N�����{x�8��V�z�lk�(	4T~�	���(&l�� K��<��ε��D��C�K�(]��[�Y�lf���U�.��{	�a�����^S���l��"U��[U��@j����πv���\�&;CKbe8Q9�E����Ԏ'<vR}?���To��S�Y�޳ts�K-L�L�E�y��2�����!G�!����C���X�ؕx��״ޅ�o�:+I��u����K]�ʿ$�ׂ%�Y��LΒV����m���G%�Pi��)�x��,����C(�5��J��U�̼������!|<��jT� \f��Љ.7�Ў`�Y)H�*-m�
�	%Ȕ�@�r|/t��ý6���tzV��-����}�#9=�8�B5i9�PC��n+\M�ʮ������ý}���!�l�.NHv��wmQ�xa��U�ĥ^��I;�f�U,���G;a���i_~�:�g'��
��`��Ֆ�τ�;��H��>�*
���A��K���a����u�R8*d#�Q5�]���*K��`����'�O�ʞ,Z�KqGqUW2�s���-�VO�B�.l�l��5����x���Or���(��AG�S?"בD`V�fm[�Qƨ�BhV�V�	���A�jcQ���m^+9 ,��`*�r�b����F`Nc�&�I�C<]��}�s�:�v�&���R�⁸�槢�b�O׆ �|):I��P����'	�	����
iSƓ<Cl+$f��a(�fJ�4VYH�b��,��w-�� ���C���e;�^gaj�;�%�@����÷;�|:s���ي& }w�����V�v��C�-*�"�i'{2נ�^��&Q�4Z�!˃�vEO�묿!����+o����%[�$���Z֏�Q<��K(�Dj�h�ps6�'	=m�>ɭf��S�b{�`�(�1[���ʞ�Q�R>ʼ������n�u�k�<���
� ���� Q���YVў�}F D=�fF9�բ� ��Љ���ֶ����C�xw�MW֢`P!~��t$�Vӹ�	Ŗ�śynQǪw]D%�J�q@��F�3{/�% +��N�FYͦ{AqՊIUy���?��;���u�Ȟ� ����(QϞ,��|�"-��|��J��ȱ�괨�_���6M*nFc�L�Gi1U>j]�U��� �m�G�U���ݏo���Z���vφJ����K�.�)�̒�����f%r@�(�*|���~�1|�|��s�3�|�1<X�t��t3���HEzs��0�\�t������]=X�9�1"�W�@&�C�f:<�؝٫��q��Z���3­0���g�������o4���DHy���j����\��Pm���B>h)ؼ~�Jg-��I�,:���g�%�\��z�箕U"d�N����QG.�LK�@i��J.���C�k�RJu,t�he➳��7���Ҍ/��e�[�ݗ�"ӲC��T�R��#�${�QZ*=��b�nt^l��>��KZJR�՗,%c�|a�,	Ӊ��;[
|�.�~�����Y����`��.�Z��	�����YqV���j��6I�8\$������>]���c�XߋAߞ�4̸�Á��q��A�ծ%�:�@w���{��6�'B���$�^��(A��뿾��|��<���#��=%�t�=I��x��յ����+K��,�r7��"�N��Ҟ��1�>���N�^"�D�]�hY���-D9,Pp�g[ �i�N�� lw�m�o�ilb�)�/x̥`�i�~V�
��3�%j�>6Z�����2��Qǣ�ƍڼȄ�1�홆�}?���N���{����lHK7ᬛΧ
r�R	L���^�����r��G �s�)KhAtuV�L�ّXt&�~��\ ���]���;4�sB����{9/���ndL�.B+]�D�\j��u��#�"bN-�Tj�=�Y�����J\�u���$���^���9-Ü����7�j�̔�áaF0�v�J&!T�2�� ��tU*b@����ZG�,27�|����Y�	�y�M�F���q�1�괤;�yص�gɽ�K5-O��+E��z�A�0a�H����qB�d1(ɒ�/���?Ἢ�����I��2���d�j�k֐�0�rQ��~��f2�J�|��,hm7��"7-�>�k�+�7� ���-��>���ޝ��|\O4v��P+ui@M#��S!u,T�:��8L�mI�1oy�vT�èt���A�k���C��:�%������X���F&���rD%�;	H����X
8�F0��H	����	��[<�-�$6�m��KkoԪ$���J�d	�$(	}��OWN�hf3+���m]S��3��f�2�r����{��g���2�]}�rR���Ԁ��xD������`�z�����Ru� \����OIMN�Lݔ����G5l6�<�����|��k�������{Q8A ��|�k�/-k^��6�4*�,�vi#���륨u��O���Ŗs���4P7�t��ء�@܂�9
���JWL�4���R��"'�)A�k�ǖ|����б�Gi�ii����~��6��`!�A����N�͉-c:�o^�����vs����(�5�;�n��6v���@(3���=`Fo�Յ�	�����$30�بJ[R�c<���n
� ��"��cq�c	6��QH��(m�7
̂��TK���u"�5����-R��5b�C��8LI՚�e�z WW��z�����k�IQ�h��m2\� M�XP�B��	��,�?�J�쑆c����y���ߘm�Jų���V9֎��@M���e{�뱡�?A!��3�E�~�
�R[<sF .[P��l�ڭ4�Ё�3�3�6�Z�[;����(p7[�?\5��#_;�T/���y���+s�>��?Z�&��.�Z���A���T���E�H�Ҩv��#�e�V�	�P��u�1$�Z���؀.�d����Xi3K�Tz�%��vt��ȉ��YvsKe�.
�0$���ʕ�ߪZ��d�r5��N�G[��w�R�`b��Ր�M۴3K�&����$P�r�_���Z-��y��:�Y����#>�V)�T�}eY��6J_Rf��̻�Rv_�ʂ3!{0h�0�Θ��N~�Âp��ŕn��MI���B#��P�t�U	EX� @�H23�yS��������Ud��\T�c�Yg'�=�>[F���m$`��VAfe�O3x~��cg���! ��
8��A&N}lP��k���1;��D�m���h"ǹU�]��Z����U��j�(��PC�S��jCO'���������=�w�VUu��o|v��(b�"~��g��U1�3�5���ϼd��^s�`�@m�������!ɵ.�@�?�����ۡ�E�����击"RxȲ1B��JQ�Q�0q*�t�����ߌ,�]U7�^?l�wMm�^Z%L�|�j��DG�N(��h�ڳ<x�4�|�wl-!�Rwyҁm���`??o��ص����⾷�s?Oõ}�k�k��V(��p��	���PG�<��Pe�۞u����B�\c�L���uL�u�	�$/�Β"�-Yd�*��P�k��(H�y���H�w�_���>~�"�_rD3?|i����
���*h�.�{�O�	�
U0����-��'�O��o^���H{�3�@3��j�'�����d�e�ӏ��}���];�%4���1�@�%V����ϟ?w^;�ί/���a�Y���=�ܲ3��i�����(�%��Q�̙��;��J�3�ɯ�,�?	���֙��"ޠ����jL��
W-�/�L��7�<� �62�?�b���F���A�>c���5��5�-{dlx1�׫��o����4bI�z�݃p�=�6n�ygQ��4bn��_?��[^	���ɍ�Z��x�A+p�̥U�T�dl�>��o��^L�^�U����߳O�a�
�e[�������@�x�*]枫�C�$S7x\op��T�djH��ձ��<%�JYT�cܸ�8�^�~!��$�|V�V�=��C��@�v-�~��qqpo ��G�n�Q����c�|���*����m�XKDdB�g�wt7
�H��[�d�I�?}��D�CZa���p�<R ��V+�>t�<�Es�ҫ�E X�$>�H)g
z��JHh+ƕ=~��TPgn�8�B�B�Ƭ���"Z�e�)���B�Y+��k �e�M"��"=d�P���k[/i��ء��ׯ�o�|ƣ�pwy��$� AZ���;��ߘ�_^\���;�R�O+�JK�ɫY��d3jQ��J%�,�\M�/�z��,�u����Á���7SeVfs��T!��}Ι�I�+X��ǃ(s�����Q�l.m���]���B�d�}n,�����9z�c�J�����.��a�#�f������$���BY+HA�*��4\��=Y���1v�v��0�vaͨe׭Be!*����_n=���Dr�]]�J��Z�i��]'��3��7����;�y� ?�R�P������[վ��"�l�����������Ƿo��ŹӺ�$[Ec���^����L�f�ؽ���|��ˮU��(�߶��b-��3t;�(,�ptx��Y"���������E�2��x����X�	��ϟ�g/���?q��\��,H���
��LP����F���4j=�gK�- ��h:߅��=%5�4Ղ��up̂Č�:T��(�p�5��Fg&��oۃ���k�Ŧ���K]n�?>J웳D���S�8���FS~��,E�w%�E� �����;�t�0cɣ5aH\}/
��&9��u0��}9�jOJ=�B<�,��P���R��4K����N�!6�h|��l^�ߪ5��ٓ�w�;}���PK���[]e�+;��P�"ia�>+w��+l�,���}r*bZ>��D�;���qcьmY�'����i��Le�� ��M����@�yG�AB�:Ȧo� �
��5��"�b���%T#��KI��D&�*t�����6/���Z���&������ai�`/��0�zYE#ri
��FK�u�"^�
(#�6UYD�.���2��W�6� ~y}�C�������:����Z:��=��� G���;���	�PI��}IY��TG�j/�*��RU���%m�Y�J@�`�l)���K>�m�<����������)V����r��u�tCW�������F�>�	��\�,x�!X�R�v/���~�'Y�]^�
�z���^��i�����]�|�I
C �� ��%@�\�����S&4�l��dA��/e+�:�4fj���$?Y�=��=[�w�v�?����@-SU���G�U�m�q'��epr:��2�X���J:R�Ҟ_�C>��Y��HŧŶ��a�-�O�5��=ה���̒�Ҿ��M�T��n���Iˑ�6\�R��UȰ��]H�CSIU�x�V���>���)VU�թk��4O\�U!V�p�m�Ҋ�����þ]�WO����S��� ��7��t�Aا�����»%`���f�Ŝ�9L�<	j�}�m����Hջ�uu�8�ɫ�\�>��={�O�+�#��:ؗ��Lj���V��'���_��_�T�
�C�YU��%DU������O��r�
�A��]�N3/�ku������z�V���HO,~�fM6I��w��r/�2*�=���4f��C����$���7A��o�>T%��]7��&� \GFH3�8�@|�iR��ݫiQ��KY�N�(��]�����Z�M'%]�R���{��i��FߓlK6u������{�f����󒝝�p��E�����^����~�] ��[y�vUQ%(�H�0�G��jj��ř{R&�.��{�¯�0?�%�Z�ˈ �#|NhF�� ���0�L���F������(F+���,`�
�Ӫ�6��<���9��y��b����M�<|ba��aߪyt֥�B<�&�<�3�1SD�������(��E�f�M�:�^=}��n�Gq���W��f�J�a��cB�D�- �b��B�����p-æB�d�V����hgف���3*,Z����9`kK��W��kq$�?=������R���Ύ֟�㑱��h�!�e����Ax��e���_Kp�.h�F��k�t;� ��L"��3Sk��:^}�}D�p���*�;[��}�hl����ɤ�Q8RYs2S[���<�ϼ=����h��V?��b*[��z6�J��Z��&����S���%K����H������QD�a�(�XBw����+�[�gV��u\2��JL���RK@B�﵀CP�ʉU2v��/�&���l~�J��h.��M����B�JD[���:J��k�3u\��J4s(�v�P��k;�T�|�-YC��`��}�'Z�������JƵ�]��=~���%�N[������������n�]�h>�$��%a��! Ȍq����ӧ���_���}�oh�$:��Τ'�+�!�*`��ϟ?��?|'Q�@�> �D��"r���"���G��w�Yb� �������[r�.2B"�+v-����_�3V��COy�}�i8P��D��_{���]y�f�yb ؛]��������-�C+�aBӊ�r�ETDk�d~�M�F��[?����
?����vY=&Hގ��zD��Ts�5�8���	�ZNi.�Bkzf�w�P-jT����W(k�.�k-�������k�ח��ga��K�嗕��g��A�c��J��1��v���p�Ï?(��û�0�*�2h�j��*��A�ǌ�I<��z�������NO/$��!�.|���ܥV#�fz��� F��;���'���t��ζ"變�l�Y7�o��C���0��CE'��X�d�9
7�� �d�U����o$�`0�@.l��j��e���ԥ��#Y�1^Zu|{/z
Vi�GG����pp�/�13$�1�Ev�.#p,�y���3��W�D{�{�&tum�!c�Ks������ˆG����1F�2�Cw�t��G��[����v5�:�xx0�;!�"Z�d��k.O��**UӅ�^��㳟ݵ
�����T�s t�D��b�E%�X o��F��OG7�>K$�0�
F���A��A'�T�A7b���D��ڛ%cT��^_���K��@�6U�x�($v��\� zhWnϧ�x��h��4�B&޲�0��5��a!�a�Ug��Vi���v����'���]���'��]����~O���,
Kۀ`↧�-�}�[�s0	X�K:�v�� ��Be�;����a��pϱ��:G��@�����ӧI�*>��T����$�UҔ��=����}�|wc	�HV��U�� �$:1Ӌ��NY�;�@?}�.ܾ;յ%��Ǜ��Q����l��]���E�������������_�:/�/¥%�nz�R���F�
��`g�量
ƬK��+�͢��Z�ȼڽ����o��J�t�Q����΁�"?=f��]x��4���*,���s���Dv�[�@{>v^�z��Z��.�Jw %��h5	7�u�*]�����~��U��5�"�Ơ�(���$c[?Γ�o���Z�X8�U�Bu���3�8��'-im����c.܏<Q�0�B�G0�񖺅�p�,�Ì	�eC�jb�ƿ���­ZZ1U���i��թ�ĮJo�+� �(�}�+��[��{���2=�_��w2 �eV'8�"T�)E�B�����B�E���
	�����>3R�c�.��#�ڑ���zT{i���	�DU�������y����doW6hg�w}g{�UT�x��J��.2�I�Hɑ�v]��C(,�8� 5�bq��.�@�߀�A�{O� �N��|���I8><����v�P�l�q�cj���A��#K��(>���3�q�����3K��Rm\�a��u�. '�*A���ж��V]ׂ��{4��q����i���a���W�r��MD�j�?[�-H9PO��NO<R�3eLD��N��������p���ݶg�Zb 1p��V���y߾O`�(��ª�{[��v��C�%r�%p3O"hˉ�.��Z"��Z�q)�m<o�����XC����@��V�M^�]�s�<��8�I� ���� �T��4��Ձ����6G�ߏ�@?�`�~�p�W�piA����y+<�zr`�Ӫ���в ��y��e�I��%Ѫ`�1��=���<������lW���ّ��n�tw/����Y�+E-h:ܛ~�6��3^�n� [��B�^Jn�tE'&*eL2P��������9!0(�)\G
��3},��o�ُ?���$���G�Q�1m��#�����8:��г����c����#��z#%?�0��uh7����E�1�:�3K�y/��.�"wv��g�4�+�����|����	�$�--]����25`��??���>>����A�ŧ��D�L���`1h�>�ĭ���z��zu��L]�F��y����"F�we�x���w��;3:ծAW�r���o����V��EU]\7�GQ'M�1��@2��9��r�iL*��"��N����;r�"����6 �����s
�v�Ө��
I���N���W��y~������j-��d����Zw�!�n���fM(9;,|[|{=TF��Εy��﫽���\*�-�T��-�X�"��x)�P��XQiv���r��ǌQ��<���di�Dhc�EQb?7���H�Ti�H;7q}�R�)�8�.�J�O3tm��1���*]�9U�}6�����me=����YY�q��ٳ�\XKһ
;{{���H	�d�~x�}x��dSfM���mc�Q�!��)|MHPTe�����,�p�j&t�U�y��ӧ:im>�ymf�fa�#�1�%��h�w�N,젴����Ϭ�������N�l�����6/����	�"�
�F�i���&��6�4�bVЭla�>�{��a]:��9���u��89���w�n�Z���Ѻ�ܳ�1����J
�Wͳ4���Y�һ���'Yl��0�Aaj��f,D[qm����������D,���K�� ��l�$+��j�Q� d���c����ϥU�s�J(Bm˥���:�ۺ<��7W7����*[��%'t���K�NÐ`��n��ګR6��^:�Z�+�����c�M��Z��К��=��nHW�ʂ0^�IZ� �Ś���G-k�T���K,�����!\��������z[�2y��v���6R�	�O����> Tunm� �hYF1��n�u���7t�琧��إ}l����U��bl�9$�v�����p}�������������b�m�um/�^~V�3�=�["�A��4|������i8����ü�ϾՓ�P�������d.��"Õ��o��$�xo�^�/uFE��JR��^&?�@j�v�U��Ei��p�ߗ�����rb���y�%�)I�p�`�ަ���cE.�Ő���� ���u�]HΓ� w��]
)�|�V�nFJv$@��<Q�un�v�TG~� \�դ�S��3	P���N;� ��g����²��Pse��!xx�vʯV�g.��؆e��"EzΛ6.\��S�x��BPe�j�C�Е��R�A!I~��I��:j����@���=���h8f�����(s�o�tH>��ʝDԧ3>�j����c�z�Z��}tJacw�!�Z ��J\����u����~?W��=nmuT!ɣ��E-���Q��*���N�V��K��r7@�ARW�`~73�2uII��<��|�����G/^��ݝЅ/i���e�U#̞��O�]�	��*FIJ���W� �ܑ���*W!jÅdё�cމ:��?�Ujbj��_�0�)�$��l~_�Tx�R��!c���$MbL�@�B/�D4:B0��J�|N�T@f�P+��+����y��_a����:�����0Bu�H�TEXr��n�������*�d_H���p*��JkV�U�?�_S��x��M����9�I\��<��{*���PX��K^��U.l¡ɾ���m�9�
������U;:�-��h�^��B��Cb�@Y:71Qe_�3]�TIWQ�ΰ�u+�GPyJ�,RS���C��pkh2�wlC��B�x(K�A#�R�5=�3t�^nՎ���hq��{�%�0�C&���~i�:�[��z��@"�~Gi�}l�2�y�uX̑�q���m�H~�Q��~��ʖ$��E)�sn	:tK���/�(/��?�>ZR!�j.���[����CK���E�~}{���ӟ�~|�>�s;���a��cNړ�1����`t� [(�(dUѯ�A�r���oΙ:�-em�H�=�7������S+i�P�C�d%u�c����M��ԡj��$Y٨7f���q���]�
��hH"?�����-������U�M�:y�w�[���F\���2�9��W����Y+9gf�X�"�#�a�o�˫�����qU����?��ْٙ���=�)��P��&y�O����z=�E�<��L�9fj��n����yΘ�����G��NѬ�� P����{����jp�������´�*,
AJ�;�H�E������k3RÈ*�95R�������j_V�Q�Ӌ>��^ p����Z�D΋>dTL"�I*	�3�*RӹȀQ�!�$�d�'�_�vU�Bd�yԒ-�aL3���![h͝�hp� @rR���]����Y*�d�P\��x��0zE���H�u=��q�@��C�FU�j��+�}��L@�n�tA��O�D�������N�3
usw�-J�`0+yd/!�?�	�d�$h�up�J�v:�xxK�e泊:zT�f�(+I:��!��������@�>�����"���X�RsNT��-�l�)��s拷�4&2-p:�.d���Z��2�2�g�P���Z��c3Ҽ�4"�S�w����5`��;ڴ=T	]�g"b�G�}���2$k�bi�7Q�V��x(�C`A�Dw�� ��}����
@�]<�{.��U�����f�N'�pck��!�ّnr�7���̥2I[^�85r}'�N�}�1����	����v���
��j 8�6g�v
����po��}Z���ҍj�����'���3iZ�y�,�ph��\�����t���Px���c��-��Թ�,  �I���"�x���,�V����7F
�ɢ��v��LH�z�jϦ#�#�T&(��"X���'�_,s9׾٧����.��Y�rgvͻ�wtv�de��^���m����
�����U��Q����%�ro�On�&PR�?�E/��uE(����2��{v�U��IG����LY�]u_Y�#�=�2�	�5{��ԞI��e���jTƱ7��f,��Y�)�6lt�%�ԏ�pk�ny*�)Y�]�q<1D�CU��ڮ�;���!�����焛fEtt)��Z�G������7a2�8�:Gvg�"�mC.3ȣ�&N���zgs��*���ĉ�_|��VW���CT����H)8H��� Z��ֈs���"���Y�`�\��T���c��!`O��K�q���蘬XΣ�hP\<��Eą#&B��G6���J��,{*��K�M�n��c7�5q	�"��Z����hI�Q*R�f��N��ƈ�k����QXf8��A����#��fS=rL%i�jN|&��e=�Hv�2*cS�����'���?ܔ�����"9F�����!��蝉O�D�Γ���}�6E��"�{���[G�A�|��%�7�^��.���/����2d&}n (�Ygh��`qf�{) ��ȼ�b�X�
�'T������Qz�K\�1�X�Έ�D�ckS��*���:A�����V���1N5^"�bq{��`�V��ݪX�Ǽ/�A���0!Yc��-�4�i�v-3{N������7�ښ%a�ӗjSi ����>�\?�G�o W�n�^p�챽�D�(�͗��^.|L�����e�8��;�L�I�2�2�J�v� �5��{xtwy.�?����d�D��M�R5d��E�^���eO[���[ˢ[�����e���Rޅ#]YUZ��{jB�:8�	pp��S���p�l��L?ڹ���C�>��%*�l5�F����)���"�2U9:�o�aTcj��������~�S���G�!��K��r&����O�jj�4�>t�g[�����������[��=�]�	PE�F��\W��j��J>s�e�s�hĚ4*��/V�_���;80TϠ.c�~rZ=g�e�`k�~*-�ռe�f�[;��sjVHG9���.d��e���e����cx2L[;�h5�9�W�J3���R�Y�*:���oćy��_?�j�%ʊֳ\��ۡY��~�Fs{@��2�}f-eX�Ј� ��*}�:j��jBO�Q���;NE��HʱZ�����ʵv�����������ə�B��c�D����4Z9 PV�٦��R�\V�M��rX��R/��
e��k�2i��$�w��'g~{k�^[:ܔ�U�	A�(��Κ��q@�K���+��U�����*�#��ĭ��NG��9�~:���Y��g�3�Z����h�`V2#�xh���6��,֣�na�V��cd߹��5(1��-]G�R����>,|��J�����^�GC����x�[#1�tk��o�����ǰ�w�> �y(���ɡRP�rc�4g+ĵ���}��"l��#������"��9q�n�*P�	�'r𑰀��gG�p`izH*H����B.�~ �DJ� ��Ssg���h��J�N�M|꩞�K_k���s�dm�n���-���҈�y$s��z`ی:#Z�Ϟ?�W�q��e���������}lk��R�4����e�渚T��$wΑl%D��$�5��o|�>�|:���*V��\��!@%ȅ��D`=Y���mX=M�<k��0_m�]�/��'�����*V�8k۠yoh E�P��׶ F�q�����Ѩ}hDTF���-�O����v�p.c�!U�����d�?�ۻ;�p�������nh��6���am]������m�IOә=��0̝uO���l�t�7h�ý�ph���ˆ�]��G2ޭ���a)��l�+Dy9���g���qƻ���z�y�%:�8.��m�.?��g��A5��"f��Q�k����j��#�խ��7�,���|�����("�z쪓����t�vA��]\����lS;�+�x�v	DG ���.3i��&���CGwV�������SlLZ��<�Xt�A�W��(=-� ��_/��xrE�Y�T54>��Fh����D�R�ꗫ���W�s,#�@�pD��&e�
Ǩ�x\g�4�"�XE�'�XӬE�o��*�.�U�ቦ�6l��s�̧�3��ABWw��/��/�7����-h�*�{Tm��jR�3c9�F�Y��ة$1�e��V�	�ں�/���
,�vc�K`��K�-Ts�|6c1�2���g��!����=$fsq��*������+mdq���;-��%���P�hX�k{�^�k�ӝ��*���RС�%9�b(�Ѓ7CE俷{�d�A)3^�,��Ob	y���}��͝Ʃv�	�lvn�cwQ��, 8֠�y�"�ϑ]㈅�s@�����]�^����}��0j=���ê� J�0�-��� Qކn�ג�-�)�����1�2����خ����~�oB�s �'�<�=�S����wS�s�v_MF�sL+l�vm�3�/�V��/zk�k���'\��� ̶l��4'��4!��G*?�D�C��J���~m���@/O>���SD�i��QvO�}KB�_�4�9��+��́�ˮ[��tq��L�5Q0K�*�]�4i�ɨL�L��g������5�*��p��"(�gZ�Xf�=���L�4�'�i��y�Ã��}�ph�@������a��ǻ�?
�L�r�� ���8h��|�	����LA����U>c{/���~�,(�l��ߧ��&�EYYE�a��3J�c)'�WZx�۟�#��	;�g#E��|� :]�-'z	`H��h�$K��8�,�m6<����v~������4b^�(�y�)�y����j�c�7�����B%h�w-"�5͈IT�{�UI͗AXv����˄;���h��"
��Te�0���4�Xy9PE�V!��(j��W�)fy�f��*�E6!�y�ڦ�T�b�7�Ϣ���Iֽ?5����4��Aeom2[x�v!>�5� E2S��x�Sh��,S�hP%���B��*j�اH&�������*p 2�E�wy�N��|>����׿��sKe��f�3�#D� QQ����A�O��pg�β9��<��^hE�gK���xB�/�g�DY�?��Pw,b7ð	ےH*X�BC��P�悹����=��`�2l4h� q�J4CB)M�J�i�#���E��"��E6-��bo�{��,tp�������q��9J�k�J�+20��m�9;���FXX �����H���a"�/߯�8�^z�Y<�����.��;�1%@[��]��M�B��¢�s��	���?M�($�.BIY0͝�#f�A�}�2��X���7�������/d�	@�)`OZF��Đ,$pz���y\�0���1���0���X0��j{�v��2f���3���a{���a80���; ���bb�R)�4��me2�S���
�N4~�
�&�ex)5"Ҷ�]	K1{���sc�14�b���'L�<\T�9*W��:0�X۵�[ӏ�� �K��&<�ii8��D �!D���3�s��\�O-��}X���e֋�+!p�QP� ����'SU�(y�'�Z�|��������cנ�	>�6"(��*h��_{;�"יY�r�x
f��n帜���899q�x�\b�r��	������^��>'��J`D���;ܢ&Y" O#n���_��Q�<_WS�	�f�h��kL��$���H���Z��ՅȆ&j^�j�vwf?�0��h{�@/u��RS9���&i��L��Ns�UYo�&֬��w�ݢ�j�-+-=�c_��.̘Me0 �OʘJ�;[1�e��������yN�`�-sG��zq��6���8)���,q���2�F��/��k �`��|���T��a�!K�������H=�`����-�'%�*��?@�-�a"�/]��:Q��gHA�6A�ڽ3o��<*
�����=����~c��]"�4���Y����"�J=wƯ'3F�?<i'�8T�m�Z���;6�
����Y[0�)m3�d]�~:B#�E��K�v]]{%T+��]> �J��g�rǘ�R-���/c�@Q���\!G���vGcY��Z�fB9l���9���(� �Pr�:z���Q <�Yp�Zl�Ä? � �m�:E���$�kWѨR�^���mM�B�q?[��Ȱ���4'�Z)0@+�U{92��`D�����k�%���x���HA;
��ӧ*�,�l��T��h�9c�@�T��� āx�@�ư�%%y�ˌ*�ջ�;�}�;[0?�°3���ۗ���gtk��N����� ���O�vl����T��2�j�W���q|��|�vOm�|��
�j �l�ޜ���߿�漘�
���ԕ��$[[�>�4�{'����ߘ��sг���Pd�kf�]"�tJS2vQ���W�x��t	BXKz��.To?G0�c붽��`���of�9��W���@t�fK���Ӊ�x~Tͤ�]Ub;9?��/���ȡ8�ϊ��b34(AK�����EhMQC_
P4%��naY{�E����+zQb���O��"3���mP� F4sUX:���u�K>>+k�Sᙱ�F�i����8�y��0-��J���V _���G[�tđ%�Wa�"b\g88�@?��٦l"��a��ѳ�Y������]�~����=��WAk�ԩ�8�6���Ls-[O٤���4�����n�o"��Y��0�v��N�]6�VƳ�c�S�>������FG�k�Z4����ߋ�R�|]ZvV�B���uxx���=��ˮ&I�;����u�9��@�H�jA{�ۖE��ڞ��P�4�1�(��?��]٦Aƍ^Y�
4o�-�����6:�'=M��@�1f����z�Q��\W���U���ξ�:��O���e89�6�ԫU�g��pn�$Q�9g3�Q}wN�1l�vD���t���#�o��
�Lw����+&r�5w{>#��(��Ԗ�Q�BC���ENR��e�M��k�ɤ��jߟ�#�1ë9��񆔗$�$k����3�$�ڻ�dڌd%�q��d[E�**�Tr�m�}�}[%���1'1^��p�(�T�
#��e��8&6�K��dQ1�yN63�2b �	n�Z�*+�B��b�G�����ҳ��.ʥ,�3�eDf�	�x����ί���� �Z��u0��TC�C�礱=��6��k& �:;HgcG�o�q%3�v�(�n�GR����We���k�&Wg�bb������!�=�zas���)���L���	3{�����dLd<��?W@rwz��}
�gW��|���]�	�5�H	��&���1Oae�ײ�6�ad�i#s��v7�R,h́�d�5(��5=h�"%�4�[>(к}�����b�yyl��Wط�~P_�=���+?��4\S:��O�L��^��
�a��lM;ɶ�����8����p��{0&[=���p�1���;�BT�ٞ�b;!��Y�&�f陃DyB������hd[b8�}H�J-��k�S݅J��`�q|p޼<{���dR��l��H�2�K�����xd��x_e��Ӫ�m3�#���ZY��8.J�RE@-UŚcZ��HU�
oP���H�\�E ����x۶�djk��i����H`���fAa
�挥���F�I���6�#���rU��&�,K�F�71pc�����ݏo5�Z.ܐ�Z����.z�"9Ə��c|��Lc/���%��g&z��I&�D�:5��po��_����$cM�3�h��I�;ْ�+W�J�<�2ѳ;��Yq0�d�d9
7@��x��ut��XF��YY7���C�����ʚ�u�~���2�Z�N)����"���9�g##u.�R}�Q�BG�A���T�^��# +�5�����ZDA�(�F��h��!=(�Ke ���/��=uD�H�^2<��i��5=�{^��ep�e�kkc�^S��NsQ���R��=�O����Ϭ�j�3�eI%g*�M�J�)���s��0��~�����?��E��ر���C�m�vvv°�u����˩�$F���O���ť��e��Kg�j5;r$����xd���y�Y�F��c�\��o���x�{s� {n�/Uڄ�ϥ؞uEʈߎ}J��^PV���]�[�"|���3�D���YЃ��i9�b�y0�z'28�����<<A��C�"8`gZt��x����k߂ ���a��Z���B�A?�.���?���R���"�i9L��9~���c�;��\ƈhYd�<1��?獩5��Q�tf/p�#{��x�0��y�A�\X�nd�Ӽ�(nKo�$�8Ώ�HNnn�c��X����.����>L���<X�S@�[�.�c��SK6f�^��L*x0�!�B��A/[��fا�70LO�/VKi���C�"m�+(�'ס���Xm*D"���%J�mm[�r,��F����]Ά����G�W_��v����qN�*]=C_W��e�AL
#�\}��)GS�Rm�\��3	g�g�+9,D�f�Is��MB������-3ޗ�-\���Qh�����"��e� ���4�t@Y�rz�-6�Z�<�s�U�T���N�����B�:�P�5�׽"6)e��%=p���+��wEWY���H`)��r7��D
!���G=p`-s�6��Z>��	3pXt�0V�Z���U9\��	�!妅�A����� �j2���g�`{�8�V�ψF�\Eۑ@�C^|&=������"^5:xj���d�璋�<��Z�#M쀏��G��xD3��'	I6�5��!�G��󀩈��=K�O�֦��D,�����K[�,� +�D0��Ec�	
2m[�'���1�|�&v/�׿�&~y�ÞZH���^!܈k凨R�֫V>�PD'����DQ=@(��m������Pҧ�빹:o�K�:��"�vҶ��/{C�}��ٓV+hH�3��r�<#̻w�¹e���Jn��������9�˿����p)��T�#�:	v�P��Eb�:�]7�ω��4i��<D"�  �N�����ێ�y�D�C��C.4��D�˖dЊ2�k���m�``�)(��]`�*E�RHz:78Ƃ�gm��*���f�g�ƨ~��H��^�u���<��nP=J Z ��)�2J�s&��]ߜ��ӏ��y�R`�cv��L�c/o���w��ɀ��Mv�e����cG:��I��W]D�,Wa��##$�:��2�S�aX�����T~�$k��!�psy�>��ҏ�}�����k%/���k�s��6J4�v��S;����R��H��a���ӕð��3i�T��i�
F��Ո$7I�/�������x���*Uk Z��v�}Wz��`s~����?}�_«��N�i��������U�$���j�1��(���H.\,xk��,���������i�\��̌؍���J�n؉tx�������'m �� ���Y�]^p���Ch݀_��E��g>� �k�D�9K�J�N*J�g˅����~nD0;r7�SC"H��z����l"��u��
9^�2`�_�g�[�7^-�ؔ@�Ρ�,�<���2���4}DMM�Q`��,�xFR���,A1��
�ک�F��x�����r��
� �G�-��5{��t�]�>Gq+zn5�nq?��3�= �6�.E�@����߇�˟�����PX�E��4s�8Q2,"*��y��0D|�f�l�׆X�-�>_Y3RA�R� �Pj��ْ3>�@���GeP;{��`�E8x��F]K����9s�����a�q�bC*D�WJ�pb�j��z	� >{L�#�1J=E3�J�x�����,�S&#�>�n�̌w @�qJ�2wސ���*�5���/D"��"�(���dq8I�zϕ�^����ӳ6=K���o�2���-Vk ΄@~�/����J����#�"s勬l�h
}T{���˼ pa�����v�Z���t�B�lWJ���f�"�h��<�X����w$�C�|�tq�����Evn �-�:�p_�,%U��;7�l��\3�ː�s_��d�30"ֵu������>\߅�|/,;����C��7�o[�-�x�3a��- ��9z(F	�X�A��`��E�Z��IC�!-2�>*�0�h�V�lp���|f�Y.�4�)k'���'���kQQPM��K�TWro1���4�g���3)p�(%J6��k�'����]���,����9�)�r���U_A��YX�pq]�� ���_Gk���D}v�g���T�̄M�헿�8<{۟8@�D_V�wJt�Z������f7�����3ǥ���3ЕNk�*�8�W�d���Y�O����:5����aQF�g�Þ3�����=��:�'���v��3O0���H����<��K�7	)�g����3p�hj$a�n���se�h�z*W�,"fޯ}])Џ���.��zoƑ�"������t�m����sl�B�I�t['z,��(ۂ�+
G�3�1�~�V9
2�E�f�aP6�Q���/����ChX6c�Y�9��ǒJ�0�RB^:2��C�|2'0qr����F�2���e���w�ӧO곡B��W��4�,�j%Ks0�Q,��@�k��#H��4�ϡ��� ���b�_�2|��������@�*�;�#3�@�1�4#R��9ꅍ~'�ۍ0�b|왷��}~S� x�Wr>QD��������'�*܉P�����*�J��CtBI��OX2x�����-��J�U����^_X`���8 }���h�lBt��~�`xpÓ=a䫺g�3h:�D��S�7�O�O�_�9Ֆ��"��|>�g�[����T!������>�5�C�Α=3�ˎ�s�m_��� ��3��X:;������T�e���ՅO3];�N޻��2��(P�{���i�x)��(4]���e�N����{A��ٜjF?�!v����V�o�����9�9�j�q0���$;eVW�|��'�s�����eoX�O5~�ĽM(�=��ʯG\DҘ�� �>cH���wF�4fH"ј�Q����x_���b�JL��YD�c'7�m'~�4��	���g�xXΈ�\#9�L@�c+*Id	����askG���i��1c�udNX���0��%��R�P��٨d��82Z9#\���R!�z��v���^o6A�O���,\[����������}y,�'Q��Y�b$l�52��++���b�����g�U5����JX�n��z��@�[����T �r�&���k4:�C"sB��R�c��+U!�
��J��u)�R\��Ahv����?'��/L�V��1��?�F�f�a#K��-�������a�^���Ww�"	����O��
.T�^��R�R�֮-Z���^%����4�K��r���T_AJ=s��#6��Kb�3�O�%�:2�1
D�4�e޿K�j�Py�&�A��0��C�r�Z����<�>��G�^JkuT���r`�����z��8|��7aW������p��D�O)�ޤ���a˂|�,p?lY&|h�igW�i>����Z����'}��Y蒍�kl��̲,�!<�#iB��DJ.�:ʌS����> �9X)�o�=nkB6��q���&AT͈zJ��L\������I�fU��mѻKP�_��&����$p#%_Z����˰�1
��������������>��iT`|� y��ۍ(6T�=Ҍ#M/�u�'Oj��z����:`��Y��6\�b1�S ʽ�h��g��-�ɖ-�2u�e&�:��" �@��U��Z U�z~_�y�b[mW9���J�]��MHj�ѵ����83co��"�����^2�VtU��8�=:�?���;9����ޔ��>
X�>�NB�r�96H8��L�dv��	�A�����]��R��i��G��o�� ��X"�8���=]?�}_��������I���XP[�T��Z��k�>�3�!Pn9-(�c�/u�V��kUz��Ȉ	�CUTA"��F.Үg`�6���Hס3j������W�]zy5��2uX\qo볼�|�^�������P~���L���k����fn���Q����!ցXmK?_���kg9���p�{�*Խx��w�qM���!E�k]�N���P����$˕���4�/�%ؤ���J؅�=�S-i ��s��MM����v`�l�M:;�W�l�Ҳ���7}�,'<X�Y�inQ��2��*�0Uk�"X|p�=44yHd�D�d[��um!�ٯ,b����KI�	�M����&2����P�A�zZ���{'~b�N*t5��E�b/͖+���Z�j��,��kh�4�I����c=������xu���+k�W}��ō���)���65�N�u`׿��ڦ�Â�IHbs�fh��_���/��0�2z��)�-Ol�r��u~��6����ɇpws�1���=]{?
��#\,\� '��_��:�I^��Ӟ>���=۞9�'t����Y�/8�����"q=�̧�$#��gM%BH�<���CP��MUV�sWo��>�K�˞����U�\���j����D��x޷�Z�:
��0�ۚ���i&N��_]˨4Ĥ��vzy��(SS�\h�p�AEE��>�䒕��a2Ot$˘qy��~������7��kl�o����آA����zŌ=4\l^s�R�I-���N���� ��N�Oy2��g�}2<��h~őn�J��lF��Zw�rA�l��H�H�2
�Q����'kP��]����2'�Et�+U�R�VsۗWW���������ك�9��ZAg�BX3���Ps�K��i;����*d$�T���P�O�5�׶;?T��n�eP\-��Y�ph;[E�_�4���K��?��?i?��q�~��:Ro�I|p�³_0*W���֬�5U�J���y�W΁�F�]�����_' ͬ�Ԫ�6�^T�#*U�	~�BV��^{����	L���(�$&0��֠�:���iW1�M���F�Q�f�W?��*��{�v}&�W+�������?\K��?��J�y�
��Y��	V겳־��R���+�����໌Lrd��:G������ �Ͱ��n82��r�������b]�Z{6���8��&�����tZ�/��#����amG�%��!���p3���{uu!������T~��qj��F��E����Y��\�O��R�V�l�Y�!\-ܸ��2�a�ʣ��b,U��{1;��2F��g��ș>B�x��b�$�sr��aѷ�^�馈:i+l"8�iJ&����ێ��h#X�{`Yߛ/���^��;��Ks�7���'Zoл��{�8��6��@Y�ut�����QT�/_�"���&���_�@��Ȯ&v@w�i7Tz9��-ϰ��lK���#ef��I �<�^��JGWe���o�����u�JS��v����A�9�U�:J�cs'?�N%#Y�0�z��m=�N�!m�F�*�l/���Qx��u����J�Q�s2#�:�q�������(I�����z^zFzH����V3�%q[�ttv�x�M�J��_�{ ��٨g �J��S�Ԝ�t�������p�8A�����,�jv�XA�1� C$���DO&a
��q:H�NH]�����e�8&���ΞEy��zΊ�uyp ��{~��!��*U��)Μ����R��'�C�����L�EŲ8�F�'/�tا�s'Q�;��g�ߍ3��:���(O��?��?�f�ɚ$��E+�1� Ҍ���ʹ���ޤK�ܴO@DT	(ٷ�v��Y��FE�ŽՎ��1_�$��\�p��i�f'��y��M���5�ă�G#4?��d
 R�g�Ҍ�,{D����|�r��2s�c��ũD����no�@���m[;�N����SH�R�\s�L	��������������n�XLqd��	Hٯ����3U��Ib�@����c�;�^j-��|a,[פ)\�9���V�w��s�g���`�P߂4�
�㔼�_�,p���C�%,IA��O��or����r�^�����v�%Ѝ�,E�:��Y!�g�i5͕�b��������d��m�<��Ϟ����$�>|�(R���yÉ!\�;U-~fbzJl�njb3<��)Rk�⑭�S x(������Hr,£O�r]�<�U�D��3F��u,�FT5YiSs��xdx���$#���[�B�U��(;/�"��,��ʉl����-���3�2��Xd΋zp���*	�$S
y�=ܐa��\�М��Ʀ��D������~��������?�	c�^(� ��û�|#Y���s{{Kkh�)z��g�@| �6�=O��t�*�e;D/Y�ud���īqXA'����DN5��D�d0Mt��1^j���pO���`E������=�X�E)�|��W�섫����ݮ�ї�٤����������m[&�H$.��P6^��.�|�H���
P����/����k%�8�
��w�w�ʯE����[*�	��9�v� �Y���i�4�&D�\�� r�mS��r�K���$I������ΔP���1�����z�3W9ѝ���H>~6f�D��"d�*ն�2�:#8{J�������í��Z@!y�*�#)����X�\�A0�--slGo�k�S��g�d9��cFY�#�� �겱�k�|>�B[B�C���~��z��k�4�����@�9#e�h��mͿ��h!
���y��hbD?S8���v���T֕j쫧�Xy��+T�x�p�p$SU���6 �_PƉ=z�hŞGfAu�9��N3r?��i[=������m6����vU�A�|nv� `��0��C��#�([s�ɹ~�m�x�-�������0��+���O
v����۔طFJ��,��^��������i���x��;��9�����w�(��bw�����q��mP��͛�����T3��Ml��}rqs���;t�N˜My�-YIZ���U��-����)}u��v����I4�r�psuI��H�߷H-�MoF�Y9JM�`���c;���b�)筄:��[�2��Yİ������~l���9��őʄI+nRP�sWu
��g��$ν�qIW1��"��¼�+ku�~y��u��PIS��!�-�?�F�qh�S�M���z�[)C��ޘ��[t~�p�,x�;��]|<�߿�l�A�{��0�-R���:����9��)����=/���,�����tB�l��AƄQ�N�+����!�/�YPb�X[[��H�}��`��8}����ж��2R(���Yќ�/��Xz��x����X�Si��?�`ri��Pℚ望�h,����
7S�lN͈�,�j*�i��s/'�I< �N�<�P��H��$(;���>�^%�W�v�|-dl�Մ&����C��y��)7��]+���ɅӮ6��!_��b"f0N�P	�C���z�֘��5ok��j�B�| �L����.��0�̸H��M��mt�׳��7����,�pR'��L��7�(=��=Yʀq�tX�*��jJ��Z��X��:��iC$�3;N08<���bI[I�@����c[����gbn+=z��~��g��,�J����r��p����h�Z�AAE���g^��E@TN�u�r9ha)	�����9� �W$��`��"��-����PvK�6��\��P܎�H��\Z Op���,�\�w�� ���A�AשX#�lH_Z��T�l���NU�T���_H'��%����N3��HPiYz))�,�z-��:=7G��y�	���R���T����U�:��:(%�����`�6� ]�s��-$�%	Z9<�Э��������m��w6� �: ��p�zt̞���ݡJyd�������kؘ�&��J�U��f��N�I�������e]���uzR1/�l��u��o�zo�v6v��!Yب�L�ҫ�c��fRY�K�����b�*��Bk�h��L���-C�W�ʈ{��[=�[����y|B�M��pA�2��j���`e��x4���g�O��D��|T�I�@D�s�!�`��z[��m�nf��*��L�!�d:��������p`���`#��?��������ʨ�㩮�22s�d��A�l�����Bxs�>��Q� PF�b�A񧳉�Kkݛ��'ο��1��'PY�nt�3[�v� id�c����ޛ���\oZ��Ybױ2#1�y/8 A}de�p��9?�.�5���Y���d mf� K-�O��^���=8�'avo�Č��,L�'E�{���p���Jj(h��$��pr�)+s�����:��-�jV������n��|n�nm����Z��8@��!�b2�Q2M���w���Z h�(��;!�Q�"+h�1��C�41#<��>-�Hӹ�\�Y$��=ht 4eu����y�"�DQ�m���.6����R�ك�!��lf��`<�w�׆�����Ƶ�R�l)�	�Q�%4@@S:�K����=3���z4<#wX���Oo0�dk�X��w��sT��#p�3n��Dc-�e�`���/Te
�kd0sٟ����W��ʂ[�� �tQư�|��t�/+G�#H=��	�}�4�=G~��XP����۹��m����Yx�ڑ	��9��6��B�2�jK�豾}U�4A`���ɇ���^�a��e��d'����:#{�����j:sF��g�$���}���5VF���]�#-�D�tw+� �1W�~����_UW�0M;r�� �1C>�>j~�
��=���-��=�:*�SUH+��M��^:Rh?��%��%�V"�^5[��n6ZSۨy��Tۇ9(�>��L���F����q�XdL���9�f˙�0�z���J�_+fd�XnW��f:���@L�������a���<|~���p��{Epp w{Ͱ	U�8�y��1�f0��ߒ��w4rR;ID"Ǎ�T�T��EcD�axaQ%���ˣC��@�T%����E���ܣ9�;;܋ʉ�)[���H7ʝQ�gSp�&�T��p��k���>ybß}�R�,�Yq�5X�?/�΅�ꫯ��|��mx�L�@�׿��p���CG�^�x:֡����i'��?�2T��mQ6�{�����{��3��/���J�l<�M���?�g=H�� � �2�`H�x����r�W)�U��R��s�k�*E'�>�}8�.s�S[��b5�{>�����pj��c����|c�؅2��R�Y�>���^;���TW�>�A�zVeG��#�֌3۬/�BPD�$?D�s��"	y�x�����,��f��ϨW7��cPUK�B��䚉�].��S�ǽ���|����&c��X��O��LÜ9k�k07ʙZi$p������@3cF���,E��PK��q������B�|�5{���wtp^ �g��Ǹ �Џ�H�������ٔ9k=��p����6}ܦ)
�U���
g�碡�jgZk���:�f]y?��L����� TI��1H6诣����ρ3��3�����p����PU���O�*ӹ�Z�L*)��i1��Q��O������k�ᛳ�hVh�5mg"���G�JC�$'K�2�\�}Q�R-�}C+��fe��l({�q.�7d ���W��!x"sN�gnn*86i��sz����.��Ȕ�53�y$��ͯ~�j�\�uo�g�`� 1�]p�c�a/�q:��s��U�__�59�1A4��	I{� �1��B��%zPvJ�������س�͆�2�4mZF��?'̗�����xAY.azdf�p���
!�x��U���a�6�؁Tn��䳢!�೭��ճ3_���J��7��5ʯf�aa޼x:K[����� _�a��;�?Y�x��鈮�bc���F`0��S�%T�-T?u��1���{_��-���C�Ć�P�,r}�(D1���b��{o;�-2�)��S�S�Qa+e��P��R/K�Ll`4�zmSO��@	��o��z�7�Q�t%�Nֻ��+p�;��	��~�Oç�s��8��bP�9#�������砪E���&ڦ��1t)�[;�g�o1��襡 q	�,8Pm���zY��N��R%r�	�g�x�2Ld.>�T��AT��Se�K��W�E��вg�7cз5Û�s��[�c��$��Y�T��s��7�'��C*
Rx�ɠ@���F�)K@�ON�td��U�<�@��Јt�b��}� �����}BP��a��Lld�y���%�,��h�DJ>�p[y����5Ƃta�ֈ�c#
j �U��,f���У����5:�G<"
�ҿeG���)4��\h:��"�ɏ2KI�����z�Ke��<AQ��T��ަ�#yO���JU>��;��9�Ab��f�����l�uC�5#��� �O���dnY4��
[���MPەzt��zr���o߽��Z��T��zW>M�F��$��38x���F0h�z��Y�?�Q�Ԟ��O°���m�zq�^H�z��Eț�E�sN��5eӨ��0K��$���3RJ�$x_����s�L�[A��k�r�T�'y�۵���a��sM��&<�|a{}lA���M��);Ki��X�"<�܊۝�;�!_u���$Ī&���} ����eܶ5��\��N;iE���t5��x6V������l����_�MAz�aN�QEv:f/�m\U�*$�x��!m��ې-ř�'�HAbsv��2��Q�k�:�2���>Nx�X��8�H#}f�R�Z9B�7�'A��R�M�H�R,W:�_h�v�+��Y5U�b.PĒ_N��C�l���qx��R��O��)é�R���Ce��D��i2�m�tT��}19#�<�i��<n����{$�D���a�i	�E"h�)��p�?��}�c�Ȝ����.=(�E�c[��J�w#��^8��Kg�b� ��{����0���MX�;�{"��ڌm��ʁF��5٘�n�}���բ?���;Gw���޼�^=���1i�#�2��e�����X��g��҆LJe�M[	�@j�?�LB����#o��@�8�� t��L�;�ga��������G�3�ޱ=�����~C@�xF�P ���
Q W%?~�ޥ/�r_���g��>�����qJ���Z�p��D�h��O�����i�\�����<.��kx������7�Y�g"/�rX J��!Y�
1rg%�7#�}|ݍa�����k��Qq�7�C�Bũ̵jY�e�2�Щ�T�!�W�*8��l��C��!ґ�eA�Q�����q�Hf���-��':d�TU�LR%̈�pF��ȃk���3fCk���[�*!_G)��b�*<�(ml��v*�8�5Ug��RZBX��f�;�7Wᇷo������"�tk�:�`�@׈u��%�,�`�`�1�;�5�7k9]�����H�׶Q;��4����Was�ᝈ^V�������+�K�0����y��#A��pp6c(h<iSz�g�p�C�}p����l�����e`��J�����p
�݂�4�$T/h�\�&�m�	x綷!U��$���UC9'c͡?�һ�i\�./5��*�NU(q����z���(I2�d�xf��h�J�`$8K���ͭ����5���
d��[�Ȇ0S0�v ��ػs?��n�}ֈm4�L��E3�7|�l'l"�C�Գn^2{��)BEF�C$�o�¼;h#S9��N��Ă\�EM�bf7q����������9h)������jn�Ms������[e��[���o~l���`N��N�!����ц]�^(WЄ���͙ ��q��m�h�A��4�m7Т�n���F��3ޑYv������[i��?�����>�O(Ȧ�PU$&(c�C�3�B^*��YֵR���<4ˆf�PSs���kgC2�se%Y���A3��oa�bӐ�,}a�A��2z��7�on�`΢f2����F��:���c�(7����P�[/�Cw{ԂR"'+�h����H9%f<��L[�h��vp%>�=��}%L�@I,/u�(u���ͨ��-����B�]ˌ̰\߅���L����a��jL��^���B��<2��WB�yFI�8U� %�D��$�ўZ>��%�A���1(���,JW��'�g&��穌Yl]�Nb_��u7V�?����p&p_wBd�@|1ˏcR�_���a��v�D��D�2g�XW�R�R��s��@�7�{�Ou�0(���ѹz� �����:���0��ޚ�H,](�	���?�_��$h�H����룰��4�E�G~8�ic�L)����1PJ#��h)O��0����zr�V�A����e�_���F�w
0p��1i'��?54�z��z�̎�6Z�/���R���1�`Ks�C�*2��aOgˉ�c�\<����O���j[۹F"16�9ћmwa9�윘=������p���K��!��,$s;��Mi5�~���w�lk���!��������"�ˈ&E\��z&IKs�"�1[�$��k���R=��W�)�˄�=�.���I`L��A��hؾ�����~���?�P&fÀdi�p,>2G��6���=�ۑ\��6��u4�b�'�\��TF��jm B}����.@)�� ���� ��r��t{l��I�\];�Z3�A�}ЂU9�� dAB<�d��U��0�y7g���\%>�u[�CQ�����t�2��O�T+��S���2�Zv���K3��rmk��p���PyDZ�/.����X�"�� ��e�����r� �\�qi-d�5�C����Si��
������W�	��_��p�k�}���?�������z2����~��*��������Q�����Z�b��F�Ʈkck�����>�9�)�����c��d���� �rUK�u�{k)�$F���(��d4�J��vOdsP�!.A�4��)X�szM!ʠ�K���(G���=A����Ĩ��E�q�l��s|�$J�\$ݰ=42o���HN4�Y�B�Q�LHk唚� �<��U��\�T�"I���~(�5#=j%�7�p�Rsrg+����^�lz��ֆN&�
`�1:�d���G*}.#��(��U�"�2�����V��'3д@�s^�/�G��`A�g�<E}D�l��:�YiQ3�L�z�|�jBP/:�Q�R�!� �; ��^4�,s]e�b)[�~.���Iy��pĠ���w%���j1'����o���`����n����Ok�����������N�9=ֶ��=+��]��%���1�a��$ T<>�M`hl2���VN���Wֿ��pP��X(�no�÷-�
�M` 4��d'	�V�
F=�pi�:�)=*3&�Ng"�����+@�)̿����2s�~x���9
������7_j�_�\�?���j��-p�|V��S�ڟ�fG`)���n?�Z�P��Ǡ���O"�ȧ�N����}����4�k�m������\=g��Ԝ>�i��=A�
YY��s���G8��$��"���h��+�c}����:�\H>�ҕ��J�5�d#ɋ�O&�U)2�UgS��4ET��`���	Q��<���/��|̝9]n�H'��et�:���e7��P�m��/5Ξ��0����f�Ȫ�OOaǲ��08c+7��Ӊ�}.'f*gsg�*�z��!A��}g6
��V@KҔ�0�>LA��8r�1T�p3}��%���oZ�{>Ov��f��._yV糘�z��=g���cK�VtG�Ɨ�ᴏ��Gm��r.Vv�l�7���/�٩
��-�)����v!���a�^ ZmT�X:�,{?�� �������xvi�0S�
89��G�𿀏�tP�:L"ηW����a�KR~I/�iQZ����\(O�J�ՅD�}죊Ƥ}�̳��j���L��8Xz(g�Gۚ\�_�������2`J���lS�t��ͭ[\N�7P`$'[��Uπ,G�tmd��R9�P�$���N���\�ąLp�dp$>���@y��Hc?�/E����PZ�U7�6(yv8;�F�k����8��g�dN��)�,Yr4v�<ǎ�b�Ԗh��ۮ4��g�l�pe��D����6��H#Jr}ϞgvE(D;w�O)�A����u:�a*�v�E	��� �M�P��	82�V�폏�zO�����@G�!'ȱ@�}�(܋/_���~h��hH�[IßE� ,z����Z�9���7zo��ݝ�@���iv��qyqf�B��Ζe��03�v���U>�v�T������Bbcvjǲ޾=�wv��s8nD$h%���{8c�-h�փ��%.���mߟ=܆;��ω3�@8�Q���%Z[U�����c��*�o�}��u¯����ůG������s8�����e{޵��[U���Y|5�M	���I���!p�]�c(w�?�h�)H�g3Q-$�PϞ�F��jן��Ɡ]����J�ߥ�.��Z#�C�lX�z$L*́��]�����0M��CyH��R��<��]μj�v.op%p�<~�.��S9ڲ۟i�#�|pSc;F9Z���j�\��45t��7*^�2̉=���?YT��)Ά��Q8���@��l�t����1�33jw�-K��8���;s̖%__)m턮E�`J�n������7J"����_�����s���� ���;���hz�k�8=.Ɗ��9����ŊQ�A�,J4���%b<��TڰM,В�=a����n���`$w5���4��sy�G黕]��uC%��c,�\�۟��7]��'�僞J2�T�!�L���� !t�|��<6�3U����LYF�"��% [
,��IU�t��$t��I�2�2�8�R�_B	G:T�r�&A ѿS)�@�lʰ�P�@��Sb�GL�&.�O�gW��ә�)w�,�rz�Vϐ犳�Hy
G�����[��zΰ����Z۴&����-۟��l`x�;�ZV;��p0T=��*�{^�G9�����m3 X	F�	�k`�rl�9T_�8v�S/RgH�xJٹ��7�Le*'�_#f�e���a�"�)�%N\!��L�m&�UpK��F�هf�S�w�z��BV����B�d���Gn �y��W��:ե�*rٳ_
d��~�çS�\f�m]'�"�{{�5;?x! e��	�a����_�	��J*ԫd����?�:�j�YwQ\F�+�L�[/_�L��-��׿V����O���K��L}n�JƠ������
��b��YX�B�aB�Ӟ[oϜ��
�TA�Xq���#���ˁ6Q3Ui���vo3���?������a�?�Ϡ��m�_jrЙ����3gM�EUi��o�f�go,�z0����_^h�2`���$����^y��w�j�aOA�/�,~E���,P�f�T�^KZ0O�g�AM{�5��4mD܏O�h�@{,���VJ�6IS��aʚ܉� *ƿW&�&ٚ��6H�NV��a{�w���R�ʐ%Ν^���fH�!E�0�� x:U�S)��^����P���<

�H�ճ �E����o�N吼�{��6Ş�\Ur0�ʝ��5Z���ݻ��
���#�;���{/�"���WԈ�Bt����>G����������߆wWgB�,�M:��`�^9X(�T|͎S�q=�?Tr��@��ܘq8[Nm��m7�p�B9[4N����Qh�¹}٤���gd���kS6�X𓸪NM�N�"RƬ>����24F֮�ٴ�3�,���V����xaP��A(S~�?��*��Yаj.up{vp��qo��tЍm�}f��c{��Gs���abw�(\�ztR��"�4�TD��n)���e�N��z�r_�EH�ʞ��.x?S�O�+#��E|����*<�5��]#�O�ړ=_�� *T|��d�mҺ�V��[��H'�XK�Uѐe��zc��LGγ�d(�_��,AJuY�.O����{8Y�,c�
����g��-���S����F�k�8fS�/������/`g�7����S!��[�ȓ!Hj��F�Cp؞�xȫpg���oA��~<gS��v�+�O�����G�\�0"�E\ce[�8]�aj�-�EFh`o#��u|t���K��� ��'�g����^�}���Zu'�>�z9������]\����8V�8��X���(��ݖӇ�NZ��Ys���f��L[ݰh0ni��ר�06�G�,q��=Yt���)8�8>D�5�TrՈm*�/��W�� Q�P/f���=���T`�����U�ʟڪ�B�d���1�i��\$wX9��pgK	�`G(󳛫pg�ڃ�Ih���2m�3��Tf�����l��Q^E�Q.	�D��\��I$��̒Oӵ+�9_CO8�v�LW<D"=��x�E�0�eQt�rtw(	)YZ6�$�p�ƪT3"B�-S2��g,Nq����c@��Hc&�^���!��s���}JJd�g��"����h'��D+�ԛ���Y�|��ԜaS�$t�����L2GG�2�S�F���^okv����5�p�1�Ӊe떩��B��i�%�t�1��d"V�NJGxq��zð�M9ƥD�g*�(����wo�[cn��;�e�IS�JY��ʑ�2E��m���x`�k3�s��f�)�ƹ�r��[s �`��غv�MI��N�td�kk��:�V�3�A�h`M�%�Ele���m��Z��Z�\�,dZ���ߔeѕ�Yt����bl��<�N�}��C��K��X�����+�(�R"ʯ�<k��xn��c_���g=�HZ;gU��/n;�~�4��v3 ��@��*�A������]��`�ќ3��3屗G�P��i0Y��4k�q�#��2�_ZB���'Smii7��.Gא�o�����!$RhN8��:d����Oa����D��s�D���Fj�wK*>9.���&��g/�x��LXN���J-n }�߳h
a����pI!����MC٥O7@�`g����0�0�R�T�����2��hs�cMR �Z�$Ƣ 	ڷ3O������9�}A������>'��Թ�8"�dI;(d=f��x�9*���'�C�)t!
�n�P��,%����@�G�K��V���PU�n��>j���T�m�̆�N��M�	��!��s��ּ�*A�� �1s;� �I�
:�K����i�^76���}l����s�	�E��&b��t������e{������Hh�Fx��k���Κ�dE�ā���+@BX��F��W�8P��:��]�d5�T�qoQ��V''�H�F�Y�#�5o� �A�ڻ~>xt,=�ԣ`GS�ak�v�8߭��%��ҙr c�)�͈�3���p�����K�IƖ)�UV`�@����(w��=J#��� �^���B��#;4�ab�c"df.����Tܷ̙6�ME:��L��L���������&�}�.���,�e!7���e���ۓ��_��Q�20�n����x��jWOk�]p��C2/ႚ�Ԍ?f{5-�?�}�1L��̇v�����>C���^��B���{��D�K��;�$��8`
��\S�"�w:�-3�2������_3(���i�Uj/�1��e��F;�O֟�K|����T	p&V�  ��IDAT�rZ����}'�B�zow�z���^��Jg��<S��A�eX��ݪ�S�_>��Us���i����U���V�v K]�ƝY�zEa^���f��e���H�
3��Ҽ6_�;� 	@��`sG��w�N�-Z�� F��s8/�A';C��+�D�i!1�B9'.�����m�f��3h���^w��̰W��-E�O�i+�1�<�O�,;��aD�|�2�m'Q)�=*y�U�?1B�zw�ŝD�0@geO\��W^^M��hK=�`�l��=�@��P
@�9aH[��p�"�HD�I�� o<�zDAH�>:k���|�O �n�&Nv��{�9��4W���ed�,R�ӳ���\�`�\"x>��Mk��D��~��q�MQ�O\���,##W��<J��྄���k'k�ёF�4�-]fT`V {�L�P�9l�m�X����"L^>�*)\��y��}���VB����݉]<��Gl�]+\۔��<�<�;5[%�v�u���sgs?qTHY߮��-eM���}��X�
�݅��+a��N`}3����	�A"�eIц]+�yM����$<;_�^la�d2��2���dDx� ժb�-t.*;3��x���|`V��Z�V�� ��E�hȶ>�0Nn��H;F���0�UC����RGRr�ȏ+�V���T�7�B�f�!j7Ԑ��A�g��(�6��yS�r�;��mh�ᇓe?�����PNK� ,�Z��*�H2^�w���,tT��3���ۢ��]�6���0�-R�΢����Ζx�+�t�_��n�/�J�!x����BKV8(�R<�dڸb�aF.�,#�]��:�W(��*@n&'����;��Fǲ��*�|u�%�e[���l�n۵IC�s�R�A��p~^�(6b�= �@�t��J։|��T��
4d�鶖��ӣ��5��Z��H3s��U,a����=���$R�+Q�[����c���	�4�D�D���XS�)Js՞�܅�2����r�B3��9sUM�!
�2Y� U���_pN_��J�;ۡ�1��g�)=A|O�܌��|�
9�*l���=��n�u}��]YSIF����s��  ��
���m�q��F�h&D+A�'0��K��z�%p[Yp&r�T��%�.L���Z���ܳ
���P$p%q���Q ^"�C@���&@ߒ�a��J
xR�b���u��:N;Q;�L-�2��1�PkK����h�I��+�ԡ��U_Ɉ��>���j.��<+1Q!x �Z:r�U�`1f�c��2�Ǘ�q��Y7�.c�ƛ{e_������;"���*{^}{���XFp s��.�/�;4��Q<�
�hs+��|��!g�@��_́��桙�-l���R�|�]&�����hk�Q���_|<O����z�L��6���|��|�?έ�b-qh����i-���0 ���譩����}�����i�� ��x�	�mh{�Ck�ϕ��7�U��6�<Y��
zD$�bAu+)��wIX�|ΈWJ�V6�oʂ�&'�@y�>_��Ξ��E��yY�.�x�\I��KˍX�p>[!Ъ��[�5Ek�z(���q�a�yR*A��5 ��^��9�0�2��s�\A�\\����F��9Q$�[^���%�D�MW��H�!�GT����ot5��P����aN"�Ռka�Xc��s�C��5���>�G�#�v��aa�0�o��ʔ��>��j����rf!T/,".�����e������2e������=�,ɮ4���O�V�JWA��l��W�����
�k�q�F94�h��h�P(�:CG<������s�GVS��CGged���ޣ>����@��|w~�m72���������W�!�bP��Ϧvh;W����>�� c��,�����F@
�Y��\� ��=�+3���IҞ�uxC��l�nv���?W!\�d�穴�	d��E�W9������*��Ρ�ỵ@�S-A����ZլՅO��R���d�g��ݛ瀚'��#r-������|ik��UW꜔7.3H��x/.�ώg3_jg����F��.(@e<}d)Q�P� ���4�$~��i8�%(�\��^,��@�T-�H�s.�IW��(3��yDr*�s���<*�G����DA��o�v.�k���V�<���8+�y���~_��Z�u���j���7�Iˢ^*	e}�-�"h/cV�i?��G�T����jn�_��t�@Yk6lg�����huI4z��%x�R�+�ڴ�^-���:��?�Lƀ�l���>��4��������?����
�a��F���w��7ߧ��>�V%��� �0���V��P��g/S(5�LJxn�υp^7����U+�2����me�%g�֦^w�p��Z�.�^����KR�K��z��#�PZ�t08_wO����-	֠��~Ғt��v:��*�F!�{��M��E�+^�64�,��]���j�\�x�)���=~rV(�ra�ɲ�OUA�d˴%��y�+7�s��P�l������DuJ�L��ᙝM8d���9�ø��:�^�5�½��5\�q�j�<�C�I7�r�?�Of���I�����@�����N�$���8��Ȥ�L�A35�LNR\DX�PA�k���OON���+�O��;���S蔔	+�f&���-rjQ��M��7w�*��M�Jώ}����NZ�]*W!�� ���B�NU<�8.DN��>�@�#�0��woӥ}	]	
W�+Y�q�$Ȳ���$�h�Bh�����z.Cm�w�q�g:$�	N-�����
]���M���}��K*T��´�Ce��_������|��w����W_}�`��\�����-h�t�w�D���w.8@�A�Z<{�$�W����O����E���[�N��V�x��+��8�,0-aి|w��-�����{�r�`ӎ
�e�) ��VC�"��>�ˍ�1v �$�����X8/ea
� ԡY���n ���J{:W\mt 8�B�Q�֑Ǽ.�ex�-Q��Xu�I@�(��J�$r�i��$��k���L�O�j��:Hh��<���_�lI!��J9'T|�UW�E<d�^d$w�dk���U!�Z�˰�c|r��d�ѯ8O�Q�Ě��l��S�s:�$�T����$�Q�hw[�����3�׵p�i��gcݧ�Fb|nY��Z��<�'��3ivy��,�]�)Rk�
Q$�d \Ž��}�$T�B�w�~�wФ�S�pr���)f\k�N�hsO����~��ME��U��uR"��2��Y��`-P�J�$�v��<}�=�>��SKv�����W���;�p�"��v�����=�{J ��]\�[b��ma�A�˴ļ���G'*���W���j&l%��2�f�W�c�d��&@�I2��<4�;���V�'(���j)�4��)A���r�z��BҖ�����r����@oE���@���z:�J�n�}W��A3taC%�
+�6�.y�g�&,2u �a�y���5�`�!�#6@�!]Z�4�f�5ʢA���;@��,��p�t�=P��e^#o��	�e�r/�w�"^��O��A-f;(x�Q�3go����DS�����CT��@~{���X�r�=��:2{/s��2
p��ޖmr���F�~S��Q�ZXlf����	O����N��Q��J )���4s�jDY�~��F[�d{����x�z?:>M�}�yz������{�E���|s�����{ �&ȲO#A��vn~��,���b�±�	�5F�XȩR�����BF��9��w{Ko�Nή�m1JϏ�����v����3�����`�%(��%wQ�ֲ`���lXv�=} ֶ&����J��@�/G��1�h{�y��h����M�s�-D5]�jJ[�^����D{��+�+���H/�J{vH�^I����5�N�
ʟ˧fQ�����l���h�Xpw'f��t�)���s@)�ss?�i��2fռG*>h7+��|���c�Z	4�k�Ύ���?7vͥ4T�[L������S�3��Ź(7x��hC��ַ�,��~��e��uw�������|ѿ�*���c{_C�z�̲��4����3���	��:�u�KAΪj�|�墲�[�>��ҺQ��A��t������i�ۡ��_�����u W�6��lqr�<��Y�Z��Wě��Yg�;��[��dk�>#B���
�"D:H@��~��ϟ��O�>O;��p�r��BQO�:<=� �IQ����G=����kۓ�E���O�ȷ�sCkb�Ck�8�[06�B��o�]��Q~(ϗr%�|��|��ﵮ����nN�֡`�dr�&;��BӔ��r1�@ ��H���{����X��hO���A�=H�VA��N�5�V�e�}f=ᯂ������]�qKv/+�$�:<�r�b�M�G�I�N<��[���M����'�RNXhC���V� �ME�/ɹ�)���ɢaE���zc_�:ʄ�� �<�n*e�)M�I�aV7����[h���tR��u|��;>[�J�߿�z{�ꅃI<Њe�H+u&k?���V��������rU�Y��m,���W�[��.]O������Zd�PȖ�������hf�$�����g魃e�N�
��[��7�L۳�b�����X�D�IR���#mj��!s�!Y�ݛ���y �,k�'*o�u��T��[��Lp����ގf�t�b��y�<g��A���k���JZs1oŻ�B%� �t��N�'�1W8���]˶*��^��l�k��,�JKq�Z��%�3�K� 4�V��s�٥�(l��!A�׷ ���#�Z�/q����w�T�KѻQq�mqz�z��`���G�p�+@Hj��¯�AjۂF��t�-��ڂVΒ��!���Jg:�_��/��u���kU��xIl��U�_k��w��0]$,!AÓe-s_��H>�� �a�ʾ(x�_�J�,㻕�vR"E/�S��t$�\�R���~ e�Ƙj���}e�ٮS���������bѱ���Y3��E�����Ӂ��;s�D�_8��[�w��$�8�����Q�,��X�n����j��Y��,�'ѧ ��'�t0�&u�Ty�w��]�����'�S�˟����h�џ_��7�8�l��g)�X�0> RoT�&oy��L�}B%r���\5A�*�);\|Z��[;���E���o�o����;ڬT�^�������켍CG�Z$��Z��P7U��	�ҏZ���+aeDMX�X�f
���4�siF�y���t���qnAf]�!TP9�
$���%��^"e���֍�bK�<�$.�7�P�Hݩ���-���D�ڪkwP�\a�b?����	d�Uۢ����!4]/��D���6L�Ꮶ6�Z	�P�%d΀� �5��񇋢d&�us�Q�Y��x:�Ѐ��,�}�7������VG�;�	���CU\g	��u^8�Ta��l�Fz���y��"�5�
�r6
�"��ަ�w]x-����[�e���ew=�J���@|�εU�tw��N����+a^p������{Eb���Ѯ^(pֺ>��Qj�����h�q�%�.o����k x`D0�M��{)JR���Z��ʁ�;2�A1,i5��$թ�Ł��pk�Z��f;��](�R!�b�Y�>�:� �t]Fl��8)Ώ>�$����歨A�7����ltfl���dׅY���sK>fjQj�4@��Y{w��Z2Yr� no�,O�\���r���wqs+����:x58ьU#�p�b�@R�z��K�;��!�^_\����ݳS;OO����]a�U�(���0� �	t&|��]��Xf�)�QUvz|m�F
x���XK`��EG{tl���F|����R(��Ψhz)��2�	w�S7���}�>��|�TP߂��𽞺��\��u�,A��zg��%;W��,�k�Ҙ�]�$NI�Gs$�{����(	5��3?��W�l�-"+pT\�Y�	X���깪�,5����\Br�mh!��K&q�L_%�w�5�! (�B�-��_�F�3�����;�!� 6�n�/�--��"# �Y�FWv�������vT!��W���[0U]�}�H��K�y��Ӽb}Yܷ������"ra��j5K_�}�^ܜ�������IN�k�d[��%�-��T��h��o&��w�jUm�BP�1����*�4�6\I�'��.���{Oָ5�M����O[�yH�(@CY��ˑ��'E��_�,+<�C��#1?8bY�j��	�[�]��p��(�Ц� #5�ܘ�g�)�M���AnfR�6���.8�ö���N^a)a�L����I����g��9�g1�B;N��w�^J� �#k��<x;����Z� �����la�5��hߑ�O�<I~�Izz�&]`�������	-�\��]����#x���pM�{�57�6��T�K�N���+�5�����H��j�U�����:X7�k�ި�Zۚ�ɓ������v�~ש	$v1p��Z�\~&� �N��f���g�W���ע�P=yt*@��v�v��C"�)������6��qP�A߳�[v�������c�	���_�g�;^c�Tx0�PEok�ݥ[W�>H/��� q�Z�����R����m)/��vj^� P���D�	�b��KԦp��K4Rv�����6*���0�u\K�-���ɭ�j	k��C����o�������j�Ud���vI�h�W��#>�!i���\3�+t��lm�,���ߋ^�̱ƪ��a��]�%�4B@i������W��oiK��J��������I>�n�*�>T��oԎޔ2��}X�^F���ѝ�]�v 	0�Fi]�N�+dZמ~�K�Pƌ"�K
���k�qs``vtt�v�沠@��.0� +��M\0I�9��9z���l�R�p玆� С��>�x��p,<N�im ˔�b˷�1��Z��x��=��MG�@@N�z9���/�H_]�IgW��B���J.R�?���5�Ƣ-����}>����g���Y�����m�qr*��=;xWs߬�P˳�|y� �+�ؠ�=�[� k��̓0%c#?l�~L�����W�����L]s��Ѥ�)�IZ?G)x�9��?T��#���{S�^wVQ���xC��.ިtO8�n�/eb�z�j��o8/Dt�+�qb���G��ޮ�ൡ�1�~��pvy�6_��-
>Ĩ����7?�U#��BRR������L�������Cw��v��!�܅T�>�����ç���M�?�1�7-t%G��JU���z��e:�;H��'$Ϋ�8�7HZ�xm�cj�������z���:� ��-�퀞"8�W"��w�V儇���b�CE�p+L06�>Hl���#��~Vkt�	2z�Ⱦ�ş������Y�fmn|<F l�Ô���(����ѳ��-"8,r�h����z�\�����?�W��ֲ'���;�r�6��Z�B�=�����-3pʕ����&���O.ܻ�U�`5�Ŭ:<1��3��|/���n��'��R��K?~o����c�zv���Z�Et�6Eʑ���=8y�k�jZ]�l�҄�p�v����9ْQ��F��l�tQ+Z]�2�t�TE�;�t�۰<�+f�됖�|��縴sA$� ����wq&�&UD�/�{&Or�BQ4��H;��ɬ%_��h�C���ڜd���g~j�m,;+���7�w��V��������Bҏ;��T�����6H޾j̞�r�b֪��o߼J�W����Xl���0%���E��0�p ���,�gj
t �ɛt������� \�Y���G��Of{'C��-`|�⻵�?O��a��d���6��r����l�J���`�,�+o߷��&�2Y�����t���{㴾�*�o�*���lt�1�Ϲ@Q� ���9�Z���RhN�Zw�x�U�}�ϷMơ@���t��Q�i���j��7��C5j�z��q���x�k)����P�:6m�x�|�b�p�Q����T����1!��p����'}��xy�^��G��k򬷎CU�|9`�gܲ&���X7��Yr�"k����������5�~5w��﹭C��8@�d�f[�k�ʻ�ttԁ	D��`U�U�<�ONR���j_��+��U��Vii܍���EZ����Ī�k�ewW��F=i#��J^��^�Ģq��	�2��_m�`��RU7���O���Z�CF �Qd��*K �?~,`�-ISpQ����]�޹�b������I��.
v����;�ן}���=�?��~Mֲ.�n< s��zpf�f�q&�d�Q�6)���.|��O�}f�3�����<�J]ӻ{���Y��wu a�
ipT㍝{}����,9��	[���hфmӍ�<�i�7l�����￴ lI룣c��H�7��鲻vut3�A���{:R��x	I�8w23������>�l��e~�X���o~)Q���=�\8!ΛyU�V�
 k2�W�E|�L�C���0և���8?Rt�W^#�+Mvl�y��&��'�^�Yٛ�<l3x���C�����;��l@Ax֛�~�G��	���eZ�D A�Ȃ�Ֆ��6����Hawۨ�]&n2A���ŋ�����L����(Љ��=3��E�z�psiC�×-���UfT��meC
G��+W����ů?s>�}�N�ߥ���=ܖ�We�ד��td�M8�@��\����5<c�G�pG��,����4��v�tX-ڶ��h���g	2[�z.;׋,�-3�����T��� � ����=�p�Q˥t��'\jG�G�����x�Bb�T�u)�.H�N�!�ބͥ/\��0SqW���SAm�VH[���l�VU����8�cZϥ]��Q�E��a�%r;,��P�~��ߥ�w�شCkC�Ш4�^�G"���5�D�j�I·J^��7�m���ѡ����FR��pX�=�:J;�'��z�(�:x��q(q�2E��?WVh[t����"�;ܔJ7�Y�������/;N1�`P����y�.�7����×j�n���_�z1������%��2ڢI�a�Bఔ�u�z�3�tc*��	D��lt� &�)�]5��2z�[��;9<R�{xx�>��4��ق��)�����7����C2�,�}O��;�˴o{�h�@U0�pL�n���ξf�@��Tk΅l��LV��u��FhK��,�E�� n�����P��'�b@������@�O5cS����pAܫ�DAc�$�nɣ�4/ڵf��Y��Nm~��z]�F{� �y&���܍F�EW�x$n5F���Q�B.���u�BFW���:q4B-�����oI?�m
���qCm��{�ׅ�����vZJ�%�f$8�v���܅F�u̢����E�E�J��q����|���ڑ����>�o��䟹켏�.�܈��1�'�F[�,n��|۠��ƚ���P�$0��Y�B�IѶm 4H��P�:���-z;#�qH�;~/�P����d�,]^����s��W�V���ʹ��3
!iK�v��������~�Ĥ�G^����yP-� � ���U������N5�����w�v���3ٗe�AZ�S;�ok׎��-����A!9�]��D?J����婞��:^�vh&�!4/Ckۘ�j��Ո̿tKF��|�Y�4�Y��}kq#���_@=d�E�h/�q}5[m�ZI`��-�G%Q����6c)u���@�����K�@�����M�ȣ�>	A��Հ���k��|���:-ə�Qp��*Y'9��h�'�[
�z>4��F8xe��D,}����<���rJo�	!�p��6��ɡ�T���.��l��խa*:Dσ�x����Q*,8�7�YN_[��q�ͬ�,��T��^��gO5k�b^�{G�Jr��#>I�6�4]�~��YPb!�����z�4�!�@���;�����*��U�w�~��T0�lR'��+��4A+�߶��;�b���&��p�r(��a�'���JrG�D:Itȇ�- a���

{H���&�(�w5��H���C�t (��?�����*�u���H
�*��ˋk%$i����y}9�
�]Z؁����GR�R�ŉ���Y�?#�G7�5A�#��j(}l��ٞ�]L�sb���֨�,�H:
g`���d��R9R!G�<�N8q��5���ٚQ���м�!����_����W����~͞�)��$Y�����C���� �ʻ2+�%6
�`_t��nY�Fm(i�1	-��Q'TB ��ݿbk䒬�:���mic��H�R���I?��3�u��<�=Z��om�]�1�M;����|�m��y;��Ѹ�$�zr�^��O緷	;�%�{��J˖�����3��s䚻j���Ɇ�:�
�ǅ��n{�+R��{\�BN�n�L�W�~*W���~�&�]ԝ����~g��~u�bj���=��٠@��s�s��Z�{7��p$���ήԼ�	-[ݶ  kn�����T���&�k9�L{aY�v?mnW�dŎi9�0cAj����T���TN��+���H�B�YC��Md�1����3��{���r�$�hnՏ����+t���sr\c�����'<�e�&j|����+%�<SWOr�=��]��ɥ2���.L��ȍ��bc?g3ݤ���D����u0f��'�@ #�tBHָ\RH�
��Hx�sA��u�ڎ�Q��
<R�xu$w#<w�1
�����L~�4<z�>�7�J�x {�vP���i�Y�$�[��؈�����m���J���[���v�JW���.�H:p��k��i8�sD���6oS������Uz��u�Z��hf�$Q�{���JQ��Y��ӕ�/���뙤d{����+TM?[D˖ĎQ
i���q��m��{
u��� mzZ��;#������c��eYb/��X�*K(ґ��]�Z�7�kT����٨�Ჴm	9����?JǏN��In���=�@O�U�G�;�UK�����m�t��&s�P-3�CZ̸Y�6�&@��	#':���Щ��q�����.ܗC���.>�T���;�a��yTЭ��$̓�j2����Z7� K����K��#V	5�X�s�;��t90��粸WXLq���eXS��t���r�*I����{�r N��Z��r�tϮ�w���|ظ�&3i��H>7nJ�EܢcKQX�Xh�o�y�������i�=I'U�Ξ���T���.o�hI˦i�3?]��^�^��EH3�po!� 0�h�����{�ju�����s�p5	O�\�pұ�
S��"���� ����<�-������Awt��>9uA�9��,ח��/�����׿U~������E��ܺjL̃�&�������v0���VQ0<���M�{WW>��{m���7��Qq:�����,�^4�.��jǅ뒮˨������h��4��� ��E��`�c��7��E#��RW�7aYwc�9�OHd���|0ϸ��:��7�w��@ ������رѩ�c1�ƣj�Q&+�,�FZ�(���u���J�-T���N��ޫ[.&UĴU��o�ab�@�מ��0]�M�%�&�����n�ԝbv��q�G}�jmj��E��mwm��x_��&�'Mے�>h�E�	\���A:�J�|�#u�X�j���n��ͅD򡖠�utr��..u���O��T��u�X޼|����w�9�vDy³��	���r.kL�G�	�?nv'~p��]:!e-1���ܥ�k�������M��tĶp�?�ĭOroz���w���;;K����̗��r���V� AB��7NsD��v�2��H7|I��Щ���	�7VpM-���Q�B�m����u�A���Oh@-㤡U��E�T�^q��!�G�B�ܫd�gA�c�,��z��������9�.J�|t��旍�Z��o��6�~�J�[���$�Z{N���c��ѝ�Ɨ.=K�WX��^Q�K��%����ep��h:ܽwCY1���7�GU�8�\�ljԝ�F:��I'��id��
A��NaT��q�8z�f���a��1�N�"�b,
��#,�D?}��Q�髯���a�@�xG�JRJ9��YU�ζ��X�l��:@�Q���ĕ52��Dpj�rГ�2�6+���K{�;,ά��P(
��f��*����~:��6# ��U�h���
���?KG�>��7r�x��]�>���2c̈́�0�@FA�f8��&U�O 6���?+7Uz�T��x���(������6�<]\��?�������ÃG���� ��},�zm�ۢ߂G@P��3w�p$CĽp@��t�@��j�H�#kU��t�	�`Tv�2�3_Z�\آ�<���yH_�r�-V� <U�:	�לD@�c���+���a�X2[��8��@bg����v�ֱ�PFk{>�B��΂� �ЌM	��8�5��`S��������v4S��B�L2@��{0�,|�J�]|n]���K�:؏�ܰ�rP�%������`L�j̒�]���ܱxb�c��ª)I�h�Nӣ�C�1Z�h�v�h*a�د��^����[��dH���@�/��ʼE�q�d(����p��wgkW:�]�I����#�\Ҿ[�^��ڍ
�I�j�xe;��o�i�lK��*�=�d߼ycAr�잭[�b&��u��^큝�X��t$��B�6pc����-(�~�˽��� �
��g�ӓ�G�'g�<	�G�c�x�oAuI��#|7ugs'lA��9�3��;Bf�)$W�1Pʫw�Ô!3P��H�ei�����Q��3k���~Ï��W/�yF�c0x�5�M����2�\�^��2Nh��Z�;C9:��ɾ�r��hM�j!��*�Tz��U�{>?���2�{^#�Ë�/�D;c�wҳO>J��-�k�i�s���u:�ݦ���\q*ˁ߯��#_���=�Gn�c��k���>K����M�#���#� u`�zQ�h���N?���$Wj�u�ѡ�AVr�Q��X��\��h�of+ׄ�kF��X>��S�����(Zі�N�r,��N�� ؽ�H����A��y�a(�^K�N,E�ǖ�Vk������g��>�N�MR��KT� ��E����2x��tA���^�z�'�@��7������W_�Wo�t��G���)��P��V��Rm�V�Oᄱ��m>�L8/�����7�PuPUw��3�ף����M)�nb�|���X{�	jPx5��+�������&��R�hI�KoWo ����1�jD����M&M�hf���%7J��'<hM笙"���T`��C�Ͻ�>mlt:�<>=},���}��?{��������=U@�'�������!�F<�	)�ƻ7�J���	�H�{mJz�S)�*�|F��BSa�:T�21�5���d�k�+p�d��:=����}U�pCgv��g� �N�q��k���!d*��r^10jm�˹Ь��c�jìw�V7�4�l�R5�-
]�/�d���8�$(\j3�� gm��"�j��$�nDM���.�m��K�e�8���-�>:�\f��*,�P�S��]\I|��H"-��T�������?umt��wV��+Bҟ��4~��0�Z� k4{Ugr���쪭O릣�I' �P#�KЭӌH|d>Pރ���5*�j�ty-\�`�P�/Cm������\�y:�;��[1�v܇��W�H�s �ɸ�r)漲��ǱJ8�P�(%�Q]�5c��aydH�aCɄ�]�,�:/!.0��Ŋ��Ȳ�йܙ��/�����_�
��ZR�UH+F%_�m�����,�����xG�<�'�<A�(k�_zHM���fl��o������d�m�le\:x�#څztt��?��ftW�/�"LY:q}a\�È��J��JtؓU]�
t��U)H[2 �<`�$��S�<����4�J���{��k��8���9�r�*�?t�*ti����B*�l������ԍM����~aA�����EpfQ/�X�*����u��k;|ik��.���p����N�����+�w6P},����A��ls�[�u�P�9J=�
Y�t��
�b����V��=�
(~�\��RI������+�d��LP�	ʼ�ĵ��L���W���������7"UxUwT)U�V��!e�C��d��#��/q)�`�H����"�?{'ay�H/6g�!n��M:hl���4M��^\�p�x�V
F��K��q Q�5E���r@�T�옓����l�z�ܘĀu��:��֗���J�;��_%<BbbU4s^����E�ʿݹ�� V�{V*s�%��<�L;=��ǅ�y������D�%�v%�>w�ɾ��?����}�:�e�l�m'�� ����RvE+�Y�ފ,3��?蒱\U
 )H���|��+Q<�V-KU�vIȦ��
�9����ʒ�M�m�;��O*F�R6л��ӗa�?����ܣ��������7��)���ӂ$nFg���4�E�dtSDP� ��Gn�k}E�ݏj��F� K�����\��<R
ի�ݎ61ߕ����N�(w������v�x6�ɘoGW]7И�o���.��ga���z��TN�sW���X�I�q������N+d3��N����I��F��k�wڢ���ף'��s���G����=]׷V@A9ݵe���(nVR��$��x�ֽv����?���y��I鲔�I�	ylAc梱���҆�}<N�[�v ^�]�B�I�ށ)'�ӑU+��(ޯ����N��p�R.�)���U����2� k~��Uz�򕐲l,��]ۄ��9ܳ�o_l��tr��v	�}�[� �ℂ�mF,�_�
l���AS�S�u���(d�}d�E�v�����ttx,t#����
���m�E��о���6��~�n.C{�U�C{�C;��m\�fi�P�5ai�siٌ�RZG۰�D&6�x�T����d�� �r��;���EՑ�^̪�³{���8�Cg��y_	�P��������{ U5
�B�P���ֳ�C�p*a�Ch���9�P���;{�6��"d�0wA
0�=v}�:���y��t���H��pH:��bpX�6����p�U���	���W��<�ZT�u��D�(!��S�,�@5YW=w��~v�cW�7�}�wm ����reڄ{�n�Iڽ8}y�����.��x�W�]��%�fi�<�^M�m��}�*�
�Q�s�"������ByD��`�ֵ�N��ϼe��>ढ़�oHn�2p0�m�S�]�e��,�����@<��t���u7���p��2��TX�mT�hp�񾳾~v��U4{�s��$^tu���'�GN���Y9L~օ����C8�k_��L�C�~-�؍��YE*������"f���l��<��-��F��էR�ٺ����d�Pw�fqm9;�H�,2���@e�əNJ k�!�"���~ĺaV�*��v`��z`�Q�*Π:�qu���x �tU��ė��t=�U�G�u"B]0+#>�ړ����u����Ʀsݺu��ӧ�����6F�Py�q����'r�y��i*���:Ӎ��`�ù��@Ipf7�=)qfi�� t"־�n�1��L���裏���m�j�L[TrV�2W�(?�?��b�m�2�2?�Z'�KvW�>�(I��U�e�9�̮�����6�N���z���U6��8Ǎ�W�f���rI>Z��ᵓ����LW�̯���u$��X� 
��Ar F�k4'�\��-��V*�t�9E)����&�s��(c�i�e�"]ܹ��:���mY�n�yk6�浖��zE�ilI���+���N�J%�"Y���^j�+���;�c�	��[�_Z�L�����(�c{�^.F���h���Y�mВ:N|�ߜ}�v�����P��%�k�w�x��b#�b���ٳ��g��rh�y��9O���'��\1�l|.F��gvG����PDnX�_|��ڍ�^��́��:*�wgR @�ý��T|6�)�ݷיWP�r��J���� �Y,�
�h &� T�4�C���U����<�<���.j`�׻��U�Nsh��#w+cD�^9�Ǎw�h�R�P� T!�vhl�H8���ˑ%�G�sT�����e4���<ir���0��+�h%�h-^-3g�>?�-w�Ꮅ_m�����ῧ*4�\�"��(��
#�`]eQ3�F�/u��n�\���>=Oˬ��h<�dg��D9���)t~��+���̨��5�S�,���@G���Vׁ��b��I�EF��=+*a���k	��'O�3�'�K�K?Flet'�?3�b6���8���"X�6�����Шv�c��QNek�	~����]�Q_�-{9��Y�>���l�B�UQ>�z������Ya��/�p��Ͳ�7����E�����zd�v�s�z���)=:y�UJ�Z��ˬ���sd8�JD7�����T�rȶ	y�ą��޳�!�~���j��n�+�ޓ9��yᰡ�[��1b�j�7ns�jnY���Z�ld@',:�-�����{���5h��n҉������:�/ߦŰN��wiv�&,Ze�
��,�
n�xV���UrW�^�,m?{�V[��Ȭ��C�&s�_��g�KJ?��wk_�����iH�X�s��nX��kU�?�����Ȭc��3�\��,*�Q��m9̱�G7��jn�;�5*]��Z���4� o�V@�T�p�5h�=}t�� ��@��٥b�h㉂�' m�T����K�>�͊T�Q>��(ɿ�g��SʐA�n�x��Xpy�����_�:�X�6��җT��^�ח�����q�t0ZVt��<�q�ɥ�-F�y�'�w�'�^Њ��F�Z�p�z(��G�V�IE�~���T<�S[2 ��
VAv�`���S�oF�l�F����E�� ��<���;22���H�9�]:j[3�� 3� Hl*������Tctx�z ��:�KgFh�ݸ4g��N�����=9�8[LW��j(�+1�=�g�l.`��x��x>N5Qb�~�a��g��_��ݝ���uj���DuVu��Ȳ�r/Z��F6��Y����{ۊ@_m�,ԡyj������W�#�u��~�ZR��z���l�V���Ư�+�g"��W�\cփ�lm�]�!
]����:g;�=X��ڸ�<#���c� ٞ�ʘR7N*.����T�J�ƽm�������h��ίε���6x��}�"��@�s"��ߨm7�X[I�i*\<�m�ㄾ��lo���7��~H��D�밈ku�b,�<��Lo޼K#;HD��w��n���g�	i1x�Es���ʕF捖#�3d[l��i����f��8]��I�M̕��82=) y."����2�mU�jq�[hQ�8YlU��F��vlcL��٦���a��`�>}v�Jl0�J��K��ަ��U��j���P_���ե+*�,V�#xB�[Oi��R7�z_Z%U����4:��p�l!��ñ��p7̊�f:Ql�k��T/	��j\����?�o��	��snK�N�޶ÇyX�<R�mi������ ��J�kB��|4?����Y�)z��2f�w�~����s���8�>w�pmQ����2ߥU���\�����6�*@~h��5	��U�Ԥ2Ț�p�N�Ӯ��ބ;�%����O�Z2ٷ��h�0��?{_;vF��7��+��oIIH��@4���w3�R����I7v��ߝi�Hg-h�#�k���ѵс�H[�����1�z{���	��e�)�t��D�J��ҫ߭P�ۦ�����{�9���쒐nwH@!9��Rr?c8�����t�p�oR>�=�o)�_Z�B��ɷ��'i~;��oȖ�O� |���rյ��ҳ߸�R"y*�mߩ,ٟ�㑘+�IT�=W/����ۏ�������RV��/�./=�e�o���9'���c �t�����X�L��5x���-I=�������~v�v��d�::]x�_����o�Q�s3���B�W�@ɢ{�y�⅕�!��PI[!F	(�]�g���Tc;J0��s.�
v��Ҧ�ꥁ6@}ϒOT�@,�2:T�*E'$���R��9.�Fr4����Lg��iS{�����Pe�n6�u������Mm���U���|��@B�]�X�rE@ ��0���2������u��-�
O�h�$)�b7�O�F�3*~����Z�x���v��1ֶ�[-�f�6�+�D���&�H	����I�iC,Bv�����ךּ�M�yO�y3�8�B��g��`wh��L�\ڂ���(���A��G���0]]L����4�xus���`��j�(��`A��S���Zu�;��(���b<>HO��>����6�Z�V��V��Y���Y��0�6��a��a=FU��9�@���%�	��`�Z�O�Gل��xܴ�Q�j��[^U��/�YXHm�2u�Х̄������$ �9��������qk����6�Qd%�ql����B��5Z�|�y�����dA~#�����A�XA��/;��Q#�~�
�������ߴ!��ć~�<������=o^�L���&�lB�� 2x{�ZӼ7Xr�
d'�S@��Y��#�u2܎������&ڃ��5��?H[�;�d���c�4�Y0f��	���6�_�x	0P�a�I�c��m�wЙ����*�J�"�|m���Y]� ���f�4<�{��(K�<����w��W�3�!M�Z^���	X;�C���R��0<���R=:I���o���b�D����~d���������?}�^�=}���߈hW�<|�0�b��?ɨ�R�^�6�NV�u��<?�� �D\|�ׯ_*�?��Y��o~�>��s=/�<g�?����W_}���se�r��wZ�EI��*�����|��>�sN��:��A:�Ƌ��*�����	I �	�w�sz9(�jg��-�@�r�,�!��z�8�Z�Evdj�!wY�X�C��)���M�[�6��g<~rnBGOrF�j����z�0���l�9�ww��G�3�=ae�uW���|�}ڝM����Գ*M�,K����>O���*,�A�KU���(o	��� ���*��C;�M:��b7�J��1���R����	#���% �,l$ �k��,�K3����2{[�y�wM��`�}~���M�ޮ�>��W�f~����F�tk��Rϝ]K�l���Ȃqdgkc��&.�W��Ҋ�5�s*,�lq����>r�N��'K0�����4��F ��p�*z]�?���`,񥅌�8�T�K�x2�D����]��-g��cq���h�
Kq�3�6���L��-������-HUorZ����$3D�^����v0�� �!����E/����0�����vt�Ic���õH?�L;,T�J\�  �z�=�}�c��z�Z0���
�g�.� ���H��#0j6X�;F]+��pC�c-	����>�����Q��Y�Ⱦ@���<�L��X��uf����,�aK �EH�q>sn,���U����l��C�����ko:�]3"�����U^� |��4�����#���>��P]��H@@�M,S�{��ʥ��������G�����p��LR��΄ar��w�g�Q���/Ŭ�2�����P�^��x7WWbx0>���LP{r� -iG�3���:����Z<1K�=��8��+Z���#�ԹoETuШ���{��>��3��\o~���������?�o��֋� ���a]��x�L���E{6�'�~��ϵ�4(�;�sY���������G{���
��r]�����xv&���--!bT�`>*�䬗w=����>Em��/������܁���3�j�vhڥ������O�~m��^���[�34? 5y��m����/f�����!B�Iq�A�6���2�Z�vm6I�!Q���ɔ�C�`dA���\9z���K��w�4��K;��ڵ{�b�ǌ���7��a#p�*.c�����4\U6�X.&�!���M�E�Lw�*��il�}x��w�V[6zw�8��\��'2P���?���,C\��]����͕Ͳ�J��B�b��+k�aN�p������ۖɼ�N�b�l!WG��ɩ2�w��Q���L��)�KQ]��	0
����ݜ��C�rT4<W�9s8?p�)?0ĳݸ�C�����ބ�q�9�l�*G��f���9�c�*HE�o�VR�r�1khkw�*�Qw����Di�@���v��[|^�zPu���9��w=�
rKR���2������sV�=�����-C,�6�1>�v�v�r`�a� ���ۧ�Z����z��h�|]V��h�0����?l�-��A
�)zrK;��E��~(~�ؑ�n%��*��~��*r��q �KQ����N��<�q0n#'`��EtA��y���	N��U�����$PU�͵*KZ��)g�"Mh��!4�q���,�
�w5��wijׇ�A_��Nt���U}5.������RO+���#)<�M}�. +TlP�J�P�F����ܸ޼���c��3�<'�m�EA)NH���̬�{~q�}�̏�}���xg?���k�c�t�ϟ>U%��������˗/uN|y�$���Ɋ��������������$5���|�$�9�,��IF����G���B�{��(m Ȃx�rT������(�AnS��k>{'��4�u��c��Š&`O�4<���*ܳĖPY�͜��������������E�MU
�v1�L�.�U#s�@���:ZՀD���|H��`��Y�8�ݖ��=�b#3�UE����k�ւ�K7�tP�`'��R�Z�Ұց֦�|�K;�fw���t~u�>{�<�o����2D�Y��%_����|�-2;	(�UK�v�(�DF}�ô?X������t����҉U�[����Z{a����� �4��k/0o����E!4mch���D�K(2N-�]YU7F�sk��V}�Gv���vtc��z6�I�U�L���`9�V]���8\7a����k���:/��*���SP>�����5�nP8|Q�"�J�0��G�d�ڙ+�b���xR�چS�h��E�u���[��m� Zcɑ��-�����Ȯ�2��������:SM�b��gj�Dm�C����?࣑�������Լ������֮%J#U�[�ؒ����J[Tèɥ@��=��UO���hT%)v�JzҾ�D(h�e^�?�TP�޾z�F�b��?A8+�=�Go:�����Q��������`�t�Ł
���R-��bH�2|��s�k��]�<��]9e��\&��\�k�:[��6���8�FO~hA��)IS�(+�<@���T��(|�ѭ��k��B��RB?�"$Y��i�g���� ,d'�}zٗ�A�b���6+�#�n���oi���8[$���}I���v��uo�^BM�� �se�	��~�.D�r���y����/��|x_{���	���NR���ߦ����?�)�����?��_�2݈n
�S>�+�P4�l�աI�b�*����=�W�DaL�{Q!gIk��oH��B�����u?>����`7!�K��_���,4�+F�,lK�����\�d��J!�򑚨`��6Kn�?C���[���������Ę������]���?�7��H&�3	��l3 3�J��NB������sD���=�f:;�-RQ{���I���0��u���SW�L��I*9�?:N��8h�����-���h&��ki;��_���*[D��/���N���:�M�:Bw�n(U��h�2�^����>>�NOO�ӓ�=��ýt�sS��f�b'��{�^-�W�d��/�ծC+!��A�|[2i���K�6�J�:>{��|�Iz��'��䇠4�앀p���+>f>g�t��;����؄+}�� ��lB\���-���GlW�&Wȁ�Y�AN�#' wR,�)�C�>#�f��r[Eu}q�I.���꨾��2��	��=�/U���}>��U"���q����nnId`3���:���˷���7���s�8fO_9�l%e���8��� �u�{�B�l������8yr�v��.sg���(=;},o]�}���-c�%tk��x98�����ϩb�=5#h�}��5��Mw�{(�
�D�I�E�}��B)�����աԆ�Grh{�Z�}�j�5�]� \?PT��0��l���4��L��'۽<b(~̇u̇��4Ѯ�1ya�s�$�䮷5R�}L[4�Y��du]�u}�d�7I�L#�RJ\�G����E|�rO�Q�_v
X�%����[B�p_�>�s��iź#�F�O�g�	��?�r^R�c�z�D�P�V�Wu�@�g��?��*P�J)�a(:wK�ym�(��뻫4���h�[�@_�xi��Ý� �$�Ǒ��k	�8�3�@�C���U?j�7�E����^��L�D{��(IGE�C�I��a7WJ4O~��t��bǛ;��wv_-���4��\��`�ݖ�:Te�g����sM�'	�'2M B=�mm��M*��iӫ^/��:��o�*���~��n��5;�,�Ck1_kS:	�[*��dh��g��`Ó�GV�X�\ �<�E|F�j�P5[�ƅh`�4��$;↡�L$�,S;��Oӕ��v���������j�n���L��i�7����\����l�8s�p����N:��Ǐ����N:��q@��� c�k{�ۛt�����n���%(k|[jW=�p)PVۮ���)���1�I0�;�'O��g���Ps\��i�{ ���vA?���$%+�s��/ׁv�G�:����o���W��u�V�����#�u��T���^ג7��c<ApbC�	���w��*hD v�Ӂeړ|�}�,�:��\y_����В*av�dA*[�Pr ��CZ�*��D��������s3z��-��I ���.sA�g0���"��T����<7��GOғ�Z��Ez��T�ڽ` H�G���Z�Q�r	@eb�U����Շ*Or����:�kϕT%loZ��(n�1�9v=�hp�K���&�=�(Ў�����.�_�B"���^ �T�����KByk	�t����	��,}Q�lW���y�\� �G�,/π]��g�U����>���٠u�����s�N�.�V������}νa�Z�<6�{���PcI|�{�gIp�1��@�~0��m�G��pV) ֮�EВ.	siڲ*S%]��e�  ���6t���X�!�
�����\Yu	��p��[�\{0(p�E�a�O�u̮�A+�Mg�X�N�+bKB-�Z��x%1� ��u���l�:d�sU�M���l��)b��Y���G�U?	z�u{�/�ޛ���i���b�7vN�������N�nbӔ.�J����R�zsM�&�[��n����@)z��ł�b����2|��}�XZW�;!T{�[��������7H9{��C�oU�R.�F%�y�����?t�h�Pˢ�̿�ʐfl|����ȃ�����Ӝs`���W>�Y��,�b>�s̴�J3n��������V�޺έ�7�5��nʴ;�]˸?�J��'O���g�����trb�ww���Y��Ƨ˔nI|��7��o��ާ��m ��ve�W��~0��?ÿta�lm��X9��^w�v+6����!-%��z�p*\��B.BϞ?Oϟ�k��LhS�?F	q��� $ ��bm��d��)2H��Yɫ�LQ6��A�E�Cm\ܕ�|��勶)UWOM��
����*�'���K�{�]�~i�KjQJV���}�'U1��Xo�æ�J��~��4�,Ɩ�e_d����ڒ�8T�8�qjZ/�
����nE�V./�ߨ��]��V%�)��GO��_|�I:==��L��S�nو�D����V�"F��>��j�N�z���B��;�X% ��)�ñ���[F���Mݼ���GV1"�����tu}&�D�a*��A����)��Y�ME�:Q��g� �'�E a�)��b�������wlc ��L�h#�d�mT��on��V4ma�%K�Ğ�u�K��̘CiD@JKHI���g�X򩃨��2�qR���B����
�0��K�4k6gȉJ,�DE��Ų�JI�*���%�:p��ܘF�J�*7�3Way~��+��{�����k��
���ƍ��ʲ�k��-uJKɫr�YвtV�s�x���(zT�	��.q�dJ���N3'>Flt,j��w�i��N���g��$m��̂�)�l+f�^���
݇-�;;�vGv��5���F�&��X@�F����L�=�$B�y%�69�i�����2�2�ʹ����˿I;���������~i��A�zѷEdpPl%�I�h{O���G���O�Ԥx�U١p�X�E �F�ߠ�����B�Ꝧ�u������,�*�o��Vsi?k�b�`�0�>z��]^�0�^�`Ti�'�*�U��cʓ�sZ�G����p"�vc��e�����1Xϵ(S� Hc��ާ�����Hc����8}��qz�ᓴ�o7}g�vwhu�!�������6]��H/�y����Ez��,]_ݥ��*ݭ <VCz��J��~lTD�a�,���=N{V��X�-4"�����o�w��"�	�aZ�;�⏂�Z��M�P���h�G��Q�<H�Y(ì@��-�ni�'W�s�t��N� ��@Σ.vz|��?R��T6�#
:h�P����P-<��@�ݿ=�'���,�f6�8Q2���
8�BX���ǳ���! h4V�n�#H'))� U3R�ן�E����s�:�#Xռ�Ls�Y�x��R���3�eqOmQ�l�v۲����v<U�ϕʉ�;߻��쀾�I���{�s��>ɲ��7Լ�n�:������)�󃎠X����߽t	YP���qO�� &��^��+����"ߏ�V%�4G {;e6.7�#iqn�Pcֆ�t�+��5�Me{�n���)f�'@�RuUd�X�i�]9-M�8���C�V�w�nOr|�J����wI쀖H-%���L�:�Jn?Q�y��*NeH���'�����T9?\3���'�'\Ԛ�w��`�Y�9-�JLpk
�6��6�� n�֚K)�5g%P-�ܪC\H]�Bҟ�FB������{��S��Q�f�+OX]RB'�6<�֪7v�V�R�j}��/Ա�-�؁?p]�(�,纂�`ܳ��wPET -�0�4�KO�D�n܇{��Q��|�n�lO��vV`0�o�e�-ڪ�z�(���I]�6:0�ҫo����L9m���b�:�E[����m�0��ߤ������f��חgi��e��hV%g���J�eɳ�. ����ٞ�}�X���Tvw��l�#)������\�I*M=  o��8�
�C��NyH.����9�m�!l����q�_�4��
%	���G���.o5��]˖ТIb�?� �m��!�gt3�;�O�;A��R�Y۵�[Bp��<���Mz�������[Kn�`�(T�2D�����q9�T(iac�ǅ�m�׷w�u�n��R4Slҫ��t}~�n���ZO��Z������9��3�������_V�ILe!����½sMy8��8���f��&Fm*)4e]�AF���;>:N?�P3P�͗�W⌓���>�̺'�L#�}�k������������Gif����&}��;mzYY������U��
�O/�}9(4�/�����R�nk������L�����j��Uֿ�"ñt�����JN�LT6`!-����[�a.��,����+o��V��3s=��m�nN�6>Y=�'��ڽ~H ��F(i�;+q�/N��(Wj�r �
�q�� A��w�	E4�ǥ��� n�����Us�Z�3-�W�Mx�+N����eWiI;���{W�xru6��!�0�D�U��1ʮ�[��tjgM@CO�ˠʥ�[��k��r���6����D�N[Y��i��P�x��{��_��?E�%�=�wh���HL���j�#/�c�;O���u!{ۨe��s��~�9��.� �E穊R8�V�	�<��N���_T��.#y�<P�5^�Q-�(�b�k��޽��[�=R������+ݖ�^�fL�#�]�V�DYE�Y�wO��W���[��Ϟ�>�����Ox�� ��Q����"�/�R��ǇGB�Z����s�� T���b���]��& ��{���+�;�.&�7E��C�C���2�^ڱ�x~�,���Q�L��흃<�'kӐ	z��΂�D���+���v�Owd�.�%|O�N��vP^۟7	ۄ�q�*�])͜<�
k{�z㾂o�j���wo�������cz��K�~�Ց^A��;�vq��� �:�Cvu|=}��*�qٵ���*P������̪��t��>��=����t���ٵ}��)����U�Ӆ��v0��ּ� L]��g5Ңn�/��'�0T<P%u47� � �Ȃ0V�|!5	{�z�B�*{r�v��
�$`O���?���G�}�6����7�_��i~�M���!�OCO������%�� �B k&g���f���/�j�z��8�;�:��[G�r�<� dV_�N���~`�����B��v���f݁bR�r�:f�{|t�����A�"[h����Ks��f�Ve�mˋ�!ߛ,���w�����R��p4�*�v�Y���P�Ď�ġ�<@��9�*~+w����$��ȓB�܀���"悅������HJd�!9TG����+G_OEXe�o��J�U�;�Uц���"�;��E˝u��0#�v��`Y�_^*P�	A�NG���4!��d��Hb2Xͥ|��:4�$d�;~B�V~]S�/A�}Ѯ>0�h"�1w�"��,ٛ�i���ѯh2�?f�J��_/ј�[IIYv�;V�-R��֓G�4Vʞkĸq˪�a��d{���<�+��P�eu�^��v�2�.��q�2�3傁����=�-T6{��9��'Y�)Λ���b�w�_?ZWM�S�0�1KfӴ��Պ���)��g��>�Ԫ�;�N[��	�X8/�Ѹn$�ѵ��ܫ'�G�RES��t���ic�מoa��qa��mZ,dT�B�G��}�Ɯl�s3w��ݾ���-�
9�Xv��hs�{;��Z�aZ���-��H�����% �A��������x7=~r�,Ck)�JN�!-�߽}�ξ�!���������j��.��o��&agW�r�؇W�� �V�7�����s ٷ�\®��H�%z o��Y�������*o*�T�v��.n���~����>88I�<Q[��7J���;���y�*]Mo�B�P��z$���U��Ъ�:d�b�EX|i�遮�^�Z���S���m�h�,-8IN18߹E%n1�J�n'�G���>d�|p��B�d'��H�
)2���Fy�o�?<8���`{W�
�5��Nn�_::U+JS(�}��ג�$�l�F�6�����!���j�g�Yv�u8���&�W�g�SNT�<ߩ�����x���Ik�c�G�� �j��C�a��u�ܶv��B���#��������~��4��YwJ] S�g�^����~/��$'%J��(C)�籬)��s͏���sDɸ��r��z��!�~큫߳R�?t�6�#��:yW�����&�qG���� m� ���=��W�z����`�͸wK�����?���)����Q����^��u��R��q�B�~kԵ{ݏ����tM:>�F<�46)(���޸D�TH�%]��{*�Q��et5K�����:��I��q)at�Zd�cB�d�?w�J{m�24?������Ǔ�%�=;����Kk[w���Xܮ+�L��;*��~�?�G]B�k ��:�9� ���B��b�3���W��Rf���?+/Z;�����$��U��2�Y�ju���!AK�9+��#����� |���A��V&%ZKO�ע���V�">�Y� �Z����$�]�8�u
�'�L�Rƿ^I��v�݇ZJ\�,�P��*lՂ&�Z�ʅ�ygϽ����ݭ�U*�n��0��K�Тc��i�݋�������^�����;{}��F{�9��`+ 	��m��h��]܄j����0�K4v?�:�Mg�Zoդ�RϦ+{�UsJ+p����j�>?}����_�FA(����G���Gi��ߥo�����oP�cJ[(x�~f���d�3`.D���iA���ޤG�,��{2�h����1efUe�Y�fsC������pC�pA�h W�^pI�$��:�YY�{�ln���"�߹��ZdsQ@�&,���LU��{w<��lx6UPֱ�)��v,�ەӕ�h�6����9��c���j��*�V��zED�K�Q#^8�;���������G�/���38w8��wG�*��2�@lvZH;�2�O�?I�N��T��4�����N-�3��.�%{����T!ݷ��,F���%�"�C�b{��@���u���ۃ#��{G����^/_�F�It�;v�f�6t��:1�o�h�YZ5���w6���3q~�B "�9����=Pթ�H�b\�����=�J}�u8c���֜dC)#ܫ#sK��	=�����x+wu�,�:��{�y	9�v�b�h��W��Y4~"JЍs��r;: >),E�W�J�s�����}��=ʙ��ߺR�N�n88��ө�:���OH�O�YV0#�c&;�S�ϕ���Y*9�&�u-!�^ �n�a[2p��;�P��C���b��|�׮�im$z�/��W�e��n���.�)����-~EJ�_xe
GhpI�Z@����tbw9ǩ�����Au�i�#�Җ+a�XƑ�7r���`o(��z���hTi�w�n�u,��� �����
w��+�j����(�UZi\na���H���4��������YN�,zӪ�_1�d�rP�!l՟�$%��W*�8��Q, ��d�8̑��(A4�+�E�l��rn?kN�|��R[s��+�������Ekc(01h"(��1��\^�H��T����Pg���.}�IK�llӖ���\�ڜ�NZ�{��x͡Y6�%��@@�t3QY���<���������}�:]�]�f�C����l���2H���U+!�5��ި'��^��7�@`v1׈}��f P�do��'���č�r�vۥ��`�l?����7_�E��Ͼ��n_�2�у#��k�YJ�� �ױ]�t�7��_�Ȓ�����Q.�]s��wD<��}�3Ƒ���`$)U��ɂ���Q<��R�؞=s�̐;�pٕ����\b�kC��֥��\آ��/�2���̡��9�Е�pXu�Qd0��uA$c�5��y���H=i��[�
u���`��Tzb��YPJ��pj���+�*��6[�M�^�XuBtw�<�|k�u߲�	��yܘE��e�ʘq�� �!��x0��Z�A��!=�ss}s�F���)I�#�������f^���#�-�ѢI�=���mV,i��
���:�C�ȓ���G����ޭ���pN�R�S��!:O�*@���g0Ҵ*��Pu�:�65�.ef7�Ugx3/7Z�p[k\Ezȕ�|��J���s!,~�R0k�4Hv�����FN�3��c�R外���^�
�{�x�=z�>y�Dr��O���:�i�5�^k�b+�.���db�0�����(�K�,z�Y}�(�$]n+��t=r����c�˘�Ȝ�1��d�:�~nk��#5+�fT#69��=WB?��2�ҁ��%y&� ���`v�fa�"�J[�"6l�"����:�Yt@�"�`Ϊ�͂�g�{��j�ivS{��q�;������ݼ_\��eIK���&F��ʀ[��B�gY`�n�Eg,}>"F��Y~�`wY81A)�q���91��v�Y\�wu�^Yƹ���eh�K���:]L�͹oҞE�=�}�<c��aPyz�@�f�w9XC��{i#'�_�&��������3�Ŭ�!��,h�*�4���&���1���+��('������Ʌe�ש�n����?	tun�py������a:����݃��*9a���|�N>�j�^\�(���6�玕%Å�j�v��6���	��~�o��_|�E������
z8�B!�QB��/-c��ߘS�_�����7�G��ѫ���+饁���zAK�B�Ly�`gOz�d�88 W ߠ��A�����1��#'�`�$#9�{c�6��20Sz�E�$ ��a ��Q��g�#o0[Y��	�ʌ�(QR�n��L)����je���F��F���5pg&]jx���=��se����2�"��M��#C"JE=t���}��V., �{T���۞%���j)��� �"���]��Bp��d}s���_�_��W��.;�D��9@�q5�l|F�B���Sy��F�zN:��٩4^΅��n^���-�C0Ȑ[��[�@�h���6�\����\�y�=;U@4/*ȏ��r#3�TP��?N�8Ȃ�w��G�̎dR��ŉ���N`���#�gW�H,���W�]�Y�]�q�C�e�í`��:��az �����j5��̮���6�P�2�c�p2w�鹂P�ш��X�W�=k�F�*},d�e���:����ή�C����-�{�ZI�ĥ�(T���un��?��@w�9�u��d{�%0���&�6����V��Tu��;c���?h=<иӮ����Ƕs�x?��ck���'��,'��sps���������(�(���J�ήn�2�3�c W󵢡Z���ڸ�U+�vᚥ=���-��ۢ�-������=P_�>\s���A�ަd��60�@��6õo&��G���=��k�A��z�3�T�����{���O-s@ǗL��+�f�&�o�� IZ�K�\]Y�l_�ʠ@\�:w�{�G������!�`T�C����J$�m�`lRO�6�M�?����K1wM��ZIͩ��cF bq���o�A:^zI0�Dṵ�3����_�_��eV��/�Od�eїS�@F�ϟ<S����Ԝ��H�kXpڶ-�(d"Z�Vr�1������JV��|@9��2���`����\�Dׁ��u����L��� 0B��L�h"�1h:K�'������ZUz���1'ȿS2�y6@��鸝
Pد��0Ӡ�cx�o�罼ް�/g��$Ve����P�q#.�<�M��`)T=�L��]�&!r��u�م\Uv���:�Rpm�;Zʙh>���
�E�\
fv]dՏ?y"L��_wFi���pz�����P��}[�t2"g����}��9��:��n旑�]f}r͒���*V�p$�T]> @bTs��"$S��n2 +�7�4�Y���g�j���������~���{y�z����V&�����؞6ݙh�M��#�ء�۾�>���Q�>�ǟY�G��:�n ����y������(1:'��=�=e�Ͷ'��/U�Ы��M���ߖ?<uY��)*�� �Q�N�	G;�o�|V�3�f�6�L5�uoV�#y=�3�;�%ߙϢ#���h[<����%.S����`+��I[�+��o7����~�4���gN��M��Ʉ-�]�WgkJo@. �y��m�2�#��f�tܒiNS=Y$�S�f�ƃqj7�D��8\'8���G�r�D��O������ˆO�D@�<�Qې��Pj��?����?6���Q�5ú�zWo�s�J��8���-��&'��ۓt{r���4
%���9�f�E��$��3�}�s��w 7􃴇&�9c@N���X��6��Ӟ�O��"=}�Lt�cʓ�4��:_N՟�4����3�f����w`�P�+R
:�BzUNi�X{�@v�|�<z����/��O�I��/��;�qݤ���HЇ�:����&}�٧�����U�?�����\� i9����� �@RP_�Ҟ����s��sk��GeS�����J�d����M��p�=�� ܨj����Q���U�ә�tc�1�v@�� w+����,]|<M_��b'[�3A @迠�C{xx G24�F������=9���ҋ��0;��R�E���x�}��R�ɢ�~�T�B����/͙}�씹o�=%g�$���=�p}��s��~������[��1z��R�
��x��22�A'v�g�������/��n1M��h[�������1h��t�߽�^U�O?�,�v�Ƈtg<��=�0	CI�Y���ن .��nׅ3��<V�u�*~d,	���;tF���δv�R!�E*nϾV@[�U�@T�8�&H,�,���0�A�с��]���{�|߲8exH�I!h�}L��8a��[{���*�����y��o�ԋi�Θ�k�	PT&�\�snA��zV�^6`O���͔��]=��3N�,9B��./��}�M��g��lӶ��_[E�qG��(�����tG��x�ۘ:�X~V�L/��H���
����ގ�,f
�q�s���߱h1��
�P8�6��w�J9^���%���*x{�S9�̽�>���Ev�W�� �-F�J�M�0�-`��bҝQ��S�����(f�Q�^��U5�Lز/����P;ˀ���ض���C�Y�^��P��͏r3��%�ҙL�����(���\-�)\O������?L��7����9��s#F�a=4�����B�W�Frp�y�J�\x��0}��ߧw/_�����{�C������f����`�}*�lc�j\�39���(���V��d�1�/�?M�|�<� �;L}?"�l��σG��N�w߽M�~�6��BQ���Ŏ��_B���`Ha�Y	�j�(��s���������e�8h� �ߗ�tJ�ܬ�eM�ѯ�RF�~x�V�7�	u�n�09�ѡ�8բ�ꊌ�t�z2w�^d�d\�F1vq��QpZ��8�e��Hy�G��}�wЙ��B�qm��v�a���FY�b���23} ci�����8�7��H��Yn��������>��g��知g�?p�}
�3�� �NP�8fڼћ�,J˂*��3S���7_�����w/_�j��w�����B˕���˟=��㥴9G`9���/m��������޾9����Ϟ���Ŝ����c��O�=M��_��n'm�� �,a߲@( a!��C��5��>v�\͎Wv�(k�Dx�H\@2dbA���:eИD��w�`�Q &�WϳDZT�A�T�6!�P�xI�E��o��>�Nﲽ3Ǜ%T3�1���~UT;�$� +��S�K�4/��t��/^�y\Ɂd���_oS���@�:�	y=��P~ݭdgݍ5�M׵;�����$"ɒ���&;hi7�K魢�vX�V����>�']f{�A��u�����9r��2@W)E�7eA�����#Ӎ����]��*?.?gg|7K��^�~6��ν�u��.���Ẏ�4��}��@��� �ٹ�&ŝ璱U ���^��&�	���W�۞E~#�o���|`/1':�k������ߛ��)�j�}Jon�RO&��eN����(G�y'$
9 ��@��̵&}N��fuo����>X�y+Y@z��dlv3�k�R�,���辄O*Csb��ߧ��^��o�.����t��+�Ɣ9g�"t�v/xE!�چ_�x7Ʀmz��K۰��)w��ݵ�~��Qڻ�>���ز���C���]\���o���,�}''���*��#`?�sCq�z��Ԑ\�	.����Q ����<�໎�n,��x�6��w}��P��	ӿ�숳E�͹��"��/�p�sdk�Oo�W4!�%��s h��䥡6��E�:��	�|Y��*��*��ld ��什�]����Z�r����������Azo����e����p�v �s8�6#"U�� �o��ݍp(̦3e�#�p(ہ:�������!��ߎv�bWs��@�j�q�ފ��1�dǰ`���:ؗ����Ǵ0G����SϜ���G�,7Ǩl%�Ѯ�@>������ڲ�����=%��ʊ���X��A�y	nj�׭>�r��A�I[3�GHl3��
y�ɬvn��Ց��k��e\���E&�	܌���y�VKw��#�SdbYW�
�2N� ,Ix})2������I��d3}�����d�,a�~<��j�e�f+3��R�?+'���u��|�L8o�Y�u��b
k�߳U8ɞ�UE{E�FD����&2a�j"�,���v�����vn==g�?e�)���(��k���<=����������Gi`�c���3)�/<}���)%�Z�����x�l�~��6��,����|>�u�]��JHTeo�_�\����|v�iL�E�}L�,�pIU���"`��9z�Zpg����F��ʹ����Y��L,SǇ�_��������QZ,no';��� զ�;ܵhg�2���1�lf�m�j�S�uEGS�b�*����;3�1�N�����d�2e[��q��pm̠�xc�fc�g�6Fo���y�0��X�8y�!��?H�ތ̻�o��������1?�{/ɿA[k�6�}K�ϭ��5��ڌs΄��p@4�轶�6t<�'�?KO��4�{|����-C�Ӧ�}y���}H_���O�����?|��/�0�#{���`�@QWޮ�!�Lrf���c���G�=w��aA�A�������͑�$����޷l�7�7��g�,����Mzp�a���ӕ��Uy��,` ���ʓ�3h�1�M��E��V�+n�/�2�ABw�� �>%��]�Ke�q2�#ڱ=Bf��w����B�N>x�������a���,�Ҝ+��0�H%)9�@�O�\�@
#�~e��7��,��N���;rm�j��fD	�_P�R*�C�.;��|���h��Uz�.y�F�kƟjG��]_	�Μ�ۗ����yz����Am��u!HR�I�T>�5��W )��B����s�`�]^��oΜ3{B� w���K���S��H�����S{&'u�j�\u�"ƋJO�6?����-�T.G�=�����Z&eE��,-og
��JW�����(q�s�(S��X퐯w@Q)uWAu���r���5�ke��w�F���]V���g��.�R&��&3��e6�����yvZ[��*�6��y_֑�>�U�l�ȩYC,���n<X�F{#�,2P�������T�o�����c����jS�����ҥ ��=��{��&���	ב���V����+�N!I%!m�n-�w���$�c��\�|L���D�����_w�#�|Ǹ�Ֆ���{��r��*��❞}G&��Joi����r�9�ۘm~��z�&�{E�Yi�*��$ݮ
�ؑ��JQ-�5?(~|���!��^C$`���t)�Z�(e��ŹJ�{v�����4[ߤj5�e��V\�-ЕeM�������ٰ��������ͫ�ތ����e�� <�To�,��8��D��$S�����Q�����/����>J�����^�`5B���im������|�Cz��1u��4��-��o̱��=�ü�hkǲ���x=I@e4wv���ޡ2��7L7�O�!���h_i�	��JB0NQRCp���؜ N�ܥ�g�����������ܞ3�bGi<Ļ+�-�WuN��2����tߜ&���i�{�ae����/,AB�"�<J�Q�����^��S��������R�̮3}Q,�>2'[y��ޣE�q���H�5Hz��k{��=��]{^0�h��L��Ҳ���D9�A79J�ߩ��$k�w^z6E�E;d�X�p��(�����*2��ߦwoމ�_�=c�i2+@gD�c2yw���p�\W���?y�>y��2�t��D"��L��2�~ y,S4}�`�W��gz�ひb�E�S�� O��nA
��֌~��J�0�������xw?=~�XY{K�Μ0*g�{�	�n�l��}�ֶ^��s�ṂSZ�k8#�˨)T�Yh��3�fˊE��j��Yz/K�4�_�S�ց�`�5P_�>=�O��I���3�3���N�������lb�H�H�=t֭ �i<��ћ�H��g��'VB {T:�L��M�fF��A�*,Q�i}�ׯ����3�*��"i{C��m0L�0J��u<HR(#��]�X5I�X� '{��� ����8��Ɓa������c_*�r?�^�'gm7[6A�g��G@$9�z�T� ������u��Ѩ���0�m2�Z|wZ~��۱y��O��?�	_��y�&�]%�s�;�v;�gp?z� q �, !A1� J(M�5���62���0;fF���=�i�D�ٹTfv��=�,f�>���Ň�Ԙ1����7� ��E���޲�w����$]]���	J�M��@[��v�/���qh�`�1���j���/��/�����Gi|o��I8_���w���"]�=M�^���ٛS��EfBy�Nxa_��q��C��i�df���!�����>�3'���f��R���<8�N�#jI���d��Q��z����g�ʈ98ȽQ���u��_�Helk�lSdP�C�YC��Q%��4�d����?=hթ��_�O���>cT}���=|�����W��,�##��6ٜ�|���\*O2����3�����%{��kʾ/%-i{���������� kȖm��	�%m��Rv�{_{Y��Ih
1p�.wIɻ��G\[�yn�:ҷ��]4�5����5eT����J���]Y��r��!��@��f����ˆ�1#N���+9�j�&6��)���T>ND0�`:JL �v��m��y�՛���`�jNT�(�3����\m�c�k��?zdϫ�X�k�g�{d.�o�ԂG���@���FT E�؊�-l�r��<��Ѿj����F2�nP32���lcT"@I�,h�YP�`](�C���֕kW+���i�r�9�s��؜�v�)���رu���-"�
��H��G èGۉ��@?����z�����܄`B�U���y�L������5΁h%T c]��ށ�s�n;����K`��ޡ�0 	}��.E����.�({�`HkM��<�xi��!i�B��z�>�Ys��&�7�?��a��wC֟<+�Řʨ˪��y`{y�~����V.��|1/A�B,?�\�Ҟer���,��1/�ke���C��B=�u��gXDLj����Ԩ�D�?q�>HJfȉHS�:�������w���O��0�ڳ<c���<���2�����\�^��7��,�e]ƨ� �w+�
������'��˿�E��/>O����TZ����#�-㞟���7'�������ߧ�녜o���j�~nO�G�L&���޸/�0���K��vB;�TF�Ӥ쿼��L��ft��0�m���S�c."�p0ZƔ,?|<Q�����F}�woߊ|��+jQh"�1�3{��B��2FU4oG:J���@��� nG{�*%b����g��w���Rs����2��A��^?R9GM���p�W*Je`���?:<�SB�=�\"F�4�,���ýc�B(���������C�XɱҧjD�����S�R,��Sgn\f����^�E�UY[-{��`�(]�5ã͜��Ѯ>���[����U�����d"�����W�o��G�X�y��F�P�{��@��E��3�d!XOw8=�*i��g�e�c�q���7|�M[�ȱt +�`KMI���ɳ���C[ӕ��6�q�	_�~�����|(�-�����b��K�O�����yn��1���W�)5��*Xk�{�U4��) n���O�.��`��
 *�#���3O��G��lJ��D���\9%c�yc���5")i�� i[�|9�Z�{��|�]Y�x^&��{�&�5��TT�v�@I[���e��.Dq��7\T!�w�	�GY��{����ܗ���%~+4� �Ψ��̾߬T-�K	�_wG�2S������1��f��ߗ����3n�y�q|Y*_�,؇���Er�A�r�� �?�wOHֻi��<N���M��I���D��N��p��-���"�
��G?�008!vw��rN�B�!?� �(#�*#U�͔��̘����^LJg�ަڌ��2O�`�Z��g����2*�_ͮ]�X��}ў��]�06�`P�5��ož��7�LF��{���{��O��_<�L}��4��_yY����,��y�����Y��1�ϧ��]X�b�6�lوx�`��Pn[/E�0��()l����H{o(4/���?�"��T!���gfP8��¨�ތI����~��B�.So�T����ZH^;�Hg��,'�9���}�7�x\yn�G��ɵ��nb�BQ�ʥzÈo|��H��uH��/�*������gi�������i��,ҫ�o���˗/�?��.-C����R�27�X�g4�u!F$������@ٚJsW��9�ɍ�@�7d�YW�ݛ�K��)�4������@c��Ӷ�~�P�(I
��(��r�C���1Y�d�N�9�z�e��}0[\z����(�g"V�r��*�[�K��)�q�L�,����A�`��`f�B �/p�=�^�g��p��fJ��d��0��c����B�۩�Sš��^����o�Np�G� ��y`�5l�\25X�����,@AT���L��z��m �ե$�xǑ�џ�]f5*�뺺#n���<g}Ĉ߃GilAc��/0���x/�AY@���B��J%��v���l۔�zD��
vr�ڻ��k���W����_9I���;�
��ĳ	��7�2n=����4�6����=PzI<�U�i�sR�F�:s»#�}im
e�U���n��6ۏ�K�	�}o�H���X�&S{z�
}W����rzݱ�I�������[�y+�� �9�{h����i�\?ϝ�-R��L��Fޜ �-=4(6}�C���O��x�v����-ǌ�1�i� v,����-�ihv�vE��Έ�S3֫t���As1s4������զ���X6�Z���p�˛˫4�����Ej�.�ʾ��ޘac���ReE@c��Xfu�N,>��Q�SU
���ϐq`9��'=$������	R��kS�3`�,����`3G69o��e�˙6,h؋w'iI���is3O�t�vʑʑ"ఏ���(�R���'BG1�
1܋��\m�F��Zu=�wf;�����aDA=E3gvoQ(],"G�d�d��[�?X��9��b��/�����E��쉭�N {VB�沨k62,�Ԇ���2����]�}��"����W��5|pd���в�&���7��7�4:��/<ϽC]?�ۼ���Ȭ�*��Md�^�?� ��������̐b
�h��LԦ��rcY(��
A	�fl�a8i��L�o2�y^�f !D�@J�h�����֣򠃒i�ڌM�c�ږ��:�i5����R� ��e�R)� ��R{n��N&�����^����F>�e_ � ^QQ�u��i�^�w��*h�ch�|�>� R�h
�+=w~ґRlQe�F��֜�R��[��m}A��1Me�`����Rlq�L��|nA��#7�5� 8ۏ������]1Epz�f�E�	=�s�����:�Z�{��]ẽk�ft��c�qIo)��i>�5�ʤ���8���ޞb"u�o��ƙ�؋Ȭ���uJ.�[٧�H�rK���W�B���Ȯh��:�P쇭���%e���;	�vo����c\��~�2�=#��[���W���(�J*�o\������1L+�l�s��6�Қ����@K ��U���3j��J\mZ;	tl���5U��|�*��K{F�0G�ts�(���q7�������)7�Ғ�s��^����$�=�#K�S��N.�zT�\��q'�6�A>��o{1u�R�l��yz�kt���#� c�:��"��f�ʅ����hpc�B��D�j�W�h��Q�����?�w�S�p�Y� S/�G��ۃ��/	�Y������ߧ3s�g���q�v��F��?8�x�� �%CS(+j{�����^����~��_#k���Jeę9Cp9[�G;H#����1�8�a�m.8]/o@���E�v�0�8�#s���ӓ��c����i:?��4��sp%4�0 2es�Hy��f���7f07�o�eK���Js������^!��7�k�b1fQ���v8+����B�P���ze��c�o���}���WZ����Wi��q��Н�\�o�	�!`M���$���[}�� �'�HI탵��&V1��|��CFx%�z�irq%�-�a5��k�N,0������ ����I ���kϨUwtmG�FV��&D;c�Si���3KE�#C����E	���hRj$���{�8i���̛�;�@�{y�T�����A��g<*P��5�C�akެ�:m�z+������Z����;ʆ]z/&b�H3�u#�[�eY�߻2�R,z��^_�	�����E�;JQlp`$9X�v{{��~��Zi*  J���%��ҏ2a��lT���2�(-�E&�*��V��C
�}�z�},�W�cTT12w����u��w=#�q�r�һ8�c,'g�9P�Ylv�~}���/�Y�+���̝��28������\/�M�$KZ��H�@�y�S��;1�5]0�~h��������l�+Wi��S;a�
�`�����5ќx�(�����jiY�w`�L�gA)����v�.H�Ђ�~^z֨]�h�%�&M��^���!�5TB�
���q�<2��b�2C�i�?O&l�@���|G� �-FA��X�3����P����kQu�n��5E��,�?*��)p���S����)OU�3|5m\3@��\]\j��/�M�ӌ$�B�V�έ]�'M^���7X:�g��"&ߌ3��������]��5w�wl\���,�E�Cѥy��L뚬#O	�2�'�~�������r��A�oN�($g��tbY�(O�������_�4D��o���DiӜ[9<�-&�"q\��:��Fpy�f�qfp�#Q }��� d�N*sJ��m��>L���U�r�f������'m���2����ؽ�ꅞ�ei�?h���9��@g�T-�Y�x�J�{n����R���cS9��:�`8��Y�a�.�\ Dq�������3��cϓ'Od`nfv��t��W�e�T�j|6W=��L;�0h�֝�TU�L�e� ���3�&�]�M���ɝV٣g;����#{�YQ�ӵ�8LՍ}qH[�H���Rg�φ�#\�NU�Z�f�(Ȭ�]JF��"H��z�	P�@in�9��;9kRѺ!%�)����}@VQ�	�c��]8ӏz���2z���ص�_��~�e��!;��m��w�ɯ�iSV ���'�j��"o��1˞�1����u ��CA.QYU���:�h/D.\a�����O:�q-=��W���*f��]���[ם]l���,<��FW���G�	�Jr�+'SaT�{���J��P��hX{�q��j��7���k-�BZ��X�-P �Vߣ���G�2��M[ �Nn�;��
���4�7҈�d�Y��3z�c�OO�ʜ�e�δ�����fKҭ�'�l�u�Ӯ�w��*�>$A�~�M�j׃��6�?�%���';���m�������զbјIÙR��7��0���m��S�rdX�攭��}.��#��E�f�0���ƃ�RP�k(�Z<��d��j�/'>��׭eXҿ�6(]�p���o�u�)SW��{P������+�]g+�`[40'SQ`���v�!��4��g��P�-(�0eYu�`GD�{�����ã���ͫ�Z��\ڈ8 �y��Mz����e���jz$�&� �wx�q\d�d�+	�\G�:�^FP^����,O�D�{'��,�q�4���V�@^�stg�v�)�;�0�]��g�K�g���2�����0S�@2�����r�����u(��ɬ�d,7�d�`�����zJ1�K(Bb �&�A��Ԛ�'ѻ� �&���W�]��=��{G�zD�����U���p��s̍_]��?��Ho�H��:,\��@ H����2�|s���sm2t?��2������\_=���<��q��@�A��>�1�l^OՄ��J=O���,�Ly,$2���9������;�^��=��юO#���̄=�x	7����P��a�1�Z�~�[g�����U��S#��c{y];0���Ν�]����kd]���펆�ݞ���ы�r�v��w7�7�9��6C�R}���	��n�
gr�E:�^!Ѽ�]��-�@=��y��1n�ݺI�0?���@>lK-�1o_�����@(��y�{*7��f�c\GZ��>�.�X*J��⬦�I���\��\2�.?�ai)�I��3f61�m_�>J?r4����������l�4��s�l��2k�7N�hWm�VcmI�ە��x&�E��E�,_ܸ�K-�ɦ2��lv13s��*\�Y�������	k1�%,O'Z�e0��϶N{0D�a�ƍxXUV+f閞�4�E�,6�GDt�E��i41ԾR�k��l#�E3�϶υ_��O0��Bt�(�ƙVF�>�[S>�(��Ԛ,��ӏM�A�`WѦ�:!:}�
z86���-�UKQq2��=0c~`��
"f�J9�i�\��$���~�i��?����>O���a��M.��lj*]^��������ߦ߿J/~x�&�˾9[Ѕi|pd���J��;)�3�������ԉD,R�Ӻ�/@��'�)�{����0���i�#��T�x������i< Xcrd��n>�}L��\��+��\�4*��s���P��U9ej�ڜ��z�^��N�Ҕ�#b��V��՗
���2�/��o�j�.�-�����"~�����2$���g�8g�)KЅ�N��-��Ǵb� ԙ���������O�9Л#�؀����Sm�!#0*��4��2I��Lԙ� �!��v���rN�Y+0#��!����웲��Ⱦe�%��P�3T�̋�v	ə���	��ҾZU*�J�t�P8[��m��CƧv>���W�8]�:>��t��K(���t����l��n��z���W���<�*5�<W^&�Ve�6� ��Tw_[�:)��r�� ���y��(���q4�M�;"J��*��Y�щ7no&�,)B�%�M�x6���6��pK]b���|�`� �2;~t�/t�g�E[���B{*��/��b��oo޹�X �`@�=�q舲=�V;���D����Yd��P��.�3_|�yz��~�rr�ޟ}P��Dan��tA�}ފ��@נ=',���rv�����ղ�)�ބwa��ۮW�5U�N�J�2�]�?���3�h���?,{�~�"Rʤ�v�*�|��(���/�CBi����O�ԽN��G�J�CE)E�JR�5y ��R�P�1��63���2��2�92��q~h���C�ܦ�Zmӑ��&�$��M�?��N^����r����7d��q9��/j�q����� d��+�NO��nz������O���O�ѳ���O���{�.� Jfrq�.ߝ��/ߦ�~�>�>I��f$'" ����Q���{idka'K��)�j�*	v��C���1��bp���g��Xמ�;����]�\`�"���n7�H>���J�����L0��[yu�j��Am�e-��;#M_y�a�.ҥE�(���Y�ZwlE�?�ܦ�16�yiT�����P:��JB��y� ������3���������/5���ǻ�'� �-�f�BOXd�mP
nBUH{�ea� 7k��1����h��R�7�6[*�彆�]��LOGB�����X�8��:�/���)_(���l,=���@�ʌ�ƒz"����y�/��'�gE9W:[��P~�7��]���}[�A� Z��ь����y�WQ�X��!�i;��=�<�l5�+JP ZAa%t9��3/].W�4��L��He$s;�y;Z�˺|1j����^����)�挅���[�gF|��Ld���x|�?�iݕ��p.���k\kl��?��V$9�7�� f��_]�l'm(����LA���A�/f��T4Zz�>g�y�Y�C��%�dբ��pCSt�U�������X��uv�&y>��JH�����!p��b��

Q��FqR��fNՖ��	P�j��F�-Q����K4f��D%��TǋW?(8���o�s6�F{�������\v��T	��Z�T5�"QJ��E I���N82��U(1�p�=ZE ��+O` ,��'ё�H����Y�0�O�S��Um_=J��К"��[u�oEõ���{d͐{� �(Ɂ�%� [��TO�@<��Yb0�� l&����!���U:���-#7*SØD_@���5��{���J�7@ۗ��	���AnX�(��#F>�2zEDd��Ҳ��Qڻw��?��~�4�8>y��O�Eu���ί&���<����޼x�^}�*�{s�&��2��I옑�3ݷM�s�Jˆ���-r��;��yZ� D��@�ͮԂ� �ء��#�-�J�u���j�Ԫ,�A����Z��6�Y]�0=}-��
;]����:m���2ɞYS���%��ɲR����刻�3�*�&��8��hD��]�,����̻�|��aG�W�}��z潭{�8K3rj��y�Re��g�`2�П8ae��8���9!�Z���
�lo|:��-; ��7�h�u�"�$�;�\����R�S�q�d25C��Z�S�5\��qv�[i�2&_e�L0��ٲ=�k�5m�<��u ���8���� � ���)��ѱ�n�����e }s�3�0����}7	Po?y�r:�TJ@��۫�P�z���D�S`���V8�NN�{d�v9�3 �x>Ig�jY�`��:(z=w���O��Q5c<�`�	2z.a����9���~P}��y��3#y���)�b����t��m�����W���� ]���S%�"�]do�nj=��\���\7�3;�<7�U�B�4W�:���V���Ν�{�s6��\��^�X���L���n�����'��t#nX��a�c-��,᪖3Mb��������9-����u�ݠǯɘ,��=�'S�:	�X���XUW��t�����^��2$��,�dS�agT��[�����pz�oɳyrĕ�r�B_B�ƀm��ڴR�
�I����͵�J%d���灢#R��� �o�n��Cx�Ʋ�����wv5bA`/2� ��N�������L�R9�""یY���ޠ��~w��$}��_�g�x�|�IJ�f���e#lZ��S�t���e����?�I�/-�`�n��fwv0���G�y�U�X�e�X\[�O�������'�o��
�>�"���HFKtG���NAV����J�@=xi� l{��z����|�|/c��qg�C ���|a9Z�b��:8d�"Qq>,:��
�Ta
�B�U���1�V�Z�c�%,���gs��Z����}`P~x�.�띦K��!�>%��3�,~����xGG{槔� �u!s��������#��fv�՛E������ջ�ރ���<�Yõ�ѩA�Ч{���e���;N�řZe�1Ⱦ6^&�wpNs6 �L�t�%�I�L�'	}�� }��iKy=���h��R��\��z�D�N�9_�! �\��u65N왰��c2��*0]�	�&�RY����N��a���v�=K.�q��7�{]����x%��1\����;<����].s�~ �� A�Kh�qd�:����ϒ��!�(CC��{B��0[q y]*k�����t�Kh�������΃��K�U4"x�kyw}� �������Tkw¼����۳^Jp�g���i֡�S.���X����y.���"�H�+G���u\˕%�=�[a�s2Џߗg�8Z��a;"sY��[�5�z������m��� ^�A �x���V�虉Of��Z	[�@=��?)�yR������p�<�w/�,�Zϝϗ��xB����0��<���#����1�ѦUͽr�-�*]�z�[E��:�d�{x;Ĕ�F��%�d�p��j]�m�ׯ���H9�/���d��Q1R���!�+2���z	u���q��Ɉ��ね7"�}�$'|���˯>M�}�,=��Y�{l�lZ��,���F,F8ߓ�ߤ�w����v(-5�Z�;i���"�4��2t߲���wvO�[]����j$qp�2�B�7�����.��T�]���]D�9@D5 H1"Wu�؛'�r61g51��j�Q�9�b;�N���3�IK���(˰� +\�4�G�ל!>�֕|���h�,��B�uO#P�L!�t�{� 1��M�L3�g���}"��]�����2$�[g��!��F���M��ץsJI�p��^[u4���񅲉�g��G�_�Wo^w�ګ}�kFL3� a�v�s1��۳ ��O�+��@�*�t��" K |r9�
@�J �0,0��<p��<�м�M��>(s����L	x0D����ܩG����R	�����«KK�L'3m��$�����k������g����$���d�z����/7���,w�������![yӁi�3aGO�I�rds.�V�Q�C�bM�ˮ�犋0��NU���K����֕�f��'?�zVA9*�}Qv�+_�iس��X;_����2}�'ټ��o����q�>���u �̫IPH���=a>G6�>wr����=�_Pf����y��yr^�����uhv���گ��RU�k~U$]M`5��e=`Y�5t:��1>h�si��ū��g�#~ZzUc7z�����ˊ��������;��ή�Z���yw�%�(���8�[7��r<�0��=��*l$�~tC��"���JdV8d�}����cgi��� ̨/��似7|W/cӋY.	) !rp����!�M9���[I������L�|Ak�`���/��U�Ui�B�gl|�u��
V/���x� ;w�ۆ���-6i�V2��c��6|�0}e��g��Ѿ��L)8�R�������ߤ������@�gN�^-���#����M߀�5'|k����k��kttgi�j�p�x	�j�R�Y�<���Ă!X�2 ���l{��R�4P+��H��L)�*�b����^~�e&���!�Pc�<ku2K�O��z��h��N���|d�l�����@�U�	��+Rr���s<�w?�{�(���O��o��C�5`� �U��܎�L��Շf�HQ��R��� �Q��	j>��:�K�	PUF�R�3�K�0�Iլ
Y�RA�h�5�30�1j��6���w����>u>pШ)���Z��������Q�k�H�a̦��h$�t�޻�Ի|�y���(_s�����~�h�N�c�L�e.�{�����A���C����C�`T�v���hI�����ha?e�`�b���Q	�^} �x?��U��
΁����S>�q��;�r�{"J�t����F�QM[h�;X��p����^��]8k�9IaI9�ه��(��x���X���@�U~oG�IAV��Vq��(g��������W�jC6������<��g00���@��f)H��Q�\FQ��j���n�B�h�Mt}�5�:''�Im��������0>����탡�-U ����C�ە��4�X@����g�$X�4�����ɥhpm�){��Ʊ���̯*��˲�ty�O����y�hfvx��,�E�H�\~�F��C���%	9��q��ʔ(�p8镥�����!4�>�x+*��LLTp��4�ۦޚdޒ�M��U:�x��u:}�F%h/����#e_�6����-�o�-ՋbQv�"�v. �;D����!ޞi��BO�=I�}�L>�����N.g:�8�^�H���k�f�ROZǻG�Ҟ9�j� -!��%���<�.��/.��ĳ6��ٚ���i��4h��h��SXj��iˑ�� ��t�G���v5��A��aF.P��=��k��p�UL|έd�2�럒�w�vm������m�a��ؒ���� @ￃ�&��㰐9p�z��R��Q0ƃ8��dxvo]�y+��A�eF+�08PȍB�v����@{3��;#��(S��MLZ�����!���T� ���;�Q(n2efU� 9i�n�c<����O~������S!_SP��4׎���*;a�93�.��-X]��h?Fx��B���n���v+�Wn�Ǉ�.�`�n�L
���#(�@�g�Rld1S.f'��֩;���@D��e�۪ߕ��&u�~$gb�{�2�<�|������U=L�}/Se�S�e6q$�o<�,k���b٬��5���i�W�}�.2`ߴr�ō6�yz��2�rt<�^�x��ظj�� �ϳ�#^�����U�ApL���y>��b.��޹��Gz�j̥���ĝ�>�����Yy�m#u��%��0p�`�������t�UP�EF-��;y�H��*������:�҅0��I��Lv6�
!�yd6������z�_k���V�#�97M���:a��**�uu�]Sf��l�D!B�I@z�������'v�d'l���o���(�G,�f�H��G{�K6%>X�,�^^(�B<���=S'��4�Yo�d좘��c�X_�`�7��"m��|��5/5��D+i��6ҍ��nl#�  �Bgu�P��t�N/.���uIy�������N732�n 5���} 6&M�ADv׮}w�W�cB����̎"�0��A�~��+�9���X&��z̛�ע7�Lw��͐\�}�	�V��%t('{}ט]���
2���DP��Y�I�=S�h�twd�o\�������n����k�E�����,�J8�u�*���3N��	p���4n\�P��r��?fDw�U���O�sL>>��,!��<zO�t�Y*���<|�0��?�O!|��Yb�������e��}@���;"6����v��w�bTnѹ�ep���-wr�Yޓ�a��c���g����i��VxcY±���ɧO;���`�`4Dah��qµv���I�ý�Yi�(�T�2�W����@�^��-�Z%�M̀p�E|>�A�?@>�f2wF=�r\ �/!W�)C��MV%	8�Ֆ�R�7$1�˾���J�� �No4#�,���ѝ%��<�����[�k��)�rL+��.�~��3x��g�0��
�����ێ�t@:{���\f��3~�s^��s����m(ze��~82��2�(@0��)��:�r��Z��\�ЇnCब���c���f�7HE� ����8�h��hd����tC���P��Ɯ�՞�h�s[�e#@���_xk��4l"��@���A��j'n"x�_��E�*�m;�y��RcM����k�ef+b��(���	�Y
��B4M+$���P��cT{ �A��+	W�����$���2��2��>���<�E�X��>���C8���e%��G�Fh���\Ra�����O�d�\�VT�����Zgi�t]�y�I{�9-���Y�x�>M/�EWx��Q:��O�<��2���2�k�.�:  �0|U�?���W沄����<4-w�^D�of���:a2Գ��A֮g��l:�dg� �ӹ6�ph���q�H���6�Ԃ�+s���uz;���0�A	��Y�~(��K�����Y�>['��$UZws���F��e�9��R��ZF�7�Xf�"RTi����#uQչwXJ��ޯS���pu�B��)�=�Q.]�2kP�񴂧��s
��,����ZQs�%ߢ�P2��֨)?~�$����>��3�G4�% q�����F�GU�T��۾��������Hu'{Ɇc13�8F���'�{.�������sp�����`�X ���;R]���qL���q@���cl��O�A=E���l�r�P��8�޾Q�HAX��1^�"H�,9
Z��Hhv[�jWw�B;Gg1�5�T� �f��҈�w��z�Uٕl�O_�8�ܣ��lЕ�y6[!`�p�,*��b*LK|�f�$�^�5�����rr>�*8�W�g��	�A��c�3�
�nɮRY{�t6�w��GjҀ��v��"?O6n[�NF
�Z�pO���l���u���	�M?�]�������L�2e��g�H�I��P�WuZ'�*��Rxߜr8�`����c|�1�=�����3am�iM����xy?��i�.�1c  /����'����/M� E����C<#�Գ������u�O�q�`�;*�����V�A#��a�ߗ���p�:�'7V�Z�a{�?,0�S��<_5��.�Q\�CD���Z����!����ǏB�7v��@��A���8�|�T`=����y~~iQ�sH�阡,8�k�-\]���F�[z����ϐ��Jejܜ#`����˾#W1{鈾T
�|�F|!>�R$0_��wAvi��3�����2���D��̗j$��J��POk`�����txx��X$ψ���m:��x����%"�RbV[����8�	�X2���C�(/��ZǘH�������y�q�MR;u%�Fi���V_�p�Q�N����:j7�����(φ�P�rG�)Tى�є���^j��a�(�����xS���PJ*E>P���T*��i�/���쓧)S
�SW�2Y@7ZEyu�z����d$j��~8a���Ȁ�l�t3�@<�G#/����;̜b�G�b*?)�|5�t0I�����/�� �:~��Ș�>CYC[�tlD�,o��^}A�R�Ʌ�m"k�8�Z���H��W�3W���F\�K�M�_�
!U���>�[Z11�%S$ 4D�R`���9ud�ͦjM
�4�2����n�^o&W�rD{��i�ZU�J .�l8$�ـ	��Oa�W�Z��dv&R��BPi��9�_~�<rU<�[���A�F>~�vec�`��I�Q�}R$�+r0G��2�og��X(l9��:��x��_�QA�^�8�q��.���^���.��j�֓�����?svc]9k�����絁��ŝ\y;嵑���%���t�>�-�I^��V1�B�Ku��g|JB��7W&<w����W���j�52m��Ğ?v����]�J��*�x-��}l\��,��r�Vǝ��{�#��V���p M2p����z�7�?�������R��m*��.^}�#޻�Jd�`��l��4��lrJ�G�e�vvFi�;J���~�r��ܒ��5S� ��!�`n�'7�6PbV#1����#��=������k�W>�t~�rH{d}����Xգ���н��ފ�S���X�(Go,���{�#d�@+6�8��eTf�����o�Y�(���@�xzj�{���;����y�<[��<�]���R�*h�����;\�rhN�^�c��~vNP�V�l� �y�R�W)s�آ�E����+�Yu#4��^�,��B4�=i9��9��,�t���.E��"���KvϣRnh�vY=e���Բ�K�*��)K��l3�h'd򈎰a2Qf���Ud��)��n��6��W.�i�������G�J�1ّ�z���D�v����e3j'9�ǫ�t��Z�6��<�2li�6M���Ĩ �x��2�S�W�pE�f+^½�a�Ħ��!R���wo#�o��2p��՚�n�K��D�� �m=���#/:�f1�c��#6��+�l�ό^�@kG)~�e��;:8@Hyi�B��>:׋{R���k�ɫ���r�,�,���]-�E�쐰"� klr6��Q@�cj"��g.����>�$c`,\d��V����F/����ҵ���I=B��G�dA���s?҆^0�,���ޗ��2���(=g�x޳��xY�V�$\P����u7�-�G��={!���_�2Y��j֖��rKaنC��6�+ <�K_�t4t~f��x�l?lyGfg��"���&겛X��X�'	Һ�{NA4RfF���Q{�tv3����f��A����գ����oz�����ԟ��Ԗ��G�����f�ΑEk�^��2���BFjH2Df,Q�!�{)�,?��tog7�ȏ�z��l���qp��(G�@���
�|xp��-�E�'�YcT���z��*�eQJ�� �z�{	_/90ԭ���� 6*UZ�V�l�nў�2T�@#�#^�C�%�E���
�cv�����o-��[	34B��U�F^nf-Kw���mZ'&mc��rٸ�HU�]�2פ�(�S��F���B7�+s�#'�"�D�ʄ��J��QxD�)E7^�7j/�fi�쾉�p��H@U	B
��c�����G��)�Z�}�z�a���A>H޿�@B=������1�� m�Jd�J]d�p�6Q��r����	����3���� ��x��lN?s[��Ξ:��K�:�������D9��+��s�6v�7(;�fg;�����G#����\�"��(�z��%h�þ������ڱH��<��"#n�Z1�7ٰ�����f�8@\Rx��b� 1�����T>��0��x���mctD=�;�f<��͖$F��2/t��{ 7e�w�Ÿ́<WJȦ3�Z=��P�{�^u{_��t쁏[��_��%���N�w��" I�������[ttqn��[�d�8Z2S�$>1 ̇���c+n,����MG��j���({�+�`��3��]GU��	!Eh��~��g.�:�A�z��y���c�^��U��{��B�BF�ti|�����;ͺ�WGak#��Im���R�s;-�J�K8�W����\��˦��%*{eh	t#�Ag|�.��뱵gs��g{��w�u��/�����ӟ��.�vi�1�;�Ŷb�� ���M-e�6��(Q�X�#<������w�P�UGI`�����C���ig��&��鶲M<�Ų���4&sC0a�0��˴��(�v���T�M;����qk�yc�Ԝ�z�v��0Fep��񆈑�ٺ~�z�����9���7�W�<�م���2��RgW*Gs;���?�J�Nӹ�[s��~�<�=w?�ے�Ty�����%ן�(P�-�&��)P����x��|����,�m*���dw�"�24sW*�:n����!�2�k� ��FV�@��V8ϰ�h
W�!���?ġo�(?��lX�������8ۖ�j'����7	8Ѝ��x�J��K�aL�0J�ާ��"�f�]�x��?;��g��J�nJB�o��+�	�gcΫ�'GyN���ֱx	2��"�n�'�� �6�M,�����j���BC��̟���<^Aٶp$.��z^!�ː��[����~�z� 1%��h���}lA.�{5�����lz-�aF���d��\�+Q�G��I
&�/0I�ie�j���3�fnt�e��y޴}�ʵ#�W��@4����N�N�����4�:Zg�s�;1���B	��V�k�Guyѳ�����97pk�j��|.le>�s�Ǣ
��2��Yk�a���<�/���,z�k�
N�)�D���-^<��a�}6����z�<����r�&�^���z��_w�#��v���H�9V��n���X
r�]�!s��_��_|�E�m�ϗ���Q	LE�8s��ɂ���e�Z��ǻb���"X�K}��ߥ����r�V!����Znu�	����,V�d0�ۯ���4s˄/,���9������S��Ov¿O���Ŀh��M]�S�(�J���o�7K�4��nӎ�+�(Q|�^�| �2g�!h[�����=�]
��J��EZ�{���i�����q/�������Ã�C�0r����h�Mcƶ0�:[vQ��L�P�a]G�|q�V>�!V���]f��%� +���{;��A�C�'�f���۳�tv}��' ���7e� J���^�m��T�I��Nb�)��D��kT�	}�b��t��;	3��g/lzG�{�VEiX�՘�TϪ͚��4��{�!��3b�U�iØdV-�����a(�+0״y�i��P���2�o.��?/�r��:YY�w�1��������%C�󬐠i#w�q���ro2Ӧj����L� wؕ�(��w<��'^����J/8���s���G�R�jU���TI
�y�����׻Q	!F�l���8�ֶٲ.��� ��11��6;u"���N̑��A��W��B�SLzrb����,j윏ځP�^h���" @�Ĝ�es��F����y��u<�< ����K�Aڼ*�S{�8�,vm�%������&�WULX�(M§�����@��6<8-"ku�V�΢�QL'����=�x�!*θ���	p�>��Yf=���y�F>�����s��ΫWoӕUױ�d�v/f���n^�2��ZP.��[�9
�zgvs�&3$VT%�K�Jh�����c#k3AI�m�^e��VF���e�k�71���\si�����&z/�}�Qmbn�(疽���ZVV.�3��5�u��/���o99�vM�V���>���w�s��q��������?��#�~�����/֖�4d�Uꉅh�|&�s0���`�I��a�v�V����a@��h�ym�Tn�i�8�W�\��tb9|p�z��{i=�.�����.)���ў�8
���و�R$}s뜣gW.� �m�.�T���x$r�|S��B橧�	�t�[�9f'j�3�n���2`"����<���;;K��^�ȑaH ��NT���Q�1���B�%R� �P�{H�|6ZM�%�Ȇ�T�������TWڋr�z=u�o镶�J�T�RuN)Y#�3ҹ���w�X_(�%�T�Y�xS�<qxWʎ3�L6�?�Ӄl��O�uB@d�!d ��J��z5s#P��)���fhI����P����{�N�������K��� ���{�e�}��q�޹3CEZ�-�T2;h��n�6E5r Ԝ�� I�Eп�?<F_i���� ��GQWpK��-�Vb�Ҙ���	��R(ˢ(����ܹ���g��}���>whɑhy������{�>��g�������$�ny�(>a6�G!�$dT#��f~ܴ��[<t���d��9��&�E�	�`8�����h;|^�w�H�uI�R�t���|���0窹䀈��O�����'Η�h�J&A斯!��>]o����{JO�^�'w�s��dol�� ��D,�ᇤw��e�H΅�B�Q�L�*Fǈ�ҨPU������5�P�/���ϣ��mS�,�ɽE,��t�5�i�I����C瞏D�ȇ��p%J`����܉wC:=�{a�1�wS��)�MQ�9wߧ}�|���i����E7�k���wm�C^�ͷ � @���Qr�BD�Gwܩ����v����,��{�����Z°���H��SL��WK��~�n���('�س�uSpy�zqL���SG�.X|SȲ�o)L3a?,\]���V���,n<��oo+M��hCu:�l:t�A�)hw��c=H�
ׯ<G�ܩ�'?��[�Z�&zenbw��t�C���kDċ�{�^0�se�Nh�{� ��r����N�QѺ:��(���#��k_ǧ�x �<��U"ｐ����M"O�����ˠ�t>�"�����Q�E
dѬٮ說�*�-��iN�~z��b� ���I9&��j1H/c )� ��>����¶�A�O��n��*�nD�)���'_Nk��PS�yOn�R�KW�_��Zgw86�T"�䞋��P������W1��"uY��(&�[r'���z\�D�`8�ijκ�]t<��p���'b��"GӐ�Tr���8�Ni0K�߃�'��;^E��ls(�W�������%g���k7�x�lٱ���j��t��Y�D���p�����(l�#��D6P��4jO j��|Șa��I?w6��ߑ<��ufk��ҍ{�ɇݥ���9+eq���: m��V��Փ��7e!Z�Q��m���~��o谥��V@0��@���dG"a̩6��ݺ�kq&9`}�|�=��*�soE����<6�v�>O2����l\�j��G�]jCt�T{JM��~l��W���,�\��XV2�0H���}7��L������1P�nk�cc�5(Ņ�[7�gR��5<v�Bv��]߿Z����]��>�Qh�^iK�sj���������@yʅ�p���NZ��������jA��1�*���Y�bA�I[�O�*G6ۊJz��U3�ۍYM���~��^ʷl��x[$L&�y�G� "9��̡Nًn"�����Q�^N�b��!&D�����CD�h
gV4`�]v�Z���j!�(RFg$�ק+13GE��x�jŪ4�塸�����#�7�o��8�s�m��4��� 7�Z��l1��D6F�6-�,A�w�!m�3�7�I#���:���������1�O����p5�
�>��u�#B}p��["�.�(��bc�-x1�!��i��gUe|�(��dWJnVB�j�C!��1qr�T(~_Hw:20Y�LgT�a�k�(����{{"Bz�~&A�"E��E�:����$��v�he�����(���ύN��v��T<5��7�]ٽ�[v/:�`��}�vH��bN��9�G*� ��G>F}�����\�S~[�N�wy����	�.�/\.l�<]_}nO5`&�K)>Ά���_��DVaZ!��m��lJ립���"iNUr'^��5/&� �sx��3( �L���ӡ$ú�W�5�/[�at����07:��l�c9Aǿ�eE߄��FzT���o�^ǿ
�H���ӡn]��rV��t���Q��D��C�͍�i�"����@|����14����h<HmEA4;��}�3��ʛ�P�/�_���pMzYӽG��1�B��1�s�<*91CTO�5=������(~t��H�*dJp��uއ�W{	��oQ��213G��}���Z�.�w|r��ޘ_���j��;�.|��!��)�>��_���v�M�uS9�0��
t�~5[��+|StvCOԜ�?;<4wNO��.�7n���#�b\��HX�S,R;�z�"ʄ��aԽh�8��c�~͡/���"z��|���4�oD/-w�Ņ�uD����+�qb�F�74��F����X�)m3����~8�����D�~玸}tħJ�ͧ�2�06�)E�8�!=�Z����{ts��Ɔ�3j�!�[o;��^��o1~��84]���ke�==��3��Zo��(�Vn�PaT 6��U0fg�XO��Z�*F;EL�%�'�;}MRɱ^(bt�hva˼(���Qh�g?a46�Z�ϨB��0dxq'A�P���mA�.50�t�<wbN�c�}L�Aae���Ĥ�A�H&5шDԩz�
�N��@j)beq�Cl���Rި%�����6��nX�<m��|��;޷Ή�P���E8D�Ʌ�oA�@oYy���Q��RF��)���BNb�`�(�u�eh2I�O��rEb{Qz������CtSء~/�=g|�����e~.�(��m�XN34:mk�X|D��Y	��h��z��(U�j�u��u�#$IE�Y|P3� E�#5E�9���QD%H���i�!f�Y�%@
��fH�n�.���!�|��U"�W:�]�hҿ⬾J����<H�$�[k�ނ��N�8{[���鹤���0��"�|�ѯ�N&���PTK�{7�5g(�^q%-�C��y���M��&ȍ^��z����X�>ۛ�_���to�@��:t��|����6�l&�Ch����"(:�TJ*��4�tߝuZ�b�����Si������GM��f�ҕ��w̪��W�'_x�#����>���:�R��6����#�oi�&�����E´5��i�L��4��V�s�q@rE/��Ն�Q�{Hc��i�}���*���9�Qv�>Hq��f���F�-��":�/�f�2}M+fHMC"��'�+���v���z��x��e���Lƍ�<;e�5��	cd)��K�������G��+Wy�*Y{5���+�����	��@�k�������)��R1�Vr�$XD�+�o�f����7}�l	pU��1^|C�#+�;QC$4�D"1��9�8�BZM&�Z�b ��M���,cm9j�o��X�Io���������=)�1
��-	�t����CLz�!'��pJ�
1||H�����8�^Vq9Dܚ��9~�L��1"��e�7d�ˠ�-�9EHuƚ�1%*8m��^��"V8.v��p���c��H����P6����mD�ΕJ -����zч�Q��`O`��ްʺ�V:ۇ�Ql�8���UaA�)��Ί�2�E�L�b������{�L(�Ъ-�����-~=�
�A��Z#��8Ս⨙wAX���6C8$�kp>Ӂ���!(D�\pa���#��r�n���a�O2�*�w^�e}�b���>�!�D�C��KD�Aڶ3�̚�"�c��[�0�tJ�^���rRx?�Eq�������9Ş���ډ7��ޢ��=��G���y=��C�E�rʚ����r�����4�}���Szɩ���P��ͥ=-
?CW��n������vՍ\�����t��E߫UUQ�,��dR��U���e�����/��x=*�s6[)Xt�#;�{���e�������}�[>�x��E��"aڂ�4�+>z1�|��zS2�B�( �!���ێ��lt�*m�nH���~�ĄjDˁqZ�Y����^�s�A\��b�o�����B~���k���\\���`Vs��u�v~� @J�@=�c5�Wf�+���ࠞ��q/N֜��2�����ڄ�\	[<nZ� B6��0��zKr�s�qHu���������|B�*Jq��R�"�r�b��C��v��1	�p�Ӌ�G�Ǹ�D�:�M
�% �;�f�iȉ�J�q��w��0��̈BU��K�A!�e71h�o���"_74�p#N<�n-Hy�[�t����u��M��n�mB-6>O,���HRTzߨ��vS��f���ﱐH��XpDE�x/�z����2=�9�R��O's����d����
�����*�IY8o�_�=e��gS�.{Z��@
mo��6�?sK�l!��A/m�+m`�I�qG_�q�p2�J�ɘ����"��fu�l�3���ֻR���3�?^8��������ɂػ�3�g��P���G��O�@��w�S�������y����~�u�"�S��''G'2� {"������7{3n�d��8�;z��Pj��8]��.�����q<��ӈA�s�=оI���`��c���1ESת.K�Z�%ݯu�ԡ�?5���h��Vl��֗^SU���rM���M&�~�����+&�ݻ�,�������۴�5��8�v�\j���QML�L�lo�o��窼sy6?-M��}��0/	u.�cuN7,��x�!���L߇S���Pb������E����4�ឈ#B�&G����ҍ�4�����3N[|�r�w��%�N�b��郛���ꇛ#uP��M/X����)��3ނ���\��,-�+�ר��Aa���6�/t�,9�wQU�Eq��T�G ΋)���4~�U?ՉBgo�%�)��a�pR�u�[��ЌU�>� �tf��"�Y�9�P�
c)��:����i��$e��#FQ6R�"�CA����mrº�M�L�?X EEq>]��[�.�1�s)��{�1��<��*�|9Ԡ+���8#����n"Ig���h����G�\ߵ�"�v�X��mmk:��=�od�,
r��L����O?�"�G��c�úveU�B+[U5$Zеb%x��5��c�tT��W�v{�t	y�Bc��K'�Մ�'��o�`:cL��o�X�&�S�nWM�6gD�m]k�-�ɦ<�J:Ѫ��k���^��:+7R;S9�u}okJ�t�v��xL��>�~��o�J"�l6v)eמ�uto��f��.���J��A��ӗfs���̊aD�H�x��ᑻ��n�l}�]���j=���f���V�-v���z1]�(B�cE��K�埣`�E��-z��=�>')rܛ������
Ob$�d'��GDf�|�~��^���EnD�ߒla�/����>���#?r���t;�E:�q4�m^���&�����Y�����o�W��t^�U�+�) �mb/t�yt�,d]O����[�Y�N��"�=��];���Cg��r:+�Q��"A]"ކQ�7T�s��n�9w҆)��A�*<�Ȳ��v��&� B�a�	�0#�� ?m��_���GP �K
ft7�VAH�)T*N����3	#\�\���%�Hpi��D�g�U���Ë�T�pכ�;+머.�t��7�����aJp�f6��A$���Pq��ڜ9GС1)��LN�Z'm^�(!�P��@��B�4 �5�Lp�4Wj��)��Jn�)�^3ꋸ�,(9�(���d��RǦ��>[N�f �����?���P�Ed4 �~�x��+@7�������8G��{�{-}L�v���H��'����i�S(�j�e�jM�۾����7����p��SZ:�w����t�:��>]~me6gm��X�.аT!���J~X�zZ���RGσ�C���Dj��shS�Vw~�i�qS���1�Nz�P���<�_��ž+�S_��ݹ�'��b!���w��6	`$�~�~h�Y.�o��?X7˲��ǚn�:�De��-��׋3q|t¯Ϡ��
n����=�c.vq�ɵ
�]NC��-����W��>�6�smݞݼy�Iꆸ���s�?J��;��������ihY;g��c��T�y��"˷����x��_���]ۭ���^�`�Ilց��h*�CC��{l���,��9���t�5�c&��D���=d����	_z�=��������ͦ{=�U�$-l���b�qv��5kDr�I�\��b��iJ���І�m�`�r|�Q�.~1KN�h������8 f͞�>������_Q�=ԣP�`M�.y���;w�/����$�
���k��zC7�z����2�lW"8��f
!����j:�Q���a`�)�s]ͣ�F_�!q˧K�/S���[���:���Ns����]�:3����	�����v~C|�ژ��ўk�ߢ�\�Z�t6�����G/��+�9UP7dB�{�,��z:q!2��SD�"4ZK��`1�5�u�'%Nݕ���v�^���~m�혅�n����t�Ƙ~��x �uXӹM�����Җ�ѷ���龀c3��Im�(�3�u����XWYZ�˶���"�j2�˥{eo�_���b�7
|�����'�3�k;� �E�/��(�����O�x�{��Vz=\�������fM��p����7,�+{�[��l�W� ��� ��W������+�ݛDT��5�f[�߸���ܜ_��{�~�k�R{���7� �� ��u �����}�����H�ƍ�g�Y���B���-��.M�!�a�C�.�{���k��!d��&(R � ��u.����M;2+��m���'�w��g?Aw�"����nz���B��u��� �f�cD%��bghJS��p(���lp�I��(��@�0|�Ά#A:a��ŻBj�7�^E��(v6��=1C�t�]�s�2���d&���>�������K���V��Z�2"[UO��C�O_߯i���*�� �{uIUb�^���8)�h���!��H�S���4��n�\��:�4��S����W,�Aux�������)G�q[�-_i����_k̦�W&���t:���8x2�W@b��;��'ĨsA?���ͺ9^o�;ĝw�oj�Lr�"7�Dn�g�zZ���(�,z](ԛ֥�k"H#i��􅑴����!,��-ץߛͤ���@���J+Tׅ����(�{g���[�1޹�>��M7���>�'�����Ki�SP,��������'�Ղm��ߨ��X�a�̯:��S��%cj#Qܬ����4��71aӵ_����6E����0D��|��;���ފU��j��6���ȶ�'�x�?��x7�M�Ⱦ�g�l8�����Xv���}d�w�ǲPZk���֣7��d~{~��}����O?�����
��k���(��F'�+һ+��t|���s���p
��Y�����jV���uHf{;@�����]Y�1$}ʴZQ�Uy>�J4n�Mgl�i���۴�({�^���l�S����|�=ХE;���Fe�Y�	��<��%7}��kq�\���rmWDMt\������EQ�.�������ʕr���\ �S��Έ�ά�Z�m��:2���=fʋ�Ġ9E`ҕ�+�i��_ӣ"�\"e�XxD����MGD�ߨk�am[����E��|������XX���x�i��;��[������n|i�Yܣ����<*��S�����1E�k��>��xSd�	EӶ't�kR9+� 6ɀn�i���	���ԥ��V&���:��u�W��ț�
�o��Ț���G@�{�k���m��D�������{����ݐ�(�`�h1z*��Ѫk�	z�K�qND�F�bD�P#fGЬַ��'�V��PKc��#t)%�0��m2	�Q��'���a�|�Ƨ?]�_{��z?�7���Z����F�vϮi7�8L����<6bC/��E���>���8���X����}��eE�ra��(� mJ!��rSn6�m�6��Qz��I��%�K<GW�ܥ�j�h.X#�e�D��,�����x�>���Ѣ�nyU�B��[�k��rq�����g����x�7����F��3Hcŷ��u>v��}�N�7�{F���}_���?�s^��ԗ���j��5�$��Y%�?~����ϧ�ɤ�R׵����\�����˴�?�� ��%�*���h�A��[��7�M�zQ}�_�6ә�-�����}�yR��(���@�H@E��Ƨ9k��I��o�)���w˱����t��f���-�0KI%�? D+\ﴙ).8�H$|Q;��x0p����'����o���g�UZ	[�������Mi!��뎎Oo/��/�����j�ot�~�[}�n�g�~��@gFF��It�sfc{.W��6Ϭc��q4�]]	��W����BUZ��E�.��U��	��]�"Z]aޕ"�/�V뛛��T�/���^���_�6_�e�{
�[�n7�:����8fVW5-AM	:�I�@ktFı�s�g�(�q�;0�{pg>-Z�}���|�2"a��Iܯ<��j_a�Fϴ�ؾ��qПT|G_����M��|�������Z���,^���nu���֛w���ѽ���-c�_��߽'ަJKFF�T-��l����r�dm&/X���VE�5��ѬǶ�~�H�{ꪺF�C�����✊R��us�i7�t�^��vS������V|h���Y�6�Cf���8��͕~��Lʒ	�=��|S?��4C}�	�Vid"<M+�ܻ��m�x���o���/�=f����l�'bZ�c֪�(Jݶ�;Z|�c���K��m�X�5W��N��%
�o�h|���W��=�қG'�_������o԰�����R�Gcd5�S,_�W,F�G�TY/i�֛�[ߣ�zќ�Y}��o�VM�����kEW�u�#������v�y��������7�~+k����U�Z4��m�Y1�U!zY�Sq�����zR��}?�ZS���EA���_�����e�b'�0-���nܸ�����Y����z�u��e�@	a�N!thq��M������{����GO���D'���^]�����Wˣ{w�f��7#c<(t���Gz�N� �"�v8�t+4�h�<q���Q��O?�ϖ''wh���������B�"�S����D���_����Y��/�l��d��� +F�S}3����]�*�Q#����.
4��u�\  $#IDAT�+�q]��~�g#�O�q�����&��q�����}��E�yŅ��������x�;����2)���z1�Ȱ4$�$L��օ��1�{�9��)>��@J��_�X�M�T���a���o�t:��:I ��(��*{t���ES4��H�p�K��m�eo�0�A�N���w!H8=Yu\���UJ��C@@@rIa��\���YBJ���k%w�ZJX@����NiPx������|���9gΙ��y�Kh�e��JeF����m�Vi,(:M���n�ﰴ�#C~Z⯩�l��%���6:9��Y�°NC ���J�pJ���7� <�Qɰ�����8{ƭ�ZČl�[.�O�_����u�!mN8pNrE_�Rpƾ�%wpZ^J�]��p��o>,��q��OR5|��L��X�In���g���
Y�C�g��Y$<�'m1=4�����U��s�3���*�eɌ����}6wf�d�0|?#Xҙ��ܮ�Ga[r�D?�.h���z�Uȋ��aV_�`�%�I��;����hy����ټ5�$2�̂x�a��_��3�S�=�,gOnv������������!�{���J�=�;�Xҿ� î�}T]Zd�TWj������.��|Cl�"|*����x�	������S8���*%�m�RjƎy-�������Ə$�
{�q�wVؖ�����-�p[ ���<�ӆlS�%��nk"*��$�Y"9 ?��V����d'{�(f�<�{߱�g/��%6}ElA֦ǺR&*��
��פ�Q�e�,n�dV��M�10"������J);���;���x����ѿ���,"��.�S�i r�>%�Rw���x��Jt�:��Pa}?U+p�j�Ç֭��<�!�>	�.�4<;����\��b�=l�(�iP��U���|����b��֢�%�/O�5���_W�7W'z,Fjl4��{V��k8<��.�ɣ4*b Z���ɷ"��
E�^�$}�������ۧ���q����O1_�g�d���=�	v�c�8�N��`��e���6�O�@���V��(Iz.�wӚ��Z	��|,�҃��я�[�߬|�P}J/��3�j�d2M�z:��H�8�W
W�h���O��%�>�e�w����>ȡ}�=�ԵI*mP�������`o/�$����N6��ߺ_�x�P�W����"e�=dC9E�@�*�8Z�f����i�? h������M�����A�Sm�����qSݨ�&�jy�]14��1�t��]�*G)T���io�^���o����f��3"E�:�k-t*Ⱥ�� ��5j�!�g^i�ʡ�֚f�y/�Z~5�"��λg�#?����x� ���~E��<��RZO�g��r�<�����S�X�r�d���8��G>^��͛�CL��"!5?���ed��d�l���f&����t[��C������w
$�)�1S?�CG�X��Z}�^�0$���6�}$���[���Է׳��Ș�X��'�hm��Փ~v/[�ɚT�����f���C�+�L�_U<;��BR'�R?��52�p�^��d��IdCz�ͻ����!���Qi�L�A|���"T�X���a3M�&�'��X��>^� ���>
��#ɪ�[�Ȃ�_a�.�W�9��[-5�ɮ@B'7����xe�ro�.3_ i��ܔsX�z�D&{@M���$�j��8�ش�1�M	>�c���1Z4j�|��5��0n��cUI�6���k䮽��!�7�#�7�!��+�N��\G]3�]����U=O�wǎ�.h0uYo"m� ~BC�5*�"h���-1�[6�\N5�k";#��M�����eUώ-�\="��B��%�j�U�Uf�% GN77D�	ih��>�d�A{��j2�i=�X�y��!���k��_z� _����'�l�*�\Z���CX��<���}���2A�a&�l`�2�������{��p2�V�Ϊ i4�B%â��8qI/N��_K��(��D$1[�}G�uon^�k|��6;ʱ�%��/�|�-;�Pq���	�<"ΪF*wy�Y�*@G�?"u��B
��6�Y(&J�J~��_�(k^�7�D�0*/Z1ȢQ]��n�5���~���9�FB��T�k�X,�/+J.�����[ ��n�9&t_:���Ïa�i���g�5Q�0ߎM!�wߐ�\���B���/�]��/p�B�>�P|Oz�?����/����i�N�� ���We7#i�g�xR��h��>nȱ��k�<ΐ��㋐�2��0M�W&������q3�;Z�����h1�d³a�
-<Ղ萬�QۺݾVￌ.��e�-��>��|��1n���w�w�V�������7
U4�Ll��w��M�Y,?S�l�6����P���[�&.�]%��u\$�A��=G$/7
�K13�;i���A�Π�J��L똻+1F�.z���:�����G�+h����j���F�3��+����l!� ���W��̃2���٠�rU�칏�D\�ι`{�d?n�[z��5~�ީ���~�~� #y����M/�$s�u��MyXˉ-�w�X&�=(V	l��}]�j�qvVVT�W�x��`�F�EpyQ�:,{����gР)�9�'��;�lЎ�rU�7���Úѷ�wE��-\y��n�;f�u<�w��N��P5��)}�����Y�d�|��y� �1�ᵈ�&Dm�Vm?��%��(�Z�;�N4Y��T�";C�u�C�E��MAf�1�?��aI�p�ɬ2wu�װ9V�4p�+|�_Ev����A�iugy,ߛ��_�]n�m_�HZ^��,d�lN������<���ӵ̃�����!p��.ܚQ=���dEWh�
�y��%�<��}�D<�^����f��"<%E$6?R����X�m�!�!��*��2�ZJ-�L$tq�aοo�n����(��#rhT6��.ZJK�{>���I�i���q��ܞ��Ԃ}��(�c������Ѩl�|M-O�y�Lk;()q̦���ǅs�9�j�^���7*6��e.Q�������Q|���I�l+0�bp��n�{i�8�HFm�f��p4<qq4���8����MS��mv�<���k�Y�:�U�#�-�I�?���!P߅���7�����O��=�(,_�ͷ�SY���ꍫC@C����M��i�rs9�z�{	�2�P~3�z�Q��:�X��!���fh�^����a�Etoi�.�/Ue�$n� `!�J��+���|-q$��6"�[�e�����#ccr=v���Dn�`��w��N��` pBO�q����	 ��o���U�q-��|�Fh�!���j@]w]�ŏ�'h$���	�
��)��/W�)�*�;%���k3��i�"p�WOU��f���iUR�Y��+��J˶$ζ� �3_J�"7R����a�8Y	�V��P8d5�P�����g5-��|oR<�汔&�.��ZGn�Y4���}�����VUw�������Y���Kv����|͐dY�I�S7��a7��%m�s a���m�D��qK���H���YW�X2ـkv<�80�-�@��dۉ�s}����"��%�ԉ�5�����=� �m�I���,�=�5����Z2���D��y�#՝��X^�	�냅Mg˥N�Y��I��y�>d�VgFS<� w,혍G��X��3$���Iۭ�����p�.���%�
=!���8[�_����Q0��t��VLAt�뵧a���L�L�Ϣ��N�A���I_��ǰP�v����H���FHタ��.�_��
�~$��T�5�#��� x�K�D庝��<�x��K��)�ص|/�ShM)g��Ek�M��o~"4~�)���m7t�{�gXD�-��j%�%��Oi��WΎ���O���]�5���7A�nB����y�������E��,�ڶ��x,O��x�dZH:*����#���Tr`�Zw�b�g?}�r*5ҙ�}��|��jL�ZhV��`[4�⪙�w��l'��I�Y^z�d u����2��Rj~����Q-Q���ZJP�F��A�鿌<.�`��߷��-
ܥ�����m�*[���g�M�vi(����5!�N���}p�}�lnv^���fl]R���n���ݓrH�b��uG�mۨ��M����O�j�|�]z����rX�c̳ _]\)�?���rL�$!��@�0U��
���:TW���Z��5��=e�5mj�+�0�������LlL*U��|�w�:]D��/'ڹ�<��*�aH(lN�l�%��$LG�N��s��������I=׊|�����W�	E�(6��J�zis|����b������ńVDP��,雗���T?1y��fP�1Y��v*��%��N�Φ!�/{X�	ί��|�4�󜶟_�ۘ[.���0��}��e�,z,�c��VU�����iGQf)J{��ʈ�Y�f�]��C��$�b��:"|���U��l©��{lZ�Z���^���2*Ǿ����aF�C�����~?��iIuS=��('���ѹ�N,�{�r��s竍U
�/��x�8���DH���p�+��ū�1��
)�&+��o���K�n�u�w
$���G ��� �ڬAC���|<�\G䫼D�ߜ�)��+�N�<ڋJ�+pcTg������`��I���|$�`n�k.H�4}��o5����L�0���FoT�%T^ԥ�E{������K�b��������&��~w� L9Y�]�5��Un�����D6m�9o��4/;�D��)�R�/p�;F��q|'â<9��bϣ'��E�{��҉����c��m<y,�;S�U�ٞvE���o��f��&��-
ۮ�(��eR'_	[��������|őֶ�����e�X�p��Դ�R*63÷,�.Є�|n�S� NË$�Q�it��c����*mO�W�4(����+0�Jm�я�a�tA�^��kkg��92��ʳ�5si��X�IO�nvQH�R���?�%߄���ϖ;[Zo9��U>�i�=��-L$��<̤���:�O���ES����c9YȤu����a��+��T���s�W�?�T�+o��Ǡ2rZ� ���=����P���"�%,��Cu:AJ�U��6�&��5��r�h���*@����{G����
����׮���&Z���)�d曗��5;�����<6�H�|�d\�u5r��r*˞���܈e���2���.��wV��Vw�a������\VƆ%*�7�0�2�o��LI�U��U䖌���
	O��Q��a�ۑ8_=����Y>Q��x�$\M��ET͸@�~^��z.o����Fmud��&�!�0�H(�d�c�S*-h���pMQ�7��+�,���ה������0���Ί�D����)���l���õ����&V�k3��Al���A���ϱ¿��܁��6��>:��c3�w|R�(���xYո���W�P�-'mÒ����O+�eq�U��.~,�����n��a��c~���X��4�bLYq*�DB\�o�t�K�k1_�yRt�"_��6M�%�-oI~��Tp��$)��������&)$��JeCú������Z�5EU�,"V|qO�u�����Ά�U�#w��0�(��������>�����Ѿn~a��O!U� ?{��\��i�G�S�5hN���O�J��=yn)����?I����#�Y�L�0�y"�tț����b��v(��v���~Y���:��aT�d!*Q��������~�~O��^��}X7[o#��1�j��4!7��#���Z!��p�#��ĝ=9r�剛��/��3��q���7��f,�b�O���DU�fM}(�7t�3\H><E��+��Wl���@~DiR�P4�Q��6�G�yi�ሙ��AGS���A�*��@���lzYf��yʂ��W��Byiq�3OJ��� ��V��#<�>�ڢ�������OŨ�i�N$+��]~��VQƓ\���((�M��\�%�2nA�����/��fM�[�h�Z�^.t��M��"�#�n��ӫU�Hm;ׅ*P(j���L���>�ȲӺ6���ˌ��Oݔ7/I���(T
02���`�[�O�O���	�u�u?f�}�C/������DX��N>\Z��v�/��lCA�.�+6%	���0�ޭ��>� 9�y^-N4��V&��ޤ<U��6+Px��A�Q-\�7KV�9mcp-�����K�H�I��t���W���v<2-��e�A�A�RW*�n�/V�.�sz����0J8�HB|70���]E����̸��9���5w!ww�+4�����`��<h�p���{����0����K��{�e����M߽;m\(OvsW{~�{!�O��\l@K=�2�bՈXFBt�Ҋ�k�33�'DW 8��b�����Ɍ�b�︎fV�a}�	%�a�ȶ��Ul���v\|�Z:z�	����� ��3�D��i�E�b�z��T��d��Z3�U8�gۛ��M����W/�~ͥj��k���ކ�i���o1������>�4���Y��I�)2Ɂ`}��x�(�$\��A�[�E�H��ǤDS��D�HB�2��$����/(��+�j��jNP�3�[e�4E�I�SS:����h�U�6c���:���JQ 	M�wE߻+K%�,Z��0Q��UEP�;⠵J�f�Y9v��BGF �!lB��2�]!C���b��C�M�WεN���ў`r��Ue3��s�d���K�1��>R��BXӓ.�:�ҋ�,X�Zu����]c�h�"�s��r8��DR3\8�=*WI���
cJz;�'r﫠�eH�u����A�83��,^㮢���\Y����u��ws�Nt�i����Q���U	Pn�P��1)�.��D��mY���B�#�.Xm,�q�.A�4�ڟY�SLJ��K^fK>8�r+BrP�AB��K���5�1�S�O4_
۳�=��ًt����m= {bX^�.� ��rH}\�uwf��z�a�[:%䪯�[RJe�KǀU�jVǵ��\g�X�bbCrk '�)�
`���	~�kC���n\
�+��ִ
�⃘:7�&�V��t���	,��V.x&cOra����s��;9.�W�C�� N�Ò��U�5�'`,�G�x�9��E��B0\�=B �|id�G<m��D�l�&1}�Ze%T�F���N��!�FR��3Ol}����f�H	/:~=;c��PY�_K8}Ѡi�y�㓈x�oƶ���@�ǴL��21�ꂣϞɴg���9mT^Y��{=�m���t����(<�2���ڑF�;L�}�L��g�o&�����g�d<����EGw��ΰ���0iA��8Hb��6��J���dE���=��_mBrS4� |M\M��n|0�*?fG�W��@1�z�9�̶�I��*��e��� G%�@-}�t�V�[f���4S����7)���������g��t�zt6}�L�O�
�w� 'ۂ���y\(/�d���l��D]l{n�gЖ��(��ڛ?g�\[|�{�G*bO��v�}��t���c�J��z�^Lsj����D,��}|���-���a�����kj�mG�	9�S�HVxl��"}(�iM�g{�A�QC &$�]����͟[3u=<�ؐs��?g;j��G�j��N�(&��a�Pqn�o���C'Oi
04%ck�3���ĭ�_�F����Ť��sď�W�jA .�T��Mb�k�~'�����g{��4/��o��			�
�g��&N_I� �d�^�fB�_�$��Es�#ݘ�3L�t��4�帀Ƚ�}U�q����f2Qʹ
��-���u��=Z[OJC3�= P�8���:������ͯ�����K���V>�~���w�]K&+y؊~���O�?H/+m����D�1-�� �C*��h"XL����r|�B=���CyY�zW;�&�8jU���1�Qb��|�*���������Y>� �ͨ/5�Vt%�ʙ��cd��QmtO$��s�+:A�Wcb|�����Y�aϲ7��)s���`L&�̠�ީ��r	J/��+�8�1Ɔ9��QW[�}�666��I�Y��/�H�FX#)ӻ��sI���Y��k���<T̽�m����V�&�������B3�`$��B@���`�>�}��x1����{�ݕ��Z}��襰N�����NC�u�y��<c�M{fbM��6'ޙ|ʹ�Z��ϯ��ٗ0R}�_�,�#�q|�����}�����a���>tѯ�.]�j^����p���v��[@oD2�vVG�{��u��^YM��QǙ�cGἀ��N���'[�LBow��!{��Wm?gH=��6,�E�Uם^��E�"����V;�{�ȭN�u�n>Mt�9sW���� g��&�bh����7�jn4��>^>?;{�\���w��N~����d�[��y��ǣN�P�f��I��t�&�z��(rr^?1��� �p��������H�l���7mk9ޛ�����O�[I�4�R"sߖ�:;�s4s��ϱ �}�j�;�t����v��֒���3?�gq�h����7�W�=R�%�&�������GS)T5��!K�'E�ܖ2*����޾�d�А��QN�J�����L��:1-��:������\M6�ͪ_����T���~�߮OV_}
�S@8���~�a�?��Y��j��k�<���_���EE���G��Ⱦ����߭vԡ��������1�	�烷�����v���s�es0�����3?[�ߵ��G��Ȉ[��Be�~�3�gm����Uq�7wuD��A�i6w�%95 R���� PK   l�X��� � /   images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.png���o&�����[��ֶm�v��ֶm۶m����U������I^�y'g&gf2'BQ^  �KI�*  �Y4��յ�?��^R�	 @����� � ??R�B���W=������+�O��O[���6Y��0�I��I^a����8�S���{@e�ΖxuV6Q�޸q��Mr�X�$l���$҄����vsba[!��_���%�{�����~s�ύ38������$������bz�m��x	�������^������<ý;d�ȝ�7a�����$��?$��Nu����h�Ɗ|45���IX��ˊ��>m��='*���'�_?^��<r�|��p�q@O�������f�����n����O��}P}ʯ#��y7d=t,�dE:�K~���!�����%�� �������)��q|�J&+��VKyri@]�����uQR�c�|5�{�I��au�t���Ԏ;��X.�h������K"��`�כ}e�kq�:�ŏ����a��Q��?V�~�~<Y�?
�Z�~kzH#����yZ�; ��_���������n��6���L�u���m�����DH��	�����)^J0�P8�8�cȅ;�r��y��0��o����L���{P��?<��笔���(�i���?���\r��խ�R�H9���\O	V1<���+�*�h�JY��]�6��0z[C��5�%�c�������sN�1��e��.��P��o���'e�����"������v���p
lqVh����m�[K���/��7���u�G�T&m�骦���WBԷ&��b����3Ǵ�{��^�>��	^rh-n���Ǘl��'/ė����5��C��D��@��x���"�}!���֭%�܋�el��l�J��=EQ|/�sGo�D�I%�s��� �]�+����3p~B��5�#9{^=�	�����[T΁�O�~��9Ρ���_Y��Q��$���0V̑1ˆ��M(5% x� �p�/N�,/w�@���{yDXoW�N�^��|�� =1"� ����Xª]�|uECf��O�v�)�Ȅ���
i�'
8#���P�1v���9�ٺ��͕�1y:����%��e7��5�y`��H]ݠ��LN�9�j!�ᣳҭ�V�A���t��l8ط��`��ڳ�p�����������o��' \(���P�����^���κ�����w�?��A6�iu~�Q�l��<*+�����"<��X��I�I�"������ΜR�{�^����ƭh���^l��8��3���V$_��ı��q�����k�Ke�2	�/׿e�jtO��ʅZ��D�����*oD�n)�ɉ�M��9����[/��|�W'�����N�O����e��|�s�q���!uO�U,C����a۱��\܇�c��}s��rs$$ط�A��l�,:|���;�A�Ě9�c�M����7�����tx���Uw��[m�ω�3� �^�3��Ðr(d^-dA��b�ܰ,��n�����#]���b�_V�Cn�&�V��W4 ,���J`���a�5P�R���0��/�d�o ��آ�K�Jiw5a��Y��*��)X�m���U�ZH�W���J��̇����J��g�q�j0f��E�] ��0��}�eD�	ߦ)��m`�L�xʭ&'�d��j����]\���\���[���0�t�܇����x(0ˡSC�g5�B1�V�U�f������!,����4��O$e�[���	sk�s_�"p����r�̙���|�}�`�o���]�>�gs,f�����[��n�p�GK+M��K���֞�
�E��Ɔ�Ϩ����,����`�5�y����D�Q���]�^���\��E�����H{Y�F!K�e��|���%�\)�ٵ�v� ��,?8���fK=��R!�Z��Ci��^~q����R��$��C��E����������_�l��-�df��� �S��)MG�l'� ��1�k��d{J0���������󑌽�,�X�����b���]-sg������6�Z�	b�93���n5���A}���O��2x9��%:����g*a�z��:��?�r��?�w��� �0f$�gއ��٪��
���S-����b,�#��W��Kl�����E��L������șxhV}!:�2��[��3�Tus�ke��oV���6f�(S۰���-�P�С^�$Qxy��ngp�s�>Z:�,dX�1ۧ�g��ޥ��Oa4���y���3�m���YsImS����x�sãY�
�+NJ��5�4W�q����wAyۛ����+_��q��GZ��s�#���Ǯ�'�6�J��c��P�X$��nЮO%�-���L�1��1V8�?\,�&�{W�D�ӕ�P��t��i0�3J0f�t�b
�i�p���H�R�����
ϴҭ�:v�^��֨�o,�4� ����<>l���'?���wt�=��^�����o��[��?�8g���Y/T����w��b�Gp{�������U��Y~�x�U���1|"3�AA1��d�~~*��Я��hQ���M�MpA�zY  XT~�2KR	t@�f�
��y�x�'�"���QdAn�@S6��f�����|��}QBR�ҸBN��3���ZNZ[�����S %$K�cE�_ns�x��x�X���iv���N�Mc�؋z�)���h�zA�=**.�_����K�AQ��i��pP3s�^$d��.��H}�B�ֹ���o_�@�To��!��a�h E�@L�����J�K���uL�D�<��UJ�_d�Ou@ڞ�f�H';��$�@�N�<ۺ}��no�~.gv�0Iv0��z�^m�E��"'�2PW��\oq=�<BR�ת$�u�[���p�(���6�m~Y�\�� �ʎ�(3XIo#&y[������)a�+Z(nh�qn*n@���t�Uw�B6�M���,H-,����AS�;�rc��V�o=-������1Q��&9G��w�*��i����b+%��;_�X�7>a-P��lja
a��ÂJ?G��Vro͡�l�FE�������"�=�c�[@C��Y�����Ivl�X�f�(ѡ�_�Hk�����peL)�������������Y\�h�-�x��JNF��YZ��5vx\@����^�
�F��=��������AA���Q��Q����0�^��`X<Q�[�t� ��Lk �^ސ���p�U����^��C7bZ������6���'�m�bQ	�A�l4,�@��Dq���S�t���ܶ��z�r�9��O�Û�|u�?~�>�?3~oU�X�� �|zjS���Uf�l6�]���;
It����/���E������q�1aN��շ�X�:;�%񒕞�Y�~�VcbE_�e���aGx6L�a#g�u�i�a����Be��6,���7������ਃ�j�D�Ҟ�L�����ieA*�0�Q>����a��^e�*:,��2��2�^$?���^��*3;�z����s�ky�1����r7��dB�p��q�� �@PCb�~&d <ȭ���6 �C�H&�1o�*
������~O���*(ӕ|�����>���:��̛�7�P�<}Ōi��A�v>�;d��iN�bsc������.���d!��1���K���օ��V�����=wOܼ��`��n_�h��mx����u��\=݆��w�5��댼<1]�'c��6��a��wN���+O?4܂�J�c~.����Q8N�����8�=�w�Ҵ�H��R�=\���!l[q��;��}ۑ�����ZT������H�=)4�]ؒ�����d$O�V:>�l7��V�р�@�T��A변+oǍ~Ƣ<J��T�L�R�i�A��z�R��>GI��8�� C�r PW��;t�v�~������F@�S��4�U��p��/`"c�Px���<���Xd�3�:�7�<�WTYa���}�q�����R��[L�k�*vP7/������H�S�h$��lݺ��9�^�t���b�^��
E�U5�z'�1s3b���O�g��
636o'��q^���RE�1Fo4�#V���}��'�Aq`�-�ñ��	�ev�{�78!��k#E@�L�Tp�? �b|(��q�٢��ҷ�L���b�?z�[�Y�n���v���ue[�qk�#���$9�d�����,8�T���!D��s)y��h`��V|'��6��÷���i�ZB�z�0��gW�H�3p����WV/���x*��h81���"�2�x�~�NJ�W�vg`���`����C���N1c��&/x�A��|�iRf4n�ZLvL��5��)qА�5Z39wĨ�G��;6��O�h4�J[^^��374��PPu=$n���Da�����h��� %������g͡!�����2��]�ܸ�/;�(��}Lak������_�Q&�n���R��\�~��;��y~�������4m=id� D/��,g���Ӻl�ji�]�0 ��("�.����TO�m����A�/!Zʸ�.B�J��3��X욻d�-��f�88|Vƌ�`ʹ�0�a~ݚY6�j�Eh���<vVsʫ�?�B%|Q�ЏW�e�dQ����Ʈ`ÁUXS���4* ������)� AE�P�J�tT���,�!צ=�kd�x��>��M��ӧ�Z?4�NM���r��!�,7���Vv�y*�t �����"U1�P�+���Px�,�8Y:�{,�X��c�d�W��Q��n0��E����T�����K?{u���A���B�J�p��pj�wG�r)��P[��I+9�!z��u.Zk��-A�,O,DS'���*;D77��N�(AQ@��{��H��BAV�"Φ���݊��z�?���l�b�:��U�}�#=x��0T?�1��������$�6���I��7������mlm�=T�W��)AA<4��?f���{�~�=�$.�w��n�]�eteL?�BE��&C�k8�H�ղ��5��s���"6y~��V=��[��F;{�m��|��ʘ�`�%�1�pzw�J�b>hY;D�X��!_�l̧w����hO����(N�`�XʰI�����Ȉ�7c��Z�f���#[U?����d����ǹ���n<]���5&����.굘s�7�K��_ ����Us�-.?e�e]u���]�抋bL�I&C�p�I��a�$��+��K�t���0�-��yf]� ��?#-J�]�2{�.��SI��UuЮ�(�)��z~����)�\��h�����i����,*�ܐ�e���*�~"���%XPj�U����8|�=u:#\�]�CQ{�����X��ݢ;3j���h��1��p,�h�.X�l�G@����t:Sh�`���V��2ĉ�A@C	�u�=.��B���7<��(q��2ޖ�����2��5��8�6�d��Q`�2Ŧś�̐DTһ��% 
�ڲ�tj(���d5#}kKl�J��M怣�M��A��ޝO�`�hF�t7j��;3{RÂ���(8��o�k3ғ��+����MW�z6!\�^��
u��U2�����A���x��&3��h֥?u����D��� qG�e}�9��JJ��f�ep�Dguw��0D�93�-Ջ5C��vA�~�V��4]qrw&�M^'e�Õ1��]�s���1�V�G��3����csGL[��=�o�U�Ʈxv&�R�5��g��Q��x�/��P�a+�3'9]�hlc�p�ʬQ7oؽ��ل~�֋8�5c ��E��w��[��Yq��#��v�
�:�׬�!�g�Պ��%Ng}�_b������I��+���ĺT�ߞI�qfZ��� �M
���D���j����&�J��̉I�6s��Ӓ`-ՈU]�eh��H��wĆ�5���?b88�꜕lђ;]."���"Ma�ۙu�Q���	�3���mdFc|�\c�L�y��כ�	1���,�o�m-#�S��7�ǘe�s�jCHѐ7�FA��+ơ D�Mw�=��;ѧ�Y�v�k06�������#݌�
OL�*) �F���v����Q𩇟������j��W����}Kw�'U��@���f۽�+������t�H	���Fc�$�lM�I�j��K\���o�^�e���A�}�@�3x.6�+�.7"j%� �ڭ�Et4-�Vx�UJ1唲�f�T}���#7�E5� ��l����Թ����_�Z˕%_?	�M% �q���<P9:�5:1��4m�������c���xRh|4M���|�\b$�N��>!;�����4�BZ���t,��Yg��)Ԗ̢�� �5J���f]wC�qr����T���Yʶs
�N��Z�ģ�
?)gr�s栞��[������#���"�ݖ ��D*��s�ڲh��J���/	��IL6�b4�� �!�E� b 7.CƢ��	��,~斣�#x��/�sr�Dn��#��w�w�{�
¡�8=>s�k�&�K�3ԧ��Z)��P���k����"�x�������#1�R
�+D����}L+ݾ,�ɼ��D��>���@f�wO�}�:'��~?_�1��w���U�	m3�fd i)���Ǚ����;j�%�oڧ�f��GzS�S�	m�,Ze�6��6H]sQ�c��%Nݿ�Qf-M�t�I�PU�C,?'O�?$|������W�)���"d�&:[n�9�5��#��ӀW�gQVL�1���;����-��BP���N��jJ1�ȉ�j���pǌ�������h7G��N��ȹ��U��M����)��H�t���!-�z��Kc�Lb�w��>OX�`6��O�{�V��	
٫�}��݌7��	ĸq�/> ���g���Ƕ:>�Ѝњ�_�]m�nN�b�.�� ����\���d�
<
8�:M�< X@�
#m�1QE�*#e��^�v}B B3���d����Ev��Fb�tw'l$|*��r�M9ŦR�9H�`��������2t�7WE�{��c�w0��`3�������m��:��*5?	���5�3�I�;�p,qB���{�q������ܱ[���=�Q?ٔ�_����"g�3GA���lKt�Ѻ~�-��Sxb�)��6��:.��z~�MƢd�3�]�{@oܰ_&x�%p��j�$u��G��,]�0��u|����1�H6����Vc%�����R)NΎ8���(8~���R�L�;��4�p�=lZ;觋+��S�K{�L���ʽpz@ a��~�x4Te(���C�N���Ke�r�4}�J���Q���s$J��wv@���=����:�=p��U��`��A�����!����qb�̞��U�F�x�8����˲~��җ� ��cjSŵu�b�I��X�9l�)�x���ܙ�"�ã�z�	+#���>��˼�!��2/��+q`�������H��:Z,��	%������p��yf�,�Dr����~�1�w�4GC��������%��+��X����j�E�D7����g��Ì6�5�sM³$}���I��x��8+*-�K<Ǡtɶ��	{����;�@�k��p�hH�/��B�H]
�I*�_�N��{��]߮ɑx&���x�J��]�s��R\v�ӷ�`��=!9�[�����O��A��J�����3�^��}����XK�l:��֊���B�T���t'~ą��rۙ~4��yncߥ���g�q�c�fM]�_њ�����kV���n���:K�8�Sm���e��c+���2b�\%8�[.T�GR��}^~���*��e�⢐��S�JI��S�x�\�.]�6Ӄ�ja���l)������~phQ��R���$�^=�]�*
�+*�NLI�]��z5U�F���C0�&��/�DG�RכmG��.:Q'`�Q���8��H*���F1|���:am��.ݩ��v/S�b��C;���v%gy�	��G'|��O���+�sJ�����üdn�'�e�Ry�P�Z�7N�9�80:o`�a��]�	��ICDp�m m��kW�ٖܲ��̥A�z��:�&XYMN�u����Eg}���4F\\���S�t]I��t��qI���+�C��w����"$�.ņ����[�n^�kӂSuF@zQ�Ӽ����j=�Қ�T�0.䮧@H<�ގ��_�� ����SY�C�EB��U��a�ٯ8��Z��J].�h]�,���ە}��Dӡ/�1g�E饚���Km�y�J4�5٣�4dK�rZ�y�j6sdz��a��Ԁ���
���� ���j8�o�L73�s�Y�3���i
R�g�ȥ�r����L����F(N�lx�
�����^��8�	�<���A����y�%�x1bz2l���S�5e��|R�� l�"D\���h@y�� y�RF��sSJ�H\B��lA�O/����rz^G6���>�!�����I�\Q*�@�B5Eh6�; Kˆ&�I�#��%@Q����[�s2xW�rKB-0y%���!����#�X��!#n���T�#y?%8a��6zT;��l�.��0+�#wZe9�a3G��G~N�}l%OŞ�3�w����tP5aj�.]�2$K��cˤ�=�uc�6HC�����5\�����m�F���u~JŲ3�ܢ�`��^XC..  |K[�.«�lD?��-��Z�z.W���p;�}${Tsk�ƺQ�P��{��qgV�����Ҏ��H�w1u/�g$hŖ�AܩC	��p�&vW��A}QkZ'D���d�%�a�LV��:���������iW���_���%���]$�N$�y넳 ŧ+�u����Q[��^󞠦��=�Y�˗!�bQ�d��8��z�֢%M"	O��˷j���z� ��?GSELg,�h��V���Y�-��X��5�ݳ�FU��Y�SUW�-4c�����0p�!3V_T	�!�fu�0�4Q^��g�?��/)��B�1���֛��P\���P]IOgN9d�A�Y�:i����,5� ���gw�%c�{Ư)<u�b��ψ���lf|�f��$ ���ꃄ�R�<����g���3=s�Lq)T��D<�k�l|�O��ˍsiF�c�t)b9��ԑ,����CO��a@W���l�4q$՞^���M��5�][ЬJ����������I(T�.D�'ڑ1{��qIg)�/A/G��
��B¿X7�?��w�;�o�����T�"�1^�� �n4Jg��/�~�U
�A�@?�[�JO�*��{������e��\�x/w�q!�~<=-��X�E���qCb�\Mg�m�<R:�|�ˬ��[�K�[��i��xO�᝹'Vq��������[}����UO��5�ꃘn���� ���_��nEfj4]χt�{m'�}��D���?>���հ`��S%�V$]W|��B�����[��H��_��iYO��H�_+��|#���ɕΓV�A�i��W�I��h��k���9��v�Ӄ�t6Sj�08� .i���I�9�ܢ���t��n����."d�]Tg��<�jK
���\�/F��yJJъ,Vy���+2%���oD'W4�h��f��2�l�>p�R|���9�L.��x�/Λ{�:(05�����S�qeG�Rl����iHo,����7��ϱI�i�m�����#�9uPz��>�c�O��n��G�@>J�E�ʴ�]�R�2R/jU@k��ƌ+��:07=�|�]�@�R�N������~		OLٴ�WYUu��S/W�a�JLnRxg�$��;d^�U�J�x�;�,�vBi��7ٖVw��i�O(Sbcۢ��}n��E�Ol���������u��>�վ[�0�Uk��&I��\�ZBMe�&WS�rbY��Kn?Ş�����#8�%Mn�O$��<BR&��wU�$���lG�
T�%|u �����*{`�\`�w�^ S�G�J+�
|�����G�l�d���ʜ�
z�&��ɷ�!�i��B�qztG~�U��w��x����\vߥ?�j|�X�|n;��� M#�&FT�I�`B}5;��Wgh{`�p���Y��?��wv���Tip��j*�CA�xPS��?������������|�bg䱡�V	����9�;�p:�9i_9�����I<�>�9'��(���4��N%|�V��s?Olo��61����1��2����*�rN�X�Ӫ�@�:N���M�|_�=)Q�$nu
�A��O4w9ĉF����P��|ϴ�V�׹��ҋָڶ��Ͻ(�*�9�ҜK��ʭe\m�����'W]�J�F\����>d�!�T(!��`��A��b���I��JoeH8k�q��N����-�����ԍ<��NB��-�E����yt0��Ի�+��;ӄ"e�0y*Nd#�3����>ꗾ�l� v�;i�?D�����T�3��9	h�xB���9�:'�d^�4���b�~`�~����j�GD�p,
�j\���]&����Ԣ�x�{����%�y'�Y�ypf�Y<R��@��
��:t%#L��j�L�\)�u�(��V߶
���c٢�>�ME�e�jFV� �
��y��tJ���B�!� Mg�h�X�bMe->0d�a��c��%?����I^ �$[�ǃ86�ڙ%<��{r*�be|�H?�O����6VT
��;���Y6[����c�*���B��fk9J&�pp�@>ߋ\�q(��>�*W�Sr�c�s���r�7���L�/�@g�,ŕ����6��[�Oe&���A��hNM+��V-f���A,���QRV�_?�cY�
��
�#��y�]	�x��-2M�w��F�p��0�}�JP�R)�B���&�xP񨡧���}E+p��l�pvT�.L���Lǆ�b�n[v�����!'=�p���N�޻Yr0a��,,��lvs��i�޾f��i6H��b���3��h`�p=�]zZ.v�6���:Z���=dB��4�4��4���r����q�j��s֐k�eZ��0'kh�>���YG*W����?\��l.b5�H~�:+;&:S����yG;*@B�_A����V�8mK�5
�@C�K�����ۯ;�rF��i��+��Y�#��3������=C����84�Ą|
�Y���:<Mi�+������`��o�	�u�E{5��+n�g��	A�L(��v��+�;�� .�����-M�ݦkI=shra�9�^�(x�;i�2P'�y��Rt����;�W�cC��K�,��{�ƚ4�X5
�>�Y|Dh\�'X􅙆�s��s|���i�|�����x�����VFH�
��c�㎪���1F� n��ͩ���V��OYV��{x�2
���L��y����_��G�@|<�GZ���&a{�rv�=��6G�o�&�*�[�m鱰X��[^�Ld��!���js��{�" ���5��W��͐����4�ر�rf�f�O<�����O'�}�� ��D|�l����Ee�scg�\C��S��.�YAI��I�i���c;��p�RZ0���ɕ��z��~
M�1�u�#�b��w�"�Q$;^M�L�l����S�����BD�Yު�$B�;��E^�1��O�4���.�q
G����Ɂ��8�y��EL��O�4SO�z��%�Z�LI�	�'*ln3gR���S�S�6�=Ň �a��rTIF���Q~��"� >���'���r���QcˁX���S�sc�y�v�����UcAex2�	2�_y�h��Mf�������Sb��&�����6Kx��6�9g�Kґ�%`��؆m���.5sR�L�D x������7���Qb骭��b���*<�����V)�9����Ԓ�	���Y��1���.�/1(,f�p�U�Z��ջ��@!���3s��P{1��'rf�w}�)o�&����3��u7ϝ��#w]<�]Z��1¦�O)m-Km���+�� �.�p�!�\���;ݠ17��@�0�A��ܒ�9aXy�dA9�w��4?�!�#�v�_+vGkudt��I�ۤ-�&=eޣ�Z���2B5M�j+x��V�%�C��U�� ɠ^1KS;h��ϧ��F���G2�ss���N�Q�{�s�Y�f����ȺÄ����k�Mt'e36���6	pg ޮ�Z��"<�1����:�_��1���9���}�ETM���o2��GE���:	N)��_�e@䝾���`;<����(0���hqQ��T[����>���')U�'����d<\��K���}��R���fm������qL*j|&ZX��ie̸
���p�~Y��I�w-�O�`N u�I�Gu�uװ��h�ȗZr
�Q�/�j��u�
�VT����gt-h������p������=.ܡRQ�Y�k��G��f5~P�	�U�����4F�x���5��H��n���v����kt-T��u��5���݋@���cy|�wa��G���v�.D�'��� �����W��ιּ�=�޺ؠق����77Ej�Ts��ϱ6ȅDΡ���rlȷt�y�e��d�X��RyO$W�,�q5�%������������� ��7�ŏw9�}�z=���j����`+I�B���~�3ԧ2�x�~���K@��u[s�?�2Tuy�|^�8S�$����u>���a���:ņ�i�
�-��U�tj�,()�]O8����唎㪣��L��M��ִ���;D�69��>O6�5fm/�4�?c�H��`�oħ`fg�<k0��~�l	����jfiA���հ>��L�2��VS�J�����ݖ�=�*�Pwt��QU�'=�
�r��(qqf��-��H(�m
�a�ENS[wt}L�A�%B��Y4v,����8�O�K΅�a�.u�ЀoI�>�j�v�ky�F chލVTx��2RoW��D��d�߮N���oi�圎ow�6D���2��� K��I�S+8+� %� =��T�{I_ڛ�]���z�}_#��b�5&?��h�Q1窛5(�;v���։M���Y�>qّ��h��l��r�^l�c�g'�Fٞ��ZX
��Y�߮�?��U���A*@��=f�H��Hlƈ�����\=8�w���txj��D3��p�(B'�$��Q�S�,iE"���T�ČM7/�A�ƴ�f��8�u(j<w�5%9يE�#��u�9,�7�e���Q��ׂ�����@�*=��i����C�:@���>�Ǭ;�������Ҙ�x�N�}��E�ّ2<s�=�s-��q��]��ܫ멏ut�%E�5i��vU�������SI����h4������Mh�%{J"�7�Y*�\bs'� ��7$��b�;��*^J}0[����WP>� ˶k"�vy�j�x�A��m��GG��_+m�����I�s#!�ƞ��~�E��1��ZvxA��O1�9��fN�B'�Jn�z���M,?s���AR~u����0�-C���M��x*Ӱp\�Aq�E0������c^y�r$�9i\~��p�zdEJyܾ�>�ء5���G}?�#<JO.�����:�.4c��t�Q������yɹ���ޤ�;��KM�6/+��Wz�IUZ��)lѐ���o�I�x���l�=��L���#��n�ڂ�^�9O��QDL�Axv��u��2�d��R��0&ri�O�.sjí�������<������F����gL�̲�!E[O֮l���U�HEA�Cp�
oIͳ�t��!� ���jW���.V[p��h�߿�3�KrV����f���$��7Ym��[�nɭe�W���XQLcCt�Cc��A��sU�jK�@�Ƽ�]Oק����P{O�n+����Z9��B��r��0�ӧOT�����闚4F�]#P��G��Rʠq���r�k	�EW� �Om�*��j�Z�~������7Y{�%��q׏�h�N/y���r���[{ڕ��5Z�ŀpFe�s�UQ��^�2��N���� N�N��)z�-�0e��>7'{��ST�qZ�߱E��X�J��x���"7?�ْ���rC�d�C�ٹNa�#0M��}�,3��Q�T�Rr��]Fl�-��pl1��Z��0���X��<��ؙz{� ]��VT����GE�������T(��bH�C���?�ۯ��?U�=���׈U���q npp���4��:����I$_��΅?�w�q?s,�Q�� 8����c�x�r�{͉Hn��[4*�ϻ�퓄r����{��M{};�*`ls������ă �y.��qIZ�ҍϳ�I	���C�Ͱ��ZX��;(�
�~����C�Ϭ�@�ܩB����N:��?K]@���g�Ɲnŉ�b�F܆�El�o�A���b�S��ܣ���ΰ(:mQg�����y�����2t�h���Kzy�T��5>S�b"���c
+t�:G��p�������0�(I-/)�Ė;�6Ab\5�Ś�oNg�B��%W3e,4�8->� �� ��όƒ�?y������c[�k�7T�;D�k��V�� �E.H�!!�Ǩ�� r]��~�~z�|Xi8�`���Kk3��l��Q�{��Kkm3�]J/�
�~�+������u*�a0�J�����T/�3�H۲w�~�Q�ZZ����^����+ͺ�4�0�Nh �Ǘx�r�w{�ʯ���N��ǧq�Qly�])�wm���ޝ<&��$""b-�Ji��n}���sѝn'��u���F�w����Gn�6�(�K�k�������WB�z�W����?��D����JY����1��)w�s���	�6�#�~~�G�p�\��Ž8��X�X��W�������p�b�E��w J����^/;T]R��C���'�j/�T�7M��e�g�y��;���O��-����B���>q[��v͙n`+OP��[����yS���Ļ��,�y�D�:����7�T��G��S���t�����}m��&�0{��+�2������$Ojc9dj��	U���w)�V�K�&7��;�^�6ւ�)t�9w�AQI"���y��s���\�-L��P~359�k�<�hwч��N�^PM�d��S��z5�r0"�'��y��
_6yל�ڜ0��p_�%6��3�L|�lO4��^@�I��]ă�+�xyz,dV	�
0,3�����&C/'>��^߿U��>����"Xe��XNKC4V��87�����V�>˶��ϑ֦훐j7�Ԉ��<y�s���|��c���͖n�,�++��y����j���!�3��_k���15�-7K�d�x����Ŀ�sVܖ9�fZysQ"��d��5/u0�'�M�mqef"��� �<H�.4�z\h�뤰� s#�z���"��bF�qA��;S������d�g-���|<�)\9%H����V�ёK� <:�r��s����iDr��@�l����k���r'"<ۀ#��'� ����:��dnb�ǟ�+�ȃ$I�j�"}�rb����>�)ጯ�F�m��b��Xu�G�}� (�R	�7�G7�9��!=���at�>��(3���I���*w�9r�2I���7�4HSՅ�J����p����j��[E���ֻ�2�A�kh�2jN�ZB�m�1�Ě	��N������7)q���4^L���I��$���Q/4:�����:�:�W(����9]�/��m���w<�@c5���sh�ʎ߯�h�	�M�L�ɷ��lz\d�������O�w�~+Zm�FX1\�j{��:�]))Z�]�t�|z7�6/幕�ਝ���:$2A!U�,���eL��.��E�N�l�(��MZ���?0����v~�R�Lp#mn^��t���Zsݠ����Z8:�N����%��*|�'|���9�����H�#D�p3^-S��ra[��{��%g�~F[��=xA��}���X�~bzR�}��I<ࡢ&����6�s/�V�Mn��|�X�uR�$]�͖�zy�`�9K�����h�:Iʜ�	�)_1B�+�7o�T�������?b�O�>X$m�����T��VT��g=�� �&	��_ɒ�>�l� f���ˉ������:~��ǝ���<�?���:�k7�!b\����U��� @���!\��A��w��΁풉xkevp+��"	��dq�^��5.��4�����NÍ���D���~������8n���O�C����e� ��yB�/���n�j����V��a ;f}�+y<Y�TVQS�GZ�`5�:�y���vε��	�Y@̑�{]_ �<��qM�W��I�:"�_�s��أ�m_&�il�g("�CϮҳ���<��%f2�abSc*�ɂ+��bKn֍���	ٻ��N�!#�jebW&v�,Ԗ�@���R6��}��`S4g�sy����٘�g@o��S�lOV�,���^��R]�������k�Pt��[g�8t� `n�.���h;�a��p�����֮�<TJ��i����{a��(�n�u�a���I�͝T���C�H�����G]D`��\$"���*`�Jt�CnR_\�W�pE/89�]�y���߫��(��i�s���;G&Ғ��^�uG[K��u��)���8����JJ.�xz<��ǌn0�G�V��l�����fm�e�D�bϋ�����Q�0�qR�j��`�ώ5�ʒ&gj�.�%�Y,���ȏ
Z`m`Sh�cԍ��w?�ɪ�[eV
>�Q1&L��

a
\��:�A����� �ӍQ������J�'�G|Lz����
E߶6xi����`_m6���������w-#<��Χk5�?��ɕ���z�{5T���qi��C�i� [�OV���K�m�3����_߭��g���bśU�Q���'����J��V�B:�A�Yf���eS~e/�����/���a����h,�5�b����}���2��2��LfV��z�iU�fk���o��-���`����:�o_KӞ��Z�cg�\l������k��l�����A�i{��{�U^u�x��@�9JUC���O�M�M�-V��tFc?� �e�#.c�72H��<����0����+���^�2e��X%td݊�ZX���oq�S��l�T?�.@n�\_��`j��eǈ�>�-�^@-����c������*)��da�٫Z���|ر���X0>�5z��"�*	���L8Bz�l�
���}k'��UW�G�@�����Χ멆���Z��e�kem��\�Ϗ؎R��L�;�0�����>��;�k7�F��;3���لm�{��7�	����Y,P\��G�m��]�)�ޯϤ�l1�۰0^�VSj���XuiƊ����u�T��6݇�R-�ՈM�ثP�l�qh�o&̈́���*w?��Ƕ�=�.j�g�s�n��:Uk����¢(�������jKO������:��j�o��jK�0�7��1�ꨖ�>[�=��AU�k�:Z+0,V&(�A+��i���z܏LC6h��s��UYbZȂ՗�L��Y��9[k+@b
z�n���\���w��k@�Y�cfQ���L�
��6��]*s�֜���+<�T��gU�L��Zb<�
e	���q72�[+$�0Ȋq�r��vKA4�	n%7��������:�I�{��XL}2�9�pŻѓ��}��\^�3S��*D�^�	�R!�����k�b�wZ��$f�	�k���>C8 U@�d�e���bw�V ���T:���;u�w5Sx��C+mJ��yE����G�ڨ�e�w�_c֘�mF�D �^=�eRF�.�w��{�Ge�[7L��n]���	ƍ�?����!m@��|�GQ�IuO5�Yg����=l;O��0B�1gcb�{����*O$׀�=*�+{a�m�[�$ �2A�D�녺��=��o�zcPZ��!Z�W 2�Io�>��h�4�8¨GK"b��V����G٩ׄD51����s�v�g�jb�3�xգ;׸W6}M��AZY\:�.;�V0�	��ES@&����@,�%8����
��I�=�z˰�o��x�%[A�҃�u�e�$��͘�D����}����O�Qp ���~e%4X�p�	"����o��Z������+���Q'>bheBbOh~2ʷCYl�19B.�a��_���^�rr1W�E�Ƴɕ2�'���d�@>_ks�ҤVR{븢�{1:�;���h�u�K̶��;��1>�L�
��`�mQ{z�0;���"��l�g�Gl�`;��?>2��V��`���^��;�#X��+�`�2�����c6�Z���Ⱦ�Q8 �սC��3v;t��p^�;��9QN��@�e݌�J�*�<���~j�	5�keL�bRl��؀�^��F@�n�>� ��s,�៬�1���1/&#J��e3�F�֩���2��Z6ױ�V��3�l�ِ�5�F�w�Y�V��Mq<�Mc��P]�� -YSX&:��+���k��>p�a��[5�����d���w����4<^�an��_�-�L�Lk6I"���� 
�1ȯ�0����ٽ5���kNNU��n-bn!�:i����]6
�=sڗ���eX+��{���`�������~�V�b�X��?��I���Ý�_�ɍ�����-�Y���D���lw�^_˭�c6����MV1���t73�\�
r�� ��o{Z�DVcT���.�g}�Y'-+�C�z���b��
l�������(C��XSP�Q;�b��H����I�O��]T ���-dpV|���������0���:�6�s=X1�^ �.{� ��>����-�`(q��g\#���0E����}c��F�^�����B���W��K�@�花�d�#�7��3)�\_I_X�+3>hSZ2�m^�B�
H�H���tc�60p� �����(�-U;ۖd�K<�����XOr����0�/�/��S��|���5W:t��d���o=�^St��B�b�G
*�Ω$
��@6�6�*#>9�����!&�� �Ί�4)6z��F�vf'�2;;e<���Z~ү��v�=xH��k=���#-��R����-v;�4�J�صn�([��1���%���[$���"�ϟ`d5ݵle�v��ǁ2 �w~앵5�6�l98�g2����t4��єeIY�b���?�I�ƅ>��W�
���P�[��K̯���h������)m��3cR`�c0E�p)���1"���2�d���a�(�ؓ�7��1#+BaX��� ?3�Њ�� ��e�<��2`F��D�)�u��fw��K{�A7k����E��i��ى���Q�G���ʬ,�X���4�`��J��+�+`l��Y���HCjT��j�'��Gv�I ��-6+i�E�1�_%�5e��on��D'��ϲ�����٘�F����� do���?�z몂�~ce�����,w�~��4��e<���"��]�"�|q�*�@˚*���(c��K�� Y�&յF�/�s��K��t��5�Tй�w����,�zez��ɜ�F��x���FxV8%��4J`����ۿ����{�V���F�ʺ��n��"�%2l�H�$n����lp{�^��6q�8TA�˧�c�5X9<���t^�<CE���>���gv/-����l�y�mVr�md�*6>�� �bM����|�:�8�v����n9U-��L�v���<�}T�")����@wL �:2&�{�X���šNq�^���������K$<!�=&�Xti
�Р�ި<j"���M,h��[Ϟ�!���`0J�P$>g�B��aѰ)8��Y*�����5v�j�����~#��s� Ys��;��z:ޯ՘,��^�-�7�� �Ǖ�j�s �h>�s5:(����Fb�Fw�8.�lF����R�o�~��(�:�cPɲ�Y�׼�k�[�vDGcS6b+	,�;?�hu<��0ϏS&ǌkhQ%O	�q����^��:�w������k�_��hp/J�"���챋3��k��g��`-�N������S�H��h���y�F�������V����浯.e����d#��a����zA7`3e�1t?S��ÿ�W)����OV���<yX��P?;A�A�61�ٽ��`}���l����El���QۦoX#c�ɇ�bA��\���^F�6��Ɔ���0X�t��e�<\ 
!"Ļ�K;�""��m����4��J� ��ũ衵��x�i�v�'���䢗z�=�D��am��<��Q$s�R`���{��!V֌����욲� ����(BM�6�x=?gK%�ù��374!�+�0/g�0 �Ѽx������ ��N��FY���ZCun��PU#�^m���d��e�ǥ��s����n��<���j���!X!`q�ݵM�`u;}�eS���H!r���d�,��$R2���uU{�#�� �Jr�[�����d��$��>q�v�Th<���y�k���]���d+�3-X�o��%ť��������:��a����� P���:�ҧ���Bqy] �Y�V��j���[3�N	4`�(�����|��������3$Iӥ25�(� ���|����'}�����?���Q�l�f�K�*�EH�7\T���z��)�Gl�n��<�ҏ:6��jŅ)!���ʉ��7��\���}xJ>��9����8&R؞��U<@t� e�(�fg*jL����т���t7L-�&��H-̫J�ji���?�n���քV���B��KtQ�8B\����k��:Y��Gl����y7���R�Fj��o~V�7o��)�� Gd_��tq�ȶA��]I�ݖ.P��6xQ��z���� �V,�B��;�~�K}�_|�+�[pX��Z[�)$xnɌFM��cRBB�u�
2(}S&�s����jbٿ�	�����)R� ���e}{'�?����(�z��3t����[�Z+��(��~��Z�k�3
��~yJA(�	{%B_:~x�<�]�Anp�^Z�8X�u	��a۶s�c�c�F��k�}�ƈF��'�E���G��5��ve�ʑZ�c����'��
��N.[M����7����Q+�1���+#-��<H�Ǿ&�}�t��~�4�c�<j�Jr���6����O����p/?-��z�����ѹ��[�&C�(��b�u�
�	m��<��3lL~�u���*��V�FK��*���*��S�|����@'���`�=�:+9Q�YיԶ���MZ�1pmq)<zX$0t:=�6���zγ�>H8���>��C��Q! �BݫW������v�x�/.�"n�]����Z?����J~���'�@��p Nv�P��%X�m­yL�Y=ȏ�k�_<�d7e���s�j�����֛�/tQ���R��F�TA���yzfȖj]7	�Bk9W�6����X�%��ۡŵZӇՒɓY�����1�n���q�Gs��a�y��t7z���@�\�R�����:P�ʐ�+�Sp���w���c?0E0�ӳ�\���D�[E�)b3�Ģ��Q��lD�&�L��I�秮P�s��Q`�RZ��Z���>�Lg��ց�d0!��Y	�C��{�"�~�x.̔�K\vZ��kǔ�$�ŷ	�&�+\�d:�x=�mc���"v'E�]ڞ��-��ҳ���R�������1���vk;�A�./�F�H��Kit�L�n�B���	�&�6D�[l�������N�'�cc솪7���ӡ�go�&�<n�ֱ����h��uN�^R���T�y*�V`�r?(�p+$eo`(R�B��!�sR� T@��}�M��n �>P5[��Ko8�O��CA�T�h���!�l�Ԗ4�z�ߨ�y�	5z���阌�Zj���v�L`���!�c���������e�t�3lBw��y�l�����ޭ�����h��.Vo.��:�3Jg�e�
���v)�o:l�Tw��N#�]=��pe����e�uFb��ny/WՅ���%v�X�
j+����L@kne�jPv��ѫ�e���Ο1�7�����㹮���Vr���앭)J)��Xneį�^�]>Ah�k3�W̙����umn���ѥB��!י���y�0>��k.�C��:	���.�~��k. �,o��.�����~�zH��8�\:��m�$�V�K>�}9���i<͈D: �'��4�g�6�m��lL�9�L�������j��� ��s�H�RvZ�܂�qk�PX#��nа,:c�#�妎Buek�f�m�0b��VΘ�Z=�'���f�(0�Ȥ��E�-嘸�u�9m4W�p_|v9<l��/{S���{�vj*1��D2u��u=�B*ix��P"�Q%���U����Ԏ������zA��o��m'�O��Z(!pK������k.(D����t�bU��G��[((���a�Hw,��]=��U
x�_��r1�31f}E�R:~����o>Ȼ�k�е#��J�x��) ���.zkI`;n��*[�̏�G��F�x�o�R7/}d���w�brn�f�߅/<�k�4�w�������J���J����V'c8?��nAa�XeV+<zC�����-������ K�E�g�\���l��2�tMQP{�����ה��ul�ܚ�Ȝ�Ţd���L.�����G��~T�Hٜ��[�1���٫+�Q���$��dG�S��?��޽��C���U���^܍�74.,셉?'�Ltp����.�'�XWa��1�y��woso�țk��%��HK�L���R�1㙅t	��]�q�m�i�=tF�o�E�L�z'�U�u�)���_J�FVŰ� ��s	�%�H@԰a�0{��;��۟L/�����r2��(�?m���K�-���-=��9���A$<��[ñ�:(̓�&{�e�
}��=��a���C7k�Z��w��rC
d:�yă���H2�@�%0 Pe0��oj7����ڞ?�Y*����?Y��L�M���ƁUAl�M�ƞ�ȧ�[@~Z?��v,
��MJ��td�%;J���
,�4��%ܕ���7�NG���K�����wj!�=���D���ƑUm�F����Uw#�-.��FhI�����ݘ�����,t�vˁ��xʓ�w���A�z�`��}�p8�NX������+�T0��çz-���}�����o�g/�Ե�W�����R�x���B8�~Q���~���q�E�D�N�;�'��O����������%�H)1��1<Tz�!co�>]oMܻ^��+�h��]�!AV�,�gB�J��.p��|V�c&g���Z��۟2�!.:�Is�{O�0=S�FK�lA� �y�<�fе%EVH�`S�d�Z�*6i�M��W6�8�V�s�̟�w<l�o�Lp��� �_��_���毕����|Jŏ�p������taC�a�X	(�Q<XUn<��K�+��,���tf�L�-�؈	'Q� �(�x�1�=�#�^F
tu����%`���VL��{U���{{�gL��]�
4+n,����C�:���xE���mh�'�u:�S��*Y�F�#۠�h��ܮ�V�Q�#�� l�v���� ~ j5����^��kT|�4V[���AA�����P��­�����]�$iQ���'|>��/� M�����B�Z#��.��2&6eޭ�hnt��,�zP�C��͛��g�|-/�.����{���S�0�\N`�8��7�d:��K}�m,�r��bAp[+�@�b5S�=�eM{siNr 67�GI��6[&C_��B�<�Q��֖0���B8*O���ۓ)O��8ؕ�ĝ�Q���䰙uʶv:�=(�r��xy��~P����|٫���'��? SgI#�m5�Hbw��Ƥf�A��:� ��}���'�gC��&�G�Ŷ촦�ѓ:>g�ťG�c�Xu���榈�z��)_ 5��Q»%;5�[�bI0���S�]�=L�
%�nY=r�7�/yѴ�u'5���[� �5���C 8��N�=i�L��V�O$Zra�	Bϸ[�]�馘� �����G�㞺2
}Q]��h�>���CG4�h�lE�;��5kSˋ�Q��ޢz]yL����"�O�+�f��2(�v�@�bg�b���LV�>�z��(cfJ��_��l ��^�CR`Y�)�����h�^� x���eG$h
��Υ��o^��+lw��[�����[�*H�WV����VX��3�v�楌fc��d\�56�QV�]��z��2�Ll|�XK����`s˥�!�w�M.�F�0]6�ʳ���h��5z2�Oſ�3�1�S�2��{����x�o��r~��D�$��g��O�'絏�59(J6(���ڴ>o���h�i�E�Nx4�ʰf�}����{��0?�;\��SMR{� ���]$̊�_v?c���U�kz����;򘙢Xט��'<N���3���,��f)����q&K��:۟n�~צ'J���`L����$.d=�/�w�[��Y��)�"-V��Pp�P���2�U6���E�
�f�#Q�HԔ끥+,zG�$���u�`�q���{ۼ:�n�=��:Y ��{c�;�>�Is����6QM�m��C��L��z#���Z�l�F�a�2����hx��|�:LP4E����.�N�Bn���YT��J����pn��Yt���ɍ׭^}�F�&{l\2;���٠�Aߋ,t��E52�*gj%�k�$/K)f�0�c���U	���D���N���\��g0�*Ȯ3c�,��Tdx�Y�Q/�%��:��Nr.��m#e���U��ak"�{�����j�X_M��P$ds����$ْk1�!Rg�VG�̅�A3����_��v��F#`����Ӣt���k�{DVc`�6C�P}��"#���|��>�T���a�,�"����p]�a�����ɠ�ԗ�V6ޝ�=zoqi|J��w�o��� $��or���6�-�!�kF*�/�g27�9�:�V����҆���},Fw+R�O� &��
g�[� ,{;V�?�I��W6$ۈei�ś�v]�϶͛/�X��4���v���`"��{�/B�#o�J{���;�7b�']a�w�_��jz7�6�Z##�{,ͣ��� �[�lWX�3�hH��}��Ҩa�kL���Aeaw�nS����dq|�#}p��{k}�*�*�#�XJ4?�puH��B4����|A,��~'��7�kx*MO������������>��k�/hW���gTm�4���"����#E�E�h�M��5!ѝ�0�N� �W�c�cd1B�%ڊtAbF��a�W�]���~�?���F//{a���"
����K,.�}��/Ch��#����x�w�-�S�n� pQ��#�ʍ����E�#���K㢲���H�:|�!�б|�떉��V��P@��!��4����O/Ӑ�_T3��d��e�t}�`�|9R.���"�9�*���=V_��p�YFŁ�	��+\a��e_�م���3���\I"�P��
ύ�\e_̽m*z5b���!m#" ?�|}�L
sϋ�
�il����<޶�R��4�$�X�\I���ޫ�jh~VS�j���
w��'>�[�/B�Sa�h�b��<t4<@���im(]�G�����G���r�R�g5h5X[�j�{���%I�4pA]�\�V��-��*����
����v;�])�&*�Ɇ�(@�a�b�Ë�����I6T��{�i��/��g�π7�>���q�B��<��|��x�L#�)��K/`0�2��k���4���5�r<�f�(%�\���nD��ҟ �o���@,ئ��j�;QJIh�5�Y��֠�Vz�4���ʍz�L��RIѱ\CX�z��^�F���r'��,rYJ5`��� >Y��_]/;K�F��KL��Y��V�Q��1.wɽ���hÈ@�EI'����dA��;�Qc�7q,����<n����,��:�XPё�:�����d~��)�3 ���EO�K�ɇ�qPx��ֿ�Ȉ��=��r���Y��2^b�4�	0��&u4�eQ	�q˝g�c�o�X��|e/?r�;��EA��*CX{I����?�t9���ٌ�B�h.U���gA
Fs��@�Uf��Z�i��}VC�6�f�i1�uY���Q��y����xo찖�kw���#�ɈpJ�9�β�<�|N�H��^�p�<Y@)}�lȁ���P3n�U�ٽ9dU��>����>�H��(�J������}���	��x�	�:�R�SK�J�H����nT?�iܻCgk#yBEB�6�����������v�?c��`%��N���h������&�L]��Sķ��1,s�#����0��(��{)@�S0j$|�0�����x�v�o�d'	O���4���}u�	�°�����d�P�&�'%qV�:Y��ul �Xlx �p@ �2�<�9�n����� �F趘�s�FD(ނ���J�����d�A
R���9�$Q��<����P�a��X�1�����9
�Oۍ��g:Ѓ��E�����q�t��̃C�3�����ŔY94x���vd�jP�]�r�6YAKFH�%8ܳ���4�&��A�;SFqx���i��1DK=�5��V��̰
��n�҅�������0r�e1���\�R��aL�UC����e3�*�i4�)l}��G��[2y.b�>�����°�H������.��0�����L��t&�O#�)����vŖ��fK3��M��p>����:|��3nu��\���[Y3c��ʦ�]�������)��&�y�9�lr,��	����g+y'���O��q��Q���:�����M�M����P�h����@҅.�D%�E�PFȆ���#H���w�>��7��|���$v�c�|�{ �˭�\ch��^�;�^�3Oʳanĸ9�> �!̈��syؗ�K��4���C������v���f{�O��G�Mz3H=�zjHB�5��P���L�maMC����d�X�P����޷���Qs��^��*7X���<g)(��4Q����qϵ�q|>:5!��^���ŃnNvwε�b�������r���e�Ww� #8"�HHr�\�?ֽM��<'{kC{�%�x��f�y���1�Ҽa+x�~Ș���#��]&*��4���u#�ӻq�'(�k���q�A�1*� ���㘺�Mj#���&㦳
����qS3��������|�/�Y2k.2��uI9����d��j�%n ���s���牏q��c����1��˿+"Tͣ��%hٯұ�x�>�K� ��
�X`�JisR�����|g� r�.�P�H~�.�,#�_�7��Z�9O?@���K�b�z�N^��n�[�?�`�Ы!�ACb��'KY]]�Ww��n��|$�g�ɠ_�(���\����~�7�?pfЏt�;�z�����"6C�\;�����y=V���4��2��Ƭu���)!����}��/�U�����;�ƍS�|HZ��k7I$\��{�b��r�bT���A��u�b/��"L�.ݔ<ꡎ[ʞ�3/1�ђo������XL�\H[���{(�в�>��W(����;�p�zb��M�#�-
ީ~�S�N���R����$Bp��S� �)g�'
�����+eT\�|��Ќ�����h����04�ga؊"�c�i��>�΋���t�'�k�ׯ��q�<������m��1�|z�0f�y�l,�e�<&[\8����f��4�u��2ϙ�kg����ć��Ê�wQ�C��Kc=�����i���Z�ٮ$^���h�� H��[�I�u�z	}|��ۙ,���y�R2~��;��wW�g�렶qZ���[��_��V�;l��兒�������b|G�f��͇g�,;��J����j�A��W�]W*�j6�nZrY��>*m������ׇl���u��d��H��3�f��`CÝ<���ݠٿ�+�a�AɌh��=�A�k���o*�������=��A�ϻtN"�[��SHlm4�P�F$����;���C�pѵ�Ѹu=TAt�~u���r"�cX�����i8��[r��Et8�^dH�j�E�b�����5]��b\�A,[i�M�4�v�x:�ߛ��?u���j���ar6o���q`�F��L
�� g7%R-֟;��a���r�8c��I��'�1EHM�a����#����5�<̻x�j�"L�Le��LV+�=�������;Y/�r;����kzzO��8A�K���w�Ï?����F�W�,пx��_�����%hI��	T`gSv\?�
E؅�2s�
���xd#L�!kF���6�T9��LJ�iΫ��LB89m��l^rU�����:�}�l4���9������<�9��W	��ܚ�c��:�!}�s7�_|Syeڨ[����	�_h���E5J����evx�W��u-L���
x����p/�Vg���a"��Tm8]W��ߩ�������iM\:ϕ�6�-���tÿc�.������)Ӏbą^��_����&�� ***���gj'yش�������w�Vɠ���%3�Y�聫����
��H�3���g����ϖ��t:��dO�~(�d-�Sr�/��2��^��1I!G���a��0���h�G��B����R�˕��n�"���Y�HqS��z�A��Tn~x+G$N�L�0���O��ݭ\ݼ�]n��w�ϟ��>��;������Y�f���u��k�l�«��\�"���[�aa�,?�&�����B�����v̸)ޑ),f���@ǱRK�����i�]�̚�>N:�^��ü�������0�[���x|�, OTx�0PYҨ���}�����zv�y��q�r��:>{��ݸ�6#�6�y��h��˺{	y���d���շ��j�6�\��NW�'3���uq!3�nx��6��$>J�q�a���H�Q�$ٯ�����߯��i�F\�J���0��F4����541�;`�'Y�(b�F��h8�y�8!Q?
yn�d�A�5�+Ak�ܜx�l��F�����)D~�$ǋ� wx�\��p��b!=?f��Y�/y-�F��6�.9�=�������^��f�~���j����ie��7K?���@W	� P	��~�����N����_��G����l(�3�^�q��Q��ƞϞ�8�f�s.�H�k�mM����V����Vs�=a1�j�,=�� Fi�n�|rhƼ�J?���~��.W��6{倭��p3"'�[�k�L4�k��9鼶��$�!vHڔ�
>G�+^ms��D�S�̥a�e4��#i8��q�&Cb)�Ƥ.MN��RG�9�Q_��HY`?ϭ.��,�Hw��^z.v�F{��Ɂ(׺�rxm>(1H~�����\<����	�?��!�2����&a�V��������<S�_��xJz>��TE8����dtL������nԫ�i^�H��+=�dV�iᡕ���\D���aUx���0��E�f+y,c�mm�5�C+C?չ�iX*�����/w��5�{���(�k���@M�/w���dj�lX��Q^��>??���_�|�_�R��zsK��j9�����(%��-K���)�ea���J�� Xr��%�Q����ҙnP��f�ַӊ����X�g��%�� \ЋB�_|�z7���G �������(($h�i��<SxD8�����%lx�2��N����Ȁ�����=J��qZB��%BP�;.���#��6�+�:�Lc'�Va�E�<~���V<_�r�_��&�V�Z����]D^��r1�EX�� %N��V�W�G�'�CQ����?^���{K�[���W�j�S���&��|:$�d� p�u������<|N$��h�g�r4>їr:�m�3O*�O�3��hM�q�h��[��_��>b��(m���$��z���1���Sk�c�^`v���T2���7O����T}��D���J^���&WW��r>�Y	��կcùJ&��,�ޒ,P9AU%�ݙ_g��SG����\da�j�Y�o�UQJw�=hm
�«A�$��TA��B�"�b�'RT����osg�#cPG8^Tg�2�֖0��l1�k0���=�2uxY<�`t���C/����xI����qK�A{�55�1�浡b �l�I:�s�q ��z4t�-�|��͆�qX�s��2zi����vT I�� ^Za*�qH�����������-,�a���0��C�0VA��-m��qaY(ֿ2��C�"]`7��H&D���3t��~�@9��ھ�.���ōn�p����uC5$�㳼���dJ�(�����!����Bi48�j��P�_���]��+���ƸN���l��`�ċs�1�J���!������DQ ��H}��1g���q�v��!Q�\�A�75Ps�~��� �ܪpi)5vF�md���sxU�=��=g(��a�xf�����y�¨���P1�`�60E�����m=��[	K�8o�*[���̮]�f%��RL�v���XK� b���'6�*��M�WKI���B�5�!�3f�+�x��ۡ_Y�߄���$Wϵ�vxsֳĈ��`0l�v<��L{�T���9e��8��O��ŐA����8|�c���M�!���J���iJ��p�\T��
�Y�P�꿣禋8!�7��"^Q�.�q�m`�<n>�n}��~C
Ɔ��P��D���͸���vd�F�.B��<���OD96R��XC8��w1�sO�������h+V�����Jօ)�M���~8�MUD���5ngj����n�X�޳7QS��}F�n�]��uC��0��üE����2����9�>�]x���A�,��`�C���do�a�3�徑)2�A]�{].�$3n%��d�c�g�04"�W�&ǄA���Y�D3rn�9�;K�V���{�H��S�z�%v/�r84��UE��Əʳ�WR����?S�~6�29��жe~�lT#\���ʥ��h=�	�"��������:7VѰ	�HER��Ll��C��>!�������b��I���g~}��K°8�W
矇ia�W�C����<�
!�wNR�����o2nM:�̌�����͜dld5����!��{�1(y���'#a�d���S.��WY�ˁ��ϣ����W�0f��p
�����\��C����,0ʃ�^.?o�v��bɗ3M���p�U�O�/�YZ<�o�s����W"��#\�6�ĐJ��g�
n�*��fir;x���W<��ys�{��������IYy��n"�
�F�a���^�¢�ݳ�n�ck���bcR���~^c���!є���zHJ���X��<�r~����t����g7�+y�n͎i�ɂE���{ު����([����;;��ᓤՌ\��%]x$��L����<��<�ތ�u�3�8�PB�F���ލ{f�G�/�l�@n��p	�� G#%j~�u���R�Hn���dې-��{�v��~ˬ>/8��!a����86)��u���Q��:�_���\D
ظb}��ES���5,���&N$�a�H.��L.5�?�{�3p9��:����$�&�^[�]N���;$�-��8�}��CB�Q��5e���;-�~� Y6�r`=�H�)*�˽$���F�D���O$2d�4�g��o�(M맹��R1x��4B�4��dPK��j5��p�����P6N�Q�����|�D8)����
!�[,Y�vq�W{��U��Q���������������B��=�B7|�=J��"��'���ܨg���[����߽�Q�^_��0&S9�'GY&��Ѹ���Y�7��_�g��_?�g@y��%(-�2������&� ���m�S�����Ρ���+
�
��C �3�ǗA�/����̨�ƹ��e���v&C�Dҧ���uԈ�����<�1,m�u�x����͞�,���LP��t� #]Y�����D)_�� f2��|�Δ^2��U���ԏ�[x�"� 9`fn�x�H`'� @鿿�w�����^%=J�u-�v�]�'[������&i�y<�<�������i��C�T����AW2<4��h� �����̀�.�Co��
I*q�
���+3R�m��yF����W�C��7/5 ��u�)�p������/�c��\�(�NFi�U�!�g�0@�k!J�r�ҔQx��Ϛʱf�3[� ċ�Lw�+��CU�1R/���,�Ӌ�ۓ�N�������������7+�n��z�B?������NGyz�#I�_?}���_���^����<��4������c�,�7����pt�B�����7��
��N"��R�c�(1���N �\��pY����Z���5�[�-a2��K�i���J��h�;��UZ��~(��?�a9Q�"������!�Pߩ)3^��̓Rm�\�|�a���O��������D^�����E� �� exp�q�u)'U�r�M_�������]lg��w�V6jJ+�w�f�n���<Lo=����J�N�'m�),`0-�%�VR^a+��q��P��S�Q:tA$�.��0l(��^�ΐ1n�l�a��0��P��/X�̓��J�"kZ9�"��Pz�$�v^�$�\yP��.c������Z�)֑{k2�Hq{�+�P�ڟ�y�H���u�����?��[��~����r[�%mO��ye8�Ԑ���^��IZh�:�~����������/��i����@��~s+�Ŕк=uN"7W�*P��u��l� �er��m�(�b�#��(�&��F3nT=α7l��2������mq�<'�Z�T�PE��zuu����Z;��u��/����$cȥ�)y����+�H�u"d���3��!k"���#ri���<^z�����2���v��̏�\�y4>q��J㤉�N�!���չ"��jx~#4{��7���w�Uf��1ݟ�/+N0�zQ�!(D'E!g
$",�=��g8E�iH%Q��N���W�Ie=em8��=(&�B����}�Ѱ����=J��r@��fh hZ!zg$�T��M�I^�}�,��ʚ*�Q]�l�tgWo͔��6}C
�v"QdwBjP6��2�ټl%?�d�F�7�~����'����gy�\�����v���e}Y6�9@:l+�q.�:eo8�(n4D����ӽ4z�\�9'��R������o�,��vuB����0<��rZ?����C"f�CqBI)�J�;[��J�NT�z|.�i�9���6�ͱnz�Vmc������փ٣7�͎��9%#����%�Tx�b]�V��� ���ɸM,���6�����i�b]����ݼYZd�}v�.]>���Uv˚Қv�hL��S7��5��H������Y�/|x$�hj��(1�ώ��5�Vr���c$i�?��gC}�<z$��.���x6�3�l���{��	 `��No���Yi�zϧ�z[���O��~ ��٭��e _�����(&Et��U拾�JO�=o=Nmo����K�+l�b̈[7�D���b�3D<G6�s��h���l�K5��Y`8�n��5�c�?�q淪����ҲX/ZD�5c"A����0�m]�����@}����k+y������/��������[~���}'6�Y,Wl�]�W���cɊ��r�_�56C�X���3���qK��j���֬�r,[�5l-�����^��������5�f��`�lU2,�s����z�e�/04���B��h����Sم�$��R�_]k�d�ȀAG�c͕�D���{Y�*��A��}�j�	1�����̿�q�Ӝ�mW0�m���x�C��)�<��w7�sq�x���R@♕X|"޼䫐½��t������]�{�bT8-�SR؉ǲ�&.H���R��8F�0�)&�;��R���j��;�t���� bc�#�D��2�b���w���{'x��dy�_LjYe3`��eW� �A�8��Fb��Z�!�gY�m�����b���Nu��Y� ��I'�ֆ!�0�����Q��aa��g�kا{�����kK�|�O1N�	B]Xқ�}��XGs�d ��I��b�N//�gA���o��� k݀�W�����35X'����VL٥˕y�8�ը�ԫ{�\���A�P���ey��s�s�# ]j�
x��;�I�*�z��֤eԷ��4��0�j+�
a�DI��zb�p���'/��P���Cq��T�a�0�Xc�𜖩F����D��w��K��׎bxYԣ�¡�b��8����zT� T���ϠzY�{@؟}[�T�e0��>���66$۵��X��C��eb��.N�������J^P,�\j�e\���,> -�j��Lo�+� U:�;#Z2S��G��ش\P�T�N�Z��tF���Rb?�&Eax���P/�؇X��e�j����G��r���L7����4���]MW|>�B�O�X�
f}Ox��Bd�9uf�I�<Y+D���a��s�o��C��<S�S^�M#�b9K<�����L�A+��k���4�׽+3��m3�$��%���ϱ��&���!�=�N ��{�8� �h%x��E���������r�0���^�ܩ'V�&{�����T3T��޶��r��e�X]��������1W=;}=�d_�h�Ax�KfųeD�lj��S�z�<�0�:WS��Oe�0P�9���X����}���]��o�o`Tz�q"�8��pbW��~���TO��FKT|�zr	T��ƭ,Gޫ��(�O+q<� �L.��=av���鉱��5�J��1�t��6��a��0���8������@1�s��RFn������z�!�a����T��5���H]��A����3�{���QaA �D���`f-����uk�	��K�qd|N��dYT����2��N�+�D��.�����7���.iA;���xtX��������~l���;��N��?=�[�g84Gك�_Mt�ZC]���ݤ(�b,���1��L���r����<{�O|9��s���5�.�;��G�B�ƉU4@6�1���>יִ;��0_os޻�����*R�O��0�h:��To�������3族����G6�.��rVCUV6�,{s�¹�ɋ����� /�O��������_�Goqx�v)B��R&�! �g��(��i��`m�g�)�[�P�*�?b>�RQx1���-���:�gCh/Y�3T�Ѵ�p��h�[*��������c�׈_7:W�W���hh���5��&*���skm*��v �0'op������7�s�!F4ϖ�'#9�ج�[�!��+�o�+�8�r4,�@`�M�@��a
/�Y�lӋ
O�!a��������l[Y���|���x�-��ϵE_���*	�L�G��8��s`�R>����.2:!g���r�a�ՉB{����~��%
�j/4T�/
�7��X����,L<�͒��g�͉�����Y8������%i�"��rv�FL�� {+�v%���(��u�;]���$r�,|E�Z�3맵u����E+����'0�j����P6�nx�Ȁ�PK���x�$ �44�Iv�`�'����mN��1|LrlQ�n����0"B�	G k�Ѓ}�������z���/��t� O�찅g�A���//�j|��
���&�_�y||��v+��Gyy���n��|2��0�eMl��s�[� 19�a�����`U���ߗF��W2;�d�׻��&NV����0PC����/�#��*�Z�)�r*�xV%d�Y׆����N����n���N@��ݔ�9���?���A/�6��p��N[o)�g�S&=�Zjhߑ,��]7x�}_v-X����
�m����^��1X�z ���M����^Y0��4���l�3JyR���Qv��UX�d$�8.��ƹ�4��,�B��-V���c��9�P��x��!���Y�����w�k5<�<=<����7Ǔ�2���l&+]0t���O_�><(ƂZPN����s>S�N�M�Ps���3O��`�!��U���O�6��F
'��M���x�0��}�PR�I��vl|�]���l�֙]|��k����@���L*m����K�z4�-�G�gHK�{������������*\�y�(��C�L��=�/z��<�N�1-ۖ^5����>��&��3����٤{���i8��^]��vC�����OT����j�Ow�l�Sc`��ӂ�f�^�a��F���Rm�Q#��s�����-Ԭ,�F)U�6�ֹ��6�1�wF�.#��,�YN@�d�X����0�,��W��ګ��Dn�n��Uo�H�� ��T�d�����Ŝɔ���E�{�Px�>'��P���?6�ӼIOi�G88�G�Xo6f�k۟�sn���6��r��8GC1��C�=�i y��͐ѴT�Ճi�xd%/�8�2U�ޕ+��1:1��?~�M�c���λ�D���ٔ�DÏTz+3��]!�xĀdlT(F�a�.��zd�\�Q�W˻\�ݞt�\�Gp{s#+��u�Vr��E�h'�uCSl��ޛy ���i����Ȭ7U	|>z��'�4i����
�zv�tj]p����I���5�Ȓ�@�!��M�}S/���V���=��9��
%h��EP7�gq�q��$��J�q�lDh��]P����,�*j����r��+HX���ʊ�"�
 ,-�@� ���0�=SW8�2㑹G���/��77�H=����9�N  ��ڂ"����M��p�Ǐ�~oƭo�k�`�тg
B�Վ6rF�
��z���J'$���S,Q�J��&+�Yզ��^�z�U�]��ӓ�u>n��]�4T]���Z���TKf��Hb^z�䣪0�7�������i�O���7[9?��cY����!��:���D&�%�C�l*�r*��Z�~�J���������6lMY��N[���˚�[R�I��;bnM��l��F.[�9�R~�ʞ`�N��6=�y �YO+
��W'2��8��<Q�f7�KO=�����m��b���h���t���� O^Z�p�Z��u�Kw�?�-�j(�򮜳����ZOW����Lx��#p��ky׻�H�A��XS6�$,pF3EȤF�N�����׃.�s��N l��r�1t��x5�/��ł �8�4Ԃ���B��bv��z.�l!��E}䓾w�F�<:<xt�ֳ��[��Д�$��hԯ��G��`��ֿ���;dI�k�ޢ/8����VYay��q�%�|�6גX����γ��񿽾ᚂ��A7eRc߮^ޛ)�Z���>5`8�`���u��A�Q���ƷfL�0��	��`U gf­-��/Be�^;�|������	N�U�>��:�lW��v������պ����2J��L�Vk�J`�������ck�=�w����Eԃ^�����˞��roQ4�F+Dqaܦ���5;_/��>Qe��!��1��Yg�YW2�l�V���̔��2.�M�R��ɸM�sӍ��	�r]�Õ�݀k�^"r0#�W̋+Bƨ	��7$.,c(R1���$6��Z����oo����
�#{[�xQ��%��$������	�N-�#���ɰ�ڱ�����漗+5P�+y_��'��ޖ˘u�V^	�F��'4ew�﵅��r1�`a ��u�x�A=h��F߷��gѱ�*��uwE�M�;��W��)�,�_?�V�[F�w]���	��∧!�9gy;Y�Y��;��~#O�QO{.�F+h0~4X���2fz�������%�p��u�;Y���xo���k����%��� f�P�aiL�c��r����&��ï��ԏU1�ߝA:	jjDw��ul�h�	� ��'P�R7-����pX�p4�}V�W�����0���Ğ�.H�`E	��#15T��Jƙ��<B�$5& �= w�C�*�W�dB!���:��'�����3?�x,Aҹ\�gr��(s��!T��oNj���=���L(� krA�{�k���볍щ^�u==���P=���C|5Wc:���odv�RCw%|_�t�u�*3�O$i��	��U� a�y�Fo;��7.�#�� M"O+OYG?Ğ"{�u�� ��βq�Ntv<n���?���R-E�<��{����a0c�驐$��7�%h�Zy�P���!�غ��x �R_�NW,�B��_zk��J��;��`��M԰���t8�����%�r`D���ú��L0�x,��-���xsE�EPK7��A�r��2��lʽ1��vt�(0?��FNj6�'�����ƛ',�)u=�Y	c�뵞�����G����r�A���I>nɶ��[D�w.�� �AR���<z�:� �D���A���������ȼGf�;;�B�"�e+19�����;��;&D�Fױ✕~��C+��qA�V=��z=���������x�޼�poI��^C������n�G�<롱�ɗ�/���d�|��'O��馅aQ����D	�&4�F��2���Jㄤ�̂zB��*n��ab�0O0T$HN�.�����:,i��!�B-�#����~���=��0�<5z���w|�����c�er"��Uc��ګǷ���9Jq�Qȍ>�#DB����������T��HpI������"{1��nMW��� ��(u��h�̺[�e�L�E�g貅�J��1fK��A+���<}���L��`��،O�1\�5�h졃��?~�v�_d�*Ȯ����.�4\y��B��F�~����J����j!K��ۃdu�'�^"������G���e9���
��3߽^�4�a���{֌�\>YDd-l0<+�q)y�٣��:3�B��1�5�������	�RÍ�����^�=y�]�/�72��|P���A�'0JZ�� �p��^2e�3F�3�`? � ��� T;]�����6Ι%f�0,a�}�ec��@SW��`�C����hkw	j0Md�4U�~^i8�d�����blZ��0L�@>]7�5�ww��net�O����B��/Q��u�!d�J�,�&�h���O�Dbמ���g]�B7�jL&�(2=:Te�� �Y0����{$ԒZ�Y
Qc5���H"a}��OP`rR8�d�[�_��V�9-V��i�uOL�L�k5����h)&��6zg��(;���{����X�����t�!,.����*`��
���+�)e��l,9,䡟@��b��F`_���b�4�O9�%b��^��^%H��wS����W���b��+]P��[6-��q�g�~�^�9�SG���a�Эe@=-��亞�[���M�n2W�6#�C��I���8�@�}��<�
�Kr`�5�a�+��U�dL�.����~����� 𰢹K��;�AC� ���!�4bXQO�������k=I�f�` {���T7�n���?J	=�7k����zl+]��^�<�pdQ4՝ #
��0�ʏ{u��/4�tl���J�Y�P1C���	ei�g{�&�����d���ьĺ���Bћ���{��Vu,47/x��pu2�{����]
��4�0n�x���a���6[9��̎�0w�y��A�l�C^��(�9S������z�$�j@�ׂ�]Y5B[����@�	�]���'��ٌ0b�6�6i~��bJ������)�l�7��{/��$��%+�����dD*�����%���P��e�E��W5�}�ެ"��Yߋ�G�V<'����\z���3nxQ�!W9�0!���Q�Q���[�S`�ul�^Y�G	Lz��Do�*!xOa�"qAc*𰄡#�rpB�uS,�p,Q梋e�%Z�z_�]-������]�����'=��v/�A&(�4:e��z0j0n��n���0Y��vM�����x2����J�.ƥ�~:1� �$J�BޚY��y|�n�������ɾ����X3��7���� ���[�YHK=�s�K�"=[�m���x�d���lj�ԺU��Z
�@�b�&'������_�{|�+}���R�\�%w���}�,/H8 \�{@�~�/���쬔
O��"@��'fq;��^@>�k��dU�VI=;����Aui�����m��:�H�ueee����ذ� fx,UM�8*�b�������W�x6�*ɘ3�&8l�y�r"x���
���q/�s=\?��\�����C!z�k��;���M��e�������<Y��Z^�um$5�(�_p��>��AL���=��t�����:z�a��p*]W���%6�·�D�d&�
����U��M� ;�������'��\u4jp���O���;Oz]?�j�����O���qs�κ�?[��c��"����z�W_���xS`T7Jf��i0�T�,�i����[5,0D��k��w��	
��������J'o

�n�Jnr-W
�����ƫ�'%�޷��ota"};[�B�zх|��"LR�6���4�n���jmiw�Rb�_�`�0!�'7|c�� Wh|�w��)@�I�%4 ���� �֍��ނ�tE^��A���Ga|�s=���B��?���Y6�ϒk]�7�z27r�C\ȾT�Zy��cj��%�U*L��X��D6���4�e�ĺ>	,�l�D� =���ES���eWz�Sr�v#�f���;[m%_������$��J~�}'ǻG9������ֈ�E�1ʳu�F�6�!߲NX������5�oO�Cޚ��lFϘ�x $�|��0F���4�p��{��+��6�S6�:nb��Z#��u�!�pF�"��h*/��u#"x�Cz��+ԡ����g�a���vZ�p�� �|=G낉Ʃ��s�n�N�op�@'���L&'�A��> o<��z�hE�n���h�tse���JjHȧQBh|J7ݭ.�ܡ9'(���j�F���X��L�V%�G��z-�� E���D�J͇�J~Ұ�.�_�ߒ��fE�~~#t����:��n�y���ڲK3� �iQ�:!3<ǒ�\���a��NI���9��[�Y}������I_�^(1�l���y!х�ԅ�N�%;���5�Z��>ox$�L�rx���1)�W�xk������ E,ks��4E���[]��Q�%]�E6Y�L!�i:I�v��@�\�d}{-�j��ۻo�j ����Rr�B{s�ӻ��<0//�<���H,��Jf��I'��:�X=�B�%_���ŀs�<.HF\����{,��Ի6�l�[B�H��a��_c���3���k8'�O���͛e�؛�gL�S_��:cO���=���
�':7v�\�5�[���<zA�B�{���,f�r���|�C|YMI���\5�l�c�ըmv�LO�T�z�v�����T����FB�u�0v�U㋵ Fő���q�� #�_��B8���&IUÛ'�sFCo{�m�j�ɘG*S��}���
�֍}�
�1����<[V��l)�h؂������Z�o�Gg���ʡiG4�Eh���;xna�_�H��3C�w:��Q��7�ky���;���8��=��]x���yB�w��`q��n��u���}z�\2�`3n���U�԰��m���*&�j�g�N\�"����߁��G6IM	�A0Ҡz1��-ԃ��F��g��a��A���LtN��g����J7�X�(Ga70S�b!�ą���x���5�Ԑ��n�`�����nʵn�:^��-c�U;݌��[��c�IA]4��E��s#����$���F�i�v��/,��P����^"6�T,�f�oK01��u�2�IÒ�'�����P����T%���!)ݜ�l��"*���ѹУ~ޕ����`\��Xo�������1�5��A���s�؞axO��3,F	�J�jH�nO�L��k����Z��!s�^�kV��L�J?��!�#��%�l����C�f�;����P���NwP~�x�	ɢ��ǭ���t"��߽�!p���Y��#1ɉ���A��w�`�4s�p�"=�%�V�Ђ��G�*��/���m���y΍�_z�a�"W�';	��Lo�w�-���_�~�)�i��
\��xNNzBr�Ϧ����),)���9p��cT����
Lq��?��/�@~@���3`9̚B���|rz�� X���J�	�X���Yo�7t�H§�r/'6.�ՠ�'?u�
�	-�y�.d=	�Gè��wd��!;7�`�����Jne�F����ozWเ5_V�U��(9>4�q\ϓV]�4����0-A�t�ql>l��zq�Ylܛa��'�P�dψ,S}���$�_�(�z�7K=X��{�dyX�t�'�ھ]^� �|��L��5��X�ٛZ�΢��ܻN7�n,$O,I�0C�P���2�-Ў 8�d;������J-�����:?۳\���I��O��j�xD����`�4���[�?�m�5D��E!a�]� ��)u�&f����u�W�NM(ݪ�f�_�[�����jDO��^��UT��iy�D�FG�Y�Éa�kx>�e	�L�ª@Ͳz�S��+�wY�bp����U�%�S(�Ld?��a�p^Q���8U#�A��m�Pb⇆�g@b	 �|��j�#Z`��ut�L�D���0NM����A�	���3��w��^���������+ݠ�u��8�1����C�$�dV���d�OP�d*�0~�ۼEp�\ZǺ;Y�}��_�<�9BJ���.�Z7�l��I�j�L�� gѵ<��RO��.p��B����
�0(����N �_�]+X,\��ɣv-�~CCgN�g6�&`,Z��7���E�������s���}h��L
���h����D�R��$�]/�D�«p��.C�'O�ǀ������,A�7;����H#+
�ڌ0
Y.�;6aƺ@#�0�s}���Nvj0�@��P�v�!?/�|�ֽ |��B5�A��䰈+�yZR��%/�/)�m�9�	J�����R=�j#wꝽ�Y4�}e�B�`���VȽ'�]s:�Q/�5�"����q�Z��A�-�����'�?!d=譟ڣe��_�ԋ6�a�֍x'�B�AwS�FC�	�i��:Z��?�\�պ���0Cb__�u�)�:ڽ�7�UA¨E�
4�3��B�gJr);fqX.�p���i43e�0p<�T�8B%��[��1��bz��J�6���>�����an�t�O���-慑o�00���Wt7��]�4X-EϮ8��[�y��<���0�=>���2E��p��ܳNH��6��}y~${�˗/�j��^���ݏ����,2�
��F��F	KE������o/��PL|�#{3/jL����&(	um�R�0��Q lB-�i!�X��A�Bh����P��
/���z0P�<Of2>��R26L��f4��
�5��Pǅ6Yi�E#�,ױ_���@���d���F[5�z��:޿�~�k�s/����"PM4,d�p���
Y���-m�(l��z^Qd�r�'-�b�eHM�?yØD/ tB�CK�YG0�W���,y�Њ�>�~f�gk�E��n������:���)V#	���,�Ʈ4t���p�ko����������y��Kb�E�#�{fn�T͂{]{�/|e&�ڂj"	�7Q��2���F~�{G&�"T�9x��"�7V��R+�(@�R�g�d�vf�V�����V��-�h?�OБX΃�AS��="��fFi�Yߐ=ab˴�ʚs:N}mN�����8� ˦��}��gsY|Ǆ�,��l�Ɩh��R^[L�|��'�ӡq���T��E�B`C�D���$�B�.�:.%�r�b$W2�&E�2���,t=���@���a�Dnn�X�7�5���͌�`?�$3���q�(������Z7d�A�Xܨ��&�G��fOp٠0hfZ�R��,W��[�ή�l~\�����qg�R'|ރ����є9�7��j8����G����X�cy�<5:~���µ�!��o++�A�������e�R$a���1��=���^G��2?���F�<[�:���xfu.Xĭ����(W7k�R����>��L�H̺��pHӳLk;�ȳ�Ȇ?�@��Y�V^L���LO�e����O%��f���E�.Rjq����>�Y�\�D�wI�@���D�����Nc���Χ��YQ�c�o=�Ԙ�:�' Pu�����|�nHZ�<���� <'�Kr-u�Y*G���~@��~{v�V��^�1*�j����O����[�|` ��t<z��Jz��)P�Vsd�W\S3]X�3�\ջCV}��g$��Q����{�U�_�T��L�?۸�s�ꏡb����T��Ȃ�@cj���Z'��Ȃ��ɳ�0t<��z�̲X����ΐ�a�V26>i��P�Z��4��~����I=�B>���굮`b�Pm���0 9��:�i��ߐ؈&�gd� ��0���9� ����0�˚��rC�1Jq �c�������&,E�$�������JSsF����5a�B�(�t�͓�[eQ�[iH���f�<�i�J�u=���1�ձ����7����~w-���Z��y;Ȑ�jy��}EM.��� ��'�s~ܐ=����
U�3�̌���\2��H�agR�-8h=[�;�G��{~��%|����lW�ި�R{UJ�9B�D|�g�<0�G����j���GHA�Q�,���p���SgeR��&�d��7��B�Wy�i
�b��)k ��ÞXqw6܎
"��jIN�w�m����`�a� w��ek�����![�'9�Fϒ��@���O�aqO�w;#Л�ߙU/Viҩ�WoU<�/EȈ���h�H�ݹ,�%Q�����	㻘�y����`�Y��Q�L���b"8�R8a�h�����6n�~5 �)�������`��ehXI�o�샞�X{px��H��^Ð�5���9s0Q�UO�]Q���Y*��d����9,"�BX������1غ?R���^�Y�S��j	(*��}~��:MO���¤c`dq*1s���:�ZP�x�M�!"i$���@��b�o����4f�9��"g8����www����%�In�􋅈争X���$>��u���,)B��~>�3��w8����	�����::��0$��?������^�R���X�Kc@�y���S!n����w�|�{����]�)/g/�kf�9ƺ�q+�d;_��Ê��W�/n�.Z(!:s�p��F5`�T%t�RE�* t��: Ƴ��5��#�� �b��Vg��Om:dSB#��
}N*�h ʀ�m��l)1t���'k���?�Ia�cPY��m�,-s�L�0��O�Ճ|ɮ�b:o��B��Ϊ|��j�@��a>�a���Z�1o�gSn����J+��qQ,]|��[_���-bu��=u�?��X:۞=�������3Fa)z������L%�n�݌�4��N2���N+1�Y�B�V� xD�Qț�r�'bdDM����`�׺�����P��p������G��<k�#���ŀ����(�����/���͵K�$6Å��f��	��.�3�����z��T ��zƙ��-��G5�,��yV����0d�|��1�*�c�։.�3|����===9�h;xnы��L��x8���p��>�(.���!�$��˙��{%C^�|��@O��d����:���@M~[$t���T~X_�1o5������zS�-ʞ�B���b��y̯��V7)���O�mxo�ct��0u�^��#@l ��v09l�PK�������'T> <M�93�s��z�;)�]����1<����9�h��$�q�"!p:�xh�ڢ�~�IB�I��	y��]��[G�CXZs%xJ��:v�!b= Q�5TGD�l>��U9�$f�䚗(�������0�	Z�L?��f䭖���.�ɲ��AeY�@AR'�{T��qa�k�L��a~�g��[����S��{��O���
�	��
���P�x';��
�Xɍ��g֘Lt��湯=\��^^�S�e6Y�z;���a��t1 �8S\7г�d	�g�H�L��'���.4����O?I9]qcn5��[�\�	���[�uN@s�)t�6�����V(������4�=5�s�1E�Y\�RèA��-��w��e�"�V��u�K��K��0zq��]�u� �6���G�߽Q���eCc�Ul�քI(���\k�Z=_R�ꊌ�)3|-�n�i~X_�T~O{�FQ���ck��'�m4��ֶY��\�����o������ѷjH�T��)��C���P"������Ǌ���|�<���S��\v^��R�4ަ
#���ai`ΕU? ���ۂ${:�tֵ>�V�ޙ��l�,��E��a��ؘ��
�E�9��$:(M�`��6AAJ!�a���u�35n��\7�mVԎ{�k�����Iu�d,�|�M���snd��m�:����õTY��\5�z˺^"��Hq�>FL�]h��zi��h59Y.\�	�y����Q��?Ӹu�\?r3l�x���-'-U0l������S%t=,�߻VH�dK�\����zV�T����B�k������	�̾�g=�����N>t�N�޾�w�ox�H��\���)�ȁL�^*�ۡe+}A%�e+{k��4�]�g����ֲZ�N����x{�v�����pzY��gݐ0l��"��v,�j�S��-�>jW损�X��l�ˑ$	#�ր�ya}29��	�4�H��x��>�!Ah5s�]X��V#�<B��S_m��g��T3V�d"��t�͐`I�%^�T=�:O�������`�%��uޯW���ݿ�� �ݪ�TO��w?�R��TVV�o�������&��N�e�+sbҿ�͊5��A[��	�R�8�I�N�\{���X_��ԆvOSc��O��`3�̨sqM���2i�[��o���4Ww��23Ľ	W��$c�gu�/ڐRH�^]ɭ�,�̚%n��В=;е�:�>�9���B��K�K��L,0����-�p�	�'JY�\���Z�_�!g�7˴`��9H!�6=<c�W���R$�/>�Ÿ۷�_�.Ov��#��5 K��F��3E�6���|^��t ��y��:ܥ�^����!ˁ�?�":%c�����>\���N��~���~��(���1@Tԁ.�ؼ���%�Y�&
4���&@U��U=x-�2z�r>�6����s9�����5�@��Qc$���q���yi�c�b��*jD�REAe ������y4���po����$�l֩�9� �IG0j�����!ݪ�"�ίË�g�AWkf�9�V�V�0�(�nu��	2J'�\�w�`�Q�tN<c��R����g)���!�P���O&���V�'T;9���l�y<b�Cc	,R~F�sMb_l��t��ܘy�c�s�7i/Jp!z���u�lO}���]T3��?AB���=q�U=e�-;��RQ�MQ�pN�l/�klz驅�;Cs!}�B����^��ǫI�A�5웬g�������Y�[s�޷�����afY��3�z��jY��ST��y�wv�.$������L�M$�p�!�X���]��N99u��Y
'����sWKS�R�m翽�T�[�n|���Ԩ��46�e�<[=57���ڤ��Aʮ�b�[�U��m?�L��ڵ�t�����蕞��x>��8AfH�r�$���Iz���ݫ�k=�:fY����'`.�9��"]q}  ��Z�`� ����F�]5j0hu�>.�mہ���~~���ɂ ��KS ��0T�P�Ǥ������|����^e鵽��A:�;q���,DĂ#�Kl�7�Bw�'wl���:[��
 @�C��!B"��uCLuu�c�$������Go|�#��{�����롪��ՍՀ̐}�k��?���}��j��s��Ut\7F<��'�t!+����%���e�:�s� |j�l��e�3�FxEԂ5�=ꀖL�dkx6�ɕ!S�H4��.��0h��R���#Ja�u�lE��a�Zx�ꡡl��9Vsyw���+=��3�RϸZN��r�a��߁��ʲ�$��,�G��~w��8`���F>=>�="�ѐ�nFm>���I��Hc�:��+�����nt/^���"���Y:�d��y�dk�#�9�#�����Ը(�j;*<���FxP����]�)o����G������7����m��K�z#�V�i�A[��H�L�ٽ�N��L�1��,�_D�V��ga��:	/��_�<�O?�d}���=�p³.(��t	��<3�Il��3�q��_�k{f�Gd���QC8�-�O�d6�`+���?�L���ȟ��㢶2 ��	�������;z�q�,�tx2���H$4.,:�r2&p'��7TM�^�X���4Q��F�����@2���T��KD2�t�\��2eKAh�]��E��t5��n��|���@/#dw��ҰQr9���� ��>��O4Vg4qy4���q"nC1�r�p	J$_���dYY�k�J�k8p���=)A���Q]��s����UN ��0���y�M�����~�}AR;�R����r���J��(4h�b��q �O��YrӲڢ4�t��%�%�[����3�*�o��<����nK�B�[k�5�sb}���P}w�߿<?���Z/O�q� ����@��։�p��G[�r����2a��$`z�����~�ð��4��[2���b��ɸM�7�FH�Y��'�"��S���>�8iw�A6�HS<�,B�K1+�^. O�wd�[a�e`��NQJ��t�uZ�+V��<�{:Hu����� T� �i�t��ǭ�yײ̈,j4e����c	ӧAg�jYM�X�e�0�����nff��`<#Dzx�Q�|�ʱ�����P�����_�CZ�:�٧�BLzi���΂2���H�qCb�T��`�{]jH���
E�{`q~- �xsܿ�����O�)��  'P��0��w����q��������r}=��zۛbG�Z�[�6��Ywh*S���B�e��,�ߟ��-�<��{�8��?�����;�ײZ_Y�]î#MKW�g��]�kU��N�k�!���E�u*��h�ބH�6j�1]�y8JeV����s��I����-{��Z"J�~pL�ɸdb2鬿��=.����~����=t�ZθO`�kd~Y!P0�����ߘT�}i�J�=����v��|�kL6��t9:�ف%z�"�=9��:ƱRG�s����WbB�hۊ�Ԝ/�,-���ξ�{�&���y�m�����!N,8_����	��a�~<N�G; ��Vj�G��1�t��"m��M��l�[x/+���f՘qk�wRw��B�:!���K}ӄ�mL�Ck'*?Y\/^�l�z���Pl�ݱ�
7-�DI]�0j���
��FL$������*���+[���VZ�Ɏp�5���֥�q?��� ��ˆ>��O��P��ᆘ_j��2��z{D!�m��xꂣTٸQ��x������n@�A6��p,�t��nٝn��)[�y*5����u)
2 �� �wA;�ȠGm(�n��O�~���&ơ����i�C�� �8�J��e�j�ݚA�c�vX��50l�5�yZm�;㣣β�umz�����6[)N�y]Ty4��)����3�P�َ�W�ǠNW,�Hg"X�NV��zg;}��H����Z����fR�`Ѓ��5VyU:�-O�/@	������X[��P~����GO�����J>�X{q:II%d@<0�(G��	�0x�\���VLф^{a�A��E��m����:�6��|?�N]�l�~���g�/�io2�"2~�������A0�e_Z�%���ϐ=�-�ș)k���λʎ�$�&GS߅N�Lm:5�b��f��'�|��wo?ȇ�7o�I�FL�V�N�L&$i5��f:�\0���p�3�D��y���@d�w�X�� ;��^v�����?ȧO��ݾ�齮��)zA��j��#v��p�2��&�v���}�ԕ�)u�D!c�cw�FUC��WYX��$t������u[�ۖ��i)�κ�SC���d.�J{��z�P�`�G�b��b%VȺn����k�`���Uz'K5�� >}�J���=0 w5���E��o(�OyG6��7����t�α�a�,�Op�!�� ټ-4j�����Y�2��T�S�7�<�A/�k��4[o��;u%E/	�ª�Q/�\O|���������{�
��O�+�K��~I�EeʪX��G*X�u�7=n�4r�A�M`�����{��Ǿ0�HfsY�g�εXH��4ͤҽs�{���T?O��5Y�$�K�Ӧ��i��d��`}�q[�Q{VK��q�2g5����I:�-��:n��z#��\v�z�z��8�u�4���Y�P䨨��^01E���LY3���?�8vtp�,\���;������w�����������uf�z+%Ib[(M��Æ�io��A�Y�F�����Ef��(]��g`l�����p��JLC@{�|�{ʶ{=���������W�5��
�U�}0>rA�q�7c��l���`�b	ɮ���3�j�L[�#9�%�+3�bU�[T�t"���8�"����d+;��S#��r�	 �N7g�vo�y颈h��S��� ��Ԕ�QO�9ORx�1���T�Qʑ��3[6`�qo�</p����|a����tgR̬5�u�,Qo��O���Y
��Em5���~��C�I�-��
 ��ࢉ'fr����t6sr4��+aM(
�Q�pD�&��)�U�Ƥ�� �un2�Ǯa/T���v�P�s�QV�2�^̰y��'y�):�fx��d�0~X?�:���7�"���&B)�r���t$������.Y��t;��}� ' 4e	��̊5j(M��c��8Z�c{��/�T�����z{u��֛��i� ��)x�7O:d�fݸg��.z�e�ă�<,.��80�AZ�^�o��7������F��Wj8����V����񧟙Uv��D��U����cbqƊ?��Y�3�];�\x*�Սܨ�>��tN��`�A��	��?r�FV]��Q�������lY�޷�	i�+��#�#@� ��'�yA#� B��������k҇�c�~�Z�Dd����F!qo��s��k/����No�MA1b�B����O��xd�,�ǝzW�h>��m���)�u#)��=�y/���˼���}Fw�J�=k���D;<���/ǂ΄�*�6Sj��%˕|:�q2ңKd	*c�D�m>�ƶ~��\��������ɢ�䥖7ɸ��>h�k��9�Z$o�K�yH�О���B���M���٦K2��*�DXFX0+[O^D�j���$����:�H�$nu�0�����3i��V� �y�M�C�>�V���v�2/	ܻN�m����=z�ʔR�w<k��w�er�E�AabY�Ģ�8Ⱦ�-�,P&�y���wV�C��B�I���'�F95t��XB}�O
qY�9k�*"��޸�K +�)��(����g�E��Y�pYxK q�����v��n�22in�<�U_)s���`闼D��z�R5������+e.�����>�����"S�u�:O35�>����M��3�k>����6}�<�Ϗ_Dw���ח�t�����������Nȱ2�~�!�{�N�I�#�Gm�rj��m6<'�����&c꫐��f�eh*:V��{FIa�3��ϖm�3yzq�T0�΋+yV����9+�b�ZGƤ,�i�dC~7Rl=�뜭eX��Z02�a�bK�s,�X���jѪ�L[�ѹ�SӜ����:WW)����\n�ȥz���s�%f�e��A��7}1��i�_Z��c���sjP��]�Õ��j�<*x�L�&�8��5��ѯa:{�����{��c��f%8˔�7���@��e����Û�����l@��!�E&/RX�Йޙ����������;x���(�	%aϸ�r^��	�ۅ�s�Vi�Շy_A�״�PGS-�8�.�Y��ϬV��f'0u���)������L� ��lHm�N��ѯ��$�"�LY�������Ȱ�tB1D�6�j�{�P&0����j�y���}��6�����OG�x�A��w�7�tg������Twm���b�(�6pKbZ3���v�Ho/���ޥK;M�|J���]��v�fp�W� �V>n^���Jo~�&]�b����(~��ߥ�}2�V4�G��l�p:w�F}e��G�[+E����ӓJ�I�	�/6�"��bX�k;����_��FcwRD.> "��\L�M�D�^K�K�}���O����F}��,�(]s�̀����B�̇�$9���J����W�̳�5�a��?��?>C�δ!��/���5�'Y�vT�c����W`%���u*�c�f��I�=��r3��;�>\��j!g��������}�d� ܭ���rfe��^o����@+w�N3j]@�)�yϒr�
HP&8#���}ɑe��L�"��G���g����g�Iw�]��n�]1l��>'X�:k�dNĄl�,���*�S��k�,������u�w�H?�Q�|!���{ჹ:��>���b>;�;���Rib��%b��u��y52�*̣S�>�҅ ?��x�3��B�,B@�:�h4$�$���oӇ��� i<X�%�^�P�,@8F��f~%#�o�n�;+]��$Yd��;j�z�=���>V��e1����������I���eXY5���n��A�RE����'Һ��4���:�#3ğ*L
���?���h�M�RQ�(k�tʏL�����Ґm�Z���E�s��]7�U������y ������6TfŬ��4v;����/VB��3f��9��<����l��t!���CArC]#f����>�<�'Tf�z��{��ש����>�Ab\��LyB�{�-��҂\=u��gp���ەL�V
�no4Y�y�����Y�Y�A<WAs^T
ݗ�=�!�����0=����rQ0��U�CIW��"G���wqOa�����s��k@�u�|Xs&�������R[p<��I�|���o\��>�!J��t��1�|I���~`��џ�0��T1�g���|�FIܫQ�@�4E�^�+'��5�g�H���,����G��ܾ��tm�(��"����ǩ�G��� я���m:���l	�Nm&ZPGf�&�`��e���[��������H(�RX�I1U�xXl���J�{+�Oi|{!�	8��r����,�n/nR��r��B�f�+Ed����$Z��|Q_�L D���tuycY���|&�đ�c�K�ԃ�e��� D��n��!H�R��^��yum��|k��9p�S ���\�w�s�0��d�A#yFFc[ezs�=�Tr��,]�a���G�(��f�ń���s ؈�RE���~�g¾����-�$G���������.Mn��\��%��_"�4���|l���>7v �$�d�괹���ݧ;e﷨RX����U�u��d�yVI�)@��y�ON>��v�:�$JZ�Iަ  �	?�����=*8H�ߍF��|�d1���Y�]Z�$�YL�'Y��ݑˌkY ąOm�v�=מ����h��_m? 3���S�΍���z�d�Ay�Q� :��V������v��uh�iB��6�L��"��R}Ad��#�-aU5.����W���6��ͦ���wN�q�">D𐁁h��cGYi����ǅ-(����en7�\�E�l��v��\���tm_<7��ŕD��'5�8q����(�K�~�J��zds��N*`r�A���S9���<�b>�Q�-�r�Ȝ��J���$5X��p��L��)��I�rC�`!�"�d��ܷ������呕tٰ�"G���v���e��W~�K�B���4�}%m^/����� %e�����g_3,�7gv�g����^�}�FK�<�j�b(�l�Ц�Œ� �_6��U��`V��ӟ�\�"I�]���o�h��`����Y�b�TdM�~*�e�����U?��d��D��G�~��R�������~-9����p�d�W<�i(�hT;A�ʀ���=�bM��,;�*��e��r�Lo�`}w}�?��_ν�S��lhF�6U�������}�❢�J�Zp�h��Ad�/�2@�L�q�OS�|�%��:�a�~]��K�J[��m�i{}�sM!Ћ���Z�l�C�ݧO�����ܺ8]*ɫ���Ԑ\*�F
]�4 -�������Q�i4M�(&O�ĳ�۬�yH?=}�bZ�Z����ΐJ^����
��SX�d�"j|:�i�SQ'j��;Ґ�G#R7�CWV���|��K��u�8��xO9�pq��UM������el�B�P��z"@�=���x6	��6�x� �;�|Å"�M�G�s�}�1�l��ѿyp��I���+i#�W1S�(c<a?'(C��SY���	DL9U�Y�K��v��&u�\��-B��@)���E��(���e���`�����rI�e��y+�vsi��r��k�����+��lr�<�MA|t���ʳ�7�j��Ѷ_>��x��EF�׷�����\>��^�J�����{�8ɒ�9}J2��Wt��wr%j��&}����!�}i�Ke�F��0�>�_��tx `gvPJ�LU�|�)���>c��/�O^d����WO@��I��On�+`�./,����j+��g�_O���(<�R��:�n�ұ9��m���;"	B��w�`>��|W[�Q1� �������Ϻo�����V��\�yE5�y�>��F Ք���G���e���2 R�no.���O���yI���~z��>�_t��'�\�vͦ���o���2��3�bN�k�>?�l��q��5�P��9E8�l�!'.	#;���6�M�#`6u˾t�z��蚉y��ǡ�E//�g n�QR�M���|�^dW���H�/�~��<MZs��e�$b��,�?���9��_z�9O�3��]�����5�ػa[���)C��n�g���Z�W�u��@΍+ܒq�~_�l�ٽ�ܦѲ�K�X�Ȁ�A�ݹth���V�$S��7���=�_t��Yp� �k���/��j>�C�A��N�0�����
��٪���ݧƧ��3O�ѷ,�Vn[��P���E��
ư.f㴰̔��x&�LY�S���0��Nٍxؘ9s���4^��=a�v��Ǥ��q���ah�����F�2�&7Ԏh�^�[c Wr���>���ПӾ��2��(2o�g�~��3��'z���-RI��yn!��E  ��D$�����?3L�vd)�چS�����e��Y
<=ֻ<
 өP[�W���Ս��i�����C�M��H��c+!�-�{ss+�r�:_v��[	�[:>���(��%#�����{a�� ¯�a�5����<��>e(T�F(�I:XzN����1}���5{���<�<m줲M��,����%$�A�CǢ���9#��Y����0] �5�������QX�Ss��$���gI������nP���4 ��I��������DM�&�CT����8�2͝��b��'C����W_��w)F���*}�����KQ�����(�-`0��F��g�d��R�,n�[; �>6�������©1���IĢ� V�T����3�'�@D�Ү��p;d�N���o�M��S:~yR�!���J���%@�G�1@����ɟ|fJ����-�ݯvy_&V6Zp~�{N���q6S��;_W���ɴ�l�W�R�pL��%�Qa�F�V϶酇[�<QY#ǅ�*�l��2���>d��l�4�hG�n8��~��8��;F�Vϝ�B��X;��̝��maYx5�ZPt����� ��ƭm��-��]�d<2p�m�E_�^���w�+zT�rl瘥���+���kO�{�*pЫU��a�j����x�>�.��EZ�fRcpw��y��O1���Yf�ڸ�v�g�����i��}ƻ����K*.U����a/����/O�⼔i#�ʯw� H�r��jXș͐U@��r.ys��Y��p!�=g|}VQ�~���H���X5��������͇��yv��I���vVEx>L���a�]YФ%qX��@�2�B��ͦC�ݫ!�ngj� l�D8=8K�4�`����TЛ,;G�˵cd[31�|N_��`kBs'<�.��I�w�xן�����t �X{��m����}h�@Z`#C,�!KZ�[�dlG{}��ݞ�:&1i��JbA8�T���t;�6�:�,�g"��҂�8],3��[b�m�lݺ�Vzn]�춍X[��j�:����ލcrp��:d�}x�g�u��0{��d����Bz�`��G@����Ӭ�un婵��bY��_ZL-�.oJ�z�_�-ل�)�.��Si�r��H~�L��Q�����Ý�_X�L�Pz�k6��\�O#��R\���<��5hn*;� ��}��G�L����<�)��Ǆ����$��3_�՛�_�M||N��Oµ1�lm�L���+����#b�GD@&�]��Uy�y��v'������Yw�MHjO>7�郓s"5�\�+C�F�Y�����N]��	����\�����*�vM���S	�:�ڇ~��L6k��ళl�͂i@OJ�D��3ɶ
N��þ�$z��m���+1=����͡w:V�2���(%&>Wӷ��F���=J��5|e����Q���j}��G�'W[1
�[]��)���&���H��)d}[O���v�is��Ȃ��t۝�RU(�d~){�܉I2t
��h%�=�@g�v¤��2Ԑ�$�� �����ԓ��q*�^Ӯ;O���v���~���h�S���ߣ.A��ն@�x�K��F�GɈ�u�,Ȏhg�ч��+ڮ��!�thG��2����ùI��@uT}��[y�e	�k��S�ą@6����(�>�*8gm̵����	T?�N���ʰ�X� �0��υ�T�٥�`�*�)Y^ 2qn<=#�Z�0FJ����U�L�N����T)i-�v����?����?�!=��e,�8��d�������K��3�gQX�P)��!�y����!��b�=S"(e��sw,�j�������9oT�KuB���t}�޿�{�I�t�	���s�O�9h�99����JX�g+l;�EoC-��:J ;���malW������l-����Ӛ8	�A�ƭ�dCɰ�썍I���l��m�d-��Z{.iA�|gȵJx���t�����g5�a��a�~X��+�~w���ƲL,c"\=YPK�l�����M����,�Da^>`�  ��AY���C�H%��ﴆ��o��ihZ��sL��d6���ɥ��h1qhʒ/��撫�>�Y�*?h�a����D;��_M\H�
':p��>���#A	 s��37[�V�7=��
��G-��Q�Ue���m���2=W�3���}�̋�W+�"dn�r�P�.�B/�3J3�����9�z�Ʊߟ��A��n��ۻ�R*2́�l^�?�ot�p���z���,���L� t������A9��@c�x�!R���q�	��M�Sԉ��A$�
QbR�t!C�YS+�ma�Ɠ�|��4�3 ��!pe*V�g�d���A/�\�fX�лKΦ@�k0� 
�FL��x�q=���ӕ?WU� �:�
�l��#pgd,��م�{����8���5��Z@P��\���Ɩq�6����}�!M1*%��/��e�o��JZϓT��\,�5O��Q�6�g�鬡G���C���z	�0���*���Ԛ��hj���~��y�J��8X��&n�M���?e�6���ڊS��JC�j�R	�B�W
v2j�k	��G;ZSp+�`(8�<N�Q[�
�:�*;Y�A�j��D��ZA�{IH�YJ�yT�E"�_>�5v�'v]��D��{ݹ%L� �W��ZA�h���1�������7�޻�ޤ]P��]��ұ-�pLY����.���7�-h�U�n��8�pHQ|���~��}���J.n�5#�By6O#/�	b��8[�'���#��7m�4���x��Qv	`Z�*�G�2ĩVV3����Uv�ޞ������S��AGjvͰ�s�JF�2�8au=#���*/SF�ZT=�<-c��ӿ�	m�|�߯c��
��ɛ�Ǚ\Ƥ�|�z��9���}�Y��_�'�Ge���I��K�b(d��32ZĴ�ı_�L��NϏ��(�]|9���F��'�|�&��/�J�X߿��(��c�R6:�{=��5��gv8�I�v���E�b,B��~�M/�i��Z��ϢC�bp}T�:��5#�g�9Jf	����l@î�� '5�&d��]�Q�.Y
pjwVQII'L�x]�6�9��A騁��`��"�2Lb�s���n1��Ժ��hZ����a�����IHŵ��6ɨJ��H�|�{`@�L�b)��Wj�IO~�~��[��dne��MyJF�Yz�\7�v l�%+'A7n���)��:�z~������J�;|H	\��"ρ��ڳ���FP ����̂�7�&�R����qw�*
��QC��43�U=[ֶY�h��aB���}�F�� % %.�?�������^Y[�['MK���\
	�Hʩo�pST5��Ќ!H�B�S�j�J�����^�W�z]���� �{P��$��=f��\���9�y��M0��7��mA������^�d쥛E���U&�F�\ؑM�>4�AΡ�#��F%�u�"ZG���u������^vO��~<��	B���b���bV6'�3�����M���7�ߥk��w/ϒ>��B���0�e�\vW���ػ�%�	�.F�V�Y㪁z�V��ə$TI�K ��QL��r���f�2��~ѿ�{  �҂ǒ����*�;�1,�,`�,�b<T-�ow���vr�o�����[3��ǳ�_��{k��L�?���U]�y���%�Z�?�s��8���"gLi��(0��о�l�����lK�B
�R�P��q�R4rb��}q�&.ox����%"�2�v+˵�O����Y%)��)\>)�2��RI����y��ҁ�>*n�"����O@�G;wm�OD����W�Oߕ� ��&f�N�pK�<?=��~�I��}���f��QZlC��<�:�Րiz�V�
(��ޅW��d�^����G�,i|fS�X ��)�_e��2��0�z��9��V�́�1t�L��ɟ�����!#���>�'9+~�^a�Z�c��3.Om�I!B��\T:���ٚ����Nk#ː�/�R�]�����S��������7�ٮ,ȝ+K�2Ⱥ��t����5,���Š�'���,��D�r��3�@Y�p��|x�NY�>�^\��WV�XV�����J_�F�r����	�K]�$\j�8fA��d���%A���tR+ �~`b�Ϭ�e�d6��\�O���ݡs�Jl�1X�}D4�B��i�w�2���������5������.��(R��L��7vK�3v���}��^pk7�N�Lhwq�P�d#H?zT��٭$O�s�JGw�s'�Hyn D��XP���OOǝ����:�R	EＺ+]y^q�Py�����GRr+e�nhl���� $I6��p�����KܻL'^�]��pQ��?z�?��s���:���Wui ��.��$��Xd 7����p츳>$�r��S�A=�(U�g�d��[��'�U��n�Ȯ^��Ԅ2��3'�l��Z���C	���� j6���+��+\�U	�#,PJ��d	�ᔞ���s�
�!}T�����u{YW�(����.{��{��[o^�<��P�_�A���њ�ؒ�OSe��p��^V�4ۼI��.қ�����%�1��lh>u�2���4�*d��|�}��e�:����С 3���wmZ\X�j ��m��TZ%��������6!`�ǋIzo��?�����U$��sZ_^��gX�1Y,�a������>*A��?2Z�c� ����0/ҷoo���WK
��M�˂5>-b������aׇ����]{|jw�3����y�hrl�l}t�2:�7�b� ��P�����yR~)��9t����q:G��RfI�@M'��8;Ț������6�P؜@��n")'������}ɷ�����mh'1������dA���6T�1�㴴sy}ez��v���˟e����D� 7s�Lf?�J�ESR�e��
G�3���I�gq��짘L/��##��g��Eߏ����jI���Wy���V挊�R.sphuWMw2��"�$�T�a(��
<��~3dG93�qyq=pM]�n��|���e�����Q^���b���0\,�Gb�՜�d� W;ç䞙e��iЃ�}T9�5��-�[\+2^�ͧ���� x��V������.�lwO۴�%0;lţ�ܿ�uyP�F#^�t����X�cuV.-8�pl�
Ң��b��	Ӗ����������v�jm��b*�R ���\k&ˢC�ͻZZ� �h�Ii}ܹP%�$�NsA|FQ:7R�A��+M����L�������&A�L�d�C���s��v�����"�k�:��j����%��p��*gD��ӴG�6e���vN���2������=�Y.:�'GT�k �{z|��
p���F�qiY��]����܊���h�PDvo򍻴�t}y�Ϳ}y��.#d�X�	��(Mil�0���ςI�E���:�O��y�O㶓�Li���L%�����.���GsR��f�V�
���ġ|��b�M-W-���T�>�EY��I��}I��GPxU22�\��م|�Fv� ��B����s����F2�A���~���p�z{���U���u5c���M���H���k�{l���3ȸ� �ϰQoo���d{�>��:�-��y3�5k�	�;���J�)>c6��B�@sPV0�}�K��k��r��������{I_[
��Mske���B������xP �A蓸�-��げ�����R�s���/�(g�'R�U���V���2*h�޽MvS���-��~)� �#u��1^�Ā-q��͇���ٳ��n˅��
!��K��#�?���݉�?b�S+Y��YB��a��ϓ!��Uw%fya���^V�����-_�/��Bo.*��P�]�w��U~��:C�3�h ����;�<w���|�0)ި�>����$��	��WǪ�>-�̭,kVG���=��"I�u���[+	��V�O�����/O�0�(��շn6@(Jw�i�=�E~�gBˋ	Sod�]�l��d��+SJϼ�IF���J8��*Nn�L�Hi������!Y��3�/56+ЏC蚱�x�c�7`s&2`�β7�犻}d<y��1f93�P�s���\��L��L��m�W�O̐�����à�N]Ri��d�N�lAR��,��I�T���&�^V�wח��Oݹ$S��d��>`/.jp���{�f�>h[}TtMA�Ogi�ڲ�[��"L��l�ҋ��[+wn�{].�e1kb�l��K�����>�	�ni�T�B;t7�/is�(E�_���E�����:�����Rk?�Z�G���2eA#I�2�S}�����@�Ͱ^tPr`�./�"��T2�]��ut��M��Jj4ܮ�.�Ȅ�s�T�����% ��/��a~PaG���X@!�y�����fgAm���YL��P��CR"�d�~�=-�@8i���̙���3�Ãk��C��Ju gb
�s��[5�/�M��2���q��Ke���<>Hl^�| y��5���'�����q>�$�,��d�i�+i<�iJ���Nb��t���]���|�|��S�A:]��	���p\��2��0kQ�$w)�&�p��_Ʀfa����g����W &�]����8�i�Ut��Z� T$��\W.6�Q��(r�)�4ٹ	sT1�Y��-W�I=X��޳�����7�a����)g��O9u��VkϨ�"y3��ʿ{�>U�H��!�e���|9(����U���P���N�b��I ���b�m��V^�i2N�0*$��k/��i1N/�v_>��l���*ɖ�;���O~��S�:�k� B��]�����˜ϖi7�u�vAR����C�qp.m��Y\��Y��0�/8��\��jUa��0��^��*�\�rXg]�C
��P2p�,�M+| ,���G�v�G�$ie�7eZ*|�o��~7P�T�zkS�n��9v~5a���\/�	��S�DTA���3�f��[+�/��mv�./��>&�Y`��6��k@?C` �`�Tr@�i�������ʣLp}�r0#���5�8e�ѷ�鐾֥xj���ɠ8�A	����^٢��0��{�yZj��Q̭�<�E٩���F'9���Ƃ�U)O첏湴�8�h��0����/ه�p������"c�	�I���� ��+۽Q5���S�������|�y�Ƒ����M'@&��2� 7X�@�:���{<�Yf������zdbdB<..��Xdݶzb2e��e0��|ڛ��~����}�����<?}�sm{<Y�IW��t�����:��<�ɏ�>[ ZK��|i�u-<Ze����Y
�
`Clf�#ê�n�uSI�K���p(˰����2j
��3�c�y�>�ւ|�S9�2���%W[I$�P�v��[��<�N���٭+��\8�X�R��N $���A)e\�{��ZKUy�
p��麆�j�}���>�J�=t!��}�I��m�|��������A��E	�k��|����c)12�oV�6d���;�ٕ͟��?mӯ|��̭�Z�Ȍ=�/;Ep�#�v�;��V��=byr�ƞ�l����S��G{��ЏSY
����lT*�=����b;{�	���2KG�K�h�UOp4>hQo�<�¢���f�H�.J�w�v�3�������-��/^ɡ�=��?@����r�SO���O)4#��P�������D46<�� A���߳2,?��:r�v^V�@<+*�,� ��We�̒k�4kw�Q��>�93�ku.x����E�t�-�.�������Bb��Go�dN�t�����\ۼ^�����6w*�����8]�ޤw��=�>�d�O/�e�����K���Щ�^��j���w�> K��g��j�~_��U0�wi{���l�ʂ`����û�ʬã�����zC=��e`dNR2�z$(H��F?�d�.T�g���w�T+�q��;)�tM����E,]�<d̳@��Z��EE�g�P��lX):�cY�ŝ{�R���f�9����SR&՗K���}(HJ/e�c�>N�@������3~������'����������2V���V�#�"�-B�K^#ƺ��8��*�q0\;�d�^H��"M^]^{�8 �.�5�\'0��v�.X�t5�--N�E	C�~W�S'onWڤ>�:�d��gJ���bcCP�[���l��!XfZIބ�QT��_yZX�L,�2F����ܗ��u���E��(�٫��E/����}��rN���:p'Y$�^��C���Y�){����9��������KH�9DP����SS�!�qv#�vS�9��I�)Lf��M�@�DnWV�q��p?!�_��N����ߨ�����=�Dմ  ��IDAT����V
!e��sK�c\��Zzr`6k+E�[��|4���7�
Ȼ;�D6�Ւ�A��R�!�]���X��a�0�����HT��llh_ @�GUNi}(�� S�{r�]�Ve�up�{2�^��֤ۮ�x���7a��%�\�?}��?��P���>������H�j%�D/���M$�ϫ����c�8f
�E,
���5�W$��;���Z�pA�0�'��U���m���r�m��$Ⱦ�(7��+��"y'�8�T��gy3K����\1�.̎`�M_紖�;EY8�{�-2���+ 1N��%��!Ӏ�޸����{'cS��-���&�H�<�tŏ?��'�1�*N\�S	���w��9�)0\M��뭞_����@}g��u��� c��¥б����(�(�L��3�̓L�,7��% �"�I��@���T+@�`�����$}1��u}*b|R]FpMC����\��du�8�k��x~Ѱ���8jޕ�k�<��`a�B��B���5�c��v��'��o�'�����xg�(H��J��^sz~1v`z�Z����+m�>���R=I��C�ru}�൵�0�ѩs�\&(���jJ�d��j���䛰Ɗ�ь�rV�?	��=5thQR��N�Af�F7rҺb�������)��l�~S�wI��¶/���%׼��,;�iS*����nh��&l��Z�
����9/l�ҳ�8�*'"�!	n���r�P�����(�~�ߥ��L��1��*H/E�x{M��>��έ�Dx�g"5RW�~�EӔ�m�z�1	}�K�M�_��4=�S����-`S,��r�B.��S��}��L�둸��/
$®Un�A����.t�#�i��zG��ɟ~��M_>�,$zO�*._^hڔ�`)�����{@�l�Qߜ�.�/����2;�<��~9��u3f��:G���`R����/7����=����!1�d \�yh�C��� pb���B���x��l�=��Ͻ�|m~�X;K;ܖ��6�9�	�j����ݠkН��y�f�=��
�J����R�C������H�,�[N�8/S�{�y��cz��`���;e}b�*eF�Ui��� �_�~- �����OS�A�*D�S_6<I�=dx978@i8�T���상ѵ�<)]�&�(],C�v�Q����S�K�H��)�BA�"�zfB��+�:I�ڹBuU���g�ItF��TV�QQ���G�� 	������s4.��F��1��ށ����[0�N{
�ĩ������ wί�:��)RC/5Z7�/�
'�^�U~�#�1j���f���F���C���LB����T8e %��ΐO����E�wrk�r<��ce��6\#��L8��}T9�A���.\�M��sa?�}����m�G,�����m4_=�sG"�A�zV���v�s�fCZ��8�����O9LjVP�����RD�p e6��i�C�z!! z	�A�@��P>sΆ2ؘ����{I���JϷz�P�:7�FJ�(����gPjxE� eTD^V;R>��!)����U"��Tw��d-��[73q��.˥K�H�iK{��Yښ򰚏��[��ӯw�U�>[ư�H���޼fܦ����أ�\9g�2�Z�GD���M���$���JO`"��i��f���	��c�{
.m�y�JPi/�F$Ƣ����R�Po�hv��Ҟ�N:��h�t�{�G*2��%���sG��!!KEw�d��� y�5ѯ| ����:�¨�d�n{�X����X���AG�p��+Q_A;q2�� �,���1���z��]Y��mQG0z8�,����`$iw�Bkaa����}fW��y{�;��Z�Y	Z�.wbA���2�l��,�ny��B��S3|����+��2'�1<3����;W�̆�=�IQ��P�xfdD��&�}�]�������Ч:W�8F/���id,DJM~/{�ff�����`b��2�V�<���OI����JA���ݦx�u��nvqJ�_z)d�q�����x>���g�6ׯ8)�d��4�������1iG�����/���)]]�{��uA ��#+��U��$�ͭ��|ӡ���K0*�y<��6\�*�Q���F�4�lD�ڂ��6�̟����鰲�a1IWdy�3#�b�Դ����jy�,�����.�l��Y�Cu�̔���#�Ry��#�pvm��0 a�W�Ր�l<���&�[��R�vV����� G%�l�=1OJw��Δ^�5�HS:l.�Є脘'��eLl���Č�D#Y![-��\,����r�ꂛ�=�W��2��:{p�׌�6���{.r@�^U$�P:6����W�����ƣ�]@���u���\)6xN�<ꝡ�M�7z]�f-)�7�l�j�s�-��4ѿ���h���|,\uޏˊ茉^����G��U���߹ЀUi�6�B}����D��\�L�d|��;I`����h:dA��L\S��+7��9v�b���+��
�l�㤆1��-G�/T*��4H�0j�1ܺ������+#�	��"�����i���3���[rI���<�)B������ ��=���Qӧ����I=��y���6(��e�vbH�)��[
 �<^Ǵ]��7��DV9�/�dd���m?��, �3ʗ�2���ez�@�~���2]֓����Z���tc��ś�����RL�̏�����{X!kE�< ɮSk�j}p+[���n)X�s�#�����S�?���8���������G�Ŵ;�N��l㚉9@�� �x��ߝ&�!k�D��V9�A�ރ����+r�d�͈v�T�x2Ӏpj���������)�|��t<VЇ®�]�M��hJW�C���X֎`
�n2{/�Au�>{��J��� %�N.�r�;oXk�!
��[lݶu:�#�E�v�L3�v������\�o�n&���9��`i������.����m��C/lKW��B��l=>�ۃ��u�e�V��,�M�6x��ѽ��G�-c�������(_{�����������s9���0W�i�n�,�j�Kmf����9ϱx�=�o��##̘3����NeiƤ��ʺo!d�N�&cs�։Y#��:W/�b:|>1��W>�eP�������uUk�W�D��1qS��t�שt/��-wz�֒2/��4m�/�i�|A#0��R)׻b�
�KJ���n�s�<�);��4�����=�ϖB�C��6��ڮ��&uv(τķ`3�:eǍ �U�!�x�{4�'T�ۃW;ɝ��v:�
�5�:'�I��T�4p�Qx��P��Npܤv�)��Ҵu��"�����&�D1B|5y�IS�ҡ+������d�L��H�پ�-ӷ�_+ʠ���%|2j;�n�\�w�v�!Ǵ�ؾ�Z�����٫�?��p}Ⱦ`|��[�¾ȃPo��&�DقE�'K���n,�q��d�*o�iR�����[���R�SkFdG�.��!N��Ӆ}R<Ke��s�>�X9+�k�#0f�RT���j�'D�v��)�V&��AQ�=2��\�	Xػ��γ�}�vYH�3�J���D�`�<U���v��^�qI�D�-7��#�^^�
:��~wԬ�Ѓˁ(����|o���E��:��� 0���~�!��୚�dp�f��\Y�w}kϽ�;�el6kW@ə�h:h��\i��~�yY�ۮH��4�|
���ʝj$(�K��['�saPB����(�ki����Ȣӛ�\�S������w��<Pg�s�=�GM9�R/zj�gzL/G�@�0�$�W���ޱtOR?��ʱx�J*��)���Vb6���mI3��Zr*�"#�̖�^:&��\���gyH?�1��W���Q�Z�!���Z��ԓso]I���r����]�pg��v��h[i�����>���&]��~��V�o	0�Eid#�H���y���_��J���8iW����'nQ�@�#g���L-;s�x6�{X����S:�uH�����,�FJ�v*ӣx|N��wi�?�+[D㢎f|�Sp,?��2��nn��x�V�&n�FD6�Mח.��ޮ>2����MB��s�k������O͌�:)�z?o�o`�r���<]��q����$��9Ȁ�"�䩤~7�O�Du~'CpCL ��O��+-|zZ�̨,��:��hW��>4���Nߛ�b���=V�5��d<��p&��%�n%˓�+I�c�'��� ɥ����!s�OP�?��z�� ���a7R�[=����w���>O�XV�N�?���S{�+�,����u���
Hw��>m>������lm�uY�r]�Rm̄,�]�z����Ծ���⺞I�g_�CO���g
��:q�\h��)dr�v%%Yߥ�&<Z�#�!Q�xj��(`U���&������u�8'�@!�~O�ʅ�ݪ�V�:��[1�1P�J5d��,��PT!��y��W�}E��5z�닐��]�-,��'n3��}���|����2�Cs��_p�Z7��--��Rc�sU�D<u-�J�r�H'i�<�9<H���&��SL��c�����kMGi�S��8#���	`lz ��N]�J�/�;�%����AS�4�
,���y�&��[���J��/>2�y0�B��3��=�����y]
���P�-}*�l�Ϥpl��"4k��ɲ��V��ߥ�\^.$��ͻ��ρêPA��f���n/��:K�7l���&��G�,� ����f<}��=^��}uc���r�
u��I�A�凲H2w.�������O �Bq�}��j��>%�޼7�gU,������Kr2{�Yji��|�V��,qt��S5�<KA���k�dz���c�&zo����������Ó������>�tU�ڳ�����`J�}��E����By�Oo~�!���R��?TP�saJ��aIDW)�����ߡۧ쉪âO���ó��ݫ:)T��SL<���&$T��%%���E&@7짪p�tl���/W΍`���,i�o��QwV���1㹆���i�ؿ=���3�*�zv��VE+<��J��؛�'���>��
n�ΒpK��k�i#�jK]�ߤO�'	��B�6�)�%}
�a�;�%Oq��V�Ӈ|6��&�q���F��b���|/��2��O~��H��۟����@#F�S��Mg�Te9x/Ҝ��@�E�&u��V�
[�W����z�%��s%��!@���"�\ʊ�e�6pM�s���Qf+��!o���$p�l����M2���� ��`�c7�����
FC�>��x t�{���֚�z��\B�¼yg奦�![Ł7�Ϯ�Bteb�%���_�28��T��z��-B�qR�4{�]ZНK;���.g�ց���^;���C�%��9ey�K-�z��ve�Ƈ�2��|��Y^�s�}�F@�߼��ǟ-�AtG�`��=>�d���,Ó8�ŉ���>�+�/��ot�0Y n�Q4Dn}`���`%+�vE��.��g�,��7�M�^e�	h�C�}�,�^d��3���2`^�'t���p��Ku>�uK�� ��LECn=���YT��t�b���ge�����nRFpw-U�J���~;��:�ѹ{�itͩHLo�n������f��(���<��BË�|�{i�1u�w��'�'��Fo���N9�!y#�r�)�sY�Q�9��%c�+�G�Y�k<�Ԭ�ք
Hw�y�YX&�g����`��-c�����@.�8�y���;�y��p)_^)��Kx�f��lڥ��,��E���Btdr}�x�ȸ�>@�y �� �ȡ�p�b�YFQfg�G�x�B��͟?� ���ˠ���t��ǗiV��A��wi|���yc��բ��m�L��!�� �������$K߯�o�����_���̷����}�M��ǔ��ͭ&�?|�>�łڿ���:��?���כo��7�l��{����m��5��괾	�oy���vR}�V����I���Ł�(#q�QIA-�y�8��\T8�#�k@�_�C��eq�3s]��R�Lz6�qfH1`"3���X�沸�L��y��͕����V�-,9XX%��C��N���j�'���﷝_݉��+/(H~tQ�k����"z�YJ�x'G+dW�����O�[�4!(��@Jg�5�2�{V^�ϛ�a�H���A�����}U��̿�"I�{TI��w�۠;L_?�-]S���2DKv�4�_?/���ya�k������}2�W�*�g���E��Me���t���}�����A6����̸<-ʶ{���`�E��RH�X�ʍ}�KO��D����Y����w���cy�z�'N�tⲎ���R4Ι����=G[C�& �H�(x����-X�p�M㗭�۷�;�X��0������*}��[������J�o���%���$���M�|{�^VOiG���`�}�/?�����af�=�9�ʽ��Њ�<� )���ý���i���=߿���2��[B����4=��{���0=������.N�x��Q�9c��[�I:��@�D
* ��~8߿�n���v=��*=����5����<�z��C������Ĺ�G��m����~����ZM:'\αX�q����鉜��GG�����E�BR}Nk�h�T��$��0��E�%���9Ť�+V6��([�㰙��y��9� ��c�p`��D�ss_�Q���a���� g��\z�LrF���'k"��'?���/��ֻw�`���U����y��Yj����� �����grӐJ��Tus���-��!�8��ӳ�d����rj�s�7Z��P��lO�(��@7�Z)>�C�^s��>Gm����?�Ò�eAeoץ_�sUv���F&��l�u`����ҿ���g�<���3onoӷ���.��: �`�a=p(Q�M�|��6�]�}�F�xD>���3L1�� �!��@��`'z��}��÷��ͻQ�'�bѾ��"\.EOY�~l{� ����-R�W/;�֡)�k�'����mg��O���6u���e���$�̅o޽OWon-�&-�ޤڮ�
�ƞ�uq
2oJ>0�žm~i^�#��G�6��ߪCitu�lErMuɆ���S�p�ڕ��I׏�^u==�iii���Q�`�2 �m�1m��b*���gQl A3����@��b��m�Ep;F��G랁�bE΢�Q�b�(���T4����2����!j3U� r��e9��s�Ld���mϰd����$�	7�=�ɼX��8sh�K=�����4��D2�U6�	�A�����T��L]�l�Y��N.[^>�5>응�e�/	~��N6��\�읚_��v�g.]��v��׵��a�]8��h[�u_]�P*�@p��/��FF���^��ÿ�W�:�����H?Z)�����M�����(�d����4������i� ��ڴ��Y`�?<��2֏]��C�i�t01�`�ﯡYHZB)��<�ɓ��v��<�sn��8�kD����b��59#�)?���sc���L.n��g�c06��A��e�ǡ���u�H�����9t?|�]�}�6��C��JX
h����ҨKY�w�Ԥ*�-X��W4e.��8l�"Y��P}T-�*�v��1���7~�]`C����
�i[�K8��Y���p���讗���_>i�;7���oE�B9k�ehĠ��"��k���//k��t��'��<e�A ��ڜ�S>o�
q��m.{3u+o��G�t
K�ܟ�٬JT��Ǝ�r���� ����9�<���s��uz�N4d'b89������d��=g��2�y����~��=� ���'ף��+�����r��������+^]�|Hd|`��br�#��{8� M�Nl1D�ޘ�wdQzA�6&�PWV:��β�"]�!B����?h�:��}������������SK>s�NTo"U~m�5Ss��0��Ʊ��*?U?���*ع��
��^��;�}�z�YS�FG,@{?` �-��N��o�5~�$ãZ�:Y){�,>(;�R��g_���!�F=�\�OC8��cO./��w����������	R��ԋ���hI	U1!z��G���Y�v�����kfn��*��}xIi��Φm��� 3�	�i��J$��Н$�I����Y�޼Q�\%������������m<���;+5�@{�]I��z�|�4.JIm�t*�^I�ŀ��F#|�UeU�O�";H	���ƕ4F��Й�X��}��4��?�⹴�c|F�S~�ſ�;��t�f ĝLX���9�g����Z��x�MЦ����>y�%0��\:+���p#2g=_���M�L�<���ʌ��a�r���}�s�Ã��O�&�3����n��`�3���l=�\J�����Z?��w��O�mzy~I����/u��^��U���"�'��)4���t=�I������Yغ�B�ٲ�FRݍ�����[0e8��1��Z� ���ϫgeoE� n�EТ@��mde~���0p|�]�뗂4�\��<����2L�a!'�h�ں�JW�}��Dd��B�>�lJ�T.�EX�Kd*�$��A2�\�
{�o\��\Y����.�L����qQ5>��X�����x�c۴V�*��JO2���d0 ��߻v��(����T9i�Ҿ.&����ϣ?�/S���n����X�W��t��o(Ղ���������]�OJ�!���$4��dQ��KÉ���O>������VϮ-��z��2F��Ep���M|>L��`�s<-�У�]eQH~^V��?��g�8�~���L��$��̌`�z (���7��g���A6�����b1{�� ��� u�x����R�oS��f�G��f��LCa$k��2����M���u��Vpñ�6:��f��v�N��"�y��h��<�0�&kl�1p"H�����O�������l|0�?���gA7���~0u����s 2�qn��I���HY �5�"sc�A0�y�V/��������!RNm�q��M�T���/�{m
h���ץ'�+W�
h�uڳ��K/�B�>g�j�F3\?X���@���!�%�F�71J����̋�����C�е�ߵ�H��㜑S�۳3I~���8���}�P�e���9O]ʨT^pab����A��9f�^F]r3\N5��(6 l6b�"r�c�,�sqЮ*\OJR�evti!�\�ϡӫw�U�ؚ��~�ͪMs��E�6��N����1cꆅB:eS^�ƍl`�aŹ��95����!��{ή>�{�}��{����`���)����a�ܝ5��!�����}���2=�������3M�G΢�1ȟ㗰�,F�?k.����^�������X�α�\4t�' ���Rw��m����1��?�>����a=	?t�Ni�ݯ�2P2��j��4�C�f�~	\�f�1ד:=�a`F���v�u'����jYT2`��Mҭ]��ȧ�H�H��x%}J/	�Z@���+�l�"�h?�U$�s'��fw��9��zw>�rKI	$TαF1���ڭ;��?4�z�a��P:�C��?�A�gvq)OY�F%Z��Ӈ����t��v��R�R]��I����v#�z����(��x��=�N����t��� _�S�Dzg�0�E�D�9a��)hvƂ�� 7{ܫ9���L
��m����B�7m�0}����'��
N=ɽ0ό�r/�Ap^�����נc߼�)5݉������EFf���͞-�r�JfA� ��r��Ƃ%����X�j�����!��DÒޯO���A;���y�p � _^V��t�H�]A�:wi`q��8��(��4�_^��U1[�M*�Ԑ��x�Q���tT�~X�'���d˼?��9M�/wV�>�z��i��;o4���W#�Y+l�3����f�L/�Ijոa8ЕqN_�������\[��9TY����q�n�����.�o��5i�W����Qv7���� �$@����dù��V�۝L}�i������&�<�R���d�}`�N@�s����Jnr�\�=�-/��w�����?Π/<ڮ���}�奪b(�P�uz? �3�!�������n��Q��6�|⅒C�;:j�*o�B�%3���đ��`YD1�� ��-�� ��տƞy	뙁��!����i]�A�����04���&�T����WO?�`R(SiNnV�����Ϟ�;
��C&Gvu�V�
���)/g��<ਪSV��$iH�@P)
���"�rz���\��QR��������?c�>�r����B �D��C�se���~nk�2����{t]h��|��ޣJ�f�jf����G��*���Y)����Et�欜c3m-4�$-�*�MP��G^�=��̚V�#�(im�^_,u�Q�������:���}���kJ[�dw�7�����ORߠ�Ep����Y�{��.r�aLֶ����%��p�5�8U��zy��L��]|�غ�T�����(�_�~7�8x�V]��d^�]��0��J���h ���3d��Y�ӮV��eh[�H�G����qK-E�֊~�B� K��3�e^b�GbW��.`m?3a!N���_�7:�HBh�c}����縗>���B�9N��/�拃6 c����u~��YO������v�%ET������ǖN�J�q54�	�R��NVz�P���P_X��˔,���&~H����R{_U�R���#AU��R���qVn��D)�N���/I�s�-6L���F6�s>����š��2�-��d�ݓ�C���N��\��,���g� sP�V4�ޞ�~R�
��cQ�z�ǖ�YǬ�	 #^~>@��?��[/qe��ej�[t�{'�
�UiU�*,�5��c��B����$��Ҳ��8|0�������>=�׳�zgV�.�Wj=ЄFwzdk����p&	yW�����M��m�y���&�l�����\d�����e�M�L�j�]��6DH�� �c�٪������0qe �kLgS�� �����az��72r����9�&��G�W!�G��^=Ma^��Fc>�xS��n�-�]\0��u�"��߻S�냰�3?"h"��(a�^��z���,�f����c��Jt�3^���1�,<%?�W$�6RR��TU�F}��<R���ofӶCz}�-���sy����cX;~O�ȡ��5[.;��w��`�L'�X�K�\^<��r��&ͯ�w��M%��``��5�)e�\
SBe��kf� k��� ��_��N�9��5�p���O��!5��d��L�������{�ꮣ�"�RYP*�)�t��!xqM	B≾,�C�{K�c���rk-9�-(��p��P5;���j��C��e�pv�t�µ}^��$3c��ĞI8<�[��(
�E���2 �b�#b��4���Y\_j���޸�>�o���8�@\>'���v��r�]!��hh���Z��%9	ZJ<�qni�^%"��rW7���w�*�y\�����E5�V�m�w�)�\Գ,܏#`���]����!y4���xo��;d��j)Pʩ(�N�W0��@�!��y`�X8�
�UvG�&&/;�pZ���LYB���/7�ʝ���r�!�G3[�QR8��N?��a�h�pUo��c�|0��l~?��Z�������T�S�y�0o`NnM����;?�|��r�VԖ�x�R3{s#��<���&|ؙ6�2��4Q��:ASa��r��$�j_�dD�iI8e�I�/�W�0�1�sI���r��K���ڏ��@ہR4�3�" ��K��)����{��pG��1����X�i�+!@֤�ת�z�g���G����J�>~�ݠ&��A�3q_HIfl3t�N��]����z�/fi��HW�E����s�^�U��);P"c��7�*U?a��+=�ևjEd�#Ih]+�GM��Q;��q��9�I��ڃ'(�XL^�!���{BF~
d��֮�\�o���>|󍾏�*�
��ɪ�:��>��}�<��{���w�;ږ_1�M,E�hj�H!?7� .�����*M
���p)�l|Xw�� �2&bdn���C���0���)�޻���IWKm��NNF�0S��x�%b�6Qu*Ks�4:n�E�'݅V���<r�t����,�2����4�:��>��ՃRI3l��q}��(pF����\�� ��>Qݜm1� �y����+�/�d:�h��z����^/hN�E�����5s�+U��*���/iN.�SC��f��9��G��!.�F�C�H���E[�C���XƁ����\���ļen��6tA�J��3�+e:��V�����@�Re�=���BK�+$կ WO�Q�3<��P����	���t��u�M;�E��8`	����M�T@/�3���ނr�p��+�WXGڡ�����
Ҫ�+�8�"�^,ԣ���]۽����^%��׶�T�����2.Z������0vF� ��l��I�f�>hr���SZ�!��N �B� �����f�%>���v��ґ���|��V͎@u�"Ø,���']�
C'CV�� XW��~h݃`���9�=j�A'�(���pB�:���$РUy�<��P��C���̓Y/�^&�;g���Do_%@�����ǁ�7T���j�P�t1w	8 �q����_�E1�E��K����b^0�F���l�m�4�gZ
�\rŗ+�T
��Ǧۉ��Je���v۽�ʳ@�8ZMe���r5����n�ݗWɵ�^k�ʔ�-qV�'��v�q"��y�(�"D�tp��B�[�q�F����g��>U_�&�12�l�d'���J�ɴ��JW~�P�r����Nr�XvQ��=�����F���q�:�c�g,x��zm[(H�.�^,��h�-S��C��U��l���>޾�6͖3��ia�b4����R*��ܼG�[��i�%v��ϳ�u/�.T6e�e0&�0jP<&	����Ź��Z��^@OcbkjAp����x�dl�_J��(�Wr����{[��V*
����攓(� ��W�����@�=_ٺ�3������WT�SÊ�4�l��F���J>��>=�ߥ�>'"�`�X\]㡓c�v�v�ۣJ[x�����9k�2�ɨ���W��l��~�w6�D
�þ�L+�̩��E��z0t���E�l5�h]ŕ��S����R�5r�+n.�(��bS2!̈yS����l�];^^��(3��:���׸$_�2�Nђi0��ǖaè:���y�	`H���{9@d3f�G�F}yRiȽ�\�e7)��G��,R5�d���2lf�2&�L���7/*���e�s�,���ZI�d̼��(&�F�����sw�;+k��k�jǤ�r�}Ջ́=��#�����3�Gˢ���$�۩�����a+�{!�����
����x�˰��1��a����j��֮=$VK̤Ǭ�N��²���\L|=F/�q/f��f���!m��$1����:� Tʄx_콍c����, ��7x�SX��eR�J��cZi��Bm;s:.D%C{�!	��c(��,Czg���+�v/ie�cMVb�|�n��E���×����w��J
:���7�e�K_>~J�_�|]ۺ�Y�����+�5���(��n-�R6�>����G_\;����Z���
7lYx6�nZN`O^��X�ەx�,�L���
C���nU���q[rl�A�	�{>���_h�X)������F#�V*�J"ج�v�4�s�5&G�h����~x��}�r�"�2���T �B����0kY����!#�0�� L��48 J��F�lG��)�i��g�	��@c��l7�*��� c�td%8s�!h[Y/OH������p���VJ S�_8�yz�Keqh;��Eu6��|Q'o��e�t�\|�Q����<���=qZCхaҽp.AoC��>�l\.Ǯ�q �w�.t�7�K�jn[�>+/1'X��-�6�1DW�����eS�d�H>|�b�:�|����eV��hm��#|�r>�S��-����T%dpvOX�{.(]W��:�>I}y�OO��hAy#5����C�VNC��e%�^�Rb��\�}���<][���Pݻ�8�����Ez���e��7[��a��*�e������BU��ͻ��?�'�8�Xn����C��ǟӝݧ�w_4��=�l��/��~����!��؇2�ܡ2�|]���n������qK����u����QLG�`(h�����O*�E'g @1���P��\܉�������w\} _��0J|e���ǧ����j�#I�5�Y�H EzzfeE�qE���!��d���p��5��~�nY�9�2#<��Ԕn�����i�%&t���<�T�r�6���&����?N��&��J��>�ӆ����"5���P��\0FiӦ�?�Q�R����gt�T�
qN��x9D%�M`?<x��q��L¦�ߨ��|5f������L��9Mc���G���?H��3RG��A=JY�K�2�O*O��1"Z�{�v!��B�y����s�e%�i(:vS�XgwגW�-�cJd������+7F�<hGj�d���L�_<QWse6 ��TS��f��'�˹��"�lMQIl�0L��݂ȵӫ�e�Ȣx�5�?�-�(Iw*A�&�����qj߻��Ke}hXゟ��~њ����{�LP{!3�|}���*p��ệ�\8E���>Soo���Y�4�2����w���Q���f�+C��V�%"@�~�;�<XYS�Z�p`90k�Ѫ�h��z�El�ap;5��7�Ӭ��}p H�E��=)������� �-|t, ��>�؛­�"6��B�a���Y������Α�Q)e%���m�>l�/7��I�Z�����c,�)#t'z�ޏ��X�Q{L��m���G2��@(&��`�J������iX��(ި�X���b���`�Ա�vu�$ݞ����$M��\�R��{� ��S�N��K��r6�9ȃ)��ij�������>|�둹�$&Z��;�k�D4cp��v0{A[b�<���w��a�b�?U��{��K|j���"d�<;��G��Tu.w&~�)�&��dU+ی�cٳ�#��yR
�Z#S�}���Jӳ~6��2��kˀ�oT�e�{a�hݲ���e�8��,��P�����T��ޝ�8��0-��_�����k��=�?��?�\�f� �u��Ђ����A��k%p���d�>Ђ ��`����va�}?��5�g�_������
M��n}���-�9[`�>��><�3�-c;j���ɂ��(l���S}	|�Y�QL�=�Dc�3��Я��/�����_��|��v�����H@�r�8�` ��M�X�~� �����N�~P�,Fu]u�Y}��CP��2��;`��jt��$Z��}��n�ևP��)D��[�v���8@��;N�xc����n��#1Rƕ&��k\�*k+�*��?�1!�/�~lz��n͈����{�}���A��;J��?#�I�_!�������|I2�sa�&e	l���B�z��W��G�4��d�ҽI������,3�Ч>�ϛv*u9$4���}f����}��:(3�0�4�3�Edp�0�8QN�C.���f�bmY���mZ�6��t��+FG�;8D��e�XY��ϧ�*zf��(g�FX5$��;LL%��=�^� X��O8�X ;�Tۂ ��*t;�:���Y�l��������ZmRkA9S��~~u%x	,�|�.ˎ��� i�<-,��J������͵�I���F���l�(-�T���F^�TU�I&6̫��ìP6���r�� ��z��%	�a!�uoe�*�,W���C^�~��u��+_�rp��L�/�㬇_*|Z!7�VÅp�T���;&B�D,��?m?�=L?:Q�?�Pj���JYʃ�W��)��B�r��`��zQ���f݅����l�u�� ��+�v*|rX�P%_yԲ?�ͤlc�df����=Sy��+|9k1��)IA�x<�6{W��K���_$����d}�Lmx���<T������ @�SM�4��V�T�I-�}��){���N!)}4�P�*@��A�`��"�Ɣ(p����lxv)�$���8}�Ё4���P%2�,p�m�0c�ԟ�Ϛ��ԁ+��E{'ї�w��K��v�){�������^� �$d�	,���9}�d�Ű� V��$����dzLU'�$Y�W凫��e��-���0y��a��B"0��^݄+�}�Z
��WS�ثO�^��=�ϟ­e����<����,�� ��iRd(��r�����Y����0�q�.�z'
;xv���,��^�_W�i<������5,��ۅ�+���}���vhN���__,�ެ����6���[����\��ެЦ+=@��{�Rb!H*�n��N�<@���R�G�r�',�8}��a�Q���!nzA<"�4$�ge��=g������2��n�
�����	�_SAd���������6e�˥����krRM��"���4�����!�N*��cF"L$��W���T����e �l8��̍㵤�Z�Ƣ����� (Nٛ4��� �t��U1�r����\ק��ņn�SݶI�[��Hh�Ah׾��j^���9D��|h凃�/��dl��ښ�Xִ�u8���Զ ���p����d�3%ך��W�T��<����5�R�\m'E	@>}z����ު	��שs�)�V�M�@�U!���>���,p�({��7��ւςv��I��{�
P�)NV���ꇁ��=�X:�YT�����^k�ծ}7����ýl9���0��J���xN�a�vY!��J {��J�(��(c���p��h{��~���b���1��˖��UN&���-e��;]���rM�D�m�d�jS���F%6lCx;dۦ!���K�{U��/� '�8�z��)$�'�)&*�F!�>�����N��	�N�v���	�tM �A*mA�i��?+cF�Wɒ��l�'��&�O�XB�bতSi:����r����EH���;�4|i�'�d�x� ��xj�����9��P�'�����f=�I�Sf�I���au��P&��� /�A�A���T�s���"�i�vv^��G�� ���Β*IS�{�G)x�QQVC��Z �L��ͥ�b��U��/ �:wR�9MV}>�}�4�5e��@� ���|=l-�e2o�Hن�YY�XJв�X��0_�i��?�^��v^���e�=I�l���aysnn�5�[���\����r��e�V�pw˩ ꫻+���Nx3�y.6�5�+Z$p�V3e�G��L�7�e'����,�927����Mk���fn�re�i���
p(v����ˢAL/��������\��jtŇ�{��M��E�2�
5{�+���H1յ{>��ǖ�rn�߿r@�n>E��\�W�.����7:��Y1c�L#r���2�1�9����Wj�[ �C���p.��5h(�w꼧�Ʋ��yl�;r��|�iڒ�	$l���I����*S�����m6��5��M|�n^1%N�NAM�vP�Є�{�{OR������qok^#��8�K���6bG�i�qq$�e�zʂ�����j��|�t�["��ݔ�&XI��5�G�����9ǓӁ����.NN�#�]H1e��49&t�X���׮%�:zA1�5c�î�;j��ρ<!���a�z����)x�,i��
��*�tZZ�xG��+o�}Y��ܮT�Χ�z�0
�d>i�i$���6b���觩�;��R���t�Cm�P��\5�K��,�)��\��B��͚2�Vp�	6�y�և8�7�a���u���xK�>s٨����XRh���ǘ�5�J
݋&���}�W̜$��7�������J�Ub�Ѯ�up_����n3�/���7��&s�$[5Ժ�q��"a���8ѽ��R�Z�T��ezN(80�$��i� �3O���}� [M3]͂��Cz"�m�Ž��71nN�$�OLX+"�g>`�laN$�h)�-��n+5]�W�Fƾ!AY�Y�&wt������b��5�y� ����P�����EKn���
*����,pk�}�.��.F)����:Ġ�^	x��CI��ې�M��h�<P2��E�Hte�Nq�F�X,S��O��>C�|��Jx�&I�߯>�Ѳw��m:�N�g�jf��港UZ?nh��� C��0��i".���e��/�	�ʨ�Eğ�!�����u���eQ�5dm���oa�������9���A�{����&M9&��Pz\D���ǅ������2�l����_8�q*�C�����	ٕ��dVJ.�w��%<�l�Y�z}ş��<鵧�"�R��n���Na�̠a}ڊm���x��6jd���1���JX0�a���,VL-J�e�voN�}�a�=��/��v_�%+� ���!P���!#�P���^ۿܬ�КO^�l�"�cֻ�a[؃����J�Z2+�lՂJ��ݰ8I���b�������D�����l��!�f�j'���)�&�לک&'��m;��i�2x 8,8&[�n�J#��VV�SJ�>�G�.N��F��@G���KE�N��]�r4e)�{��y���2"���(��w^�?�}�_?�7/��d�D��e=L;ǎ]�<��$���2/���Ã�gu�9��w��B���ݧ�3}�4�}���M4@H�ht��iZ�͍V��S��f�d�Y�R�d��R6��T.�1��U+(˒�&s�W��u��4��l�2+\yWX�\H�'jǗ��W3�t��LV�Z�6���[L�<�Z������_��K\N]s�F;{M~���4��e�G����S>٥���Ɛ�_�j-7VN�*��^��v�Z}�i�{$PN:���?��|>��s8l�E3��:,��tD� t��D�`#�(������7싼�E��Y6�����p#��t�'J��I����+�V4����� p]V��?>+�C��D늻�*i��v
��g�[�}��;ys9Ջ����N�+}��8au<����dh� o�u���%��I����,fpq��s0J�*A�#�����9�p/���bMHc$;�.�M��L��x�����Q�2�IXxo�"�2�ޕ�_
r1X��Oٓ8|���bF,��rȎ����Etʚ�;M]@n�"7DO���g����D�-��R M[��!B
F)�6��P��^�2��1�h����v��R5w�z#�1����:Ѹ�r@5������l��"���2}V�Ip��M1��7�{��ܒ����ʮ��K7z@���Ca��\�\�UE�k�_&�R����Z�fv?��S��޵�����>�XP��)P �\
*|0"��>�����W�>�����	�B4�%``A�����Yk�~���&���~�t�쿁L��Z��6����V�	2<MFKetMa�ik��=J&o/�:WK;Xڕ�bȰ&�B�7�WL����o.ȕl|vi���k�qb4� ��aK++w�o��;%s0G_���	��������߇���_�|�U��j�^�B�yX %˳O;g�pE[����{�=�[[�_-���/�%|�W+K__�^,��l 1���ˮ���Xt�r���P
������6<[��B9�w�ċ�EF(8�GB�[��8�+�6܅'��^���-v�d�b&�4�8��w���WM��$�5k�v�zx�tNM�15��tM�F��:2d[qg��%}�>^G�^����Ɯ�1�M������K��{��v�(��]��ߗF�#ń�?��h]����ġ�?_�L�,�c�"JPy� ��B��̣�[�:V��� N���ҿ����v��}��p���]�֨�BP+gh�Ep6ki%�v�g�7
�2G�1� �=L�'��\�\�2��V����j�	�e����d�7P�,˻����x� U��ug{�(~�n��avs��]kc	��zp�g��4U�3�\����+p���5��ƫ��U�Y�鿉��9SB�Q��#�$�pc�RW��ӷS��^�6�� I.Q�4*��t��U�>1��,���-{�X�	L�`,�!�k�j��g5�2�=��S��F��wϛ���5T�;��^�L�dtzK��v��aM�7J��&wy�rE�}.��K��{7Oa�iSEs��-��?r3�����A���C�'`7��5�T��R��
����������Qf�\I��|��dz��b�CIV(\��	���i�0�.~��|%���d��M=�DɢTM%6@P��d�Oa�ĈHS�Tަ���-2/X/I;.1Y�5\T1�t0��.��S�����H�E�g!����#�:��K�`�)gʱ׃�������U$;0K���0��'����=7L������6ac���u�oX ���w����"Њ���{�o[�v������-W��M���4\UI�%-����R�(��e�����}a�W���vX�zG@aj?_�矐 ����wYyi�f���2���+��:V�<h����5ؒlYy�d͝z R=��K��.^Д�D��nڭ�>г��p�V�o��u�$����Ӳ�ӧ���uqm8����}���p3[*�ܜ�a���ʻv�ْ
[+Ѐ�0�̍�]��YP��_���T�?g_�as؇_�=���{�vڄ����f��e+�a����E#W�xXi�蘩�7Q�=y��D��wهT���Xu6a�T����{�^���^����-٠}	t<�#�F�Oh0�.�ǅTQ��Y��G	NƚTC>/A�.)�$6A¦��u�Aύ���hА �cVF1���r.
����ڧl1���a����zp'�JN���I}֓8���-�]LC� ���?x\zI@X��c�7��FT��U�Ŋ�^�� L
��Ðk�yGjAPSg��lV���ts[w\��}|ܲ�PC�]������`�j\�ső��J�+[��:���y�2�V߷��1�b&�J�9�����ҡ����u���
C��E�8'Y��·l��a@ �P���;�6SZ�m�~�ɑL�x��r��.�B�}���j�9!_����{J\+���D6���!�,���F=m���9�k�a��~ƹpZ�F�(�-R�"d'ٗ�~�ߗ��,�R����N�b���~z�j�LQ��!��W���^n�E���R,��Y�U�Kf"?F�ix�2>f��'�p�Z��Mj�o�R�h;[8>��WY�v%�a�ng�H2�&E��)R5u|��8�1YS�Y!��s�����v�,R��
������ٚ����v}ԺBZ���Ó|v�.���N�/�,�w;[Beƛu� X<#9�E����C�F�@�*�Qb���}����i���s����5-O���2	�ީD�f1����3w.�`n���pjS
��{+�^�M���6*�n� �-2���- �p���^����m�{�-��7�hDeB�d���c8���"o���0�R�,H�Cj�S����^�RU�"~����>W�����K���װ9���k����7�˿Z��e��۰�	�'�fd�e�}l�nf�>���l�س�6���&���>�Ҫ#��wV�gK�s1���ʶ���dfdb�v�n,-���a��2�e>�_��f�Rxb�?�@8� ��i�I�O�q�;�V���+qS����"6�L��2������E�?Z�v+ua &��5d�wN'��@O��!Y!P��Ϛ>+6�2�����Y����4�}�Tv)�8���:��43�p�n���52���e�|����l�l/�!�ώ4'PM� 3��A1e�x&{PȰ<я��]���������VDx����ټ���0hpn�oJ���lz��ϟ?+�	��9�����Ի�����ڔՌ}F�ߦ����+ʭ"J6�r`��1��ƴ+�Lcjeo.�t�d��'%&}�ΠYK�ấ�{:ǌ˱p*�,����&���S���q��Ol����+{�&p��](���x��϶qNVvrMy�����$FSe$��Uՠ3����$����K'���߭w������}ƫ���|��e6T$��8갰ףW�y8��bY�u���=�q��d�!�ˍJT��gm@�����T�A圬�U�����}�H���a#��Vx;w~+��A���0���ءA��$
IL� )�>�*TM��P�����qys#&
*>��O
i� ��2�������ߙi��������e� <�)e�X	�"*xQ�K��ު ׅۄy�;%C��ڐ�I��%��D�>�/�F�Y{9[�ޯ�����<�⽻��Rބ�|�������aj���x~�m4��?sR��3;-�m�C��Us�M�<y��`�L�+�v��l����� �t��ZyF	��-p���N����-��v��z[��ɮ�t�ؔՉ�P�wB
n��P8�z:!�������hCY��H�&�p*g��_�h�4X�䩠l+��C��K�C���0�Lד�L�gMdh���T�7~N&���^��a���.��=����S�p���oK�nr���,4�2��U�>@*�9�ɓ���mX#�h�Y���el7�B��q�%O�?�u���0���LӉeʀU7˔7V�j�m��Ls(�B�:�EL�$�Z�#?W�a�3��u�U�2¦��٪�Z{��1���N?[�_�ﮎ�[�#��c�K�Tp����ͦ��܈�	j""�d���|(���1[�$x��B�X�����R��cya8�l�ĵ�.ןe�d�gy�?��:(��,ͼ��cտN�b$���}:N]M���PQ��}8��~il�=��xN�5�����J���'�<H)�N�����Qe'�f�U[HH�,M���)gO��x:�����r���<�E`��v���I�V��s�en@!��~��'��G]�8a�N.~	Q}#m��X�^9~��Xc}��>������x��(G��R��^7����2~/W�͇29��LS�~��Z
�)0�I�6Mi���.=;)��m�)��|D�KC�!@ƒZ��ާ�L����[�3��a*��5����6$e�b��C�v͠)�Y���U%�1d����J���:���������2���Lu�)�Ic�m}�^������ޝ��J�,{!��rO	\�Or�����/ANe�Nj�=�>�5w'���e�䝸lSYF-ĠRzg����^�^��ִ'���{��~'?O���i�O������詜c+�j�ue �}�b�������x3p�O�CVA��w�����������g��8��>�=Q���Q�+(����K)j��A¢\^֊3�t0�NY�w��[��Yq���>6�{tх#�;_�S��82�g̲I��/�t��y���U�n?��|���ѝJ����F��Χ�>|)���Iyު\��Kٟ��&�;�Ξ7��� G�Y	��UX�v}B)� �>~�Ӣ�EջJ�����@��c�.\)0xp��R��#/ճ�0��9�ӿ'��X�'�n�_���H�OA.)	��%�Jt��I��+��Vxa+$5�$��N�{���++�S�9�ռ_�fc8hƟ_��!A�n�<��Q���$���%��.ݻ�U����6(W�>Ŭ�>ؒx��mg�am����E�"��n>�+k+��D���@ H6k]��¼d4��6sljY���V�~}z�/knvo-�'�<0kF�T��b�����Ƃ�֓����{��ڕ/�Nʿ?~��k{�:�³p���죈����3Z/��!Tdm��VH��
��Q�ł�q�Z���B�sp_&�$����b���E�z��ăe� �9� L`#����p�!M���K�{�$��I"�G��5�D㦾�KU���$Pn��h�:#�Q�i�#O$�B�� ESs
����0�����M>����V�åC���\0ONF���]O,��M�?����|��]}6�x]fY�P�ZDw�AHK'�`(������߻��}�@��&�����S�������fr�[ҥ�iTŠz1�M�N�:�뻥��y�JR7���-ϧ 6e������2�sރ	s*Y	��,�;�M4�!���]z_�Q;���� ���ןJ�t-E\���i/��uhq00ȉ�� !	���&-�	���l��>�vSJn��U�*�{�M�]]KJ��em'[�G+��p���8E�7j%(����4�OHl�|z�����Q펒�MJ�v=v��b�O�i��7���&���g�/=;��6�}�u^�~�<���=+Q��
*�t�+ǣ1��YVH�֪�R���ޘE<�P�f>��$�'-�+�l�DJQ+e�����<+�Z�h�e��=Τ�g�V�*01x�Y��#�C�I���ic��챣�AI��wé��C��vP}�s"6��SJQ�y��y�
�0i�۰���|e�עu�&�O!��5�Dgp�O���l��ra�f����׍�Юfǰ����JM䲦-�j�oy���C)N��gR����]�=W'�t�7��� ���*�p��Y>���Ωm"��ٺ�����pOD����F:'���z�p��lM$o�jQ^N�.D����3,ʩL�}��� �d`r�cS?����s��PQ�')%;~��
�}>?z�-��K�+epcAM�<��ķ�R�:��:���
�������-�p7��>�S ��8�)R���ʂSi��:|���O{�H}�@��&�X��no��~��óZ�JS�L�-='�3��`}�,ck��e�__���.�m�x�i�^1����7-����Sk�į�Yٟ��ѽ��`HTO�a�r�&��Ӗ���,m�B�V��ճ� |�
E8X0$x,��m�:�R�OP<��������Q��H� ��
qX�l��*�γ�7�\ٝ��3�p�1�s�;6���b&ī� )��D et�RRc�c�{Ez�S��<~T�S��vt�s���lH�5R�Q�P�H�P9�֭��w���oD0�QI ����zk�����敝��� d��_^��/�����-|�oCe%��n&y����k�>`�I��DƁ�/�ē�ߥiaR�er�p��ZDHol�c	P��]����h���&z�����zl)�KƷ��J��B�;e|�Kٞ�u�D�U�%\Y�0J���9�t�2�Ϩ�͋A9E��ډ��vj@0��V���$�{�)�H�ү�<>�B�2���n��b�/�do2Pf�ù�@fzI�~�1\g��%d��8�x���%�uw�-c��ބ\�?�j	�lN^OYG#(Y�TÅ���ųel�����3~}�yCo�4����6��B!_}��	뗝��v�5�<xJ�L7�B�O�m��L�7[�t'd��8 �ΰ8P�Ҷ�ן�FC	�(f�W�� ��"�:#�y/�#qU��=�4����K�2�^��bZ���0���2L���=q� ��̠&��t�w�>?~K��|:��S_K�� i���	�)-��W��}��܇�j>�����LZ�����ׯ��5�#!���Y��$��Y���߶��y
���Sϔֶ1��� ^Z�P֮9/����
؀�f`��)��y��d
�ӟ���$;�J��A8�X���cƐ������W6�]�	*P�&�!P�BxףK&ݳTB���F����I�2����-��	��&�i���}����	�w����5��We�C$�W�KpK/�� �d+qT��D����hf�`��m�\HpQh���&&S���땤�����`��B�eFP��w�a��See�x�����1k�fɲ˨��;ze�%������ڦ�h��X����q�T9]Y����fZ*�{��:�dY���[x||�5���&����y�L����J���=`=���R�-$+w����XF <���_��Y3�c TIA��bs�b�������I�pU�P��3t��q�5;��o���R�z2�F���ت�O9?�7+���� @���ĵ2w���p�����I���^��+@�[7zn��٢�x*^�u��_4rQܬ,�#��[�@����}���*�,_�|������?�i�V�BJ�@�����}*J��@2�]cA�zi�r+OY���2Y9Da<&�խz�|�/��[=(N/~��F�	�~^F�?����_��/1��(��x$x��1�i,�=.��W�x���1�s���h>�����_{x���3e||��̇
�?d~)�%~k
�!�822W2	ț^����4�wחsz��樓V�`r��d䓘��R�O��l S�os}
���0d�������p���&T��;a�Og�ѧ�6�F��]�aK+�,�uʴ��xV>h���W���2.^[�x��Y[p��ms6�%+�Ky9��B, ��*F��&|���>��7+k�R��z�Z>I!ׁ���}�W@��^��DR�r����(c���맗��k[Ъ`�XpG�G��"
����47J���( �<�S�&v�Ww����'�u{�����Vi���ab+��		W�oW\�2@>�	FԶe�+q�Nh�u��-��Źw|��nH��&� \O5Nr7�6����"��j�Y�xs���Q���uù���χu��˗������0Fu�J�</|
����"|�=�d��[\�'�a# �Pa@�x�('��}قc���d���AL����e���d/�X��� @5�Ӿ� ��(`JN3;?O���I�"5߅�A��eY�x��+k�rZ���-܄M���$84�4�E�m�p�"���L��˟������&C�?�������Ȏ &���-q�u�ʢ�����t�K�&1�$�\�x����2��F3=�;�/�ql}�o��;��}Evg�{9W�v�K���}-�SK=c�he�Ag9�w����X3}K֞@эz�I"_rH��(��`�~����֣Ŵ�l���΂*2G�<�<��15�,�<�'�ښ�Ͳ�/pP��"��U��´v�>W&u>nãUk���.�ځN+跊���į��/__4��w?��}3�,��lxx��ӛ\�Vfc���^�B���Bwk�n���>s�ihQ�qb�R=[���;)/�!F�a9qͿ �#�y���ݨ��l�L�'�|V��W��{:2;A�.҃RM,XW�
�r3Y�ϫ��ek��o�'n��JM߷�6<[i��=�_�ïۗ�n���Fګ2�Qz�$q��LQ1�!.in�w{@�m��e&SavX\�3�8��U�F+{�����l���l:������m��G)U(ë3mt~W�Tn�{fcX�8sI},6o�Z&���[H�L���u`6�1@� &����s\�nZ��/�����
��:�|I�<y�&ǮK�6eW��*��4�F^��Mާ�WWw�0{5=�:Ρ-��mndA9�>|���Cm��6���Pm�%��S$�l=�&8���<�ۻp������7Q�%sp����CȐ1��<ׁB���<��z#��� �	��"����XS[�k�X&��>١�� q��VL�N
�����3d�_-{������~�gkM��>�q�C�fl*6}�ק��X>I�Trk���ٖ���b��<��p_�ng�$���	�x��٣퉎�B6��6�6�E$��Lb%u�Ro�Q(	WQ�����2�`��@�*�_ݬ­e�w�7v��<��_n}9ɻ�v�G?���u��*<,�ß>~�����݃2"1АW++���[�ۗ����5l�S�I�ص���D �:l�
{3�\@]J�v�꺧L��'K�1���a�K$��D�4�ɒ�$'�Oq"��d-���>��TC��w\R0	���n�h�fp��,��i)P�	����o�T�2-m���$ƃ�ԔO��k�;@P.��1l ���>d�Ț'�_
~�5��<{/6YD"�����QYT���(mӡ ���$j@ ���(��G I�&��C�4t�	eD��n�gO��8���23��Gs�ޗ�1@�/��Y-����2j$E_�Ŕ)��-�G�� �͚�Q��mO���Ꝡ���Q-!�R�lEx��~ѡ��ކ�	���O�:�jk�� ��~���߿Z�C_��KD�B̨�+Z+M�Wm���@ہ�<���G�F%}�Y��y�ځ�=h�@��$-=먢,<!�⹋���ۇނ�|z����[칃}��_4ʑ�F��Q9h��Bn��ad}�v�n8+3,8�����
n��EM{񯲨���,z%�-���[w45��v؅�^��ߟ��_ޞ���N;-کSUv��� ����eY�"\�9��I�R/x� �O���)P	]��@k�Mr>]$��Z&�
�����Y^YD*?>}��썌e���4^��Z8�o�1����n� %|�����{���Ca�?K�0��ܑJ��9�q���l���G�?�b
�L%�����o6(Ӎ4�"f�`������j���r��󚦶Mr��`��O�uo�����WOgu�~�!�\;�J��lsˈ� �~���w�v��r�9�	7>]�l�u�L��������JA&��9�x�Y �҉K��Ԭ'�e!����oည4�{�C�o��P�N27�>�k?�ϾZ����/���g�v�"]=?�N�?)����R�J��m-�#g�d�}��#i�e�>%�ڂ��U���f����=��鰣G��Q}d5PrJޫ]k�B���zvn�֮�J"3��0YDa�@'\�={&ǈ^Hb��`֮� 8�mm��]|����4�tE��s[(�6�H�����fJ[|g�Z�����翅�6�b.�s0b܈�Ng��Ɖ�PvD������'���5S9�J\�'��`�g�z�z���9���ᔶ�I�FOMp�ب&�q���
���3�d��|u�#�,Z��I1�]�A�2��#w�#�7�"�s��B��28��`V�`C�^���u���wC`��n���"x�A���Ka���I�Ә6��7ey��L�=�es/&�� ���!��)���99�^T+��ħՑ�,��<�I�+����fY��Dx������2��i8O\}��Y�1h�iCu(��@Wn[�D5I��Q�MY�7�@�0��Tx�$�@�B9s�zr>%a*$-�����'GpS9�Z	�?cM3��^��/�O���S�'��O1��>�
"�ezO/o�=vךf�1	޴m�m'3�����5 ����r��kVI�+��赶���)5q¯��,�b^�A)tY~�`����0���l��� �Zv*�7)��^�j�3L���=,����*���!TV��h~�F�2
[(;t��x<�E<�巟�_���h�RYav��r�egRPf]�q�JNգ}��"��݌�z�$�:�]J���'���*3��5�A�*�M�����e���n��ܔ�zE_A�ç�>�;�.��A������z���t聥Lk�+��&Q���N'm���SS]��)��2�=A���5�fY������X��䵽Ov��$�aʺ�n"�t��CĽ)k�.3�Y�b���Ir��Y��0D�d���-����}
�����>�,{|����V�p�k#ww&ʼs�Snт�fX���l����s��,��0x�vб��J�.����]�L)�.b�2�����
χi(
��Oڨ�{T��ޕr�;�p�n�,��[fAQ,��}$����W�^c6U)��ߓ�[�`�:h�8�uu$�����y�;9��~�C><��s�����q�Æ8�d<��d���@� �U1�l?��[��v��#k$�X����{jP�Qѩ~�T�v�\U\Kɀ-x�J�*�bb�X;��ap�˼=w�I�4w@�� ]��[��8qV�+	CΧ�z1��lľ��]�������e�>���-���?BO�O��)J�Hs���O^^v�q�W����R��2.h�l�=uj���o��I� M=2���N��~G�H?|?*N�D��R�M��P����n�q	4��J�-���R��	uT���"���Os�$�#��]�Y%i�be�8�G�UUC��AT���SoNzY�4:7w�ulT�2[Am�������Ƭt+=&�(�d�м#A�s^(qP��Qr�O&������h���ZO�� ��!XPf����{j�p���"��I;\���Y�Ķ�[B:�<f���M�A�:e``���(���d�N���W;��K� ��p��������:8��^%ӛ��s�i**vd��� ��n1 ����t����ǚ~Թ� �ğ:�+�N{�O��;�[� <W�بq�8o��Y��n�ۣ%��Y��oO�0�b���Wk��?­���XB[������׵�CxZ�Z�f�e�`S˄7��s���kKvH.a4s�ׁ��ݓ�l�������
8���6l_]��<��
��I&� =S�� [Nm;��a����V剓��wiU�F&'
a���R�t�k���ٿڃ�H�in�A��,�B���=dD��v�R���A\A���v�߶��o�C�qˉ�@3�}6vrT�\�7w���m�ia�I���5M����3$�{_�B>~�o����+z`��t8�K� {�2��U'�	m+y1�m�$�А��� ���3��Y�m�6�='���ߖ���Z�w�D�v秔!�'W��g(�Z{ax	�_�iB�^�k�/�����&L| �J��q)xp�˨+G�F)U�ݠY��k��4̿���YߋIh�W��n+�d =��䳍}�,"��6GS���T.~��,جM�ʁ*@ԁh:��Di�k�I���8i��+��l�ɫd�r��b/�w�ָ ��f#�^2Ν�7��S4ꥉ��Ȼo���_��Ƃ���vy�p������V��e�Vt����@�Hv۫'@�"ך�|�bY=@���qʒѪ��y�QԝC=�Y'��ثI�B\M��.�_�Cٸ�Ϛk��K*�38���X*s���-�J�^�n=��9�A-��z.US��Bm�'���"��ʆ��N2�	S��{��w�p�/ ��U5����������º9�����<nvk�� � ����i����\B�3�&�v#Q���E5׉ǔ�G�*��r��N�����Ox�������LAN"��m	~���_�9�����Y4����w��]v���Fʰ���ęJk]g��T�(y<�Ig3��ܹS� �>��.=7��]̏u���E�'�t�~����i���W����A��g:����J%�D$Ŵ�3M�话U6��0:��G�^���H!O�Y�s�\�Ų4�r2���CY�J&dm��P��p���a5*E�j}�'T�l>-�/�8N�E-D�D�`l�6r��3����y^㬌�����_��W��Շ>�{eҴ��l� �k�����w�:Wzϔ��]�Y� C[Q���ε��9&��c�zɺq��Ji
,��j:X�iu��s��5���������`�^��"����ǗW�E��ѭ���]x���i�]������:A87`��\i���������W��?�|s[6��<|�DO�ח������Z��E��@�on�������'Q���X^ڝ|K���=!���F���T��c��v �.��D��4�L�'驱8�F����l���iSP�7zpd���656t*q�K��S����Ry�8�*%'�qy���C�
4H�x�4�L��R|(/?��AA�yK��!�M~���!�A�k����J���Er�
I���{�� ���I�a:#���=���@��H�n���h�8�Q�X�C���^�3�)�Q�I��)@�@������B�EqY
Ǉ�k	F�gĕ��R��Z�կ���l2����yJ'�)f�yn�v��P�A����$��u��ugU1�̘�VM�z�I�Ɏ }�W��<D^ZH�t==�_���禗BU"@���]t^���X0_Z@�E��C?
��E�řU0�R�|�s�d"'�G\GgAPJ�r%m��Q �(v�۬(Y��j|AC���cҡ @��:�����.��z_�����{���~z�Ug;�&(X8a��>]�[�[�[+����(C|�.��+�G����F�W�r"�6��[����2���֘Vjs�ַ�E0pa��T���Û=��v��ŕ&��݀"�Oc�&#�=���r�`��Tds�,?S7��V�BA�f ʯ����9����fwq�� !����UXo�WSU鸴N�D���,���:L��8��̋�L.�,$a��s(���M
$ɔ�&y���)�@EJ� ��T�0r�����i8r���eG��Nz\A�y�+{�W���u��A�A�����)�=�]nk������6�A�ž`�Y�EO^� ���b�_f%�Wb+�c��(+2���˟ס�Bq�%a�Ԟ�Kv}Y6��G�,�����c�ҧ��c֣�T8�|6��%␅�V}�� +'Z3|�@"�"��r�}^��g9�嚸RZI�{� ������-����� ��9余�Hf�!Nl1��zi���:�޲:+�Eq����,��֓f��P$�#�N�V琗V�z���+�d�ә�Q/��<Bw��β���7$�W}��Fp�t"�%\ْ����p܇�ۗP~�r��M��t;_��l���\�������ه�pu�����p{/B9�+7B�oo��o?�~}~{� �z%�1ѕ�Ej�6-s����86����`ԜC���h�c[6�͖1a �/�hD�S]�a4���@K�>(����*���篏44J�Ё.��S�t�;(�҂�P#y��˼1�]E����1_S�^��.���O;���R�&E��
FY�T����E��EqN��ٺU�!����;��wp��Z�K��m�d�S�4e����5� a��b��aHe���sIf��wrNe���/�OѪ ������,C������	���X3�����Z�;M��F9n�(��fP5�&	�}�½��YK8NnF!�k�*�\�A��|��36wku8��6x�YRk�-��{.��� =9�f�J&��8�;��@�S}A�F����Z�,^[FG�Ũ�쾿j;������8�W;��(ap���,�@Y(��ZL�5F?T}@@1��2���⡓� c��̈��*��)kk��$޹>����vP�fEv���W�����a���Β�uXb�z�Q}K0��ve��흝����5<n�$U�z����`�ݡC�
���MC�ˢk�\���i���{Cd�i�,͵����1��\`�{su�����L��,=��� �&�>�~w��Q8�Ǘ'Q�$�5`��.6C@YΧ�>��i�U�qxW!����kǒAi�$aK�2�:*ݎ �c*X
�}	~z����i6�^zIRG9�����(�����KV�5��,�4�琽ϧWe����H3<�{^�
�1�8
�������Tm���_ځy�����3&���)+�l>�tϒϮ��~�f:X���k8}}	��&�N�&��z��	���ʲ�X�
3�_<5 r�@�
�����N����W�d�d��w�ƞT��3>˰����FL)��(����C/�;����	y>�RJꭡ�Q�.t�{�M�cj^��##��O���O���f� ���YZRR�7�z�!$|��q�uI-�i�5�;��V������p�R��ԝ� ����ȸ��~�cv�����{M�k���#���)&U[=���YV�5�PXz?�4�LY���^�҅�q��ܼ�
����%l�{���sB]����s�[1�=��l��T7~M��p�rx�l {�R�kKza��a-�!w%�l iX�CA�?1���_���Ls��1e�+*�:kܗ8˲�&�|M#iw��閜�\Om�܏�NeU'�m%.+������x�p�2��wK^¯]�_4�T/���]��!��T0��ˤZ|�j���1S��}q��)�;�*G�X��; �`�^]���.ј�A�6�3X�j��BnP�Ct�&��>꾌2���K��-��������$32�����p����ˤp���C�"�>n�kx���<�����#�_�:�R����]���}i	���Á`�;L$s2/e���6mL�-����.n~�eH]&[N\��e5��o(P�|~~�=>Y�;���)PM�tdm���Ya�ϸ7tF�xI���CS��{��\��y�QA�iv=�0 ��܀ay+��To��!��=�S�q�Cʴ	4�����A5u�S�����R�=7��cX�b��\��AS�eh���L},��y��������ihW.�L�����Y"�mr��W��)N���J>��!�b�t
��㐘�Y��g�v��<y`bQV�f���u��2��7��!�����u>�e�=�ݫT���Z�aDZg#	�U��۪j����IT)>E�T��y�\�$��&ҼNR�I��v�H������.,�1D��!��?y�� $���I�+;ܶ����B�w{6x���P� e��	Ы�C;-��ݡ9�I����aa����*�ȋe��E(�֗��N�_��.�X�3Rf�G�wHEi��h%�XՃm	L�ȴDh����ص��]d�d�ݸ��'�{�;D%� ��l�
����։������i}h!����'����NQ�����n#�KXo����ԕ�\\�<�t�M}�,�(� �s������ڒ��F��^9��3v�P�n���=k-�#QxS�q��/5�c
)U˭UP��=�Mxۼ���]x���,�)a_{}���TM�<�e��bc�~C(HYvy��bHc�6�4+UTe�]Y�i7z.�4|�]�n�H�t�tRFh�؜iB�Ol���޲���ߔj;
�:��H�a(\��D�?�u9N ���&w0Rߟ`�ɩ�d�@�1g����Rp���� �S���p]lN�Ys{ �.�ݫ�\?>>���d,=�=2ѭ�(u��!|�A;�t�$�c]�@f�*K��j4�����,�����ep�J��?dޣ7����G��#�%���Qooyu5x?$e�wS��j I�h�C`ui����)���r�>v��a�ԣ��pb������-l�����^�d}d%S�&���o�E��["��/PL[�&�쵯,���׭��
e��W��: D�_TY��HYv:+$1_R����lW�;5%O"��3<d��?�G�����;W���,R�
����'NO�ޟu�� '���]F5Rk�M'3i��S�XH����%z�������e��t��[=6��`�XM#y(`=dn������:jr�hR�+�@l�W=)�7nU���lo�˱��Z�\4U?�j�!�!b�a���ˠ~���ҍeN��4J��`ԲpQ��|s���l����[��^m��44�+��.[�̨�SG-��#��b�{?���[��#i�\���t�T!UЎ� 0���)<�fa�����B��c��E*� �8����no����N�ۻ����?��wW�E^���2Q
�� Ǔ?'�Av���Zܛ��iX�""(w,���.S���q�6ejͥ���A���E��oޤ�{���.FP��Ր�x�t��@��=���*�gT ���P��M�ļ����5q8�: K)�C+��dNl�	��.BI��JQz��嘤�P#QO6����`b�{{fӥ%��(�U�ѷU�j�6ZS�=,�(����7�� >��~�t�=���m�|9Z�cZ���a�@ǋ�3�O�"�-z��Y�+���G���`��0�@�T�T�=SR��5;��l�~�h����'�����R��Dy}(a;�_���a�
�da��h{��oU�5�7�`0l�#LD��r�|�>�������������H�O.����)!#vW�E�|}���?��3�nȖB#����Z���Uq��\geYb��ۛ0��_�p޾��V�ި��]�4ki>G�g��K5���(
D�T�D9
�x���,s�e--�/Y�y�~�dR����}J(�T������ p�A��������#�H'OIj��� ��b�ɣbEe2��vcSv�T_T���ܒ��!��w��o�4Dh�1!��Lk���C�&rt{ٰ����Lê���wx�&i�������U�6̣墸�t�-�'�	�F�_-�PNU�g��<j�P8�]"�� ��Q�j��J��룊p&�t�Gn����Cx��.e*A�G��o�.���/�w(ŔQ`K>$��R/4�ݾұ�����q{ �tO�x�2�v����'�������q���@ok�Z=	:��dD~:J���󎲳��~����r*qm��e��4աM�L�J�����Qy�#p1H,h-� ��C���? ?Zb�7n]!�"�;�a!�aD)n��5��Z���6�x�1|� ��-�ۆ��j��Ɔ']�2�
�۫��M�@2���WJ�t&�����l7h+3�Ȁ�A�t�2�2�^�[�!9��s+��d��&m���o�X��pc"�;ᏽh[:�#h�;���<�_��
O/�x08Ee�N�,
��(U	�X� �O&�>T�}C9/�����;(*Y����w9x6�r��->I7����,�����a*�h�Č��: ��K;��?��ݐ�)ifm^�C���]��W���eػ�t�ʖ�]�1�f�}ꁌ��?�-x%,�W��J���o�sɇK��Hlȧ^`����������v��$�,��X����@���ޠ�!mD�,Q��E�[�ķ�gbc �Y)n����)�\~ۃE�7������Et��ʳ�\����T;ʵgY�"���R��!v�>h)����B���j���M�zO"�o��9�B���ͽ��2F�TxZ}�}�����g#)��{k�(Gg0Qh��������m8�&3[D�d�m�]���b��G� �����~X^���*W���NJ�������G���B(��N�۰�����]�����J��+�W�a~{�O�/?[�l��R�IP0xI7��f�l!_N ��B�DG�SG���6�����в���?�c�'u���C^2ש�cϋEΐ �}@���I���\k�*���q*�kR�MAC�B��l��1�TH�_Reo�Ҕ�'�w2V�5q8J�����������좢ˡ�����.�Gi`�x>ꋤ��6F��-�l���bI,y"���綦��P��X0�=�������P�JW�p�ę	��P��z�l�W"ӦԷ �d1-�� wG�5� �����,�m��h�,٠��%�1��W���gC0S��8VO+%�+~��͇3�_4�)�{d�����@�ӿ��;�5�?��gRvRJ�dw�_�szN���V B���$��ϧ�@i��&X����ry�S���2�I�\�JmG�{�����	�nyQ���<���W�XZ���	�����~x�~\�;E�ٞ�5�*�O����HSѺ�-�U�*�@����J�o>�b�
��~��8��odM/�OX0��S�\��Ne)&�2�s�����hg���X�iQ,�f/,S c���!|��ѧ���K��t�S����	륖O%9�XD��V.�IY���Rϯ��*{�%���|��3UB}{�4)�*bɓN޴໨���	������w�I�lk;�޴r��[Y��$����C/*�����O�R4��_L�9�
��x
}H@C���\	���,��ώ �.�pc�w���G��S�\��U&b�q�sԫ-$�K��K�L8�3���N[�L%\���A�����HRPnUS����9y=m���ɴ�R·�ArފnU��#��9�`�8;F��_�M��8i�i����y�z2�j�$��QE�u_��4�i@�����&I�Z���`#27z�P7�^8<T�0�o1y/=��b����#�2s������ۿ��ڍ)��9p��4���+�&�--�w_۵��y}
?Yp�g�;���=I�t)r���>L� �M`ѮW��S��|�?J������~q�t��)���;%�Si����� a��n�s����F�����׏@{��؇�v����TZ��ցļ&oܶ��fSzh��zP����.ڗ������5�]�݋;�e��N&W�6\z]���>�K�R:�Ԫ��L,����w6�nV��qFy;�b�gE�/��\�K��#�@�	�!��H�k��p�k�ӟ$���y{RP8#V��go5�����ܾ��2
��G�RJ��'�L�'��ڝ;�k��-u�U�!�15
�m�]	�3���A+���
�g.]ފ�Xk"�.Um�0�q��|��� ɒ�{�<߹U9w��2�'�dВZ�z����UG%bLǽ����-{�΃�l�=ۨ��(O���V����D�����P����O��d�B����A̐d�������;���d�~�bտ���E_��Dn3'��E'��a��~/'��o$ ��j��Z$lP/�����nBѶj��H�j?�z~���+��O-<ZM�Xx��>=����)��u� ����\���s�##fp���Q��Y-�#��3zlL�l��6oZU�Z�z2]�	Äԋ�����S�H�;�<�+{��2%pSyTc�ʪ�"�Mam�B�H����`�Iy�d��0�[�����s���WYyp9C$n�y��<�ŢpdYE�o&� �!�$^�,�E�U*����U�{1��\C��Zzf�
x�n��έDZ��XL�6qu��m����0%�vvX�8��|�aI��������!C<Ἃ
,�ot�a�-��B!�L�6)�������j���S�|!~�;�O����q�٪�V9x��s.sf���d�Ro�(p}����Q^*!	�,�����2\������hBk��Cye��C�f\�,S��(e^E6�=��b&޸�h|�^�]}�Kb���)����@����o_ �����|q-����iqM\����_��(���^M��{C�y���-��lW;�v��9���E��No�]��"��X���_�Gt��g�V�.sW0)	�7�k�(˒�
��}H�\��O��ۄ/����n�L�<u�I��޿�/�:���qc`-?�1�Y�j�fV�Hf��7�3l�7���g ךXFm6ъ�Fq*Ejc����;E�:eNg���g���
�2���D�u+�;�ɝN5cE�/����k+�s}�|���40w�����RJ���q��`v�>���"
��ԋb�e���t������2e2_����{��N�!��m#��l�� ;�ҳ6��Ь(��!��WM���&x	C0��&�J��VbU�����ڏ�=˜�|�Yz-�����3%0��za\�Q�WY+������;C��2�:7���� ­-U�/#� <�0w�9�ץ����Q(��C�~ԃʽZ�$�5|�u��Y,�`��F�������@|]d>`T��5�H��A�	9��O%����Gqݷ
�z��j��z�kV)̪��hk���ev�/6���տ��72��8�gG|j�g��E��9��|9�B�b%�I���wGJ�	���7j��gz���[A�Fo/����xޅ���=�}w
��6�Y�B��k���Hե��N%j�{~���_j�ίV:=x����Yׄ�( �H�����j�P�,�e�����!���8�V'^�b:u<^l�Xp�������)y]��z%%�N�|)�D�3�X��NB�����X,v�8��[�rs{����$J���c�B-�I��_�������{]��)j*3S�3�Hmw��x��/vG�����Qr[:h� ܥed�el�}Nzh��'�F��J�`(q��6���ԃ}���2XMꢹN:hryL�/���C%�/��(H�
([���K1T��22���1�.���t3b2k*�J����.B���\�5Y�3�=���O&��"�݂e�&V.�U{�6��-�X����͑@zm�'QEG��R���.jEժ,f_��Ƃ�l�b�e��5'���:�gy�!KJ�[m�x>�k��HF����E�9��𸆼��}�
}V��$�X�؉UrS2Q�g��Je�>�O�b�HӘ �I.�T�:��է@����l�%��B�C�D�ݜ��'7��rH�%�#oz:P5D�z=+��AUp"��J*�>��$LIР*Ji���xpB�'R��(�tќ�r�$�9��\�����(����J2�Rt�p2uz�b�mqB+����HcqS��V�ci���az�~�n��Uݐ�i�EJW➦�8��M��tq����q�B��xm�=,�P��o���2�S0�DMu5�Kg��p�gB)�>��<�j���>E�Ĵ�����٦L>���؀~L,�#ր�'	���|�FA%lpY�8Y澒��N�Ke�Dx��^"	���%��	�el�k�:���9��duM����H2VY̺��ԹC?�Y�:p��)�yxN������m�/�C�(k��������(k��F�g�� ��,�=�d�h��,	���6��F��2��g�{=d��yUQ�W�g7Ϭ�M��[7ZHv'���m�v%���C;�6j�V*op�.�n7 �,C$�Z!�}g2��9[���μt9�^���Ȣx�d`�1�G�G9}2�X:H��Q��3�꺰f�������n��A��X1ݱ�1//�{��x���T��͌�����!����]�Ud���.�Z��<d7��F�9�W²������P�-, �?<8��>%!���@-jM�r-���nqr�z�
����6�%��8xӬ���Tj��E�&m,֬SƧ-�D-S�}�Qy"��<�J�����3 �?1(p�M�G��`>$_�ʧ�*K��(}LTk�����RF�ŬU�IeXA�+�K��d�K�v���R(��$/\X	�֛���uU4���v�^���T�Ƚ��1�̕��u�C�t����G�(�^fF�!x	o��~g_���d�xO��EHӴ�F��\Y[*�%��r��,e��.�Kz ��U=�r����9z �Ş�����fK�$I�����GF�uuuw�l/0���+�'�?��3?| �@�ݝ�9������������"jٵ��E�^����fj�",�,�f�[����4�H��H�r�������������#x
ɬ�x��`��[o&)z�Ӊ327������Sms�ŉ�s/�&�RHk0����ԙ���,�	n�]T	�^��jS�M"���x���"��ߜ�,��r� `|I�-�Y�Ӫ"�ɋt���w�grZD�A�����sެ��{#se@qN�Ɂ\~&���]�/��4�4�6v}�\͌�������j���\ �T�K�@:�fK���m����K\Q6�2[w[h�8���ЫW��&�혌�.#o��gt�0�Ux�&2����:Nv��X�*h��>��ls�TCOP�B��?���F<��j};�G7��Ӗ�y���[����V3m�I�ѓKWt�����&Ɇ�f��hu�ud-��z����m�E\K�G�RA�����ߺ.n޽�E��}#�>��p��5H>\MX`5�\r> �I����5��9�,�b�u+�V�YN�xoťs\7�e9`Kϑ�y<}�̍�ԧ��B; v�L��qr�0��c��0��H�K������u��iΨ֍$~LW�2gP���Gvl�$��0����gP|],��yNl*Ljb$a���ğ6��������S ��}�]=&PE��`�B���3��R��Ր�����5��L�p�`s�e���2����1��]�(k$��44��������ܝ�2:�1}]Y���Osɒe�c����������$C#�1�2�R��t���Y��z��1��D�����P� �Z�xD�7�;�b��@���	^��ѡ��5�6�3�W�p�A�� ap�`n�紣����f�;�ED���r�ԏ̌��7LV5��B�
!�Jt�b'֟�	�w���j63�pՑ�=��1<�t,rV��x������L�ח�Y4/_��߱��T���$<�04���-�~&���d3%)LO�y_I>5٩�d�����3�b4bܣ�޾�[)�jY�I�D����u^又���Е�mj:�%��fk�vv�,t�,.�ث@�ט�Y�1#[���� 쉤�A>n�͘N��W46)
��D�!��
�x��3C����\?)�+��!��j5r��S��*Q�h�`�wu~a�Ƃ�z��+��\�sr�'�go���! ��8jM��{��'��s��8��L�k�t_��e��ޟX������dn9ͳL�t���W�������gk�9�0��������@�GOx _l�9�|�V�8�^���gAPY�j(o���o���U�� ��j��=����4�7'�as��%iۻ�{5�<`�M[�A.(g��*)w:���E:��^�w���Y��rv�%i2�q1����??��t*���</��"?w��6���	�1&�����$u-��M�)�����=�\O� �4pU:� ����ؼB��Q�<�Lj���s\�jN{2=�$Y��~��J�/��tU�֑CT�55zeR��ܕ�#���a�ꍹˢ']ü[%:���Ibj3�y"EM��0�$n]�1��T�%�\�QȎ��6.�1�lp��Qt��Y�G�-;�%i�X!�V
&('��J��10��T<aS}�;��(�V�;�3ag�hݞ:�w��}p.'r{@�Y	]0��=�:6�nn^kZF��w�ʤL/Ks�$�51�R\=丙d!g��&�a��u����Q��=���hu�g�L�Y:� C]��'����B�N����L�mw����Lm�avR,�G�Qa!�\/J>��b[���e\S��sV��2�I��I%>��H�;�;�t(�����D�#�~��j�+2&eG���ɓZ�^p�_��� ʉox�]fe��>|Y_���h4@�^�>����78�u3dfxy��AvO�zb� a���i�A�I�z�����/.��������M���l8A�(Xx�cǡ��
����2_*?|v�����
�q�Z:�08Y�Q�:0���fj��v1s��R�h�̗��ƻ�~s�>AcG%w�+NH.�4R���Ld�Tk����c�يgySKU�@k������W7���3��tG�2ʃ��n���.�q�h[�h��۩.@��B�C�9�'��9W�|�w@:��y�L�$�;�V�y<���`5��x��P�M��,��?�YӨ�d��,�۸^�E��hf�����/
�-�����A�~�]}��Z\;��EP+1�$�D*�5g˭�N/�):}���
X����󨮵y�Dj��^�a�f	,��V�=�F�'M,,0}$T�t�p&q��1#��V}{���ϙ����(�D��;\�34���؃zl�����Dk�%%�m;2E_N���>=Cd�+���8��� u#~����]��o��M���4r�aäw,ϱo�=�[9<2N��[�&c�����9P���B��M�-�����Ϲ�����f<��֦��ʭ������]���\���ٖi�2sk��gr�.��̡���GP�6�jK��o��=�i��	Ǖ�8:���T�'(�lB��`�-jtZ��pz����1�,������"�L�Zwp����D�����v�0(^�&�֬5,�����6#{s�Xl�t�\̸e|�2V�KM]��u��#��Įga)/Q6��U��C5rO3n�}�l�cjA	�!۟I7o
z@j���+�f'	mV"k�i,M�IL��Ɓ��!s�#-�N����;�e�M�e&��=á>�>e+e(u~.zJ�0e���לv&u�T�5��o1���\�~{� ����mjN~BI}�յ�"�
]��3��ֿå���TJ�*B�%w�Ǽf�ܚ�p|�n�X��.���U�Z�^@��G���롑��X_O��A����w�i���@A��p\����r��cb�|{v�  -6��i<�;� �O?�r�B>&�K�*��J��h�7�����I�ғ��ȝ�P��]ۍ�Ѻ��yA>�S�=�(�Y��F�EK�x`uZ�uRP����i=PQ����G�s�Bٗ��%�Z�3�%6�B��"�']U`95�n V�[g*5�E��dZ���1�������P�|i�n�@5E�6<����Ʊ|����|<�I=C�ct�%(�PQt����;oSozȢ�9���$�v���°r+#�x2���H�0E��L�/��\h�y�p@}�LQ���@q&q��������5��:�|h���	�8fL��$z�捎��,Ae]-�)ɺ�Kƭ����}�]�(��Բ�����`B��_�� �=itaw�1ˢEz�簃��#�O��A+���q����+��IAR7��[)�fa��^��Paj8+�S�J��X�ԫ^&|Τٺ�sJ{�;!%���;����� zV�}�=@�s��.3�s:Mc����a9[��� 3;��6�bxqnc~��Me$ybVZ�~T�a��X<c��0/q�f�^�(q>Τc����I� �Xpe5*��!ȖP0�����9�	J�����27^b{���� ��Zd���'���鯘�y}��{- y:���g���22,��/?�Z\]sVkQ���f�=��<P�]ߚ��&��8�� e(��h��4�.H��L%��r�;UI��	sM*Ki�ǻ�Sn:���ȶ8r���وQsO�o�C�ה�Gh[��!���X gK�0��=�;у˯�ԟ�TE	�!)p�%���P�}�Ӫy�on���yd��Y)[��>�ߜq���Y�{{��F3m������Wp3T�z��Я4O�.��̌;SҺr�f���D���Q�<����;�4� k�y88��gord&�k4.���z��T�Z����G _���~6Ӂk��_���!�4�k�S�3�B!�.�~�)-���d2�7�(�®Z;F�S�w{J����xf�����n�2�
U�\d�X�'/Gr���i}�N��f��f@}�NmY`E$��5�T �\���*3�w�E�'	�"���@�ĂA��SY u��8K�p+wD�F\���ܸs���!�25��.(ɿ�?g�VE��Nn� ���ȵ�����fAG��D`C�;�
F�; �j�S�I�	�lf�@������^ѫ�Ό-�fd>{41���g��ѧ&Ѿ���93tgrq��tx�#�(k�����H�����W�*��I�ا��$	PE];�A@�����Y�p?�ĥu&Hտ�{{��Ng_��V[t:W�ϝ8��^�#>c�k�|�^v�n�������^o�bk�MlG���5{�I�t8��cs$������	l�}�6�\���f;l7pzd[���l���C�A��H	��:ql`Iɵ�
+�?��xn���qMr��L�&�8v�(�#�x7nt���%}靕��D��Ŏ���+Ǖ,nltKp9��*@��#��F��v1��l���t�t�"a��F_�Q�kq�A�H�+o�uA��5;��2G��y7�P2�=c�����k�(������En�Ef�3.�ˡ��w�8����O�˜\���@t7�(��Ʌ��&eV̤Pz�>F�b﵂�y�Ɍt��Kc?o6�}���Fy��Md�tA���/w2翕�?
���������	.�"�*��QY2]y�fd�|����Q<�����;��v4WD��k���Rq8�8��J�(��X�+�Np��)i�2�=�t{����p�٦��እYv��	�x1��t"�Ou	�6�ݠ/ޮ�lظ����{&\�ܢ�Np6��B�9�M��
A�P����|��]a�v�MQ��4	��v�;	�dO�D�
��s{#����������z.vRj�0�K3�^UO��ni5��+o3+��AD� �0TA��;��,�^G�D��ͥZrp�k�YD��??N)�l�eI��Sͥ�q\�T�t��L����V� 2� 1�!7(=pӣ���4dN�+(��`ef�F�����5�wS�.pL�8q�SoΒ���ٌ#i*A,@� ޅ����#B�gi��䛡�͉D*P>2P�ə${�h
c~]�3�.�919dR�8�Y]�.��7��;6��Ғ�6Bބ��7�BÂ~4�t \���)�~B[�v�F4j@w�H�2��ˍl!�yZ�w��L�<��2%�9�/	�?	�P�Y�?6:�����vG<Q^z������05wр���=f�d �c�'���&�yP�}��|��%���#���q���f�R0�	Z��Sm����H���7����� �9����l�0@	�_�E=����k��b�0�Iڣt�|�=�J��/���@�Lz��0tJ���A|1�u��lTL��č�F�ٯ��ėB�sH�V4��s8�z��2O���xl�AF����q���^q̫8�.lO��7fO)��AxOk���(+C&��[E�۝'����N򫓨)G���v��7�I��l@��x��f�?X�d��#ٌܱ�o:�\���� ����n��&��S��T�;�OY��t�nXv
��B��໒��K�)�m`���*aW��`P��s��Q:��J������`��;2s�2�Ǎ�a�Bk:Nr�.^��q�#�I��ߒ��Qjdb����(0��F�4�.i��i�AB���Ժ���%x��\�^���t����V�-�5��s�$�
��I�Q�
�cl*]O��vg7��k-��F���_=bF���햍��80g9 C>��>�M��;.P�v���A6V[f��t��=s��XF��I�%d�p��0�U���]l.��⑝]>�#��0��5�g�L���X���'�$��4"5�X�m��hrG�M�Q ަroi����/ &�SI�ZĂ�i�e���9d=��D~A���s2oZ0�$֣�8��tD���]U��Щ��c�E]G����PL��QG��M
n��*N`��-do�`uF!5��A����NA]�u'���ɛ�n�}����)�O��<���.i��'�����z���z*��'��
!�b�}r:Lav�cQ�k<�$�6#�w�'��hn�ML���]��E�ɑX���,g���d��3DGs�g�s5a̐��e��V&'ň�E�n��vu(��� fH:����푧��x���7i���ܹ��hL��&��n�M��9 ^���9q� ��h~\��6���k{{s����F�nO,�;�a<���α�pI	�B���՚�+��)���*j�N�a@��[Y��2C.8��ĵ��AY%Z;�>@���W؞���qn
����y�z�	��۪�x������Ā��^���#uk�B�����F���7�YNa�����.߅�Z�o�u+s�1ج�����%��x�,���%pJ�]�xq���rr>�e�=(1�4���vr���@]�����	J%������,�Eo,�8W ����9���Qr�^��Ar_z�����������i ܙB8�cv��#Ae��Q�(����("$��h�x�;h������2��_z��T�,� ;w�1�5���K��Ι�y�t{ח�q��:Q�	,�0pp��藇�b��TԌ D:���.��L,N��2m�7zO�x�M�M���2��:��$���-�����o޲K�Ƥ$�fZ�m�yP]�'�3�i8�U��	�3X���}�~�H`�NK!�á����f�RNJU��n�����ʅ�����P\���p�a95�=�f+�s�H8?Nui.�͝;^�4�G肺�>1��w|k�������M�������5�5����E�4��[���e�w���`sn2KNJ�-�9��+��ZS�Q��8W��{V��D,4��z&��:����m��=���!�$�Fc�(I��f���E�:W�3l��y�L:����b�B0���4Ռ��N�S\Y�ͤw�� @��N�x�%�T�3�����9gg�� p��<������$��bS#��Ӕ6�5��O��*
|'a>f�3�,������=;�:eΒ Z�8����+!��T,��Y8�ʇaGw:6}�LP2ǚ����m��	�Q�Av��'�rV���y}�������.n i�XB�C���%z��c9'�Y����Ɇ�S<O�̊�
hy{v�7�5�>�42H��7�L]4�Ҡ �j�C�;A&0�<���f��'��A�0��nI�]�<��e���Ew&vf���gk��9Q�˸V��/-�E�(nGzUb�ql��Kfn�0=8x>�(o��[��o
^67\[G�k� �	�
��|�*gp��W���ѐ�&��ÃLAn6 �c����\��1�iu�K�_��ьVH�%.fN��ݲ���%��"�jz`����Z���u��f��2+W��ۺ>7�TY�g��{ސP�U�[��6g�{�X��#��s��ś�آý���Ϭ����Xl�x_��w��2���t�&��C�Kl8Rߘw�KSZ转���l��Z��\�;娡.75S���j_�5��s���=<��p���$�{Z�'�U1Ώ`c��^ꑓ��2N�N�؄QY�9
�dlX80��Y^taJ��&�1&��h  (�L��º��v��\j��C!��s*j�����en�?EY��Z��.�>��1IzTA/2��?���̓f�:��:�2cP|�B�\����5����������ˍy�L.K�:kA��%��ݲK�X��Z̩�7)�gS�$���0��Y񛬸�K8^M�᧸Ɩ���?�ò���(��iej�+q�C���B�
@�s��V��k�����AZ����7)1�L�(;]Wf�B����V]n��iQd�h! �i"כك��(�J:(�F��9���Ö��ճ.��s{�0�4�}Sd�E� l��2��6[]��:Q�Ĝ�N��Kkv,���؍rk8բ�	+p�2X����9g"fٳK{�.�qֆO�F�	��.��6�w��Ъo��a���e��]_(v����nO$4�#/g�2Ct#V|%��-UH��~�Y�G���QW�.cY��@��'��_�t}��M��w1�5b5��@����j&�zŹ�`O&'���R{6���習�XK���	ѣLN��$edʬ�\���<����4��,]}�uo����t!��۱X�ytbq�2E���.�-�W��rO�_���2߳��K��Hʜ%�T�e/)���|�`�:�ϋ��0;bd�I3=	x׭U3�-n�;@r7h7p�鄓�c�2(���rȳ?ZO��H_q�-�X���u"�Z5�	AEy�,���b\A$��6j��yƀy"��8�D�v-�S��y�J�������}�v�]+O�k�R�$,	�V�X�#дf`.��P�]�=�L�ur8�����ɟ����p/Y����;ȹ�d�ZQ��-���!�Z65j&|�B�*��um���g6Gc˽��6��n��_�di��^�d5mnPL>����]-�{N�;E-���W��?ą�����09Z�4�7�.�ì���g�'�����A�e���y7�1�����2�wq�'��у#|��l�wY,��xY4��-Kϼ�]������g���%uGy{�&�uR��)��dE��M �:�35_���8��iY�|��ܪi66ȑݦ���c�b`S�v���nGo8�Ynw���.�5�xb۫K{����@6�a%hxt�|��YK�q��YA��ڻ�<����C[ĺ�}�n* �4�L�Rv��z�Ex��b>���D��GQ�D�620ȱ�J��]}�?���c�zJf-�L4�a��)��	s�)�Sklu�MG�d%b9)��jv5W"y����d����C3%f�whB�ƴ�bA�^5()��9#x]LF�B������J�5ЈXq�G/�v�m��䃻���t�j0��j�7���ۗ�>����!7���_��g�a��%�D4��ǔ_��O��"�h�.���N���3�1���R�d�bmW����1��n�E��qϜD���?�E)���q\��F�	�R�H8�ytB)1��J�R�����hx�G�g���c����&ޚ\��f���$8�O���q����E������C��let�$���	"�1�('t�A���ݛw��>��䃶��g���(.ף�OX�"C�_�����jH�'	�GΖն@���[���QcȄR$繩$\�DH���V&;��+R��[YPj�.~��ɚ���l]%�V=�=�</}c'Ԝ[7	�Jd�EʸQ�,'�Nf�b|����(YN0�jZ!��� ��sJ�,����Ӡ�8�ʝO�C���Q֙�t�g�4�L���)�Fr�E�����]���;ylF`D�9;���S@���$#��� '�1�浩χ%(gѺc�+��׷w��n�?޾�{��^,�9���^�6������$��&��3��e)��*�R�cE�ˁM���7��+'�a����Uf��2	zF��D��|G�Y�b�N����D���E�?�̇Sb�W�ʝ���y�ſ��KzA���4S@V�(Q��}�F~ˎ��Ϡ�����A������W�^�c敞�P�ת�~���v��2�s=nH�1�tg��?�ͳ+{|qi�Zfܲsz�����[XeY�/��!3�z��k�N�ƞ��<�dP<`Lb�s�N�6��y�y)ȍ�
�cTQgw�1��(S�=��J���I��T�n�!�g�!Gbk,Y��6&��A���Z�k�X���p�,�'|6H��N����w?� v���lM���4�!� ��斢}Ƞ:W�f))\M���k�n|����\d���t�}B\���{���5kCc����>�vU��NE%8���I����:����_�����s _�3r��z�	��`�:��gX ��ym�Lm�xIZ�	/��9�#��w��/��4S"�3yB�� �'	\����o^���⹣�r\� x��*�(�`��MH'a�z1���;���������U��f2��`�Զ4/��^�b�G���L��1����ѡ�eFi����h���>�%����v~��L�Xw�p=��{&�'��A �%6?K.�ʍ�f���$��L	�(�U�
Idc@�*p����R��w�d?E[!H�(n?6�!ƥ�҉�'���{�i���)��dۖUS`���?,�9���O���mv��7��Ec��i�M�i-+�&Y�p<8�H�Ѣ�Яxn�;eu��n�o�vwǌ%<�adn4(&������~S3y�%N�]�3��k8jsSv
��x��1nǓ�����(�!���=n=�L���Y�6�JV]7�W�<�O<~�7����#�X`j�sf^X��v�w��#-�Լ���#k�M7nP�F)��-2��%z[pю���Y��o!�E=��Bх����� b��h�L�e���0t!��!:�:�f%���M-�:ny���n�jP�{S�3��@q�����F� ��ʈp���ڃ����s���&����i�	Lǀ��j~?-2!�S뚦F�%v��F)��i��^��#�Y�� t�$R�<p��D�ۚu �ƹ9��o�v���>��G��3��	z G���w/}�� �!`T�f���nr:��+�g�IVs�-6��Y[����2�R[��<L]ɖ�2�,��'�W)aO�u�L��z/yG�w��'�q:����Xs?f��@@���a���2��
3�uQ@�Ae�,�Q���tSK��~�.���rp�z<pN��]=��g�W����ʴ�&�����y��t�-sZ�0ˋԲ)��Z��6Fw��%2�$��M���"�"���{�آ�ѳk7L���G�h
V3\/�e��sr�1�KT���='�ꈳ�y��|��
�:�-�ظN�7�2̥We1(�?��	�R��WE�q66:}���)Z�j�������yH
�(�'� �i"I�6NSG�v���4�gsqs��r�l��U�CF��wM��?7 ��D�Q��$�z �Aꎋ�sE����zc��aep5�C��8I���/�q�y��h���'�:�)���E�g�İ3��4��E%�y+lNsmy���_��y���_v)�,԰ˈ��-_�Hmz�����U/�O�O���|�bD#8I�Z����L�����O���܌l�xl2_�XǾ۲;��খ�����k�]=��
я��yU����g..l=$f۷����������@����:�>c)-	��v�x$�R�*�O�A����f�_/��d��ȎP"���R~�P���x�� :J7��
0Fw��Xl67K�����;��Klf�r�QS���F,�ZY��6I�b�-�����D��an.t�u���H�x�n8f3ѺxCWB�99.VB ��؂�3�q�P� �y)ۜ��F�י��aoID��Z�,����4�S0y^��-v�����&w5sĈ���;�z�a#���X]N���u�3��<^>z��X�;:���n1"��=�^i(c��i�q>�UŨA3�8,��F��9�:p6��ۍs�v�XZ�X���+Q�$[T9O�r6��`��Y��25�[]��p����s"��R����E'�P96�sAr��P~���l�����o�vĵ8���Y`�܍�Eb��	kt�^y��`|Ju��x
�R��R�Uk*���i���]�S��ġ́o\dlKR�dKn'��N�{�e���WmǗ����[������O)X�&�~��M 'K�Ԩ���~a�g�lM��$��r��0$J�x �%�Y�H�-z;F~u��X(eBn;=7dY�C�M]z�e�Ԡ�OeE�e��˫+��	�~&L�Z�� e�fm_������^'n4)� �U�g�U�X�]�� �;a�CL��	�_�j��E�V�#x�|�G.�eS�2k�� p��<	���"�Y`�p)�z��>o����	Ƕ��I�A	��8i;a;_��)̜�(�*�s�/$Y�R~�C2�<�U�V����_�،�%�HJ��X��s��Gk2�yTcx��hs�4"��:kͲ�,���I��4L�l�gGuB=����ڦ�{��w|����S-G/�mS�odv}�4���D�x�:��+�Ts}�!叧P�}��'U �(��k�48��l���$��V��ejI�N��,����s�0�j����)�4-K�(s����2�99}�wT�ɱ)�|E&�ٳ6b�%h(Ss6a���ɢ�G�=bf6�;��J`=�Jc�����|7~~+~��p���7���gU=�7�n���ϷW
t��N��������=}\3�z����iL�-�g7&Y��6���������n��Q`w�a=����	W�'���E �����3X��(-�yTS��K2虙%o/ӡ0=�fk��P�6���s~�}92/�GCGqTF�=�(�l��I8�1{�0i�@ީ�f�����NC�a��N~�U����������tk�ULSVxse
L/6�<k�S`��!��M��<�$�v��l�vh�{(,��B�T�I�94�����U����3c�}��I���s�P���R��Zr���z8�[̗ ��]� �@֭����8וVfd�?�{c�H��`OVΡ)K�P˦�_��n3.X"�We����<�L(	B�C⟦J/O>5v��#�O�Cq�[s�]��,s��|1�C+���O�����4Mad�Y%~�x���w!����֗U%h�ŝ�6��|���;���uA)���!�o8j,Љ8�Z��0�Pm6=�F )�E:�t��U�����|yE��������/�ps���gϞ�_|a���K���y󓬬�yrI�v}V�n~m��ojF�&��l�e�)��G�Q��KL�´�ܐ1"����m��e�oeJ�� ����9���D�e6(|��U#&G[,��݃�7
�߰�2I��G��a�))��9`s�Nta	_
������~AY��H`�����_Mĩn���k�k�/�D�Y����I��ޥh6Es)��+)��`�u�]���-;$����q����6�&ŝNj�С���C�3�2�8Aua��a�ߛO ����0gu�l��Φ~��{� ^��a���-K�R���qgW�>:�{E������/��t�d# N�(�[��##�_>O4��D�P��9�߬>h���^|��V�H����n	/�y����>x�"\$EG��<%� �4��Cb���m��M`>�d����O;�Lٹff��������,Kiit�끘I���t|Pe�1���El�24��k����r����İG��~6� �Q3��_|f�]-(j�&���ɓ'���3{�♽���fh7�_�b������8r6uY?�ӫg4*D�z�ּ�>�7�}Mu��ol7쭬4	������k3�\�yᳮ�:�h��C�h�$l����BʱE���d��Fq,߾}˹���A��S[�(��TGn��HAE	U���C�2�!^��{���?6�����Ĝ�L%1ob4h�̳z#�kY<��!Op��Q�n(���)3$�4j�y�M�C�BR�@.3=lR��#6��A�j�V_��D~&Ec�68W�zn���&�C��z͸�X�1�`��/n�d��8=z�pS�Q|r�����	ds�"�[�d������˟�Ϛ�H�H����@�xF���v^�bY���<�#.B�F�ſM�tsU�k�-�lz���D��*�� ,Jj�\F�g�� ���l���I�a���ɃhLKi~=,���%�4^j���\<���^>{n��/�q1�!ѹv�����w�={�)��N���G{smk:�${���>��S{���Q�vY���v��fP�;z�_^�	�i�f���.�o����k.��AȷG����N"�, �]l����N��>��7�;ن��7)�lr<TMNR��Ѱ[�`2�U<<szH��=)�@Hj��V���'���N�5�$��s�������Om?s ��jYܣ%����d�nZ�q+.�{��G��~��;0Xah����l�ڐ�v]��K�O��{�3m�2s
=g��>ZY���Ʈ;�7f�1ss&O�B��!0d\ ��k�8���|b��nKǀx,w;��݃�-�⇏�XZ�pX�^J��-;l�� ��E����(�37,�ز,đ�a��:�7K��2��8���/r���������x����菶��y�42��:�D�v�i1���=
O���K��W_�W_�Ʈ�����ٛ7�i}=֓�zK�����~�?�[����<޿�Og�^���4._�o~�[��~gO��p��-Agd�׵<yQ����}c������J?9{l����������|�h���ǌ���k�C=6�5�ã��Z�)2}mZ����� Ph&q�����t��i;/ͩ܌���&�ʣ0ǝ�g\�pF��}��^*���������o�c�
j�5�ȗ��5T*��<��g�)��6����ȩ��(Ɠ?����!�#$�9�O� �y��ʕ6w<Z^4�6*Ա[�ȿhbQ��Mt?0���Kؚ0�n�����'����|@L�1���Y�w	9-i\���j�<�Z��py��҇�j;���F2��(�#�u�������."���M�s���ғ������M��=w��|�R<���i-#��#6�r��M�\B<��q,��v���jC�=(�8k��2�$΂J鉊C[��P��g_|������y�.Wޮ�8�����>����_֒t��o~2{_3��~��W��_����/mU��,�.�0E|y~Uˑ�����Lv8�Wg��뗟�W���~��S��r��ښ�&���k;�Y�y����7�d��sW�fwk��}kp�!�d���Nx���Q���0���;�=���˨����p=a���u�%ů�s;q�V���4���6f�l(H^E� ɘLRg���H�5��y@N�E߮��u�4NSi��f�����g��H�#i�a$i{'��,Փ${6~�\����DH\ŉ�1 S���t����Y��� ���_<66�V���i7o����8�m�;��4�*.���r\/Yc��Y�|D�������2���4�7qr�}�A6�n��A��5'�x)#��<�Y�>�,���}z��{W��^Wȯ���l���o쬥9�]��q�������D�osPO^�S�]B�ё�GRѼP��nR��E���,9���?:�S������20�D+�����Zo/jp�w����.jv^�Dկz|m��������?�3�m.���_ٯ?�ܞ�]���X��M����<Y���v���y���f�I���z7�r���[Nu�h$��n�Y�j�]�ff�E���,�GCb����Q���wZK���͝o�gl�܍�Ԣ)5�u��@��yR�|F�y�1�:��߂_��pݤ9AG�%D4�A�F�q&�6J�F6Qr°6[Y�OĭL�AR�F��K>g�m�@19p�FFwON9?}v���󏿜
�^Mi����SK�gJ�'Or#�^�@�-�P�Ohy f��&2��ެA`)Q�x�An�{����+��Sxk�
� ���A��S�)*Sr�ߎ�4�?^RC7��X���<m<hM���^�XgLL3N�m6��z��e?���/"�&e
��q^�Q&99�/Ή���es����Hp3Ԓ��,8d9��x�G--_>������Ok������}�����1=��G5��=���}bO�<�����%���}��}��3{V۩�~��^�\3��PS����vQSK�GWW���{_��qw#���\hXʴ�\��� ���{0d:�G.^�	Na|�`?��iSY6�q�>���b�n��t}�R�Φ�?)CS��`��}=S���<�|a9[_�)��������,��\�d �_C�`=Ff�?���j=�Qd�'��'t�k�9��s��r�h`�����']��@�0��8���9����6�o<~Q�4��F��e��\�}px2���4h٥Y>?2�ef[<���������]�~wٔ�����xh�=Т����k�)vUCӟ����1��J��<8���(�3��#�QJ
*K|���l��<��ڰj� ����a.�:����k+�VM�Ґeʳ��l���Yً����ӧvwoo��ۿ������y����K;����դ2������LnS�b�1�f��ym�}�ʾy���twM[%�`������?��\K��� �,澾<�[	 ������O���JǢS��F3"��Ș�d]s},�J���~�)����u�4���DmA�=Wfy�����u>�/:���<`4����Tfj��
Pr⹎�[ 4<����̝H����[�˓rn��I��N�P�� �4`h���ᚡI���$�Kj�{�%��\|���g���/�7��aL�0�(�f����66�nh��;��&^#^��v �O?�Q�}�U��4�����JX�9^�4���.���o<���L�����>�{?n�f2�L� ��I�ߐL�Я��ÐՅeT�����V^sߛ��1�s��i� ���;JS���|,A]�X"ao���a���`����颊�[�f�ٜ�5�P��F�-�Md��5}S3���������������~S���OH+�����Ћ�����������������Ԓ���l�v��ô�g��������7�?~ϛ�ef�W�<`����R
�5y�A`6�N�KE��`�'����p��"F7h��˕���Ѹ
��?t��1��2�õF��l`�%>_hV��Q�#�k�����q��UB���<W�e��4��IW�pƅg��::Ǭ$��I�p4\�G�<�i����-
�� 	)�Pe�����T�m8;;������?���	nkݵU�
/d,�N��eP����J$�i��[R<�[�����X��K|آc�}���9�E
�SPZN��.�Ω�&�@(�{�U��9W�?��@�i��J��,��~\�.��@[aȁ�{�U��;} ����Tn��_�����[�,�����՝���[����Y�Al�#E�rn��t�����9������ˏ0,v��(��D��6\����!�����]w�o��d��}����}����I�,�4`i�#,s������G;{�31`5l"$�̾f$�bty� �\fy���:�M����0���8��UD�4N5�����1O���ݜ�k�+�]ώ̥6'�uC�F���"c���4W�h]���ZyhO��47������Y�YkjpL�W�.�K�5GXr������u>�����u*� :�d�fn��>���*��$�dq��`���9��VP�	�)J3鵔?>�X1V��_��A����SPN�n�|��� ���r��� �-�W�w�Mid��f\5���gՁ�Z�.�\,���7�%��t�gw`��mN�����\�$��(�e��/� ���	��,�v6�zF������k�vz�����9���G�Wg��
_�"Ge|������z��2��i5Յ����t�����.����)K|`1谁�^p�l4�i��S�������G+7oT�ۮ�V�l�s�Zo�b���}F]��y��2�g�)�&es��Sc�(�zE���f[e����6��t�kD��BB�c�Q���@Yj�;eP�2��Nr�Qe�k��ꛣ&�͔�1T�6qC���F΍���	�e�3W��w��N��;��L�_�g�LJ�B���6g���aN&��?���R��a��=��#}9�!��E$_\t�L�u[�������{�e�\GD�>�(C{�iQ�-�c,�F�}��c򡾱[�܋ں�� ��E)�H�Ś����-�T�K�q� ׿����(�����7��1p9|��l�Rɳ_�Z�s`/��K�9��nr2��������J��41?�����'�r��r� !�c��$T̀�IL��a��|č��͊%+V��.��Ef��4+ |I�H�ԑ3?�Rx�.θ.>�q�F�^qU�ڌbm��j8LN��~,�/-�P�t�P��n)�w���e��]Θ�+C5����S��E�l߇?�jfX�pj��� r�p,���靻Řh52��٣��)$�_��q�`��k*�\�~�m�Q.��S�c[`��÷o׏�n���_dVY?xʬ���N��)|o!�'os�Ʌi�;���s��ٖ���A��(|�k�[Yۻ��/���̙�t~
��Ǵi4E J��ͳ?S 3/�G/�3�&�lP��2�8[�A�ۙ�f�����1biI��Ì�w�E�G�N���H���_��x��F�Q�ܮ�.�q�:����=���QW��\��ʧ�p���7����C?|��k���MN��9w}��(�L�VNǅ[�`��`PɲӃ���I��D$_��s������$4O����a�8: ?�L!����3-�N�ڊ�͔���4�*����&+�'9c�6uN?��[�ײ1�A7P�1��O3J��EuZǸ�g��pɋ�i�1ɘ��I!}r��ٗ�Ϗk��>*��[!��;�m��la��	���������/��~z�3e���UN���O�S���7P8�*EH3�,m�d�����`g��g?�k/�ݥ��ߴ�g`����h�8_h��=v��ٌ�Cy��q\�M�,vn��d:N���"��_�D��?���{�Ŧ���v^b���_��^Q�ĿSPm��V>��D]����,�u����|ˁ���ޞ=N���Ǵ���̩G��y�~g��[;����>q 2�	�$@����Q$�����t�I���D��}�g�zsi�n�T���<J2
=/;�@�GI�>����� ��� �+^r��Ѱ*E�7���8�Ǥv�j~>a���f����?���Z�^^ɢ��o�h��pԌ���2���6~���{�b�(��r��oY���AA��r����1�p�{�36�ɂ�x��9�e�J�����nW{���=��J�;l�^�g׻;q�^��l��4d�>����NR ��'���dK������ Sj���.���.J�e# �H~s������Rf,`�f"���28���3�����!z��>s<��n��c������IS ���1`d&�]�z�4�l���πA���9���`6.��b��:�>�-9����
�Xx�E�����u׽�#m����~����~���x����~���٧���]4����1!��=���k�����ڤ���;��OMF��4�x�{ =c������^6:�(z9�cq��y��%69B?��lps� �D�5���T|S�	���7��\xC�|m��,&��y�LN��k�}��m�I͈֡�Z�����_ՍDλcs,Ä́i`���,��y),,��ْ��:�ͮ����T�~�l�.y>�X�n������k��'�g�v^����̮>��^߼g��nwO�ȃ��oV�IU���2�&����9��M�&�\��Kf10�)�VfH���b��ϖ��i��V�xP�I�������9޲x�ۍ�C�}�P� Ω{�1�</(x�%�ھ��^
r��l��c-߯�B�!D� �8�L�$[i.��|k�e�/a��f��r�m+�Y\v�	��*�R]�w���;{���/���%ʳ�����?������7���6����x`h�k%���G6�o��x��v�\���]]��	�[���r�J`Q�hmQ��z'bzO�-<��S�%�}�#���⚜ʢ���)@~��$Bga��&�"���XB��{Q7����A��\���?�����b�]EнĽ�T�O.Lg����v�As���`�7��Q��=ۦQf�3�p��g�a�#/?�\�,�Fj��%k���<yCe;yrIі�Y�ל[LvF�pOx����!b�Y�zsN� �dn'A f�t}m?�yMũw�ޣX����G����Ο~|N�> tY�N�z�O�!�r�O�\i�,M�O���8�XH�wm.;��#�ˎ�J�����Y�������kE��rctF�(�9,����%�/���W �R��s��3��SDi���ֱ5tm���_�F��I��=�""'�6{��޵�Ke�t�������a���Q�J��4��X=��5H|����u�]~�؞����_|eO�s{{��
��/�ԯ���<����}��[{u����E-9?�7���=�zl���K۾c��T;�� 7�/>�\Z�zc�����]��`]��w�7���v{so��{���En_}��]�xj��VJ�8���+RO8�􈛳�zP�dw�p���t$���"�zR�,�7LHi����Y��E�v����zN7��yd�8����D�6ɘ:���2�o��q�Ê���<���ļQ��x8�[�ݾ��C�W����t�|&�@o9ē�Ș�q�$A;��ʇK�o̪�䘝V�6�u�lhʮ���?���nV���O��Cg�gu���y?�{c���ov{{���L�������nz5x���,��4;���I8���mx��_PZ�w��c����"�.�Z��`���e���D&�M�V��'����Zf��O,�r����bW��Nǽ�}��s�#���7���j��֓��i���:zz�.Zɞj%�
[AGԖ��_�Yo�s46� �Ew4�����~;��V��Er�Wp4��a�]o�SMY�@�xr�Ȯj �|�E���E�y�� @c����ξ}�������[�2�8\��{�9�4�w(ek0�������=�����5S;������~�֎�����?�xd_<{I�ilD�=���������/��Փ˺�jY���^_��>�_m���L�s���-a�96��������L[2��I�a^���#V�� ��S�:6�,p�'AXw��jgӝ�������V�JxrN�S����4V�sϐ`�YN'��d��Y�g�ڊ�O�X���v�u�}�E���8I�jS�T�o��X�1\�xF��M-YߝvT�`�zN`vzB�	� }�r�����=���T���S���˗/����_ܺ��-jl�ٛV�Z��l.	Fv�Ǜ�Xk&��21yf�?�Y���{�F�������b��X����^r�F��_����x:��;��90�[�j�<��s��T��Lh��E�*�g�sT�t,��)N�s�Y#����$m�7�(�u�����%v𜖥<:�a�7"+T��1hQÀ��n��W?�P��z��L���?����k��S���pk�T������^Y��	���ƣm��|��~=(���n���lun;�s�������k�co޼a����W�$F��'��||���=���g'�������kp��+'x{�!�I�u*����$�K^���R�K�h�>�������2=R���mcg5��5p�AfpG_:��g^x�S�ٮ��,�0�����2���	I��y�x�8X�D\ead ��HV�J�A�nZ����X+��t?9�����r����X��E4�2=׎:��v�%�76*���9�M� v5�?�?�H�A��=�C���?O��맪�����O��\��>z�25����IHv����r<C?ͅ�'"�Ĵв�vs�����L02�|>c�E'�g�p��/<f�x� �w�ܰf����o����<1k �)K���H���|<�h���1�%��<��ϋ ��f��!o1�׽�)�E�/���ْnyI�Y7t͋������,����Օ_wQ�~��S���5������������y���?�1{�{����=~�=���|�� �����rc�0���޾�W�Gw�2�z̯_�fy��I���j���n�"<���ܿ����`���ݼy� �Q��;��mfa�j�P7e�����W�.n��s��xTW4��=f}!��������3�&�s,A}9�ן��ک��W$���T�c����}9D#A��J�_5'8wxd��*ɧv�wV���,�hp�7�f�\]e�u�A&f�
�f�v��uq[�_�ogo����u����=";,YkA\TبN���c�a%�����'���a��ʇ��2SX
�'Os��4�� 6Ef��f�C��d���7ϋ@D���ED�yd)���\T�	2��n���Dg�<P�G�X��&e�1{y]ڽ��w�<HM<O'� 3{���Ε�Z�����]�Ls�V�`���ZV�G������kz-���Qn�W���;�zHmJ������?����g�߾��b���=U�޽#�����dgn��"�>�@�2���޽~c?���Y27p� �T�Ⳬ��Ȃ�bt�(��лag?�������~z���I 'K"Z����D ���pm<��ܕ�����O�Mn��ǹn����(��\w�Fֆ�M�D��X7�㬆>#6l�0��˲��y#�#�>�]4":k^E���B�j>�È0��D��� k��tPe!衂Y3�9!,]���٢W�2�|�-8tJ;g:���L�_�09M	$�f�ʪ���ΆU=�^N+�z���vKw|����p w��q���o>��
s���f�byӫS�J �gP�ϰ�b���,�Y��v�1��T�#�K��/�����,4��n`a����=v�8��,P�{��b7��,cX��=ǿyr
o��r�%�)5�*�K-	�s�?:d��r�Mn��x��\-]��Qv��v�
��[���=�$�$G�et*��$<b'�f��������}��'��/[k���������3w�����3�������g�r�ן�p������L���q_3�oT`3��{bm�Z��v>�`�4�T3�׻[�����ﾶۻ��o���Ԕ  ��IDAT{:�+��\�9�}�D�q�[����@��-���\��2(d;�(�Y����b��ۮ2��<|�mFi�o59�h�'�nd�������(�~gA5a� k�46���ҿ��&X�j�o#�ztd]%O��!�} @쿳�ט&�Yۢ(�,��S����0�3�q�Nj�P��fH�c'xxkL��=��9f`�8ֵ�0fql�����GaA�g6<�r�-1jY���+>n���J�J���|�̅��e���"x���u�A`BP��C;Nn�U��8���9��������Ǡ�+�~�MS G�h����8wrwS`&%e:����i�rtn�|D7�ߕA��]��&��ߛ"�:�'~F-!^��g�@��̥w�o6-e�b�8���pm��H<6C��y_m׵�<Ыm�Fê���zo�߳�8�_����X�3�V������n#g�����\da[��#ŠS&x]��o����5�]�s3�ٹp��I�p�����}pvٲ�Ǯ
-Ӂ'�e#�s�I���y�]g	)P���H2��0D���{^��o�U;\\�=xQ�3��w�i|&�?}��=�zj;�IMm=�I�Kil�}b�+�Fc�%Ν5|�/a�!S �Z-?O�N�=�e�e-���M�fc��1����{3�͚�2ϒ��f�(�$:����Ȧ^�� $��4��Q���G��Jk�X���`�������QAF�JSL��n�V�.~� dA�����w�M��^���&S/��BV�c�̒3�s?GnR'���< wy�&P����Hcz;�ó����]|���)�#�Co懚'z.]�T���0�I'�|ɉ�97�%f�&��3 &-�p����>Sx�[d[��ye!�A�����>�뼮�{ˠJ*K�mN����1�7߱�{�F�`F���48���"�fU�I�����r[k��c��Zj�����A"����Ԟ�6��1�f;���O���@��3�׾^��?�`�w��z@�
Ru]��>�δ�42qR[9rБ�׍aE� ��AWx�9�Gg��.�e�\:�QD� ��~q(��Nן��Ts���,�"��˫�Qn8�����ގ5#=��^�C'�ų�v������Q&t\��@�	��S�6���/C[���FrBp]S�A��'ev�oj��O]��L/���~�m�Ѹ?�J�qu��m�ĽH�-g��a�	U%,����A��p�����{��'�=yl���R3<5�4S�������y�9'Ǜ7��q��F���V��돿����JǱ�zqʭ����$�����"w�51���� b�)8	�p�	��L�ewӱ+�<���vXhJ�xH���|�'b�;I>p�D�e�EV��;u��8����bb����6��QB���L���u8N^DdWuA����h���8�nTyq��ûeG���]�6*;?�T�� d��S��V�;4�,'Y�#8��7�r�^`��[;�v_of|^t!�<v��k�����
�q�eu�֟oEK(=&�k�:�[�nj������p�������ѱ�1D�o-���ݶz,c�K����� R_c���^�r�Ck��
�4����{��X��YoD4;j���5 2�;�N7'/F�<zL����]�{��i�T��}]Gh�L��-g��v#�޸?����1�	�����#��>������� ������f/?���������Ξ��������i��suyi���̞��nj�����b�~��`�']o�ݑ���^�i^֬	�	�=�$����=��P��'��̱fpw7�\��x�O����b#;�\%96E�a��dtďww
Z�z��5ڝ����Ҟ������M=ȭn��y�:�q�0ȉԣc���}����
���d�H��;�aZ���.��'s'�ق�����9؝D�P�ݽ�)���v�D�a�4�S�aс�ɛ<ͣ��5�j��fB�Mɧ��4���`�1ℯ�{T3�#>%ŒW��d���QM�d�W!�P�P��u��0	'
V��)����V3����'B����;����ʐ��j���z�s����M������Kj�	���|���z�<�ֿ��L� �b͉�42��M��k�V��'�N��>�7�xe�G���Ȉo�F�Ǒ�ӷ�k+�f���k�/d9�	G���9��9��������n��ynq�������7���[��̍�����.p�zs!�u�.j��!hj��8�Ma�#I-�kP�k���{{�����3:�؀@ƭ˩�r`_���R���3�tN�Y��\1���S���/�t��6��IL��V�\Ё����F��6�Q�78b��������/_|��}������M���r�A�F����~� !y����6�z�϶@���3{��irg����rj�YG{��qM���;�^����PM#��X��:��J!����ʤ~��'Wv������M}���n���7��bm��)��SV�N��x��O�z�����}���l:��Φ�RPA�DXR+B#� �b�\���륹�����d�!���� U�5|�N��b�8ک��;ʱ	d�B�ku������O����FQqG��[9��q�5�0/P���Dϣ+!�T`ţ9�lm�;�̀J
8h��M�����0�=���G{\���9o�c-���K|��Xք�M50M��%-�W��\���j]Iy_o&�D�Φ�cBV�F����� �R3&�}$�3X3?�H�zNj��;���[;���q�fC ���\o.d<��7�Aϳ'O�~�a@� e�-�L�D[�driB;v�Q�r�/<5hC���f�Q�:,��R�&n�+(n�q���n���C��[�x�]��w�0�5���K���yR�[h���8�;�&�5�N�O�僲�ŗ����\Šk|��޼fS���+�z��~�o~W3�������d�~���:ȿ��z6u�U���Wpx����s>}�	��o~z�n4�/dl�j)zV�'����;����z�_���
�����Φ�k��9��3�GJ�a��S-���^��;���Fϩ�E�2��zC���v���f������Z_�Hͱ�j�0�^��QZW*gR
s���y����ҝ��ރ7Xfim���ܦrK����Ж��]=e}>�"�r}*Q#���Gv)��$o1�{x���� l����ko�e���X�ǒp�#ސE�]�w����U%o�y����2�Wu�j�!�/�(//`a�'rh�ۅm���<�������]M��~S��T?�����������u-%k �wi ���_<f���Dݽb�g๯�v�n��f:�]��T3��Pb��ԃy��{ਸ਼�Z��j)�nwGg�u}��~�D	���!�C�U���O�l����m�D^]�R<�����X���
O(��odŞ�;�޾~��n� �K�<��(��8Aj���{��-�BÎ���9��(1��^�L�Vg��K�Ս.���)C�~����$y���o�F���~-u��.9|�������ԑ}��`y}Y3���u\כ�# �ۚQc=b-��^m/�/~��2x��ġ7a\���O�ۛ��MV���O��Z&�#x8���w���H�(`���̾���w S�^7�=�4�Jt����c5p!�����9���P7�}]���o�����z�j�p���}���)6�g�9����<��"�t�T���{p;!��p�g^���f��KAm�)m�Ut@#�,���fzB�$X2�b�(9h�y͞�"���m���T���f$���Ҫx�#�d���{�M	��G7@T6�)>��E�c�����a��D���"x�L��_554�A�M2hQ[����^��컛����{�����גv]��N����^K��>�E�z}]4j@@�G

�F������7%)Z���Qʠ���rcRG ��P� ��c�-3��|`w�v�!�?�rWe1剮�<kЃ�a}�D	�w����qo�:��_]���[�e�u6�\�}9�\�NUWW�I��E��� �K� ��+O�[ �� ��&��@~�	؀� B� �H�\mI�%Z"�쮮:u����5��Ƙk�jKNS�:2�=���u��k�˜c��7�O���R����*��'(��ҵd;I�O4��wf��ԠNi�#�i5_�[dȍ���<gxqh�g�>����z:�wr������_�7Vm��i^V�_H����J�g9o��,�
6��x^�MK�����0�xZ-��R��b���F��*sO�N9Wo.�8��F���#�ã"�gr�i^�ӧO���c������/����F�~t���=v��#w49f���\��ժ!�#�\C��Px��+����:��ј.=�r+�7�l��b�C�z�ܓ#V��ZtN��
�(ͩ�3�N��HگtU&"�]���n�FȌO�[#%Qk���Y�<>[�ϒՀحĴ
v�x��q�O�w�) 5�����;j*d�$�t�Ho������ܓU��آ7�y�bŇ`8*$�����p��o,�|fm[���ܖ����,�9�#	;��v���_\�R��T������|����%��X�ky�	l�+ԣ�mʞ*�<!��Ut�%�9>`��K1��a�9&����<12SٱW��,�zkY�h�O�Ȱ��s(��xJh��Q������(m���*7��,��]c�y.��Ն��`�1����G�[�y�ڞ���[V3&փx���|N�s�V�������)C.Xf�u���m��ܭ1�����22׼��pc���*�P���vc8���ӭ 8m�)�:�%,2��ps���ວ�5!?}J�uw7uc��p��bLz)`�~�ï�P�h��`��h��)�#p;�q?z����O,�c�2���ZO���q����F�����Be#ψ@�d1�ݭlXhtG�d�Q�;8
6h�bJ$UHׯ:3���k��L�4�C�-�ׁ^��qv�����-61�7����{{��f������,�E�)K�F�I�È��֔��?j�-PjG�N	<�Ukg!�A������H���)Ȩ7��ǲ���q|q������+��C㖢���p;õŶ(�����8�[���f�Q�pS61���3		+�o�5	a�97,F�P�_�v���4R{bB>�P�Bb>�b��7�F�����t:��*�x�d�K���V)^<�SH�(�!0����p�آ�-Ž�ʀ�6�n�s�)X���&�ð���)Ƒx��+O���
h!+g��s���SڿQ��jӺ����Z�����jv{���j@��W�e�;V�K%�Hݖӌ��y�?�|��o��������D����*�C]�}�0j��w-��#����]\]1��8��5J�2@!d. !$��L6����^Q*s���˅�uBQ(��G�X��}�.��C�sΨ���Y��j��Ĝ�.���������rZ��^!#�e��ԩ���g��k��mdW�?�?y7����rן�b`�؏!c���uF��5��KR�Fx:�3�sg�Ʊy^���1��ab����A?鶉|��lVՌ� e�p40m�a;F�x�u��@ZS�R�K˰,@�C����,�^�zJu�(w�!,ù`� �C�-y*����
�]��!.X*�	��u}��y	E�b�ɤ�u�x $7�=�j��}l�ǙxMHR��&Ӥ�a���y���]Є8(�����x��)�<��;-�`2��)���
�k`��dw�@*Bp[���u��p�k�F�*#�� �)0p�E������2ŴZi�����*0��,�
�~ʊ�K�
�J���n�Ua0k�/��J�/����#2�r$��<,n,֖�yV�̴	0�"�}$%(+R@�SN�f`�A^����+�3�@�80V���;���kߧN����yt���{_����������Tn�6��&����8�z\IΞx�Ԕ��E�=�~x�ȋ��p�����ڑ�G�8���d��\Z R�(ęqõPu>���+uF�չ���xeyf�d䂷]ߜ �T�a�AHD(Zkh���`Ɨ��"C�&ޅ	�!���WB��,*��1*\�ڣấ;��q�^c7��yr��#F47ԯ��Gī��c��Ҝ�d��*\����oMގR}-�Q�
�X�?5�Ͷ��@��(�BM\�&�?�5��CZ�7AoL>r,ǜ#TAn
�a�]�2���"�X����]]]�Ջ��D�1��K8�b�p��j��HK�b�V0)�l*�Dg���B�%�D�V*!�����F�B~��=�22�Eʊdkx>��:	O��r�-��P�W.2m�Au.F��6�r߱9 ?vtr�a��ً�8��z���m䂄o�\��(@3���(f������):8<C��)�%rg���FTy8��S)�Gۈ�Na�x��gh�P����l2 4���4i���4�p������T��b�'jw����i�QC���g/�k6��BBTGxϓ�Cw2<p_;��r� ���̠k!s���2(T�%e��Us���'t-�=��a��D�<Jv"H� d��(2�N=(����z�U��N�����W*7�E������H9J�l*-D���Zl��"}G97y$�����P�E�(��io���צ묈@��q��yCE <@	���;=y잝>!��#�=\�ܹWw�n-�/}N��ñ���S�lr��R�n�V�Vy���������2�z�����w���BT�|�lr�*]�����+�����X�0��xS�g�z�NF��"�e� `��b0 �:�\^�t��T]H�W��`�V͟ X�I�.Q�Oܩ\�q6�=D~gLsEZ����9}�085�0`�@N���F��H��>΅���Z	������=z������ƽ�z���$�pDm�¦Y*�"ճ���%Q��9�Q�����b�@|��
P8�����Qb��Sk	k�kbQ6=6�C��2�^[��&��K�y��"���ޕ�sE�/1~�4V��@i�Kc_i��\k�G3��Ad��h�5�n��<�h@G z���29>&�v��.^�܁�Dm)!��+ِ�S�L>|8����n3�+VN<�,l���f�ٝ�u`s>�+*�e��`TF5�_��YC nF���/�EV��!O����F����TDdi�y���jm�^���(&�W�Ż1n�B�P�d���7�������5XH��5�iQ���"��P�e�?����=s_}��v>8v��k7XW�j='6r��C�dt�"���G���<��cj6A)�����4&��f�~Փɡ;#�����nO����0}&^�d>!Ɍ^���'��~�=�s���m$�C��g��&�O>�������kF�I%����X���!�Ä^CN%{�=�G.��,�	���-�0H��t1�-��~G�ia�L���4
���w��8.�$P�B�&*N�P#y9�	P�����l=R!P?cuh��<S wD.LW�xy�����Wǉ,flH#,T��G5q���6��!�ɢ�*��i]dakLo�]d��^� �k���#Qy9�t���t�AG��3�(���"�p%#Lu�Cϔ���N�8P�+�c<۱l��a�c BɗCn*CTy�K���O��[3�v_#�&���~$�W��~]��345(�q�����:��[�d�����J0��SꢠQ�^�9b�&��U�H�hϵFw�oST�CGt�6�5ۑ���Qu��n8�	n�zA
�l�>������ФǱ����G�'?J�Q �S��N/2��ad�D�,(�>��K���X=�N�$���`�N�w �>�w��� �P\n@FĜb���!7�Q�0;�_�Z����4�C���{t<t��_z�C7�V�$�s���ʹ�����q`;�F�+�}M��\�(������.�kư���n��?���@{��A��Za	eӳ���
�V� ��*^L9[����ъ�^�z@)&8�<�!)�3z�!_C�-h�L:,��r�R�������aZ���7zD�>wZ�o���p�	�]%�[�v ���sy/���������r=w�{�ђU��H���HQ�B�*XOn41畁KN�s$��BD_'s=��$*}�l4��%*����gggntp��� ��$T��&��r��䆛��C����IP����ͽ\�rN\�)�bE	T��VF��øW𴀇{��=^6_��E���`��1� ��zْ�y�L���x��!����1G�<�M����̓��j���)�:Q��A��Y�v�k���c�=�9b�*QfcJ%aM����dS^O��P��d��ݏ?p.�Ç�wi�v��,�g�2�۶$�x!���"#WȂ�����}���10����VƂ@��`x�GC���̽��t���]��]y;���
�{:cs�Px���4�Gm���zEQ�W/_���̝H����S���_w>/��? �L@�|���B�[`$F�ā��h`?M�P��t�x>X�`�H��#0Y�j,�W=y�U�U����-�d������ڡ��x���jY�G*�N&$�!�	5�d�j[�a�a?�4�a�^�e2�3Y''G���p���J�,�HN����Yq�~F����;:;uA��������j�]<`��V�(��I�t�~]���C�da���'��i����Ʃ�z��:<<p�����ch��-��#7�0^��,rL�Ūg� �#(�::؂��f��1�nke�%[J�e-:�6�#��rw|z➼�T�Ł �3D�ڐ^��������:���fc�
jm`խmӖ�娆�x�%��z����t�U�^Ο�|��p���"�lgSzq�����Zx��>�fU��E���IC���C*�zT�n��!F����c� z��>�\�(p���jg�(<0��� t=�^�#ò&��*�.$�7������Vϟ'���l}Kn=Z�O1^^Aƅ�5��VS+&腰��	�	�ؓ��}��3�	E�&���	M*'�������yK)��x�7�\ hFN
���VN4/S�7�����K�e�pW�{z$0�>r>}�=���S���%<�2���D������^^Y��(2t�(�Ra`FrK+�� ����gt�u�B+�|�X�ͳ����Um�F����-��KO&�蝆
|Hr\�]�zG�X+-�9�g;1�i��Q�H&�x8Rqcm��}�@����D�#$��V���bHL���-�ۓ'O��~�Ξ��5e���ҽ���T �ٮ�@H�/����'	����&�I�u(=v��ɁQW�0���`������X	��4�x�f�u��V�: �dգ�,�v���IOt��a,�N�ʦ3��O�����؝����=)�dC�9ӭek6[��|��d�*c��ԑ�=�_��g����|���Pƒ����|��)L��l��x�����SLݪg�9�6CO;dک����&&ƻ����+dޏ�AE��] �[����ab�2��Lq���Y��."�a7��R�R����o�����t_ʰqݸ�a���[wc��O�P7��_�P��C��b��F��ЍT��D&�������ռ7>uc�ײ��J��i�Xn�!a��cW�u/�����?u׋)�*���3:�HP�P+��z�^JH��_|���q/��u�@<��=��}���{�O��2�VwS�`��n9�c==>3l\'�ͽ��d@9h���W≡H1[��0������}�+_��3N5�.�!����F�Ў�g����ݠp^^9�0�)rO�gs�0Ia�p�3�R��AC41Q�K �2R��MDE�pT������B&3�һ�{zl��'O�#�珤1&ށ�g�	��QX�%�<���C�vNO�zc��ěш!u�,���V>(�ȎN��o:�� �Jwz�4Jˍ;9��(E&̏���0S��
��ш�/hY���v�3,TEk# ��:e|ּ����-p��D[�x���Z�=��L���L��^��7�fSI``ۈ3D�}c�߱\?�r�iwx�PM��^!)/�֭��F(�������)ӵ<&�iY�:�7��j��,� z"�Y[�����8	<9-�;k�^h���B�N�4�j(�4}��ËN�yi8�ƺ��h��~R�Up���G�`ݍe�M��J��49z��7�[���c��ol��F2t@2C�\%|9�)U��^&ӱH=̄!���켲szx6	�}��9�h�Ah(�_��I���({#�9=>q�b�@?��t��ҽ��g���e�==gy�p0v���T��Lރ	}�������wk�Hj�'b Eb`d�Ioz#�Bd�,[�bY��G�Ne8�n�
�,ؼM"����k� A�mU�ؼ12�`p�'M,'����O� ��ʇ�<z
)!��UٴJֹ�W�xO�P�>:wK	1c�U5+�^���g��Ξu%&�ݖ�`(����������RBC���h	hw`�_���5���x1Ђ�Z֖��IR[(pS����S��.�B�3��oYŋ9���@�A��\H8<�T� �F���DKU�ЌǠfz�g�� ����'�z9�]�g<�s�'5C�������I8B�9�Yl�b��F>��Ǟ�C0t�_�v���
C�����1?�~�e:(�����1�՘V ��6���9}�^	�Y��� C�ԅ|Ϛd�����s�a+Αs�{�JG�����1s�����&��j/mzy~���~6�6X%^�yI~�:܇7�c��o���K���Y��)�c�jV����P�i��0��
�C'���QA�(!T!aM������%LIĽ��Q���|����ӫdRV1��������-�7��Zj�6�9�>��Г�;�\�Z��"�\0@e��R^��G�5�Tڴ\)�sϯk=�rM���\W�RИ�W\'���k5<�RC��8puX3���^�
���_7�Ұ����F��������he��p�Ԝ6<�Z�r6��c���t�$�?���wqqAl"&*{nb�J�k"��,�t�p��������������1��y ^�Ce��%�Z��6�mIC�`P�8U�+z����[c?�7h�SF��#0Ի^���TW��Aߪ�:Dr�MK�t"�e�7��j.�؎o'#������KH!�Z��Za9r\��ԬX�{�?٨HוAY��b�L�o��_.$
��3��o����eB�����o$D=�,�d�`j0#�L#�B�sL$�J��&}�<��Ǐ��i̦��]\�t\��ߛ�e_p�����D`̸�[q^=��:9C�FL�ຣG�1*��X���Z\����k��sM�"M��o߸U�\�ktbA��g8���#j�_��7�E��)�ෟ�BZ���t�̠M�<���YMT*~��^kw��F1т��+��"o�S�[`uBg4�ѳ�`�@s�xޘdg��gl���/nH���M�S���
T G�d���f=%�[����F��"�I��l{�Z�+�m�v[,qKpsGHL���F7L\z��!�WI|��J�r��<P�(h�BC8	0�Ĕ��կ.��]H��$>
�=�𘔘�vf���h���*�8'x� ���8q�j��_�R'a-�-�>�Vv�IdP57}$�yV4�c3Z.�U��P�c1i�q�tmU��a�>x�)'��V.?���g��<[|OS�ݰ�p(�<Z�ؾ���A���gb�h�Z����h)���T?�`�UZ��>ov?�ڃ�1���Y�{����B-����H�t\�\.���C��\��lg����;��3E�� ̽k��к��3���@�y�r�/�GT˗�kD������)vz(Y��c`���`"ψ�!��9D6��+����܆�*����=3;� ���j�wi���Hۖ"p��r��#�M�pc�`���ؼK7�H�v�����t����]O��	�Uf<�G�5�3X2y�0n(@ �7z>Ф.�1#ʹ�1�B����Q�ǁ���$��Ujs�L/�oϜ
����@��U�H'TCd;�T}�@��&dd���pF���&4d��)�D���;'�s����e0�^	
p�N��݉glx8&����H/�����a�.&|[GA���H�V�,��5,�A>d���o��hi�Z�P���m`!c�Ad�E�yT���h6=w�WW�����uƬѼA���.h�=�x�����BK�S@�o7����E�8�$4��Pq�F{��G���ح���1|E�61k���E<dc�s�2�\k���{*�zT;��;���qw]|���M7+'A�9�����x����[�ŝ��W4�h�|
��[w��%I���N�bz�b��wl[C��g�Z�F��1Mر���OgJ`�D ��Q;����Z����(�jR�N�'5��&���Bǂ�YL��w�~�b�6$�1g�v�%m�-�x�p��D��Sc�x�E�&ǃ�F����sQtl�r�f�A���cX"�7���0Y��~=;MS�����שo)l��&�t�F�,wc��ap|K,�J� �5C�V>�IRȤjY���g!`�0��Q�S�ēE�c���}���	��*+�פq�%����7O��5���*O���k&������k����Jt}۰�O����s1���oi^O�e��Ϟ-�#
�y�.��}L��	��I5$�B�&��7��kL�!Pm�U�ơ�Jwh%�g�p#���<=>$������r��bn�P�Ԙu��ځl�����$��c��y��#���xS�jƫs�h�k��a���=�g���b(=�_d��9����M9e~��(3f4_~$�'<�/��uIOo��s��P῿v�@�j$4���X��f�p��#X���Z�k���q�Z���r�.>��ymlP�De�P����Ѕ���&�1�=��긮���45+H�`}Aov"��D�!�@׳�ҫ�#��\<X�%:� �>��y_9�S[��vAm�߶q� �L�������C·~��6�A\4j;ƍkfܺ�A�T	ʜ�+e��Bw	12��V�V0ꑄ8L�w�����^�c$�w���S}r^�\�ƾi�G����4� F�)���J:���H<		�d� �O�%	���dr��ǿ����  *pf�5�kQ l�k1�k0�&S=�tp�9q�b̳�t5�U'*!���!*����b�n���ߐm[��ᭊ�
%23��� ����g�����`0bEl�0E�*?��O$\(ငs�p�5�!'ј��#|A&2x��뇧X�%VM#<�ƱSwP�>
l�(�L�'��c�X�)�g��������� ���6�N��C��C�����}T�f��� ��Y$V��:�{�ț���k��>�s~~N�m(�4�\�]�����2Wb����;��У�R�s���E)sJ"��B;p�r�n�nXd!~<۸��!���[+Q@*�>'��#u��S7}%^��k~��j��ǳ��+���'�	�w%�=)���à�0dd(����c<��
l�s����k�����p���lHz��q�����
(���#.�o��wҡ�lwۭ�o��E��L�vp;qrj�h�m@Ψ�Y��W^5��/aE*�yx�?~�)���M�&�D8?;g%	�*YW���U�~�5�%&B7p��r������=W
ptX(��$`�!d���~�'���T`A�xvp���r�2�S�e?l�|g��(H!aG��@�����p�?ǰ٧��wʎ��o����&d��)��	�5f ��3�a}�4,� �DER|��ڈYGxQ̍��Qiw	rF'�>;잞=f���z.�>��*�����+�5�1ȁ6A�z��ɺ:�'�f 
l����FJ�`�|ϗ�1�w�1�	C������b@N��ɱ�����\���D�{N�2�,9 ��3U����V��.Q�5o��NN��'�2���ўEqRC���y<РGg'�=�<{�g�|6��34E������"�A�V̈�9����c߮�+��;(��w(�b��pmLCFaceN�AF!��d+C���@��?b1���o�W�D:�t@R�)��;��Ӊ�������䇄�]c,!	[ɕ����Ȳ�������G(١��C=�"��l^�'g�@� ��>��[>�� ��}R�޾qk�M�$Q�n�<u��gV��$*��{�M%��D263ËB�0m��;**��N%��Z�ܫՔ�PLPٙ���b�5wc/�ƭQ:�����Y�9�����Ų�"��ۂw�閌�_���Q��IV\P!����X>��԰��!;R6��C�x��P-�G!s�a��8<&EJF��y��V����A�]�� 9�@�}Y0K٩���h"�!�L\W���6��-�h��F�i$�<��Ew��ȽE�ę��X�r~'G����M�ʦm���v=���6%�NŘƊz�C�CFy?�i�5+���84x|A=Mxe��Oݓ�S*�#�I���D��:o�W�=w���{yy���P����9��zLSxN��gܠ)�Z����Q��<�LÚ�U��@վ�<%�)�����7���4V��>}���o�?��'�5�;�6pm,X�;i����팻.��f6��5�b�
����k���k��4ݶ�re�T7��(�`8�q�}�yP�n�p@H�v2ə#˜IKғvD�V�kO2R5=.�oC}� 2�-[�$�#TO���b4�	��o]�!OqDʧT)�M�B����,�	+�啦�I�Ǫ��7WaA)��RLu���)�"���3��R1��&�,l�������J;�p�a2��m��ޛ߶k$���"���p��>5%�d�iddP߿�Pm*x�2hU ���F�;�X=��YΗ	��V�h��� \@� 	�à��<�MV�G�.�v�	�c�3*�Bi���xϊ�Ōy��f��!?$;4r[��&��uL�G�C+�n��
Ԑ�
Q��00-c��:5:��%ｧW�N�Ǡ��,�
�䪹Pm�,$�F|TA1.��:~�/�R����
׳�V�R;4'��X�S�/z�VG/^����NO����Z�~A�VV��X �M�>x�=:�q�������g�tD����a�u�&t�SO�a^�e�� 5����d C����RO�К�����lϋ}�!�b�k��^���ZY�Y�h����94�;��[�c�|U�Y�Pl� h�"�������$nEnӫk�o�uԳm5����k3�$��]��3m�Y���M� +M�J_�V�P%G
|F(���z�X~���q�φ�_���3��#q��s�$O�TV�r�S���ᤐ+��8 �݊ Uc�8�	$��kǕ���(�?�FN
7�2��m3Y�����cVm:w�9T��]Tqǣ��*� >2O�һ�`��U9: Vrp��kG9A�]���F�\9���dҶ�ވg�m���O�]A��'�w�Oܑ��:j@�0�)J#�r�>�y�SM���^j�>�
[��5:��S��,bfhfƽs����*`	զb��ޱ,x�n�Yb��hyE�%w�d�������'�<86L�R��,dTIs��)LdS*&����"I��R�cP?A���^��mо��@J�3#s� O�g��bˆÄF2���Z�G����Y���0H8K̟x�E�zom^
J�~D�ƾ"JRR�0���Gޤ�Mo)ϧ���3�������K��A+�RbOg}�lM�(�<���#7�
�E�p߀�k��
�n0��f.�r�+/L�b���R�P��}1$TEi4S1n���KdN�BK2M�c�����g���l7K�2��J-�ҕ��-��!!	��u��:��g��Vs��x��!���C����A�6H�I�"r� 2�5�٪�&�U��u�&^��������*jF��xR� 7����H��u�Z�
!�m�=j�� �t���=�^J��1��a @5s)u�b��B#�2 1ޏi��*]%�4њ���0�)�4�ct�m�c�'�mtl�c۶m۶m�v:��������Y�V��W��n}rX�=u�Z$�΁��-�s=c7��"}(D���'�Ή����M�z�!�y������'[i殻{i���{B0^l׈r�&�F�6��\S�Nh�T)j�F�`�(-���ʉ��� |w�Y�X6�r������c:y�uI$��1mF����y'R�e*��l��A���T��Jf!���
�>vw%Փ�� �Jw��gbFX��Kt�.i�0���2H`���2N>�z��dWq� �D�U�-�*�A͕���ç�`�8�Kڟh����6x#(�e��ty��_ڰݞwR	��}!f)�C$ĳP󗵾_V��x��PrZ�7Zp�б9������n��M|����u6�`�`�!�����ɇ/獢��WE�����<���m���Po���7�cuj���Le`�D������-���dV�d�'���tzΑiZG��`���>[�7�Io��5��c^��/���B�f,Z4,���o,�.,�C�7��`�n��aI�g���1є�jG�d��O��C��5P�"kJ�1����9��@�Z�����@��w��h����C��#��6?B��p�
�5C��}\Ļi ��:�# ���h-z҅'�Sn����28�;���	�k��~h���� �N�<�KY�r��}V;-EO�N@�؈BtsͲx��r���M��2�;g=>b4�FL|�z�_���5��� �^���x#��3b�#4|01#��;7w����m*W߉���U�Zb:�P�NJ���X���O�^Pi{RB�W^`")����3�|�vQ��y�/Hj���K��+��-�E��)x074�
�;�mbX�G���1�x�%	��4����r/�}:�����V<�/�ll�a��R*�Qr��WH�i���E�(&�0�������7�ӄ�Q�u�v�q8;��X������2���Y�㑣z�||��5��u\�#'���|^����<Q\���N+��F�l�m\�{���X��)h�(񖏏M���Fn�����Se�&���(����M��I=d�Dxy�	�@޿]5w��ڐi�U<';	`�<G*@m}<��)1��\��gD���GǛ�vr'7ڭ��ʤ�����G��v+m�zī=x�1u:����,I�#L��b2�C�Ea��EgӑuU�y��*'�H5�aL�3�6�u�;��{^����"o�Rw2u�����H��.ĸ�ѹ���B:���C��S���X�0� S���h��o�� ��nd�� �&4��"�spB��W<m �W���?���"�������s�<H:�\c0������)x.����a�[�jv�J7<�e������b�vť�E�t��U궥��u-=-j����~O�]L| @��鷤!�
��XYp�X�����"{燴-� �!����Z�"��IAYW.�O�n������]���}���4���M�>�t�~͑$#���bg�$�F������!V���~d�s$��3�.��8h�;X,n�'��w!炕O%��ZHK��G��&�4¼~f��`�}?խ�c��*_����V��y6���-S�Nť_��e�]%�M_ԃ�4�Y�*e��|�Y���g��{���0q�Kˍ����3O�~{0sz��%�������M�5x2f����s���Ef ���b�l5l��������k$��tg�&1(_�J�?F�t����'Ý��V�/w��e�>�h�_����PD7�A27}X(�����jhPU���!�O9P�Z��*sD�r\[��NfR��2O��G-�}���aw/��I�A�Bp��
'���)�xMѯ��������z��&Y��$�nN�ļ|4@�G'��CAB���o"�Z�
�nL���}��E^�$�v�|�l���6�����ÜTǜ�ţ��!״�]=�>W��I�m������j88BG���o�x��[�L�-6�Z8�1���tb=R2x��/Sn/D�7\�|ŭ;c�A
�9\9�*��<���$'`�*��$��E��m�M@|o�lݽ/������9$y#9�ڪ���#x�rZ��:Uu� ��]�۝������D/�����8����L�qF=m@�A���2)ј��Du/n���L�zq�k���&)�l�H�#���b�t���ֳ��"�e��j���u�fe9��5�-v���o����f�b�1��X�j�>�Te��1}Ϫ)�T��K��A�&�]ļRD�SE�����O�l�\Έ|�Ouoq�`@�gޯ�_I�#l�4Z�W�%�O4P�Y�����OOM��nD�D''&'���/s�J����eq�Le�ڝe(�T�v*U{D&hm�=*��Br���85�1��B۲����@�n�����x%Uz�q��G�Ke=x�*��LYLV|)���W%���Fl^14�1Z+� G�� �u���H"���a��Z��(}c�o����#�I�S7ȓ�(��q�ܹ��Fz�x��>�P;d�gm��t�M5�q�@Ցv�ܓ+�!�]HF����v��P#|�]&��D$Vw0iUT��P��6���Є�@��)<0Q|BZ���y��*��PQ�"�9���c�������em������%��'!Cأ-c�8B�`L{'�v��"'�1+�/����`�k�(1)z !9��F�q�R��l�;RKA�7J�6оjc[#a>>^�h��b���j$���~���<}�Eu���+��1�TRA�y��V��r,&�g2-U��],N���j��K���g:�q�;��Ȫ�����Lx6"�G�T��ԛ���%� ������Jwh"leeR~�sg��tm�5h�Y�k��#a��_|��H(�P�ʏ�j�@kXܹ���
s('��~@A�K����V��V����^�����XIH����IR^8�{���k(��a����@ͺ8$t����q)�{�l�b'������yԐq�&�G��.�A�F7�!��C���,�l�":��BR�5�Qx�|q��`�1�0����+�jA	1�#O�s���G�����;����#�d:gX���J� F�}���1)�眊�?n��*����UxM#�ۢ���ፑ ����e�%@�//Jn.���]���I�?�����MW�@!`?��%qQ�����]|:[����}�}�a�3�v������m����XW �OAr19B��#o��a��9�u�G�:;J�j�ي�����!V�S�Cc�*��W�)�X�zf���0�Ub��t�uۮ�.#�̐|��Ky�+�˨gI�'Bw����&d���+�wQ��u� R.5~�6_9��Mz�{$�&�#;�Uj������J�~y�@��� ox�Q"���ۼ��@;� ,xL/#�E<Y��e�Ĉ��o�Ӷb	�R_�0��i�Г�X�%dP��k���Z��O��c�6H���׈���г�'4E��Rd&�u�8��!-���)��D��`��`ZTq>8�d��B Iy��$�Ǆ�U#���wO��!�MI��\rE<��c�� b���� ��Ȍ`?zF"��5��%ܜ��!b�N�#`_zq�DF�Y��b����0�雋��y{tO�z��lȈ�a��|��-���t�k��={�y�}�俍�6Uc�4�\^�e0K1[s��L���#
��<�	[�!S0B�2S���CZAa����'�>��m����I��I�y�'Y�E��v��v��o5P>�(6S+��\��qYZh�5�U�{�2;�ŹI���,[�*#�Y^Q�&,I���E����"���;~��������h��-��F?4Z�z57��4*�`�k�0'�	���=+^�'Ƙ(�.#�ã�#��
=��t�݁c����,�ϑ<C��K��7?�
�r�PnҼ��wZ�Q ��iӬ��w������7��pbe͸��V���T%&�0F�����8WZ�8��Z���'#b����Bq��}�2WEp��݀�{�B�Q�x%_�p��P;�In6l)���Ҙ�i~HwS"Qm�_�ge�x�q�O0�5�T�M�@�3e89�8e�����?�Y5V�����0�'���	�����!;���:������@�����*��#n��R���>`
2x��	��E�S_��l�"̚c�' �oW<I��C� ɀ��t}PH�X,α��Q�Q���lMa"�!�l9>O`�p��F����v���D|# �������K1�z��tܽ^e� j$�Mv$%Q�7"�Z���P���+ .>�R�o�V�4މ~A3Z�x����vJ+D�Լ�����
�!���AQ&�]�`^���@�7���z�a�O}#��-4��>�k6v!(���Ч�R;y`�-Lt��m�_P���䰗�?L�@��U��v���X��)d�p�\���ӄJΉ4{n���J%��U��t77+,oPɶ>WrG2.J���l��$[;��W���U���=q�R��_��Aoȩ)�r��~��{�l�{�Xc�c�IS���!�� �5ґ�~bz�q� �����cDƁ�,`��{�
�@����U�0]u>Z���N��B?���,|Y���W�|[��k4> ���̘4�/��G\�<`Z�9P(�<��V����E����ϓ���U��&# ���ZLAw/D��Eض�G�B˧F,�|C����"��;šR�i��e*�(�"G�=����o��
I2�k ݎ'Y���aLm�����.@/묩�5�V��SXh:�����&�&Zê�*�X�����b�(X�W�$e;�����U�\��dEI$(ߌ�����q*J�R�I���/�Z���۠�Rk����mЩ��d�T��۔NC!,8fQ��/0��kJBh��"����z���fi���'�[,�^�?-ީG{�*��<ҷq��G�����2T�9¨�X���4�*��T9��x֡�fY3x���� 5����e�Xɫ��8������v�U�Br��PD�~	>κ�k�����/yjv\�����9����z��b����r�|�������6v��GڌFY��hdT*?�*�(�XX���+�;��;��&��Br%���l�l��JO����� F����X��R§�A»�����8������x�Lw����;�4X�Ҟ9��\B�w%n?�AE-T�^G�?���h;�nA
��_�.��F��,IrfY��؅e:l������������T ����mĸ�pxnu���ߺh�Z���Ǫ��ǫ�v�xs��UËM����3��7%�
��
�P�����!�6ȔR�c���%�.å��^�i��
�T��0A��m%�*d�|f�0�^��D�7�d&{Je�Rv�W��� �X���]ү��+��kΉ>X���ս�?�/K����'��Y#�5�B֐���ks�l����}�s��gw��9�v�e�)H�f!��Y�T�D�E�Pa2�ƫf�뱜�t���;}���Z$�q����3}�iw�(C�2]��<+?�'�;���h�cT0���l��A��IK���/���D�]�pFI�y7��i��ܸ��H;��D�(!��)���ё�!�����:�Ĥ��EY,�M
n]N��q8#�3_*��%2zPH��.�lb�N^0P���@�Q"�T]�N3��+j�G�����t�p��&����e�&�ٞ.�)�wZΌ��M�LC�h��a�7��>W����h�C;�C6B\+���MpG�.5�v���SЋ���n��V�n�GE�.�rl"Wb�|�����&?9צ�.0g	4�&�q��������i|�!�dY�b��4;�	�n�x�(Ŧw�����b��f^�yy��}�d����6�,�RJ�O����R��|%9y⥵ZOs.�D�X��`POH�W.�x
I��N6�6�+\f�	6ot�jY�����!��Ӹ��tX@;��W;K�¥�Y{��Y9h�k�[�u��j۴��a[VW�m���n�x��D'q7�)_���ǋ�]��bp|���=ޑ�^�hve��#���Bh�O���W	�1�}��|0��"�/�9}L���z�.�E��N���4"N2ľ���QT�<t��{���l*��K@��1�-(���i2���o��x��<;���Pߑ�a�'�)ޤ�t����T��Ԙ��_�=���a�QL���8����f�BB(�ݕ�P�Z�v���#�	q��{��-B	�5Wg��ĳX��c�beR�h	�]�\�t˩�����5!%�7�V*4t��&�� ��&�p���<ZwRo_�r{�]aM:9�i�0�j+��q�k '�-3B�/{��5g��(U�y	�؂�?�bA�zߛP0��6�QE����[��g*'d�D1�~6iN�W�@Kej�J��,��H���P0G-���,����U������6Ht |�AnaX�HTf���@��?WOZ� ���]߷͟G��[18�W��G>$P���|J������*nt`�opv�W�6�e�9U��SJ�W	�xĬ�Vs�Z���ri��e4��զ�9[
��b)会�����+Җ�ӿT"f�~�fKl�͌A�g�R	��J��H�d��՛Lr��n�=��(�G�8����+7���f��a��A�`Yk�-� _��R������~蠴��1���0�11�2�]c-�q�o�ȫ��g\2��j]�����d��7q�$Г~���]_� ��Hs���/a��̾nu�2H���:�[z�bU�rne��
6��`��I���/bU3�R�������;�#���l�i�G�&���b�
o�i�i�� HQ9O���b���$Y��{9�td|� BH]�u��V*��J�4F]匧zE�%5崛=,Ⱦ�a�$�����G�*[n���f�~L9��&����m���F�H���v�}�xr��AΤr�_�`���b�����]���g��&7�k|��b���2�j>�cpFj���.F�N���7�*�dzSݮ3��WX�	^� ����j|�h��$�W���l^���|v��;�[���(.�[�I@��S&U�D�.�ai�C��3�CY����y�%� �y��eM��E��Uu�~�;ب9LWe���M�3�; �S���mY�������s|��]m�RM�<]DZH-R"}�rP�l1�͉�` ��
��{�ciE���P�����wq�η����~�F�G�$qTԾ��[�2˳Ɛԩ19���=�++-��̳Ty�lo���
�!S榵-��I�F�<� [���%f��"R;�rXQS��M��$���^4�$:�>pE`&�%�����N��4�l�.-�[&�7Zf���'�b�%���D]�X��s�aPٳ�����b�@XaTk�>Є��l�� 1&�bZ]��7Vܨ(�7;b4O}?}U��]WH.M�>���`̿8)��!x�� #�9���i�i87��o�\R��&��
�p9o�����[{�����';������VM�g�ȕ�@ֻ��C�1 �T,5�����rϐ�F�(�u�V8aN�T=����d�������H�L.[�j���k������3W�~�7ic���} Y���D��"�@��/��j�6���|��$qma�
3�YIMB�
�F��ԨX��d�7Qq-mt������5��b��r

�Ds�oI�]���-f���Ӄ;tJ�E9D�����\����,ǷV��1�Z�5��ꡂBNe�ㅈ�UH"��;f5���<���~�=�ƌ<��^6m���Ϛ�v�4iHOJ�|���%x����:T�^m�j��M�8�Wޖ0��e�Wh�UP俰ίb�ێ���.x�P��W�jA��x #*�3���C�+��+�(�^�]�~�A?Wo�A���NU�t�sy,��u1f|��䷾�Q���!b%̶Cp@1�Ə�N���4��p�!�̽��u�#�S;1ʭ���J�F�Y�����[������5Gф��lج��K[��6��J�����b���G-�m[^nt �7�����w�g�q߷��?Oޞi��Si��qe�Hv��椕F�;�kaԄf*i�k�wՀ�A=N��f#�40�E쑊��`�¦�La����F.���8���(��NPT�	�"P����X��i�P�>V�x���a�HH�y���M��;*�-�&��>�?@̭(h�ᗰTx^���.�tϡ��Q�!�����":�X4V��ͪ3M���L���.+Cgn��4L�	0qR��,*X���ieҢ]�'�� ��r�e�A����`�c�\f��yk6T���]�;��<�>e�K�v��I����=�=GT���'=1�M�ab����h���O3�'��+�En���xgr���:��������SD��P�����籸�4P7���X�]Z'�E(���R����Y���:b�k�x�I퓠A���%P����z�˨4eL��	�o}���<D0�iT�vcg��q�dڻ���ғs7�&�7qrE ib
R5�)������1s�;B�K�?��ɷ'4 Y��� ��_t4�ڇ�p<�q,����z6[�j�M/����ʕv8��mAuHXZ�Y�a�9�qw�:��;��-A܈|?��=\l�㕍<fަ��Y�g��{^�!����J-�Us'��%-3�T��1���d�(�>��J�J	Z ��p��0��6v��V3����C�@�S5�JZu�Q�0m�_��U�����9L�#�J Nȍ1&Vi����i�I2fŅ#�[w)&���b�<��5ssca�7�R14 s�/E��A��w^D󺧌����:={j�J���3���� ����izq"��L-��3]���=�P#�.L|��׆w�����:e+�^�U�9
 ��'���5��a�������ŪSv9�ѡ���b�H-΢I�f!�����^��d�Lz`Cs�Ą�hg:6=��X+���D��<Y�f�&I�t@,��⠄��\cJF���I���#���A�V�)��<))��,E3��Q+�c�͋G(d|�z
>f�H��Qָ�-?u��/!D� ��.v�Ř���ԅ�&;В�%b(�)(�=�N����V��rRBIV�q5UD��R�L�0�e���V�
ycy�hV>c'���B�;���ո��jt@[p���
ue�g~���{?��LOm5���t7��=
Ԉ*�6����4�o䁰������uq*��N���7]�c5S��#�׊�}ӯ�k��%h�����c�����k����� ;�9������!�wr֞?,�]��c�%��m0*Jn����+E�-%g0sp��-���s���m�6�����˘*���A�8�S�A�n��� -����pL���^��C^�`W:����	U`f(�h��O4Y���N�t�����L�4(�(V���8|��3?��u��>6�N2e<�d�M8ҝ��1�81D��m�aBvlWM�.O�����ȑ0�"=���M"Y���T��p��J�T��2 �������*nV�}z\�8E��OI�L!�1�g��V�)F�E�j�& ��ԣ9=�l�;�4�\#!�R�5��,����v�oC>�Yd5l�UQ�H�ٜ8Lo���8��Mh5 �����5�
����3��8ր�I�.�.�����p�~۫Q��=<��E�	���=ng8������a��S빍\�DY����?lߎ�{���Ld�:�
=ј�G�,�U��;����RJ�$���~���;M �,;w|;{��%i�3Q�F�}� ��k��!�{��+��a�����j�od�������0�g����ȅ����.:�������V�a�T�([|q����a����v�A=|��^&l�e���i����������cǯ���/~�L�� ;fcp)�x6�X�n�hW7ԵZ�'f�J�$�C���c:�(W*|��i� F���Ya�&�S�J8_�OY�\?��Dd�����Q��^��w��ܙ�K_W:�����8���[�'h;,,M��&X��a�ݜb�������{��rj�v\h��[�l�4�W��hD_��!�N�}B���Ƣ���}]�ɧF�*?���V@�ʿ��-��dѹy¼���~A�����tr0�x˂Y��R�-��Fj�I���u� \���jAc�˾��g��;�ױV_���M�(�	U%��-��4�@�)J7;�����vdz�^����%�~����r�F�q}��pԇ��1Ch�kOԚ���6X+�J�#���k��Τ�~͸I��D�j>?��}W���>s��C�<�7*�����շF����x`��n[��c����z���l34'}s�R�]��=��eN�%q��	6N<���YȬ��n���e����>`�dՆ�}j�A��U�|f��4\TΘ�6 ����ϝ7�G]y2�_iw8p"n��U}��+���7̇��oZ��ēRȄ�]����귭&35~��=��|���_}/c��8_3�b��Y�>[��C��t�5�����ٱ�r���Xo�K~�������������������D؏��-X<�I��y�@*�mŔ����3X��rn���Ա)���uxh�������'S;��ň*�]R�=�%dBw��N#�J��ty[U�䯉�����2��d�'�����<�ڷ`T��*��a!��xu(걑zr�+@�d9rK��$?8��&�+�]��w����}v�B1±���'���ߕUW�W��Fb*ɽ��c�:1�$�e{,�~�#$�����c>.��Q� `����Q=#��:ִ�xC�����g�D�#'��t��֘j�΂F�/�����\��qi���Rr;ɀ�{�l
��b�5�����s!�!nbǊj<~��쫲m�x฿���x��a�n��3����*� +TY薑>�[�z��17����-P��QA�$�H�K9 M4��w��om��khJD�D�����u<Fr<�?Dq��p�ߓ�R�P�C����3��!�H/����&*+��e�QY��O�q��N.w�J.����
��ǎF� BB
���Y�{e40��	�qdNc%��3j��.��Ook2k$�c��Q��7�b��hL�߱�Q��9�?�h����ǈ�dƿ3�b{�s����ο>mxgdw1��"�{'��cP�;s-FQ#E���P��Ȳ|��u���];s��P((q��`�2��a�O� �F.�U���f��tܸ)��g��uR��a�"�T�)�HW�o�M�,�mg������t��kP���E�8�����@�Hy8�n<�#6����+|�v��	���o*�����`z�!��+N����������Ԁ�����D�Y�,p�n��vᵡ�������87���t��c�H��e_}�G���+i��0Cp�u���f�]�ң��X��j]�ĺ���?"ۃC'�����E��E��������}d@�gW���Vr�>D9�'�}���3�Q���g��z� �8q�?]��T�:����i�H��bc�dU|�s>�EY�����N�a�����f	�*�uAb+>7��S0��TW�Ji
��y��PQ��G.���hwl.�b)��q���#�V�%X@�=ڵY�V��(J�	t�R�i�y٨��Q��#�<@�4��*C�; =�C��V_A*d�B����,�����6�Ō�.��~y�5�/`Ѹe[�`��Z���"a�&&��w��;mW�a ��SQj~��T�c��AV�%�z��&D��!�p�J��ʂ@�����F<(2��~=4HBR<8���ؚ�JN�0Ƥ��7��Agd��j�SP( ��J�#��\M
]-�9�nk��Lnڹ	�'v�cCz���J�pH� �h{K�*V��OȖ��z�ݪ��Jp�}��kO�����J9NH�\��_�iO�^��I^��P�h'7��x�4Z��X�q'i�G0��fSF�ޱj{�"�C��0a�R�����~�?+)���L���]R,um�[���0�|T��=����[��V+���1�AZ�;z���Q�U\�ukk��0ij<.�ǠD��G�Tt.[�\�� 2��Dc���Ѹ�j���h�y���t����#S�l�t�76>������6=~w'��vrl��n�Lu�[����^s���Q(���
[9?v�O�k�#dTf+^���``�/��w��|�>h�O��O9˂i-c��L��ȘyB�{c�=�oq3�`�e���@�W�-��H�?�u�A�����'	�m�Ҏ3�	{7�"�� +,ZJ.��Gf�[&�A����T_�$b�v� �|	 �c��jit��_���!K3d#�],Vh6G�v�0���{����x��⸲��(�W
k����^�w/*�'�|�=rI�Їd��(�aY�����~�o�S=ϐI�V9�@ݢ�u�؎@ͭ���o|���|���l���q?G��O蚤o�˲k�R�9U�R����������d6y6m���gŋ�Fb
-��v�$5���J؟�"3���8����K�0���`F��J��R��@�3Z\���%<|�� �́_BaB�漬�;�A=P"yx �d#�>�?�?��N��>���=��hB�&��|����TZdL�JL����Gp�{:�1� ���6U�!"�;R��f�åxa�e�J<)�� 0�,fF�=���xG�kN���'5?�BYy����[[f��~�{a�#!7����������%v����A]�N�1.F�="���#�����ы��$���
�1�˩��(�q��q�l�t=�Z���I5��9EuH��}��}�no���Y�Ì��g`����=���UD�L1�fl�<k^�f�t��e̛�Ⱦ�����q�����ma��B��w3(s����'-�:��A�5T���8L�恌�l}
�R=/�7�eh���,�����<�ˇ�.�=�u�F���W=��j�V��3�u��Z3�|��n]#o���_�h�C*�o81آ:��a.N6_����=��sO0
f�o�e\�jd�W��QR�q�a��D5��b���N`�KZ9�lפ���|3�)#2-�=H�-�V�^�3I��w3��R�Eq�����V��]ԨZ_FQ�+WrC��Q���?��G�Z-$T������}�L� �b�/��.AR��m������o��=��{ ���vs�س�$'ԇ�ҁ��x���~�"�	�IE�0Č�e�c>���2j�wC��cm.
�f�	/�g�x�g���s���7�G��M6пw�Ax�����ST��?�.۬�kJ4H�$��ȸt
o___At�\6q#��T۶�l~��`�����I]�3~��+_��S����ȭ��Ն�A|I?�Ӆ�5�v��O����G�C>2�;_���}�]������z�-P���7Q?�{%	�:F� ��1�f���a�/P�%��=U��z�ŵ|���W)����7�o'�#�.�UB�5�'4Rc����ט�3����0n^H�k(x������&�]3�̜ӝ>���<�`Wj99Z�=���lr�ޓ��3�{���/��c?x�3zO[��������"�_f姅s�F=�ăA�zσW�̽���@�OJ4a�n����T�~zz
�J�M�1��\	��g��\dD�a�ڡ=�)Å�Uq����y2p��������7�߂�H�<���7���y�϶�^�Wӗ��C��
���0�U	�CaA/�fBE�6�>bB ���(���1E����$B�s��w�l���-��}�iz��\s�,�SV�X}U]t�,�,��Y]5��E�9����v�ϐ�f%�����V���Dr����~�vL������J;=Z[�����j�P(�D禍���;��=��tXX�b�+�m��f�N5p��?�갡ͪw</��~	9c���ɡ T�N�9��"��`y�������r�}7JU�����D=ح���|j�mW� �-���ui����'��@K&������{Fu��#?a�������v�����gGV�j��\��VN:�����M���CQ�`ۺ�5DVX�I^�ԕ 'gl�T�Vk� �JM�7V����WO�z�oA�s�hQ^�M�UP���!|�E��j���4ￏ(3A�lB����Ũm�%���o����w�4bh����Էұno���N�&nTpD�Ɓ��O��A����ҋx�	<ad�4c��|�����PH�3��t�/(�o�&F�>��umL,Uʲh����؅��� �͔gw	n��j���3��W	'�ͣ	��xE������^�!H��h��_o���kn��z�]a�.��P$yT�"�f�Ig����� ���l}�T�1�Uut�f��15�26ʇ�������(��)U���XLk�_w�g��S�y
�967��m}Ё^�ok`�Qi�(�l)K���]]]�DE���`�0�Jl�J��U�A�im�ଆ-V�K�5׽ٴ����D�mKo�^��Rl�Gh����� J��XM;v�E�Y�&^�(t�����@C�s�6���(�������d��(]`��T2n�K;�pb����rD�6�M�V���5�m��'�TA�-���Ҥ;�d[��i)i�낽�Z{{�	��E夣nS����>L�o{LH�c�`��~�.b���8���Y�\��n��n�0!rj�L��!����G�<-l�f�2�X�%��h'����o�����k�"(�8����j�SH��XmZ��c)���{(����D澄���S	Q�r�S��ݦU���zI����dS�h.��f6z��t0�o�C����6�+n����H4�x��c��!q4A�e��"�@�擓3XFJ��	�qC+N�E�\�fE����͕��7/=	��U��$M�/�:�vu"a��Na)��=t�M��I��� ]4��b�? 	v�0�%uu�q������tk3�"�	7F].x��}���.����?\
�$���j��D�+��}���p[C"���^6ONZuɝf�p�$�Ռ�
�w02u�A7�T�X욞�B�����W��T"��r�14��71�ǖ���XQ��pk�iC��B=��M�=�!P�.��-A
��OJ����m�F��ȚX���%^�i�ʩq�'�~�enrc�嶒v��(8�@��\����2�M������5t��S]K�t�g��ؕ�c�hMb���ԏ#�;���kR���"��S����U�a�?���W7j��#8�dY������'ŷ$�1���y�-�ʽ^��l��*Y��^|)���8�=�D!xv��q���p�p_^����O'��ͷ��YI�ʶ�U._g��Y
��lgt	k֨�X>-^�k����'��E�笑E���?��5��
Wh�K�l�Ң��C�j
���$����J�b>>�DPY��.�ǆ@�r�Ǹz8ʹ���r�ЀCH�0��@��udg'�ߗr嶅aw0�۹����U��N}n=Zx�D"�`���"�b�>|ܯ��)j�[ɤ5�yx�L�z|���|OC��_�O�y<�����5��2Lכ�.ţ�r����tG��2��
�8�P�k$$٥	��5C>ep���ӭ7���[���o�;a|�s�WRt��v��}�0����ʩ�������;���a �\qd�[t��F����7����tU�,_RNW~��p��P���lU��ѨBY�|U�5�_��R��TP�����d����d��o�����x���촶�mΩ�i=02�icQ�J4���;Yr���jE��ow����U��1�=:�f��#e�.�u��X���:1�YƩ��L�rݟo�s�Y%��] ��$�y�����s�;ۭ<�J�7V���ݔ���i�s8�X�K�V��n)�6u2��W�E: �7�Vyy�E�!�HJ���>mZ �,�2	�Y��Y��J��܁��7,Ld�s���� �E�6�˟��2LX^R����ժM�z)<���tÎE%P5��Ā����s�]��300�2<�$�{�tX7�TR�d���>Fk<fr����_���k�V��F�C��Sg��3��q���:�4�Q��`v�riB�K1��j�%�s�/C����4����b��$%Ͱ�Kr��=���������������|ߟ��v� ��PEW�aJ��xs�B#��s���� �ED;���r���WH5��yo8Z⡫S�We�/�p�m�l�eQȜ;?�	���mǀ{G����?�\����l]�y4�kʋF�j�~O|��mV<р�mO�Lِ�d-?�uy�o�1mEʑ��f�E����Ӎ��{ �
Be�{�k@�M��4��k��O����o7�~�N��ŭ"ۖJ�F��o%[��6�a軸��z�bSOtr�\�r�����F-3����XìԻ�=�������ɐ������̨�Xizȯ���N��b״[�4*�Ս8�[ȓ�ٻ{��{h-)ܓ5�q0x�9�f����:�37�y��3ﭚ���ZPM��i�5���a0[�:9�!��IU�5ə�I�^���c�Lx�$5a�m����{���\�ܵ�B�����!8��r	��ۗ`��#���!�Ꞥj`B�&	�	oU5P�����G�H��`�iL]�a�,���s���d�,RT��s�W-kn���5X��`��,�YX`oH��[i��%����-FԠ4�a�PZqH�Y�����Z5]*맱_9G`^��h��jV��e7���"%�!�N���e$��d��ܫ٬k�SP��3X�vC���O��*>��5��)$X�M�9���=�9{�۫"N�_zd�G��,��	uRL�ꁸ@�Tb%�r��4I=�ˉ>渪߈�p5���*K��������M�U)r���~����6��=��T$�#~1���z�J�=�����:)G�Zr�6e���=������8v?�"n�`uT`	uT�Wz���B�HB���ڔcb5V\A&���5)/�?H��ˉ2Ϥ��N�Ey�
�Q��l�H_Ҧ&b�0W(��$��¯�a��w���h$ش^Y׋?���>���>i�}�֥��d.�')>�X����l���_-s�'�䅍s����.
H�<x�D��|�����=d�����Xl^�2i�H��e���֞�w��ܩ�Wg����cEC�J���O�J9�C���|m����\����dr:`�T���2�m�G�ȁ��<�(;���B?����j�l@\:OqgN��֐G`|������SI��')���V�n/y_����kDs�
܇�f'Q��Z�"NV��AW�����M�C�K9$��R�w3�"c�Krp,Y�gDφu�e*��n��XqF��3]��q�a?��Um�5�ˮ��w���v��k.�� G(���	��z� u�nƗ�,qە:g�'wU'�}��z�������.AA-�0c�o)qn��_'ԅn��F22�'I��|��<�%��d[|	7v3K��ߙ��x�
���{qyd���-��Q1����K�T����!c���o��Q�?�aD�v��[eJw��d��3���������\㒁�0�p��t�G���=��։fѿ$�Xހ�ߟ.x�[(6��ݺgϋCaO��0��~��n'N@緶h��[!(�k�,��i�͎�kG����tO�{���>�F,~}B'/���
Z�z��Lw�*�������±�Ʊ'��b�U9����\��>�Ǽ �$�!}�m�Je+�c�^�#�l���ZNxWs-`V5��r����2y�����K�3 X��V~8���GDݟ���p8���կ[�[�� ~و����nnG�D��Y��C�0��3
+��8m7��P=ҕŅ5�u�?Z�������ھ��{�ŝ��ѩЩ�d˥��<pzh��l��p�U�d:�8����h��~X��	�����&/_O}�$/��͆D���^ع쨄e�S34&�-,��?O�y_UKxy����7wr'ؼ��h��6�vSd~qz� ��;�+̊�x9֏�y"��^s���h���H"lG������i3=<�0��"�0��
����H���u�����%��۟��P"�h�Pv��>�D"&
�>
	��5[�����PK   ��Xq�q�  i�  /   images/963eb574-430e-4d09-a29d-074ae2ef552b.png4zcte]�퉝�m۶m�<�m�c��$��m�Îm�7�{Ƿ������Z���=V���$,,  @��S�^�  4���Q�u���")���; � �b�j��]P�9�n��O�F�<B ��roLit���������ANNjڏö�6qw�=37実)RѹbW�XF�!�rW�o� ��Y�E;:YͿ�3���x;ҋPE
+Ã�.1�i�uW�kTj_:h�om`�Ue�&f&�lO��>�R$WV���`���jk%����|d�`[�cnV�~yk.��R�f�\Qpx�bRj�['���OWs�$�ZN]�]U��"����S�9���D�! `뮎�蟯�"lحt��+wK��� �pX��V�ar��W�"�����|�~M����kYù ���Ϊ��+f��?SN�&ٺ%��G#��W�S���}�{q��fS�Tt�󓬄�*e��z1��?ą��k��'�.a}2��+��KW�n���#A[���._���c��(�����Μs�e��´�tI������r  ��)ո��`���vi�3\oy��v��A�4��h�'6QPG]=�#�&�@w�v6��͸�v_�lVi�~g����-."Wa�Ŷ����y�ǀi�77�ez��/A9N�r1u�P�
��r(��{��2�=m�����#�yB���A�������SQ|�U�7��o17�C���v��v���槇\_��e�J5�4)9��z�������Y%QIͭ���S�4qu����E�����}!���87��E�:p���ֿ� i��n��4�o�/W_q:<X^6�A����y�N��7����+�ܯ%2��0�j|�x-<�Olj��z��h�.�U�6_3ER�.�.�K���=4C�`��}��	"��g�Y����+Z��zn�9�	��ٞ�c�����τ�y�W�&��J������Q>l8�lŋ���5��=h��݇�JG�;s;���K���Ե��o��5s���?�W�=�s��f!qx�?ٴ�M]`��ی����>.O��՝�����׵����#
UJH�� g�H�R�I�זKKh�c�>K�p6��;���`�v����y����{|���ή�OMC~Y��k���jd��,�r|���p��G>�9����V�ʫ�����7�J��z�O33{b$Ls��U�T*K�L��N��wD��^���_GzP�v��]_�-��*5g� ����|ojl8�����O�����h��˓Gwяu�[3a�-�tf+�����uJن�	��-��)-�G+�T�T�N�I^Z�t<��mU�]	�4�n��Ǆ(��c�>�Y-��ܸ�9�o�V��s�<�:���f��7�4�3u{�yOo�^/G��ǎ;D�q��Ī��;8x�#vX�`֤�R�H�������C������O�� ���(`�мZc�×w��tE(DR^WbĲ;7r�iߙ[��v�W��?�*Hb�^,_�۪ɪ��t��5��1�B��d�G���f���%fBi�G�jaP������
����cؙB���uY��}�{p��_��9*��;�w�$T<7u�6������{�ǌ�XOC�4u�U���s������xe����5F����s�tE8���o������� T�&_�m¯���J�����%,	\������I@�a:}�׫�̩$�C]>�_��aU����� �AjG�f֓@���i�Nb�h��ϝE�+�F��tUUY��$ԟg��J�j�Y彽�����7�溤���f��q���u�E�_|��:d���ȆO%:����o���/w��o���o����~��H�3�o͕�_Ą��gPSs	M���a��g_W�N�P�B��ع����[:*�_nTl���b�����=?̴R�����"��AՇ��Wy�CsJ��?u�"׽#���ܦ
h����35wK�����Y�zQf���d��EU��ۓ;�KϷ/nՙ$;��ICíx��	q��\x^555�,��>U�OA<�����:-|�z2a�
��H�(3��dusZ����k� �H{�\�{&Ξ
��өm�ګ��.�}��<ߧ|ҝ�lx�cy����iUg� �+�C�Y#T�b�R�5ۿ�����P������l94MT!��]���Uv���L/��/.��"���b�Ʈ0��4L���!�m�|��{��]����r?���%�hWlǅ����ݣJ�S��99�Ro�ڥ�ˇ���Sю��Gӭ��#A���ה����f���o�DpX⒨��tg�f�� �*�]��Ny����r�X��}���Wm)�T>�{ta2�U;���o,oݤ���͝���TE,.'d�)�Mˡx�:�;��7'%�������G]�Ms�J��8��鬕kT�W���|12���-A��'��&3�Ͼ�^&�ݸM���#/��٥�aǖ%]Ί�L�汸@�ϸx�����GYt@�?B�\h}W�i.K�E(��q=Ц7�Wj�(�=�N�<���VF�@�j��&�dȐk��+Ѥr��<�������q=���r7,���������ܿ�}:U
����A-C�����/�E|w5�R�����[�������6�I#Q<�59=�Ň@N
ƾ�1%��ަS{M,Y��dW�������&h{>��Ͽ!XYU�N�VU�j�S����T]��P���BQ�Y̯�������&HH��چ����{�.{;i١��v,��g'�|7�{���o�?<���̸����1%""�����dJ� ��ӗu�w'���x}���&S�55�G�2���449�J���(��%����nϤ3JW��kT��j�*�����i���N���~� ���������ՓBd^۽�f
w�{���9&75
��=���A����+F��ӤFS{�=΅i)�mWU���WVF�sLٰ��4����+�r�̠M�H�׌-�+~,L���0ЅO���Jzb� D�A0?�CF�%+7���.�9UVV�tos줒pfz� �n���}U������s�?�k��k0ߋ�������۝�RW#�N TD
5�Cqz:���JWC�3m��w�����[6>���Nn��ET�b�4�y\o)����������C 6l�������._>--��((;��͉ӵ[��)4x�)A�����i"X�DyW��Z :�]8������?ZA������kS_f@�HrV�캧��^�ҡ�Cz4Q+��وB�7F�=N������}�"�j�[����]�h�7?�CzP/]��^���b{e���d3>�
��#�k����-�&�"�8ܑ��v����9fؙ��Z�.��Ӄ3Y�W�ݷ��bFJ�1��	q{�!E|���ڥ�^I�o)~3B�΋��|�M̒]Cj�T�ot1nG��N������?[�b0~�������N��/�t��Tz�[ķR�[$x'X��/��������%+���aU���9�r��� G�h�`����ͶrI]��m��Գ���eG�hGTr[Q�����lI_y>-{3��ͻ# ��-�{��n�̑K�{_o�8؄�D\v�J��[ͼuS�q��v�D��r|;[:�tiRe�L_<.�=��2�Ӿ'�Wut\4�}N��c��;�de��8�;�M��.{�|t�ݡ���T���hhhF�-�6�mO�|yV�y=����uq��s|q����T��~�k�Y�춡T	�/����R��	l޽�w���=���.T*���A���NGo|�O.N���	�
��ާ����,�<�믛���刋Lic�كBk�t=����S)h���]ww|*"���J�:����T�������PYYY�	h��H��{�WR�@������{��$FE2e�A��Ƈ���a���Y�}�KY�ݖ�a�~�;R�kqqq�E�_+�*1�B}�\�6�f�der��R>�X;��D)2�L9Ȱd/s�ty3V�0� �	/kGu�R�қ�#T�Z�0R|4Xq�b7oH^��~�ՋY�u��U�v�Ʀ��[�}Z�q����egg�C2����:�~�Dsbe+�N�)�:3�z��c.O��G��B�"�Փ�.jZ���U&yla�CЪj&Y$�C�<�֫T$S�:E;N#Y�R�M'v�d
(}��.& I���c̆���S��P���)�ܺ��K�]==�����5P��'_Β�ȓ�R�]�C]2H6�����F��I��b��C� ��`eK�(+/�L�*܄Y�.�<)��Q$Ѷd�/dU��38��/bf���s8V�>�N�6|�.T�&�"�O�������Դ�t�þܕg�����aaeE_�"�5�f�:�P�[�Zǔ��5��߯��{*��5�0����SUJ�ËS�>>����1㟗j���D�<�E�{�y)�#"���hǌ���
%�HH[���-�,��t���R^� k��K�����͕���Y0,���;\��e��O]^6���2�7���{��S���Z=�`
��F�j��Q;pB0��g̺�ɋ��5���s9�vp��naoo�v|���u��Y�|���71FLvD��i�����T�LiEGGv�r5D�4��s��^�TyF��M�x��Ac�Z�/���Kg�La��@"�g�#F��Wh?Aj�*[���s������q�����q��S����Q���u�Y�H���S4�����4���n��һ�YW�+.^�$,��*��E��<JZ�MLN���EK���,D�-��;��ח�e��>�B.XD��Jgco|���G'��T�Ԕ<��H�) ���9"��F3vIL��:�3	 r3��A#?����wڠͩgp)��gm�z����w�"jEee�ֈ�ϔ�:<!,�y�$P��y��\x<�W� C���	�5i{n�͂im?ؽ�/� ������l�o6��:�_|����G|>ϟÔڜ\�
9;d�˲���P��&
�H<P_k���&�������F��Q��3���L�g��Z�Sz_�A| �v�
4Lb�H�����	Z)1NQT󒛺�z'��]��;G��i�~>��1�z���񍖮����d'���q��fUU�T3��[Ǻ!���Ѓ�|��t�����}�'Kۘ�����Ǉ��5,dH�Y���N�8���!ZKG��L*%V��\�@���i�q�h�#��&.��wT�o� ��W�v�\r�!0��r�W{6ș�~�O^̺I�k�9oz�]�:���HΨ���������.���8
9Jf\>fJKc8�I�5#��Ê�_���.pD�FA�o�	��q�-��~7)xeg8���������s�Ζ�%8�w�qŒH;�C�!��N�Ӂ�759ym�Ԍ3��Y�W�_,%��6Us|c4+$�2�@��(�s'��~`��gd�L�
�&�'���zlU��W13!�\vV��d���E����Rvn���C�wt8iʸ�'i������3G�>�ޚ	�C3�݋�Y{�Vk��R=��ڿ���b�M2Vk�Ɵ�
�F�LLL�<Ң�.)d4�8H�E�� *:�u0x�`9#@Xv�R&[%:�ؠ:E�j�I�����5�q��xߒ<�("��s���YbĄ=�]Q+c�^��`<���排"��
8��S(G1�{�_6�ni��)X���,�J��K`v`�dvVv��֛�|���xP�!.�-9��19o�Ș����2c�яW[���yd�"SSSf-Z�UYp�Бp��0~�L���0�{"asʗ�㪢��ީ�=�M�1G}%��S;ƃkvSNy�x�祖,	�PI�cb�^B�B]����w�:��aU��E������!�����K�㠇Z>�R��}���5{Q�F�ql������ޫ4�M�(�`_!F"��ߠ������U�HoF��q�_�1�Ԣ��<�qLd����+������+����f��,(��S�jأ�u�V�O٦y�L*B�
����������+Ϡ�B"�_����I�@���0�6s1c���c0lK�B&
�(P��Ĭt��Vl�X��Ѩչ9|E�����ܭ�z��;:�ާt�*��x��D��/!!���"?�jƂ;z�����P��-=1f1��a�s�u���� ;��<����\�f(?��!_�bN�,��y�������DV��&��:]k���A�:8~��ب�#ћB8B�&�I�b�n�W�����[�kx����Y��l!��+�5k�M�֨}F���8x�sU.�d�(ny����h�>Ǣ�-B�b�av.O����^FYN�?�� d��o� L]�qvv��W[W*|Q��d)R���<.1�˲Y��$�Qsg�@Ca`�@{L�!���U9�X��"i��)�<wb��S�8?!��[^�
lHd�^�"�#w� ��=�ي�ʮkh��r�5���P�H=��S�|��e �H�^�����Y]�a_�����(�^ʻ�
p�5Y�;�Hm@�<��c?����/����9� m�6G�<#!��`Ì��'f���<,�N���@�@z9����CF�t����K�8Ux�I��x����R4��Rf�Yt,?*��H��-d�*"�_ߤ��'Ӧ}��w(;6��~Q[�,��vk�j�S�����1����R���d�y��-�&���{�u�6p�^��1�n�]�{#���hy���Z�zim�x���w2t��t��<�Tq��E�4]F��*[���N!�\7�*�A\p�}�Fɂ>
�ύdL Q����T�j*0��a��*�� .@{��R2�+�5�J�VX�	��AL�c���:��vG������x�	�������7c3����N/�@�q����R���7SN~����p� ����<�SE��~8'�g���@��� w� �;
x�(O���p���$8�#@䙫?=i:�e��S��V���z<�/�`�#
��$�e>&���[Q'A/'J�����Y����k� -�����c�Z?��`���~��$�C�в���>�h��S�a�!��Ǿ�>��74,)i�	H��_��.Mt�J�wj�������9���P?����4k��i��uL�2�+�tid7��.�M�c Ѿ+O�%��S
o[?��g��R�~?��y4T"��;�6�+)�V>G��|Xb�i�����*a \|X��<q2�ŁV�n�_�	�>m[&�r���QBh�-Ya����Z��s�?��5��򲺣
7b�&Q\����zp��@�;��_ŵ&8��M����m�7�[���1��t�)��O�_�ɔ�L���!F,j���H���dD����=\5���H}u}OB�w�b?nWᯀ��T�z7m&1���'�;�\���,�#Bd�h�5�k�
7]BtU�2,ر%*p�|�2b�DK�e0�DU$f,�X�$ū���:�����q#����liD1S2:!����N*�A5�/|4�X�К�\�)^C�������pOF��)��s�_���3
P��R��ĉZ+�,l!��B p��?��
m��Oؾ�V�g�n�yk�%̅�FgvxK���DP��(Q�QٷMHQ�_�u�+�b"G!]�4��~���A?+CC|�+M��?]�C ���!Ņ�Q=�-qNH��d]�s�}��l+���
�J��w�O�+<�Y[>L�Hd?y!@)l3
tΤ�F�\��iN����u��h�9��F;���Ώ�gr>����h�X�@�QO�WG155טBX�ئ`g!kDI��ДA�'d=�.\RDlu�Q���=+��5���x�Bt ˹
�m�r���e/?�P�^��a�܄�+5>a,�)1.<��B��Q�7��6����K��
�h���QD�O���x��*`����:��D��VS��'^~��R8M���# ܻ�zFj�Y��gs�Q�w?�x�Y��0��yE$�]d������Ge��U�%ZrZ$�`��1�P�1}�!��G �&g��VWW{SBJ}�wy��mEY��1s�!�HgS0Ӓ��&���Uc�*6銐G>��\1sǴ
|y�٣�"���,�:�.��J�wji�Ip�F���G!<����ַ���t�@�c
M����g�k��(2��<3,./Φɗu��]���>>��1�{@9<^�]�����(TH�P�;e����`B�8�9j�:͑��U���xn�\�(�/�x��G�Z�E����47+3�[*@@J	kk�T.�� ����7G��oW!�r���(����_�H�G�1P\�:t�Yc�yNѰ�i��O�T��O���]�y��S�b�k��}�����o���ܱ���nf%����O�.�)VQ��.���t�T��ed��k�[�4�q/9G�uD9��:��ߓ	�	��
@4c��	F�Vyn�_�aㅽ�pl��a�;b��>�����h5ꋚm�o�#�߆��OA�����Y$��EL���^m+a�ͦn#Ɠc�ߵb2�!%^�n��XE��X!)�2)��a{��{l�-t�KZ�Ϭ�p�y};�1��aofk��f�g:KL�J�bQb���8^�����6qq�`� \^���/d�݂	#��Ѓ_%�oD�ﾂYJ#v'h�Ƹ����1'�
Y�b�I�S��}�	e��/���Tu�G��l��ŖJ���c.ۡ[~�5��c��iv�m�+�W�"cb|"�~/��0�f�a����Y���|G�v7]���A��u{Z�Zcn�0 ����Z;�l5�y��G�Ŷ�^�O�33�� �aE	�>��U�Z\�m>g��GX+L==����Vm�b����
�ϒ�)a�I�p�+��!�<
YB�Б�裟��"��K�%M�8$K�o�G�j,�_<�&���{A4 �2J��߼`z���������\�5oJ�KԬ=[dC�)��Ƿ����0�
>��8.M7@Q��Cc��{��m��᜖>����������zᶌ,i��j���=��NJ��6�L��l���G��@##������O�^��d��mNɀd��.,-�7,�xj���h�Q���jkk�Zm�@4dɁd���_����0#�	��������}0ȉQC�����H��4�������v-*��_�w��u���H�_�q�^��� ��~b��{ů��I�^E0N���+iT|A�$��=»͞�W�������-�з�'a�c]�|�Tym�iͽ�ӂ�����"<v�ō�W_gn{<<�ǈ�^���ެ���cY���o�K��f+R�pC�sӭ�X�+^H�H�R�R��LNvH(�}c�Z:,�w;��ȉ`\z-;�s;8Z��h���"����{{P[p��;��o�]�n�W��}��qP�<�o���Gq��s����3Jv~`1��#OW��Z�&�|b��˕�L�͘����_E&oƞ����*�Ƥ�^���@IJ�2$a�h�R�=ˊ� q+PR&��6��t����	R�u'�+#����C����$�����w���K���s�@�oG��_kw;[*�D¥�xg�_�|�>���`��o?_����@��������᭮mIZ�j5��5��MDlg��p0����'l��������F�tmh�3V|��8y�;�g��^?TVR�ۋ�ӆ��
��n�f�)���G�C�˄Z��E�'���;%���$	� �`������+��*"2��K5���U�D/{�Y���8��uѼ�5�XƬ*u���7��45+Y��=c��� i���\ԙӷ��6il��}B�`B[$�6I��2}?��j���Z
�zK��[P�@W�������(��M��R����3]�!�GV�l[T6#��n�z�bB)���
���cF�_?JQ�J�����8O��Gխ({"R���#d�N�{3ǜ�8y��:۠��D�g�Qp+%&wݥ�(�������M��dƶY� f�3�~ŕCћTD��}EۖD+{BU�-�F����ϰF�jZ�S��O�&9q,��O����Ҁ������a��6U[�����*��vF����� �{�'.	\�)Uh�xN��<����4&�I�
Jhj�\@4T񔸘8�6�J��p��F�P?I�i8zH��
@��%g��V��=�~5�\M_W�V���E+e;��D�p�IKN �YN�>����e�~���Ǣ�ŖF�	�_��"hWM���2���L������Y��1{���3��1�'��z߳b/�=e���
��^}v�V�������"F���Ĉ�^��� �?�)DSD�dr�ôl�@c�*V,��*[�U@I�=�n�O�j
,$-o��_f�'#6�O��K1Ӌ�Vm+���i��Ә#���rPZsm��ɍ|��TK�(w0��zÈ1����V�h�~Ý$��>���&����+��d������#KD_nc������і��g����@����U���Ȯ��o�y��0Q�Ρ;�0��|tb�����9<�"����EMvzo�&V���޾>�b+��1I��{˯�E����T�]D������_#�#-����-N
�Z&h/I)ɭQQ�D!��m]{8��43�����"w���{�\�En�>�9��?Z��l=��cx5��eBoW�]	-d����$!�0C=�(z���!�,�H|�nfg%8<�
��]�N�n�^�8HǓ�r�A�v=4֠X�,�M@���?M�AX�W���/ypT��ܚ�2��
-U��|K�^�� ���$<�@.ѕW#�1F�}��<�:w㌉��ږ�������^"�!tBU�N��>��ə䟺_a�E�h�L�]�����������A̯ѩ��j	�ک��$%e~F!��:2�H�>\�\�X,��K��w\���=��v��"#S�袂g9vۮU���O?%��~�B��?=~���0LZ�`d�塔�P��J4�&/�)��<K�Ψ�t�?��"��n�lJq����˙P�⥂���C�zB�ӕk�x��ESk�D�
3�is�*�I<�b5ɲ� )��4,@W=�Y�1 [��9��Q�#O���njnn ���K�`a����QX���Ĵ��'���u�n�P������X��25��O��&<Wc�q!��4�*D͍@�cV�t�������o���pu�n� \/�e� ��D�9f�:$�c�I�`��ch��#��}4g�7c���cT�tt����$��i��Gx���/
��(z�$ǣ�z�0L�ǚE�ڎ����Z�C��AK#��8c���Q�si����M'~���1�KcB���=&��`�H����#��(��<<�	Z��h([�!q(��Bq
r~�
��f��~*����m�����.qj����V�$���=XT�cQC�f,HZ<5J�%���f��-g]��Gnp��s�̕�9�'�	_���U�\����97&��Լ�E�x@ɴY .|����l�+�D�S�G�[���rx_����\�]`~j��!n�[�^�n��`n�JӘ�G`�J�o�U�tY.&ࠀ�����}.q�s�A�� ���ZD��0��C:��[u׃�ee��]+��x4ʸ�,5���&
�b���Eum���(Z6��T;Ǖ����3Y�����d�䏫�Hڌn�5[0b8`"���Q�C�#�w���c^�Ba�}o,K���Nu�l �'��㴈k��f��ծ�J.'�	�ÂC*+]�j�l��t��ڬb�*�����#uT��K�������C"�E���(s*�lh�2���ǀ��C�m��0&��ۂ
5����������L`��~�n�`.�v����,�RJ�{�n:�ZP�����\�HɈ̘�-H����[Z�:�w`t�֒TH)�\ԣ�۪�S�h�z±$�Rq�DӺ��`p���dhik*;#R*���<�~h6 ��X�~'���vFC��=-��MwEp�o�;�&����4oE�,k�h�ǈԡ��d��������L�*�e4�^#�����3�?�ѹV�pü���;8���pj�y܍@�B�F,�f��ߐT���u��
�+^�6i�̞ݺPS_A�B|)�s�0�����y��Ϊ��P��8�qń�����+:0��8Y�K�K�
�
�Kڕ�Lc�ݭO��-Twf..\A��٭r nb�άdu(T�0������\n5~U����-����j��;�w,y�zK����3�g�>\����^�qL��x���_�n�~KPx�$u9x�� �kަ���`������%nHx	��:���Qe��ݢz\\��Ǖ_P��!������]�R��;f\�8짯i��ج23�Ԅm��n�Ib�t��޶�7��k|-Gy�o�rh�a����m��X��'��ȁ[�.wv�]Ԅ[��M��.k�0�@�%2�FhcAqTi����?�=������Ap���8��&��#񪚒P��N�^�.�k=c���6M��x؁U����W�[N'YWp�ǳ�AA���Sr���E�h�(����н%͚9UF
�Y���4��b��b������Iwn��ٻ��p����������S���v-
��kO'�s�l�Ў��ik��v�'��� 3����@������a�	�WV��YRFͬ7��۽��5�X��o��N��g̥���Y��zm����!O��tއֶ��i0���g�Y2���}ꣃ��pσw�#4Q$tp�XX<�Ã����*W�eD'�2|����F`��T�7dN��#)`�E�ڼ��_Lk�^T�V��P<�cN�TCV+у�$�Ձ�N;VQV�W׳��e���'�����beO�Kס#�����#:��mZ�����|W��Pu|����{�f�ә�N�X��wB�T��5�}~���������f���7����2�����Z9�Z�k͍�	pzh��k����V| xE8`��,#�NA
����e�l�q7`U� N�Ih���{)/���#�����FC�o9�C�\�|�P�	���VH�4\�u��uk!:�u%���h9p.�&�-#	�{�#) D��s��-2͂ōae��[���q�6�(��1st�@��?�Gς�j����������d����4�C�˜�o����!!�s�A�7Z���NƲ϶�)T��f<z�qr~�#���s�Zv9.�ZtT�PTm��"i�\����Z�ѻBN�ݨ5�!-�g�Hш"��h����R�9]�e�=��%��#�6������_ ?��I����8l�ɜqڕ:�M+0UUm���Y,�}~\�hc����_Q|����x/;lu瞡#H� ���R,ml��`�V0=�`՞f���:\ŝ�mٜ�̪�BOp`�F�Zg���#>I�`����>ئ���C�`C�u�&IT#�w�*���ʀ�0vu���i���I}L
�Vu�ld7_��H�� ��!T6^ܒ?����Rt(���r��v�*H��ef|Å�0��������Y��)$0��s�u����֐!���:����Vڋޚm"�mf���i����0�\�±A��t����q���}.|%ɺx܌��,}m ��u�+Nq�1h�	s���<n�h!��)�j�?_�>�`ya��2a;�Y,�tJ��b4J�`nF��b�JK�ߍ�bO���BXO�f��Ό�t���ץ��:�Ma��#�Ĉ�[���4��	��&��݋?k��эΛF� !����:�Omz�o��,�3{��)�tx5̀������&a]fI�s�U�@|��+-4�(zV4��"t�h!H��ɲ���t����6����p�����>�cW�eVj�9{��%�ѵlįbA��d )����i��9&Kb՘�m�Ab���j"w77�0P6����[Qb��(������7ݳzP�Y���Q}������Bv���i5n߬�����H�E
�f�J�,>vv����oE�~1��yy}n����1�_[�j�^��Ȩ�2��W�_y%0pJīK�ݢ��P��t&�H�cA����=}]�c`K�o���� !_Wd�d*B�؊��ǵ��J�3M�-�Kt�va�n��(\�'H�-�c��.6t��ߟV�Ϯ����6��W��լ-��ԓW_lfcgm�"H��q]����s�����3ɾ}Gb)�b<쀓iAQS�	B�e��/a �Q�ܮ�l�E�vb�Q����xe�T��*P�Ō��N{P*h��� Rb
���P'�M�h�U�*�d������$M����a���E�MO+da�V��d!ȱj�/�r1�ij ak;��/�/V{�h���B�C�ry�);O�(rv]����S�(ɵ�j�ڭ{Ch��'DS]#�3��1I	~�$d�)���{0���<,麞NJ�M��y��V��i̖��{,�sa�'�9���xh>�����A�!sȒ��2H�Fz��s���������z̓uo�@�jf�h#��ĝJ����[WIxh�T�������@pA��� ��QrcHjw�m�����U#b�̋�*��['iQ����d�"0^�%>�<p��f��^�wxYM����s���>����%�����}S�G�Pô$��c�OT!|ߟ徛>_~a���5�u>:��O���3`�z�AI�bK�%���iͮa�HHa����Tj��P���9�&�H(xw<iR7�G,tyf���c����vZ=QYY�'�6ud�*�����M��>�%��.Q%�#|�\�|m}x�2�����+9b�����	s-�2�	�eW~o|6�R88�@�%��^�ޅ&��٠~D^��D���۾�m/�yCJLI3� E��֫�qu�f<�#�/O|fʻG�O��7r�Kw�.)�}�<���HC�(Tcn�xg?���5���K���&Þ�z���L��;Q����$׸Ń�Z�J�X�\+k�ٙ#�D�Ĝ�u�R01h�´KFH�������%�^?��?!y����_1UH��$���d
�B;�i�������8P
���~[�YY�[����9���>�B]BB*��{\���`կ[��Һ�=�Y$���kή�H�pg�I����c��ӄek5`�N�r3�-��?��������j���n���(��b�-?*�F���nC�W�Q������1m�p�N���d1�!Y	ǚ��]H�t�s��X���pk/I�|�jV�Z���*�?^f]����T;!�O��+Ⱦ�@#�mJd�t�_���y�}�f]�G�?�����O1�M/�G
mxHg�S{��iH��YȪ�� uCū��AغN6T����h-f3փi\��������^�aI��m���'@+��DvX���yN�]K�_=�����G˽N�bHL8B������ȣO5D��p'��_utZ��=l�L���1�al��YS��x���2���w��=j�X�����SsӀ\���xl�/�q����#��ww\���rX�$NX���u�
BK>���]ac�;ʿq�j;��*���C���(]=q��>KeU��Xi��i�q�[r�u&����e������`x�}��Ir�S+�;�MWj�lD�T#d%s!)�=�U꿓[�;�$��9�W�_��Z���VF&J�3e���*�����gPլ]նf��.�"���la��AV�s�,��MI)�E�\�H�AR6l!�P���,?����d�^_�_���lP�b=����c��n�eG�$ѡlJ���7�!;�-�~�d���+EtE�0�ъkG�����P�(T��*�F�/�u��ZsǱx*�7��J��v�z:�|�'xl6�gba,�`���Gϓ�~�׼�=t!F�0��ᘷr�Ud2�� ������d��S����ma8Tt�(��������6�y�_H)3����HC��$���ݨ�m�|�F+����zW��[�	["�0a�B������<*;9��'��9�t�D�IE| �m��%�i|�L|�~䝦clå�M+�x0��o�g��#S�{O���n�ʠ.o��'PH�i�<��Z�`���N ��8뿝��ə�P2��2z�_�ܦ����T��{\�N���]�+2�ѵ����Vhs�ς����G��ɬ=Tܴ4����H��iu;q9l��& �����$�N]�����(�E$��"r'V�|:���^�VI�;0����bj����S�5kՌw&�Y��}<'I�H���*�?nvHDӠ O���UUE���r�y�ά%Ӓ&'�'�� �ɷo��8����b<�Vh��;c���Q@��Ĉ�� ��ϥ�T\�PB���`dϯ$$�n9�0�%Wh�
'�	Z����a�i	E.
-2�9�$O�!���e�=����P��6�<�IԌg�bt8V���]��Oɜ�b�g���f�B36��tZ�s�(��!,H$AU
�x��f�)��h��v�@���.��{gz:P.9J��J��[n
@I��82!�H��s����q>��ys�Ie=�F��|���#��\�G��exM�c�j1$�>��M� ��)8��B���` ��b1�c��#z)1������"ow��]�vQ*��x*���:QB�M�#*d�*���bvO���rZ�A���@k���Tg�;��,�l���"'.s�6U t�	�X�� �(�	,�%YP/� 
*H�E���8��*����a��}a�8�<՘q��� �R��2O�߸Y�����?�.�z�	C>tj���ЉG98���H�D���Ô���TVA1����[$��Fs0�#�-fM��T�*+�=��� @���.���=�V� �yaˈ�4 T�q!���+A*�,��cǗ�
a( \#�ۂ/�s�d�7��@��p��}I9�B��xh�ƍ�~�&���#��ȃ|y�E�a2����1C�n��倓�'N�1���a(|n��t^I��!.i)l؅ɝ���Z(��g��+��b��Y����������Q���]�������4J�Nrn��"�'9G�M�y������������ �C�A�,Ģ�dB�����g԰����3��Mܚ�HPCK]uݵ�t��?�MO��dF $qJ$ŉ9�?��=��y���vz��gI��tf-e�Dy�f�t��{I�7Q�0�ra5mCw
!-"%��]y��<��YZ�y����{ ���P��0$�u���~���G�B�ALs	?��
@��/�T��b&�ܗJs��o����G�	Z�~�\����O|�{\��x��<�S(E�Pz1� �1����ͺ����曯s��ϩ(���N�s�n���"�F�ǩ�Y�9�#+m�������@=}�@uvv���C^��ED��S��ZZ�b]t���OF�}x�)�6��<#o���K��8�n�� �	Ӝ���O�铧hf�����Ό�B�*��.���7q�^���!����s�M�%�����`"_Ժl)��vsafOO'��jJ���U�����%d3��F� ��	$G�@�X*�0K֢3 ��2���fo��T�@G]o� 8�w�������s�I��l��Y~xi8��︑���a�#c�|���
<0�
�����{f���3z��'ibl�;* ��4B�����V�YM�S(��brY6�ug�h�$i�rp*�yL%����_}�z�{�q ]���H�59��t�}�S^��ha��pC�*��YG���y�	)��0ؘ��a1�9l�&����j�{���*	T17�ھ�bJ.�BF��eB7�f�����H:x�0>|��zqH�J-v(�w~$������˩�������cv���<,?�r����j�Zr�\���x4[��x�,&��,�
Q��������0e�V�V�x�9������t8J�9ǘ��+λI��i��B++D"lS��Lv�����S���s ��s��b?�XGIv�2�E[�ii�l��CNY�����8z\�HY/K��ɺn[����+�閛n�rW=��3<_�9� ��M�ޢ��	�J�i͊iى�j����)���H��Xa��nx�U��D;��Cy�����4�F<��l�� %p���2ir�z�b�sڭ7yʟ�d����U�=����BdB��R?qekBXk�r�(Y����4U^榛n���j׿uw�
���y.�*8���d����m7�B5Օ������Mg�{Q�Qs�c��!�ȣ�u�Z"��uj�(��F��k�u��Q�t�g�I����2P��ڵ�c�U���P����ˡ�gQs��X��s����d7�B������۽�]C�L��CH2a(CH���-�b�\r�4$�� �L!D�(p���N���E�A�T�e�8iIc]{��42<H��z��f�z磊PǀRh�S�9]���9�|�@!u!|@Q�Y���<t�)"sd��xV�?:7t�CS���S�@d�3+R ����u��S��kГN�V߬�by���5c�@I��xV/.-���M�b�O���pNƷ�\8�p�ҖV6*P����n��X��Q��$y�՗id�_��\-���`�d!D,���Mb%>�q���A͞��Ĺ�7]=���FG�9e���i7��`����C�Q�(�Α@I�
����X�y2�����ìLF8j�a��F@ퟙ	6s�K*}	���s`� ������ΉL,�R�TIbz������O౦C�8%�@�f�4?��R�
�(
b��ۯ���ߠ�B�shgg����Դ�]��n�.{�&蛯���sp*q6 ����D����eS7 ��Fst�1�Z-�!���.�:;;}=C�����M2�'g�r�#)����b@I܁�qsH# E�1VMGna�Y5.�&���h���,r3"g�ֆ%�|ͺ�x�2�DHvZ
3fN���Qoo?uvw�|x���O�Sl����kt�gg��ϓ�椻v�f�O-�Y�qJ1�=�q�38wŊV��*��n��BN�����a_�@۾�@�7̉C8��C��;�H������K�8���D\�ؓ�JZ�\��Ř��6�Qd�%w���γ���&QC�f��Pr&�7x͵;�a��9	��rB��5�]�>��?C�O��#��㙰��1J����7ߢ�Ǐ���:��E	��Ew��Mi��±�B�t��qL��E���CM�!r��~�Z��`��n6jC����*�s�l�1P����@=,>C��Z *g��A-�����@f�E�$��\�z��Gk�K� K�23\�3�Q
j���8�A����뮿����t{=��/�ф�,NIQ��5ki���TSSG㓓t��Q�w�~�O��}Qt#Z���3�
��
7�s���P���#��AX��L�|��׹���j�$��9y���j�H�ɠ�-�Y�Ի�/}P��:	��,�
V���-�.�����,$It��ݠ��Ǔb�$,7� #2Q���F����Iͥх(5�Oe����ʫh�ڵ����c.�\lc���Z������a��9s�)1z���#�܆ÔQY��p�����]��(F��sl\#׀dY��ˇ���ޣm�D1���81w�y;����TL
9��G�<�K��$G����C���*	��͋��b�$�}*DTϱ����������/�`�
D�% F`�����laDN�"���X\�す,�︩e)݈��%|� �D�ڌ_�ʣ3�\�r�_�b�Q�,f���|��2��CP6�'*/��[4#�
�� ���vx���̕S����k����Y�MMO2��[��*}^.��(sa�����j�//������Ý �bu1��{�fs��!� <��c���p$БcGEѽ�DK������ʝ.6,�Y�Q�9�4�E"(i6�H�DQ�=2����u6r�����(<������`2dg^I�2[e�ë�y�ā#��@�hSU�8͑U(Y��z���K�H�DR��&!��������e�-l���D|�J����[�a��NMsv�����K�����R8�ؘ8(.+N��\_�җ8Ŏ��}������ۯ���Edr.⟁��� ��B��8�����yr�ʩyi+��5pY�5�AY�c ��K$ENT���Rpf���(4� bBK2��G�w�w?���YGa(>;�8c��f���H(��P8BVBY.�5�V���Mv�a�n6?��]|����]]�]0&�Q"� �K�5*�E��ָP���*�\~�_d"�~����Xy�w7�jr����k���;���t��;J�S㬯�<_��������Z�RdЛ�P���g�qA��}�`k�e��`�&�l4���P(�c��j�뭢]�?@!�BB]_T4�m6�z�N�3=Z[�q�!��� �]]�(���:��t�V�u��o\2G!�������ؘ��#I���SX��8��g>��������|��_fpp�ց��08ص|����;����x�u>�7��ʱ`1��I�s|Nt!�s|�h)E�M�ZH>�)ǾΣ�.�&3�Gp�W̯	@�rU�ݻ�T�gl�>�3Y-�e��Ƃ�o���W�!�Q��-p�4�����Z�ԍW8\;��l��$��yG_�> �C�x���16��*����9Z�HE�b� �Ų�r���?�b������"��`8�۷�˃E��𵠴���~��_y� sB?<ӕO����a��N�nD���)�rg:��)������q���@����H!a�Ru�t��܄E�s�ԷX,N{����-[7�Q��0�ĹX�]o�x��|��*o�]�v��K�P}�pqnŅ�:���������D��D�	E�d4��Z˖�2ѐ����lǮ���E'���^G����Gޣ��,G��k�Ő)��@F�7j9{kЊ��}�X�N�8ΟũrF:�ƭ������q�$Q�Rs>�SYI��q'���u��G��K���F��n-�s(�#��
�韜 �FK��U#uU�W;��.��������} 
�P��K
}P ��譅8+w{N��bF(;9v��jjl$���ā�������R�RU�4<e|�&�]q���רU�rD�AXёH���u�ѝw��;���a� �s�ё��;������9R*��}��W8��b�Jί�'��\}�@a���h�`�L,�f�KZn��,�1P}����G�Dh���h�u!�;SS�~���6����U��KK��t @�d�0�'x��+��/����5��	
 �m@9��H��l壃P�@p�%��*}>�ۭ\sq��1.#�UG#��{vR[�����451Ʈ8�,̓�VVs�zU�H�|�0��O��7.Y�4OfŹ#b����*q�-֊5��124��˚o��Z�.���������@D��T|�L<Y(5>ט(�(�G���
iuit@�����HKpS���Q��AT
��a�CX�M0��A�B$�q�n��	}�bL�ٴy+�56ҡC�xr����T��|[6m�t�������m��5������k��̖��`ꨦ���g'1���Ç��ɓ'ٴ�d����V�-"�HyX=�m�&���"˜�onn���j���@��s��Ύ�&�)7�:�8'��=��-3�g�bw�O2E߫^�J��H��aA��4��.��Ur�����C���b������*<����1�_���lq4mc}3mٺ�CB��y�[k[7o���!z��YG�x"(�X��Z5-mYA7�~+����ګt��^Ӎ���-��](@�8J�9è�u4ܩIOJ8�M�u��ʬ��e@�m>O6�,��%�狷�>	��â+$�51����֪�
�~N��.w�%ǉ?q�$��������Do��&�w�=6�JԸ��{>����u�6PM]�h��F���ǹ�W_z�����$PkVo��v\K3� x����ssZ��<{���(�Yւ����{��J��<�܊�.p�{/l�\����-YRdQ�EJO�����%�������'�lى=r�(E�b[n咔�-܎��m�� nI�����w/�%&�3��`�ny����)�yw	[a:��)P����U����6�H������E�Ό]��Qn��(mk�P�����) 	�#kg;�'�ڀӥ�j�^����&CwŌ�P�\˥"(��-Dc\b���Gd�����]�.#�CAn�������=+�8�x�er��۬��ɇ|
rsx�n�W���%{<*o��M�>��a�-���݁�
�4^@�nx�:9]����WRR�;RY���|��7뫋��8=53m��Y댚�7#��a|?a�-�ײ.m��ښ�g{kD��7������(�9g���^mޡԃ���	Q#0��@%��;gHQƎ^M�ux�z�JOw��ݷ��y��_���{_�cf�7It�H9t���%�W&9�� mhj�k��`��kZy��#�������졆��+��o�ʮodd���������L�K���G�����U�L�֪V(X�y-����=iQаQ-	l9��ɼE�����+�ȥ̤�����fQ�cJA^.�������f��N�)UYUK�T�;�7��L���
52�z1�S��ZB�"2*����fݨ��{�ڗsgC@���
OF�(2�8�Hb"�R��jU
�^<��LKI[�e%���/z=�^(r"�y+�4S^V�<e)	"��P�}bt_h���-���0�ߑR$��t8����_l#�e�����0��h�2�=R�A���T\�6�]l���F����l��#��<o\���4n/��eFwj=����q���_����{�8��Q��LL�C~��C��8�J��*;C �Cr���ʺ�!���O��lhc-�ҷu���r�&Ϣ�<3a�1�ʕ��]�n,S1�s�e ����sޯ���LeAA��5������9m��#?;�O�[S��=;�l=kJ'�E]����3ȖچtXN	�ʽ@���r�b0�YZ	6��:Z���I @��������zRڐ�Q.��e��"�[Y� 0�wXQ�X,�>�8I u������YO�����ç#����( "ct1mQ��e �>���	�Z������$�0��NM[�(Z�E#�S��}��hDC`U��	���2�|$�q�T|]}�re岛�ka�a�@1ǳt]֖���5�aQ9�Z��ϗ����5>֏���6��?395U�3
@��,�̪�ES)X������ү�c?��.��z��z��l<��,k��e��k�d7��27&0(�̐��I ��� �k6���ðo�vٱ{�Ė�T��II}\-�Md
�Or�fqa�J�k�e�_��3j�V��բ���K�������5��O����D�H����H�ٖvw�}S�� y��4���@�g2`�bH��x.K
n��������xYCܶs��E��ypG�{��a�%=/e:��{:�d���I�������e���χ�O��a�>h�ځ�-�*�H �6�y;�e-�ֺ�v 2�
���5ClK�~MW�������c b��"0a��zL2��6��vxezn�y�����G�������4�����g*'�H��}F}YY�!7����~������E����ȩ`$�
��ZH�Qk���V��-�ެ�L���n=����z@�%�-���S ś�������V�y���7K���%;�@�=�4�u�Bl��4TD Zx~�4����c��@�u?�Un��:�� �/kۚ�v�ñ��*�=�{F)P�p������d���,%L�(J�ыi��ݥe�]�Q晦���[��#>��fF�iK�E�L�
\��E�ݿ_[:(��N5^�n4 ����t\)Sk���A��D�r����鷪SY������p���Z�p��b]+]o3D|�+�@���/�K%3�0�:�M=��e��>��A��5�P��<#�',��0}^Q���w@ZZ���X�)E�s���@���\�̡nvÔ=�;���������49F�t@�R��/FOH����&
������V������o�������vNe�O;P�(�&LB�*	V�*PЦeu,�[�c1)*-�=����f�!h� �T�'��AF�MV@(�cd� >BX�Ǚ��"�    IDAT����8��umd�d(jKv����[K��~�
��Le�^��̏>	P
���������\X���2��Ok��҃��"�F��B�U��t����r^��D��-�#Ci62(�Wg�	���3JV�9��EAұ�(�_nki�g�����U,
��7GO���V�>X)�@��ir��V%2]��<k����QW�B䏼�$�Y��c0��4�����'��W��1e��i�5��TZ|�J����ih����E�f�YR��sq��^Z����FR�2�I����[[~wC�9���߾��ԢX�C⻰(+V����\���E!�_+�M�EI	�o�E_����eZ@����jdh�$L4�с:d��JPh�[�#f��oZ@?���Ҋ
ٽ�Q��o���E�>P��y�K_\��K=T���G\�D�S咢������_8��R��&\�ԮߺU5<4t2uL!<�Yf���|�V�͢쁃�?�ͨ����p8S��A\�J� U"�.%�iA1�WT�q�"`39����'� *���pX-:J������H0�}�x�L������đ����+/����2�,b��1[%	�Hs &�R�1��J]m-�}}���Uy])���-m-�r����n޼Yyex�D8�����F-
@��j}��x�;T���h)�&14�����:@A���E�yL��������/@�l##A���"J��5~�>w}`}+��Y���J<�г�m@�VTq8���'�+	*�0��f��l	��"ifW,Uf���L(�pe�RRZX���t�~k=�x�����ъ�#� ���(�Ei�/(��
.�Fq
��钐��_����0�d.Y�?!Z�pp��A|�X�o�ii,A׵^6��q���[o���,'x��P��zL��F`�!�Sʫk�~<��H�c�2;?��܊��"��w����{T����2��	�9aT�O����m-�z�@]>
�{4�Xˢ�e?�4D��?$2|3?�֎��������{��\kk�#�� ����׿�v8&���H� ��j��O>-M����+�J&0`�4��t
@
@��ZzY�'a�HU]�<��Ӓ��O��/d��eT�P�q�
���a`?/,{bb����*��O�������!�����oܾy<mZ��3J-G���T�	iڊ�A���Ӌ��^N�3M#<�cz�g�����WV�W��U.��W_�����9iii�C����Ŀ��oS�;˃�� ��9ga�nCi����Y�|�nXH$9)�-��8����^`Pq�gU;� Y��A"o�]������Z7�:ohh�?x��ہ`��a@����(�nM�sHݟ~O'ӡ{Z����cX`�����
N*�k�K_��x��28�9Z��(H���c�����wI�.1FQٚ���3
[�qv�OR?����@	vWa Գ"='-�sr��e���}�%����A��H�ih0_��K
��^_k�mȢ ����ǂ����3
�F}
������&��ڬ�&({�4��C�t�Ǌ�x�;�Qijh�5��󶴵���EJ����z�c}�d�N������_s��|�E���V�@;���EA�������b����JR�.��W*'O��C/}��=�pf���{7���Il�R˾�¿�����j��c
�9�nP�����3J[jQv7��c�������'
� �a��������o�Ɨ�M/_����C����#~y��WY�C���!�޿{O�c���$
�
�	��Zڻ8m�ٮe|�uL:J����~�-��G��`Q����);PYnY��sSSӟm������{w߆EMbq����@a��(3˻*^�d�$;3I������\x�#3�nF����$&��%Y��O��Q�fcmї��2'�1�7e	�C��_X,u�524p���8��ʖ��\y��7���+J_\DJ����p�kvq�	36`0��b}��-�������() (������u�b�~��;��bC@���B
Su(�jx��D���3J-j���@���ޖ���;��%�0d̚=R�h��R�D$�A%7K�J��.(\��hm���"�4�"��!JC�/;/[�f&)y*47��k��5�4�@�4�/���M�~�9j (��T��V8}�$W�a$�珤'���MAX�(\�,�,V���fG}��T@����GP���}L��ي��]��2�)騅i���K����nnk���#0AJ2xv�Ch�VЭ�͝b��çf�4��\^Y� C��c/���$ ]������u
S����L��ŕf+^ON.}�0��L�0�[@ee����3j���C 
���U��@űl�,T��~�����n(D}�H�@M��f=� L@��ث�d��鹳�;���Q޹HQ���̿��,Aq6ڔ� ��u�t���������(591*j(�X�,���c��K@����9�8�ͅ�_Wo�<tX��IYBg[\��?~�3U�{�L���p"���ں:���r����/wԯ/]��b=5<W���-E?R��r�ݢ�g����ϥ��3\J:�]tX��U$2%��n1i�]8?;˺�G�.G��0ZyV��;/W�p*kʝn�� �z�$��$�|Q�ЪE�rs%�J(8�
8����"ٴe+wPE&�%73]x~ z����Ӏg�y�7��� &7��� ��H�U��_YWJ�c��s�x$�U�GH-������e��gZ��<{�`����%Ώ��"ini�,)������q����-lvz��$�P𐚀�Ƈ�+��1��,x�&>v���M@�fZ`q\�ͼ6��_7�ԙi��
�|�R\�=��e���d��F��N�;]��[o��:���?q���M���G�>�%sU~ߗ;��7*��o�=55��DҮO��̣֣4ۭ�nQ
ȋ�n.� $�U5���*y����߹yK��Sye*2IIj�,�P-��)�Z���h�Emݾ��Gu���G���b��4 ����9y���s�4�C�p��h��;��lZ�YLZ
Y�(��>�ԓ|۰( ��PH�	�35[Q��rWCͺ:H�(e�GG�M�L�R�p��+�c7h��je"�k&��0*\�2*
��R���9ҳ|X�ZZ*�uĮ,����!u=p�*�x�&\`;��O�D/&1�*�U\I^\���=���"/��� ����ClÃ��!P��M ��UU���%��l���I*����ky��I	C����q\��v�(��H�T��~���n�u���&''�"�S�Ɉ��M��[�H��7�LY'�����zIf�����2.r!���f ����G��T�k��5B��o�)C�|M�E�
5�v �C�S(hc x��ɚb�&�C����|�+_���R.]��!�"�� ����/]�ze˶�܏A���ɜ%E����c\_  m�����RL&�JE��FB2���3>]�/�\Gm�+�
\���[�"S�}��im�f�Z�LR�,;�'���=�[4��P���Vtf�

	R^aU�0*�_�+6���d3�P� �`�����;���L���	B�(���`-%i�Gw:�r[���g���Ξ��\')���D�쯨���wK�-�K�77?+�,@�3'[�|�����K�~�ި������ȣ��UHɤ产�J}/��խ���c��q���k��f�� �Z�Y
�@���n�Z`�[��V��LZ[�9����P���9dJ���99<�!�;35%c��� �F�Ά��zQ+��{=�Q�����3��SP}Fm�hy�_�]�J����ܼ}W��T���������W� 狍E��x���{���ef2�cO����/C�äP�2a�"�َHE��3�g7�G��Gn_{+�l!S���	7b�(d����<�
�s���@z��g�	1r6��P�.Q��{��0�>��)�+ԒE������	��F1 ���"]]=�/,B�1K����p�%Pv�ɑؒY҂a���Eʹ�?Q�]��Ko�f�[4�ofv�EY�({��	�h6�4�SO=�J��;w�J}>Ȋ<n�#RQ^�bgMͻ�K��+��F� ������В��hkk��c�	B0&@Б�)xJ����K���"k�ިѠM�Ca���*/�Pv��%{����\*���.(xi��m�t3���|t�28RC0��aSs�lٱ[ZZ�djn��8�S�,(7ai����z�j#�=�OH��4��`pT2��d���׺6�����n^�~,<9��(5����W(�������2��5�U���Zd��ZL�k�A�޵"���Z,I��� ݞU2:�SCs�*2"D�8ySЅ͛A�x|%��P9WY�d���d��G���S���xF��!�B�2?/GF������q~a��Î;(	k��Ch�{]�H��Ӹ��q�����g�(��(X���w��e��vW���Z���}P:A`�d�T�\`�`��b'��C�nBY��(1�},k���dҌ�X[�p������9Īv�{����f{ejf�d9�ܞ�}��-�?v��y$����0*�9^������������`u�z��ȴ�(�Ë�3��Bb�Q�6G&wB�B����^�ex٦�g����A��}
�@��i��l\�U�������<�a;!��(�b���%�A�>��u�2@u^\NHCs����'	T|�֘Z62A�����#�@�ڸ�HX��R�m�g��n>Jŗ��-P^Rp����܆Ψ����C�oá�Ȫq��+Pp} S��Ŵwy��=oJ��,��4/k�Eyqfֈ���,��kk_�R(��-�(�b ͍&B��|ߴ*�[�͕᠗X�4�P�!Pb�R��-m�u��mh��3g=0�jmE��כ��"�m��c֓��l\)�c�V��T��6Խ{�JFF����(\<]��@iԧ	�=,�[�Z�O#3uc�|�n���왂���ʏ�<�pb(Z���u�˻3˾��B������<������
G?�Nތ����8���/�e+	�k��ݲm�^�������-�0{d˲,��48�N����c��H+P�9�@���Hku��Y��9iQx�@+2��z	�Z�z@�LA ���bi�.��y�sv  ��pT.�:�����	uCT��:�)���d�@��L0�A^���Ys��	�{_ff�������6|g�fٶk/��0{[�5��Z;Q�e-Z$�Y&QG�$�^�Sr�\�ʲ�#-UUl(�Qw��M[�d��(XJHƊ��Y�zn�5���֒~ pQ����;����r	��-�dg��r���;8�N�tv�����(��u�h�#�3U�l���NҾ��>h ���Sg^�Y_�w����E,�(� �1P44q�Bg7�;��!ms�A��I�F�+�\��������&��%$���
rP���TfNeoq��,e�\!��J�w�'�ɇ��%�Y0Z�c�n��w�.�zM�	��fg�sG����n�wﾜ}�=�I�YnN+(�F�g-qk�f���o�-�H��y�1T�S)�ۺC6o�%��<���K�on��g-E�X�iz�(�$�t}^���������*+�!�P��7ߚ��k}v�L]�tQ����4�S+�y��$x]� ˲ઐH�̚j����H��	����-)N�׌�@���/|�7���I^}�u�L�M�*<�v���jy^�SxR4.?�(���gNK`|�{<8�Z�w��<ota��Ǡ��>J���
m�� �sz]�k4�T���"�~����o`t���@ }Fiԧ��p�M�|�~�z�R��)��/���y��/ 855�(����PS^X0�s؎6�m���E���P���xd%��C�����;6F��ё[FY�e�S���%&5+���E2Lߦ9�曔���&#���`�CJ6�DAv;E���*PL�S���Cp��)e���N2侳���lϧs}�������cぉ�L (]A���P̝�i{ۭ0Y]�=4W�V`��4�uʑ�/е�Ѫ[Dq��4Gށ�C3��P  ׮\���W%?/��&$�r�_�>ڶ}���ԚV�̼LN�>���3��b������'����~A"��_P ���{����)��� S�:8���Ԓ��w��A�����QB^�0����l8���(�=8�v0��a���B����8�(F|��^]�gMX
��Yj_���7��Zۺ��_���:uF�9{V���[JC��q��\XX`��G�em���{�u�KV�����PO���E���0���O#Jp����|}��$����ߗ嘑H�ېX��lߵW����B H���Q�9�H��d�7�u��S��~E�셮�� ;�:�~��3
@�:�6(��)P(f�z,1�t��E�"Q�*�
/Hkk��#ϑ����J J�F�*  �p�b���g?�Yٳg�D�f�?}�/d)����EX���� n��\NS��ԑ+�P� f\k��z!F�+����P��S�f��@���Ԧ-�I�P)��-M%X)�Y�R�7�j�Z3,'h!�`�y^�;\U�{n�����D������px��Ҫ,�P�(�r{��T$JW>�ժ����"\%�Cb%іm[�f`p��,����h���Zq�3�>EJ��Ę��_�'�3�HV��h���y��
y�JZ#�Ѫ���"o���YbSh��C̵掔�4�͑�{v˦�ۨ���������bg�WNC�y.S�uqފ󻜍JHa~��|�X�� *��I��<(W��p�T'�~N\ �8 �RUU�u��41`�� b�䊯���jf� `���o��ی�*�"TLȹ��b�Zj��=* y��A�[[S�ј��9^�+�o�޹��w��C�+�"sSLtA���	Ւ�����xܜ�� ���e��� +R^����,�2~@�Ba����*�N�4KU�Q�m?������\�p��:���5�ո9X/�~]ÿ��.C�K^��b��c-��� ������W0G�f��m��� �%�,�X��#Pyd�>y���αC�������͓m{���h��G E��07�� ��Flw-
�l��x-خ�<
Բ��|����"���Zkj���5T�<1t�� P�Q�C��h����'
��E$����R)*)�PZ�3-������Q�6�s���_Q)AU�����yuu� U��>4eA�F�?>v�y��/z�����@.���d� �o��c�>5;�H���1:Ùd��C 
����O���0݈-�Kia1��,	W���o��`�{3��=0pb"�2Q�"�n�<�G�&Ʌ�-�R���ř�;gZ��[ �լ9_���0RC�\ϷV{�B�Fq8����
���?���wt�e4|s�b)���hre���y��m�8+_8��|���\�]�̥Ɛ���K8L����ճYf�Q�r�)�f��n�Q0V��o������Iݶu�4�4Iqa�'��\��<O�_Rvt�Q�8;LԷ`*����Q����^�����	e�k]��cX��`���Y\���E���@T���fq�+���H��u����{���30��e���L��1���bp���=�|�{.��G�z�sz����!P�k8��.6`�#�+��K�6Er�k���7n�և݉�]\w���<YY^��,+�x��V(Tugp��xp��X�F}���ϛ�:f�(��t�F�ݑ4c����=�C�U����\�_���\�O���踳%k���ŝ@m�^ *X����'���S�͠�0��N�cXȜO<�T�VqI��x����?��\�t��EXJ+��8�
v�? }[vHpr�c�J	�fm�Hd�a��)G�(УmߺE�+��(_Q�xu��Hcy���Qw�ܩ�u�Ι�P��Ttބ�
\�����	����Lf�~��$)�8    IDATš�`L�� �msT�n`aSԻ���;
�TXI
%��o�}Z ������ `ൠ
���,_�¯��91�����O~�CĪ�[��C���WJ�6�m����|���`�D���r�T��dRx�N�X<~ks��l�/��ؐ����l"��,?�T^�ᆀ�w�^��3��d�bN�M7�2��%��n����Z��In��L%�+j��G8;444�7cH���P]M�}T�Q���A~�Y)USF9�0M;��K�!��h>v� �n��pp޳����::�����{��O~"�FG�;H~���S�/������-��#�-{��I������
N�,l=�Y���ae��y�g�.)+.2��,�(�<�V�A���~��͡3�P���V��@i�g'�ث�{�<��оOĩ�7~��\�p��;�6��ˮ�;�_YA(�%���ϝ;'C��@h��(�p�I�Rτ��f�ۘ<��oȥ?d�z,}/�Ě:T.j؏��ϞyG�߽��S�W���Rv��/=}���R=���"��z�da~�����d�歴X�X@�����V���$S67�1^YV���;� j`t�@0�`�2Q�2y�YA�Us͡�۫�.]B�	��0:N����.������9yJ�|����?(G���7n���Qz�x���Y�����S�ddhP���t_aQ\�lf9��%���s�H
B;��2�ʬMlx�ȥp�aJ7A���|d�*�������ahj�HZ�и�I1:�˩o��� ;��v�`2�t7*)��#̷|�E�\�k����R�F�Q#cc�����N�uv�pX�*P�����M���"kщ���X�T[O�|��_�S�NqSeE7�����o}��w9�q�.������^�������I88A�=�	�Qpi။Fp�뀸1'א:�iE�ADMN�T�Q�Zт���� ^+,j��Ǥ�{�"�t}+�1������ܴ���?�_w�&iln���M�� �be"pO|B
�s$?������XQ���wl�����P�g,�0���^���keB�%X�(ܥ}�wɑ_$m
+�:�k��ϯ��
S|�B�`���Ȃ���/șǸ�"�����{��5���X)�(�#A��~�A61I���p����9�EU˞�KGO����\���TAA�,��ɅȽ;wd�N#��$\�e{I#�{�4��IU�_��}�J_�g+J��P0q;p�yx`�P8\�ʶZ$ʹ(����������-.-KmS�|�o�,9ٹ�*ʥ��G~���������&\���XL��oв�(���~��|@q�	�C��u�V6����͛�=@p�t���//�d�7�` Q(jx�q����*+e��sS���,�U��y�߸��}}-�4��Xu�f�8�-h�����$~�:[���|G��uW�2�\Żw���	�C����o��0Ns�FE����빅�N'�V�Z�u��an�O}�qijj�G0��2m#7G�՟���	bfuu#6tb�X�z��9�ĩT�9�.��5�Tt;H\�zc�r�樄C!VP���:����?� ^+'>����چٽ�i��$�I�ڞ%wnޤ��D(��5��঑
��ȩ�7����)+)���w;���~�6��u�֭����S�ɩr>u���Cr�m�Z�a���H�%�N	;� ���Kk{��Ta"zz�L_�u� ]kS�<s�9vTѱ���9��?�����at�K�r,�͓O?-=�����D��9	r	�	�\�t��#]^s>��@����ܹ5��Z�BLj��o�ili%k@�����r��-ijm�;w�}b%����@����3�A`|\�+1�nn��ly���r�%_j��H���ᓑ��RXSz�ׂ��PTiV�����A��5��̥�DHY�&�����zGy����E9��g�<��!~}��y�1(��rA[��;�^.+���|��+W�1�N���Y�x�q����]��ҕ�W�0lh2���[������ ����iÎ=����E�IS�:}�ܹ}�����'I�FΉ�_���{�|�d|�.�0��	i�*��j}���z�%_jtt��x���E��Y�>p���,�����ڴ���f/#��
���NV�$��*ܑ��(�͊|��b_	���dDV��e1�B;@���deK{G���o|��̉���p��#ee<�0��y��E�x�"��aN�^��~�ZFpY� ZTt�:�<��4�u�x $���ٳ<׶�������qZ���	�.g��b<��<3H��hhSK����R5���0�� *<9�S�؏�Y,+(=��%#��^��l�����\�1���p\L
�2ca�B,��[ha S2:�;+�5om됯|�k<���:���������]�7�Hum=���E����[�������������{�il�_~p^N�9M�
EKLj���B��U��QV�(rC�aXa6*��J_�P{Ká��5x������d��\��
�b����Y[��*�ԯ4�t8L7j�:Ȇ����F@���Am���ጢބK�kk��|Ub++,�|���Z���*Gb��VX�SO?�@�
��?��?��H���ˉ���l��g���������{?�%	��	_RV����a0%f��r�QT��ըP+��T�u�6>Y��m��m�:��.�[��D@d�3�^-רO�I-I�R"@����(�o�5�G���F6>�t�0<>����2�?����#���cǎIt���w���n߱��sQn�ELG��O��
YlE��?��J�=�0 ��_�gq�<r��!VM�Zp�rr���K�RzL����D
C干8?#���C]����G����S3��
�[�e��� ����EeZ�^���jYhw#�@�;� g���2qE�A�0&�(�2�@n�k#ΫP�����ԉ�.���^cЀ��
z|�A
FD[�:��b?��閟��U������N'w˶�R[�(�Ȕ�>��y�E�TX>@`ڂ=���\���
^�Kǰ>�͞��������ΖC����6tF��>8�����В�~�����=���~>eZ����%fg���i�#7_�	B�>β��A>H�r�
�^M%4�j	�#�M���!9\SL@S�,��z%%2=��a����a��x�Ɠ�&x|��Tc	�G�H[[o�Ĝ��� w����z�ݍ������B�Q�Q���m(L_��oi�!�FL�N[]��wg�q�߰��
.\���ץ �粶�"�s��e}��s�5g�Q���g3��ԩ78<Z���Q��z��Uâ�5n��ɐ��]omkz���"�a��q��=�˴({�k���YT&P� �U��oD���j26��;�z��G�]�pik$�� 0�3q%��ʚzV�Z����B� aQ���5�M�u .�p8H P%W75����6��|����~}�xdj� �ή�g�6���Mz�2AZ���)���?��<<�R�@�-,}g��;ݸfk����3����]����p<��%*U�uһu��44K����A:�0o�@i�o,ɸ`�$��
�ZTEI����'jkk#������oG����@��iW7Ӓ>)P��j�⾖E=�� ӿ����E^(�樿��H����k�X�����w뎝�m�>�����D�L^�ֵFTY���0�X���� 9Z�&��y�3����ÞƚCuuu������ ő[0����(�?���~�vwg?sp��_k�`) z׃�oR�x5��5iU�������{dˎ]RX\&���K�}���;P�� ��Y\���QF
�ƥ�����}���xjC@]�qc��@����t�Z���iH���|qi��n\��A�k�<
�
�j[E�@��*�{�$��p�(Q{U.,��9$�n7��[w�ޭ�%��'�&&���H.�:i��Z-�U+�E_ 
`*Y@}о��p�Ϸ�^�d�x�����oMNN�jԧg����^�P+[�"?{��߳4a���
�=3ߋ+�e+;P���Ԋ�Q!��\F���x��l�I�iM}�wH^��,$j�fg�ԉ�����Ʀ��IL"�U��|�	�IMy���-Ow��s���/?:04����lF4�}��2a�J$VV��L�ʼ��ї��x�z�<��V�s�4��h%@k��$�z ��Z�hf�l[۬�aV5Y��<��<��(�Ba ��'Q�[n��0��N��@$�@q�ōҳ&�xl3�aH������줔�������Ɓ�t����૑�lUm��8=��,�J�Q偮�U�P+�_3�Z/�=�6����C�K�4- P��G�*����8s���&�CY'��C�L�e�r�����+Yy�M�P�� �SL�R��]o�)E�:am,��:����lOy���,�����,<5����ڲ(��Tf��\�Uژ����J�����@፻�%����v��?2U�zt��Ja7;Ba[��T���K���I4J����ĕ�%P l�`,�<y�&�wg�he/�Ō��@	����̶���*++�]���3�W.�������\�Z�C�X�&�j=v[�z���[�������E۵��fhړ�{f�v�UeX�I�(�5+P�T,��ֽ��nr�~�	�a�#���E�����p�y�%��5��犥2OE3j�E�G����u����^wY�C�:w�Ҷ�7����g�\�r%���B}sF�^p�E٭G/����H�>C���+���AK�<ܹ����j���BkrLL�cJ���F�Z�8e,
@=��$]�LͲH�V��y�J�Qu9)P���f�a�'q^a.+K��ߗ�Jߙ=�z6nQ�._�q�ک���
V���n�L���)P�d�<���{kY����5���aoz���y��UC��)MY]�~F�D�����HDײ(LÃ�	���/JK{�R�/,��m�P�$g�.-�܇�FC����V|�b�k��*0q_���ۿ����KC�j�_8��nʴ(r&��6��-J�Rקo>���s.���̝�g��)PjQ�~k�J[�>9 a��VA`�&i�I���~�>�3j��3��
��� X�|���p�+8�x^�X�[@-�4U�C�fg�b��/�p��iS7�n@)`�rK(0.��eg��v?�a�w��5ߵ��7���N�Y��T1`|P�hJ]�'���P����!km�����Ɏ];�4�� ���6
܂�f	�Vr���ek�(�K�+d��K����9��l��|���WT$�SS���������҂��6��TTPH�r��ĸ4�՞���r���i�=�=����������������eS�����x\l(`j�d/������y��qm��o����BR��_{ԧ�� +������ ��B��r��	NU�t�ɇ��;�ns��P�2�5�K
@E���qF�7�0\W�MD{)*,��B�v�*��8"j목l����"��m������dD���^אָ}���m�=�
?<�Ω�]�|�ggg�`M����C��0�L��氃�@�f}��7��c�P�\k�o�<
9��.@tu?��_��Ǐ�����jK|�_� ����彳�����S��I(1�� \zQv������IM}��0�a��aQ�� /_���<~BbKfΪ���cC��^&��$�-���N:d���RS��Oԕ+W��?�'�H�U�p혪�FzvK�,�>V[� ����0�JT�wW����І#�[X@������ӟ�L��8N�BK����}�n�֋��S�a�&�Hz���ʕ��-C<��g_8*�-\>���
Ɔ��Hx" ?�����v2������y�N����HwW��.��)���~sU��ܰ�Í-��x��޾}�+�#tc,�:zԪ3wcf���y�r�Š��V��`o��o4�H[�͢��=|�PL5�	�8���K����t1U�� @�]\4=C �+F��T*L��ׇ�C�t� �pz�����V�_%�|	rG�6	�L'O��C�?F����H=�f&)�����3����U���ǚR���T@�ͽ��>;<2��'&&�`U�O[�*��	�=�S�Ҳ��Mj�T�{{��� �s0�+qa�P�T����������s���B�r���_���p� ���h�Y�`�0"+�;$_�:7���*��B��F!�**̗٩iy����O6),.d�{��IY�EyF�5��p7��e�ꪫ�Ş-��?��jT�uN<�z���ҥ����¡�B�����Y[��v����<H�j\h��tX�[5%��P+�`B]�!�F׷��	E����",Go(�aP�G��ò`Qh�An ;5���ܥk��~-��(�8=r��	Tt�,����$�b4*�f�؛oq��(��~����I��BCm=\n���^c]�o���>�>�o�����o����;�~ofzj��| S���VE�֬�i�i]	*��Q����u�,�8�U�s�ǀٶ0��m�v�~�]�Bs/�J�
�h�����^\THkBB#�큵���:!U:�rgɑϼ �-i���܁���̬?��LOF�}��&��6غ(q!�(��D4�0=��P��������zx�c�>��ɓ�ᛟ��_Dv�\.f��w�Cֳ({�OUk�� >"j�Eŝ�dK�wH�W���۫��r�A"%�-J|E�p����ok ��H�3S�4h��<����Y=�^8����[@a���#G�����),N��!ˋ	���w��bt^z�,Dv���^�v� �Yh"لTW������>�y�C�8�OdQ����/�Ö�Wn��Rl�ɂ��\\�H(L^6\� S<M'�ܭaH ��m4W�m�)����]�!jLj`���J�H{Z��)Ћ1�c���
�7yy�ᗒ��<.?с6<'vq`G#�A*P��>�ꩃt�ׯz�3�M��E\�Tlnyo ��a3����<� Φ.S��ϱ�Ji9��y��������@O�Ci�v��+�?��w��r����w9���E)Ƅ���:�a�@,H��J��!�/���vKO�&�z(�@n`��(=�G���<r�T��>k'�i�ItaY˳�Kpt�v������D0XÀ��\�혶��8��x/ǩ��+)�]��S�;Ρ9S$΂vl*��`�2��wt�K��&�f)LpB|%%`�N�+��j�o��n��q�ҧ
����7r����נޙJ%i0�k�<�е=�c�L\�[�O�r�1�E%<r�B`N����Y��@�	yݔ5��Z�(�x]��fo��k��<�5n�+�6aC)��px���Cf��c:Th-A����^���-yy�
J1|�X��(�����kWHU�JE�rP]R_S{����O��k�|wW�C�ak�+[��A^y������E"�����y�yE8����C�8#���=+.5�r������3�/���r%t ԝ[79��ݿP4�gmo0?�U*3��q� ����� &
�ǉQ���	���3�<<��Ό��<� (xlݾs��Xv�ձ�Ȥ��!�ò/F�^�E*��'�[�������*V��-�� ����]�_�����mrj汢¢���B_vvv�I^��������p�y��U\�p �䙘�ƹ�0wK_-g	���B��t9..�[�-(���"4�!���-�7o6�a�K1��EDVTR�h�W\�H��~�`B��x�x] �o�f)*)������S�[W(���Ay�ź����//��3��=���q ~*��|�����i����ڕHĻ�W[n~���v�Tg���dH�S�g�y9bc�����a���ZB����i�Ғb9s��U��A�-��3�4�5��"�}��\�g��k_{���;�OтՍ�U�|k׮=����a�PdR�>��Pr}n�w�����_z��W�jCc݉�;v<���q m(������|�
����������cK+�T��p8
�Ng6[�n�d��H)��$b  �IDAThn2�+	\N�4D���XX��!��C���~eC�*A1:��S"���C*��C2��.Z[ss#����Q,�-	�q--m<���R��8$>U��w����ryyٛU����[[�﫫[�������T�Z�	���ogMLL����
}х�X,֜H&�R�?+++�������э��/�����\	��v\>C�o���Ӑ���DXr��Rg����X��H��M���J�j���������A^T��Ņ�x<>���	�r�������T�/o�����)}@�����@e>1δs���ދD|���u�h�=+?wwnN~���N��e�D"_RN���t���{���\�"ٛB%�	Ij�$�_R�t1G�K ���_F+0x ���c�A#ѥ��幙ٕh4K�R�n�{���x";'g��� ��Wp����BNI�xuNs���w<���i���ۿr��z��JN(�L�-���V/,,6/,D�cK�x<^�_)L�$��T������qa�֙r&qW2�p�ەr�=�DBQx.�����^��$S�x<���W �rNV����ʲ��X��=�YY�hvV�LQqa���?\����g����<hfr�7}�� ���;������zV�a��Ғ7���H"�]L$�R���T*�r���d2�t�xa�qg
����7��$�w�r~�;���/Ap�Jd����"�k��PM��_����@��^�?�H����8�    IEND�B`�PK   �<�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   �<�Xp&�[  �  /   images/9d6941e9-aeed-488e-a8c8-e310224fd4af.png��g8���X1�v�J5���� ���"FkoJBQ�F��Ԉ]�f�Hmj5bרYT�Z--b^�Ž�����9��<�����wF���Fzz222FmM�+:\y)-�*r�=ʺ��6EF����N��jb|%r�j��?w���E:����K�z���m�%�#��v��]���y�$ {�:(�d���im7hƑ�y妝����&vq�nv:Y<�j-��*�TrbF�:zl�m.�j<�
ee��y�2�����f�����MG@���Ã9M4/C��2N�ϓB�O�2��b�9*��	|*.�I�آ5�9�����VHadeQw����a���6���#6����j�Қ����ǈM0\���k�ݡ�����ݴ��: H�΁lggg�a�����c��_RȪLJĪ�K�<[���m��OKfQ��ڦ�̍�KӒ5�n�v�Xy�e� �����O���m����f<��<��:���1�|�x�>�	$~�g^%�fǗQx�A#xK#�Ky�Sp��[�3�qFy?*".Ȝ�h`+ߏ���9{G`��4�?�HOڀOv��3���_p�:<��Ŕ#.0[^���?d�!ڎ�@����`l�-!�w�����ݭ�]o�����
%듨:M�����z�?��ܹ�M����;�,F3o*��^�:^*\$�I�44�g]��ЌA�
���7<�30X������h��	Y���*�&�7�s-�Rz��nЏTe���B�E�E*��ח!�U�� �b
8Bļ����BĤ���L�7n���
R7��
�.Ѯ�$�%�@�pێJ�"�,�i
C�:-@k,����`�m*䲫Iǥ477���2�]V����/�W�̰�b�\6^ą{��h�˞�CtY;�,+�g�5�T���<��)�Ճ�s�����5Y�����	���bt��8޸@�.
$���E=��𓲟�_�Q�g�tg�� ��;(�d�//N?%(z|�Q�۽o�u6oC"'�i�H�y�6"��5��u~���p�g��/弁ߖ$D��x/�kp��÷��0גo���M# G󉏃R����'�$����=�..����i w-��O��z]T�O|��7qg�Z=.�M��U2Qb��I�Oگ���������jo���P���Zo�9l^��}�A��}�`a���n~Sy��z�ߖ6�U��h/O���Ǿ���.�Id�"�5}-�w��^����#t��Ÿ���P��FLt��L�E9��9�C��AAZ�Ӛi�AV�b�'!8Q_�Ҟa��ի8::Z6�e�2�4�:�g��;���cc{{��.N��{���|]�I�'��J�����?LQV��$u�I�FU6�h�Dd��ɼn��<��L=�F!���B�zPN����鼚6�R�!ۭ�t�_a҃���42���9H"fƒ��V�[�Em�YAc/FIñ8�Z���N^�Z���K�%�UW侷s����Z��T�[�h&l�o�~`�6��Qg\�
��d_{N>�@�����r� F�3�����j,�������"аS�� sXK=����qs���)gbz:�ܨ��A�s��ݗ��V+�TX��W,���m5s����2��Wd��&����t������VZY��r�r��#�E��:�jΨ%E�Jq�3�����+�nW��<֧��l[��;4I#z�ޙ{��J�����!���N�h*t�qC%$u��~����x��{��# P�W���=GÇ�(�&�����n,�ѡZL@���|��H���S��h���y17�E�˒�/_�9��ta�nf���S�Xo�k�WS�%�uk#A���y+,�׍ �z�%����X���S��)�"���mr𳤛jB��ml�Y8�3�wW��"_'ɱGc�x��P��/��Qh,��;�7~GFm�W�=�3������caїԋ�E��i�#�� %�9��#3z��*�.?ol��U�������V��Oehث�X0f����=�������r=H��:�����Q��h�����Wwj�b��qUU�8�܅p��}�/0��1P�z>����=�Jm�z���~N$�,�<-k�б%*<�����3} Է9?��r�}�Q����}LG�aޝ[þ��a�Շ�A[��jd��"7v���k%1�k�2�t���8�e%� �	Ϯ��
����ƹ�K��gɅKr `��X��rC`R;�%�6ʡ �e�,ts�5f���p$�������Ya��Ga����l�.��W�+�k�Iڏ���R����e(|�aRۉ-��Ì
�F�&���}��B|�E�v�I����D���ADQ@�roc���/��g�E��#�ϖ����G��o%)�F/��k �r�1�Ya�jx�,|3փ�t�(A_!vX�O�k���ᑾ":����6ɣ>.�9>��g}�8�6� ���'R�U"�"ϧ8p.�|BU�Cp$�(u��9ea��K��j����2����H�{CGz�ʷ�������G��i�
շ�g�S�fU�h;5�}vN���&��V�q�?�׳���%ސ��e�d��Ld�M�~Sjm�y��'J��p���h�9��d��G����s�R��0�W^��#�p��p#���H��d�P@�X �-X� ����Lup�Vg�b/�������p���F���?�b�ǖ~�J�`Z�lp���t
��k�?*%I�
'�+�P�B�E0�mF�w9Q�T�����g��0��_'�/�n�\��&x{��rE��[)Ũ2W�FɏvJfα�l���he�R�M���ٺ.�:�6��;�����T�i�Ⱦa����8��b(�c�H��wõa���Nc������x���~�4����F�6�.���T.��/O^I��ՅaqE�����N 8g}��[�Wt�na[���g��-2���ـ*S�GҖ��=>� ٣�@�x���E�N����^Y!���7_��|�{Q�_�%����Gf���A+�o<>���EA(
ɝ��@Fv@e͡2���Z��\a�jYTC�b��epC�H�Se�gn�!�~+����>Y����X�*R�E����gda(Ta\QC��QɈg����l��06m�b0�c�9�[��]ܦ5H)��{��*�=.h��͖���JO!��6�1������;+q#����?�R�WJ�B1��p�]���,L����z��XG=�&��O�H�#�N���/%a9c����aw�-��F��g��'ݱh�=xC�g��2>��3ˡƦA�J�"J�
l�r����:��hl���)��5e�W���숕v�K��Ѯ�49�5�v⬑�S.F�]�ꈡ�M�y^��Vz�G C!�ch�����OR���X�cͦw���3�y��U�a��O?]�l#W`hhHNAa��OK������c.�\��RC�(�b�N?sY�q�I9�g�Y ���wl��g��~�S���e$��C�B+�{C\��ԖF7>t�L��m:77�f��(lH+n��㠦W�)�ך��K��̴a(Ư�������puw�ibl�%5�̻�H&Q�pkǽ/I�%��7�[h�p�|����t����o@�y�t^#![žʺw\��g��E�da	�|��&M��z��D��Pr���q5��6�#~Aa�T�X^�ޚAݮ}t�)M�Ͼ.-	��Վ�=r�-�,٩�f�ܿ�$�*��ާ$K*�Դ���]	��� ����ES��^���b�����pe���9f����u�4?�U+Ӆ�O#]��Oh/�k`�����c��ن蓓�f��ߎ���*Ǹ1M圐�����Uuu��N������^�̾?<<�	�XQ��"̶�~+v����999�+던�׉�Y��rV�lo�Ajfr���o�V�r�v�+,)��͛�h�g�I��י����6��1 ؍��rJ/..V0��V��?��⿗ ��-�p{�XXg]����Hnb��T�&��[�%���Dpr@̗��H�CR���ÊN�n1�,�6"�l}���z���?s��
�Ѧ�2��D�
a`�>܉�������z)���*E?u�p'uA��S�C�6b�s����§N�мvM�DI�bXT8����-���m�WG�?~���_�xIGC-F��c� �F:������L����=w��yH?���\R<��np*�u�>뜝���������Ɵ{�wD��"��L'�m��]���#W�g�������G8��[N?B��q!�/O�衉J�!�s�����
=��~�Дq��b_���z�e6�?8��p���
&�_I�b#O$���
�'���CJCqx,H�V���C)EK^ҽP�LL!�o=e�
:��H��ޤ�WB���sSg�њ,�_м>/!�Mح"�2-}�*�M�PK   ���X�V�4sE  iE  /   images/b14b5b74-4377-48a9-90a5-00abeaecdcc5.png *@տ�PNG

   IHDR   f   �   ,M�{   sRGB ���    IDATx^�}�]e��s��u��^2�tB�ЋA�eQ��*º�bQPi�uu]v���"��� !� !$!�L��~���~�9���3)#/�0�{����������r�7�U��<o���6�Sļ-1 �x1'�"$Y�),[f������T�x�'a�a�nԴs��*폤2�Dv<Y6��,ɧrqЁ�d���eeL���p�h���t"Z�D#����f�g����?����<!�s�ݞ��͏.ʌ�-�M�7�F��v��i�u#��ͼ�����DH.��Ù$�eEOI�:)iڐ	wF�{�p�����W)���7HoX`�vl��}��������UɁ�S�ɱz'5Q�O�8�lHp��J� � <� ��f�.<�V�`\�&)�顤��#ZQ�-\R�l���xIUWQ�~�l���?�70^�梁��ʁ]���t��3�նԘ�����:lU�\��Ep!�D�n�%h z.�y����\ׅ �E�$1�L׃�I�X>�1i�U��D���y�Yt����$@o`��zWwoc�Η�h�ybn��I�NT�='.�9v�gCU<h�Y B�k�`6�	���%� ��(�� �ua�6,�0\�Ux��Z�6a
�O�=)�{��n�3'~����yC ӽ������V�67�[���h{|�B5ґ�k &	�"Dׂed�
6��
Y��dO��I���E��T�'
���'��$r�<��\����฀#H�ۘϻÞkQJj�V�����5=Ǯ�<7� �C�!����k�<���:w���L.S�	��"!y�� �.�6\�ↄ$E���
�\Ra|��L����1�E@����>BG�s8� @�z�6ٮ��dlq2+h�99�)T�pky��|���s�?o�uO�3K_z����{[N6��B���%1�c����g���p/KT��Z�U]��tw h������[x�-��$@��҇��]�c�X�`�������I)tG�d�=����Zs�ϭ��?�΍+j�ut۳?jvo?&b��UE@H�J6Tх$Xp,�I�$�,C�����:��v_Tآ3�! |�&#��s�D8�W�I� �����J�ݓ������?5.�}��?�Lp�������m��S^���tW��J/���tM���bXD�g�q-�l�K̻q/ �
��A}��ux_|��H*�3��0��$J�C﻾c H�w�8��T�밿��\�P�1S����P�E��_Z��?4�zN�����'9�g���c�+bNN-�,���q`dlfOdY��(lW�M��L+A`�$E$�O�|ﭐ@�/Pg�3dg�i�����!���a��s�=+ϵ!�-)�9����;i)m)򓒕k���֟'���0=O�V�����k���|��Yw�4�""�=.lH���`�5�(����|Z4zI�E��W�֎Î��rI1UEƝ� i���`$K�$�x�����\�g�;Ǽ���,�!���s�C��i8�o�}�@�3'�t<~[e�KO]��ܦ����BQ'���0�K��T�(��TZ�kC�Tئ	�l�%Tʪ1Xg��cv���c�[d����$1~F�/2�Ì��c�$��-��x*Q�`�K.��D�'°���{~B����n�#����t`&w�W���M�m~��O�z�,+W�j���"��04=�5��eZ,�eB���E *\�1W��dL�r��Y�U��t�
}���n��ȼ0��ˤ�>kZr�OT�@@ư!k:<WD�4 	"�r���a���*�[z�߿���{��;_����Ζ�BvQ�A�*�PS��6h<��pY"�����A,��+��'I,�b���s��sS$p�/���s�)O- ���Ԛ H>I���� >=r����tN�n&��ޱ6���Gu+�{䴯��!Ю���A����9f�{�3��|��WT	axK"""�Fx��R#�c�n�zP΋�`;��+E�,e�UR��\*����������?#A )q\�/>��c�������s���D	H�	��� #)#�����Xџ�e��x����O\|)�߳��Ϸo����M�}=���{��~Ewm�e��@��L7m�Si�����6��)"�(��m#�e^	WF��{t:mo����>PZ{m?��sq`IJi"oo|C�����f�*�.r=9k�U�pSӱ'���K�׿?�zP$ft�S��w}hצ��
�ǫ5#.4~�B�R-*�'���#��W!�4)����|��)�x��%(�-,�I^�o��Br�J��گ�09e�I ���3s�ɶ	ț�l��.�m�3Zlk>Z��e��y��|a|_�9(���'G6o��{c�/Sa2��R�"e��]@�!(�-q� 00��T���[�Y�;�"����s��~n�I�(���)���,S/f[Xj���Wk,vb���c�
����0,OB&���pdc�<�5�<[����?�}/,[�~�J���-�U����e][7}LI�
�",��!���T�\D�?\H��<!I�{)ӃE�ߢ�h����-a��;DV ��9��%	rd�@ʸgGbx}�Gcꊤ��[Re\J(4m�-!�Kã��$"��ǭ�P��4u���p����P`(1��s�_׵u�7쁖#JDQ8P���J2{��It!���łE���-&_�@�O庸��#��Bs�#O.p�}�[Ej��cDr�|�G?��r;���mT aL*�~�甹��Q�d�cBV�-3�2�fM�p�X��'���5\12[p(0�]T=��]�lۺ>j$�J5��@�n\e�c���� 
ONR��mMj�2Я0��؞�#ENI�^P)a	~R;��L�-�EF���a��U���� ҵp�7�F�I��xlK@�v )�c[�s6$� �c�d&Z�T���Γ>�YX����0ޖ-J���#����~���U17��k!")P"%"%RK. 9�HF_�"�0�$lG�b11�c���W1���*$�D��腭;��X<Cq�M�7��d%��D
�+|����-��:���/��;�B��]�l�I�B֖1`I����=���a�9��;CL�)��|��8�lK��?;��ɋ���°��j[�h!%�&/�le�%�:��1��$��$,X���[@���
��"z�^�`8�T�z�
����X�����sK��f���H&IP����Uf`�(M$R�g��R�HB�qa�-�&��:��1G��)�-�G�v�)��<)�_�K3x0���������_d�d��{&$r���+$^!U�c7�bx��M�T�7�b`�}+�d��3��)��d�W�2�T�|�������A��T�ȓ����ç�0�5%Ẻv}g���լ	x	)O�e��t!Q��t��$�)ݩ������e74w��09p�oH�<����u�*�LUĜ�Ni{�hE|i`|�@]P:E���0{A��w*]I -S-�vw�4pC�})��	,��]�l�-~b��d�p�L[^V��!'�<��)�"ï�_mn�Xc{�JvR���5�/�Gޑ`DJ�톶��>v���|fۜ3��wM{�z�;�<|V����M&)`��b�pI!¢|�/�js�����N��$e���n!�%��=C�N��+KHf*�$(¦�X�ҁ��P!@�n,������d��AH``8R��1!w�ua樠ǁqE� �aAș�mi!�>[�������w�_����L��oUF��=w����͏|?ߵcI��D�ν*����s�"
.[��%A�W$����d�0ڶ���I��d��'F/f����2?	Y�\mn�8��( ﺰX�M�"лRCy�t�(�Z�n��ц�W&`�A.��A��c�,�F�iK�ej�T	H$$�Rr�/=�7M������^�57��<T���w^:���ψ#�E�0��(`
.\E�KYc�R���T�Q�90��E�B�c�6yP���'(��i�rȪ��
��t��M���
Y�)JLZ��i�dL$�,#��uH��lz��c&��)onZn��4�IJ���>e�e���X��b�O�3� 3/!�0P�`C���Z��럙`����=���������X�P��+$*~�2L2�䶲��À�IjHb(�� 
 %�
`�[�R��PcŘ̻͠g`��id@� �1�7��HP�ː%	�-a�p0�t0�ͣ�o�E�T��@M����(/� �H�B��^���\�����av���5���vf{̜�R0jx��v%[��]��[��c_���_���<q�����n޶*�Umh*��T�$��������������eȑY��ɛ�<jD��j����:��-�1�< �>�ꊀ#K��FGYT�#)�՟Ķ^O�A6�h�8&P�͋bՂ�k(�RP����B�Ar��@8��/O�E�[ǁC�'�$Ǥ��b_elY)<T���?�}���Y����<�0Ûb]�?��Ǯ�:ګ��@�(�7�&TN�B��(HU��������K*S1�g��Tlt�ضQ�n��@A����`x0���r�5	�YP��'��M;���C�8�(��"&'\�� �E�q�c8uU��I�N�]#�AQ��KLP�	�`�Tʛ�{�����h�u�T��p�w�dc�7�=�_�������Sg����*�=z���;���<��IdՀ(Y,�Dޒ"�S��2�����rC�j'�U JI�2��nWÃ�S��&c`^��#�T��� �Cx��!lip��*�_و�¯o�� a8�e	JD������<��7 �}[#V���Y�C�p�'e�h_�L�+d I@$��D�D09���#"e�ZQ�⢓�媆w�� �v�f���o�����F��w���B��`R�B���󪤳���t�1��Ea��G�eA&�N��,"���<ޒ�#� !X��k�FABG��86��ş� ���k"�8�~��C@E	��3+P[�"�F�����C�x��Հ��nr*eD4'�0�^�g���pwpX�K,������3⨉�,�#b�����V�Y��U���+a���I{�/`F���e����y���%QɅ#f�g�)9��aʻ0ϊ��(�'�@�~C������1��!`Ҵ�=�GK���PSQ����=�66��ݛF��=G�8zI	"����փ����5ub/���m� z�,,>pZ5��LĽ4��<֢�ƽ���A��3��s���LI����yi�0[��֣�xߗ^���0�O�x�3����H��R��3pe������+��)��Qv�%�x�]�`�����f"o�X�9?�AD
C�`3ƨ�Ʈ,6�؇^�Q�Y%��(�"�L�0$�uq�@���c����2x��,(�]� x�I���LD�+�_���wT�8��ӥ���r���WC� �S��J�6N.�R�B٢{�;��s~�kٙ}��n�z�9~����qx�wi�  �Pז�2�,%�yPe��I�HB���K�%\Q�-(�0�!�1��9�f
!�{D�!�j��h7tܽc��N$�,����8�)�"1�X�C�#��Etf<��b��hi6P�y��s��%��J��',o,�9�3��.5I��m%�d^�s����<�C
Q/����.�Tٱl98�to�ly�=m��#c=�E���/�h�ܳQu*�H�0�$3w��$(����H���gN�3�H8���p^��c9<ߗ�c�$3@� ��6��ư�T�2��q!�qL ��H)m�C����(��'���2�U�P�:;��|
+-x�������S7$� ��8��UM)�F6��@HjD�m�, c�H�Q�k��{�|�d�E�
0c��l����6�����p$bX�(Ѩ��T��L�ǣy��lr.)���j��Da���$C�b,���<\ׄ�J�"�h��tk�w��3T '.�[Z����́����H[��5<=l��ݽ�q�䀕�N\R���2
�$�(�Ep��
LVCu��3-;�WWN ��z�������=�b�Ԍ�q��|���g_���3>�� C˶�����'n�bq~<3]�dY�E#cϵ$��A� C�~0wY Ec����<T-Q�����Y��5g
�BU�1���$���A�P�]��e	�+��Z�+C�4`K*zRvy�kK� =,�NZZ��:ʣt/ǁ��o�R/��O��X� �͏���O��ԕ�}`,[�D�Ř��Mk�9��g}�L�凊w=u����r;�[9����b\Jz���Q3�˘�̬$���e���d�k1`!��A�E�����ї�pϓ�x�eCi �Y^���ceQ�yUv^@���Q�Y�v�q�(�z ]�7�X��k"����$ �$�|q���v�u��VR��J�Ⱥ`��Ĥ�u�d1�7"�Č0��#՛V�����A�/�;6����ﹼ�ͅ��R{��AP�t�#� j�:*�ĸD��4X��� k*L)�޴���<�u mC6
�/nĊ�
Th��c(���%7�<�3�G�Sش5ÊW�kKp����*�{e�D*0ϊ(�/���nZh^ƶ��4\b�6`�K����G�GGet��(�LJ�3j�N:Z�q�9~b�;�*����������g��|���%<���z&��D;��IKVǗ^���g^��j"��l��fY�`NƋ#
�z�;���,�/����T7��;
)3���T!#i�wK���&��+���
Dj>�I�*�\X�"���ڌ���Ęs""�5^#��	�@%<�$�;0t����T1`8"Se�v�J�?���}r�9��?����Go�x�{�+u2�Od�ߑ<8�3F�ͣX��ʙ�P�٧�r`�`�,��t�a�Z��k�Ľ/�q� �cI���p�ht6� )��X}X#&�>ԁ燩H���@D��XV����
Y�'o��|4F`�����U+�95�X1$M>O��/��j�*���0,�9������֜��Oמ��.��������O���b3YV�Q�D���^��,[���l�CD9���@%^�ĺ�H���2��a���ܷ���/�M�lA|�����Q�X.c٢L�Rx��Q��r<�۔�eE7JR�@B����aEe	ņ���F�n5�9Rm�i�:Lj�'��>s�d�nO�.�A��<�70��
rV���V�u���.:H�[�_z�잍��O";Zw��"APD^��j%݀M �]vTJ���L�O-RX�\���,p�Q��͑��j�5�Eޡ
��=#����,*��,�ԗ"��IN$1a��Z�IVYvA�T�r�5���QT����tPV܁"K�²��ض�v���9�Jc��g�L��Tee�`�򦀤) ���Ŋ�]}��W���5�L��{B�_�rr�#�!4ٽ(!�H�Tv�y�">"�(<+���&�����J��c�*H�)0=	�IeZ�Ia ���%#�R�Fq�M�X|C��,��)aV����ɖQ'��ɵ�����hR\��i��,<3��h��;�5�� !j�"��BQ�{f$y��DY�D�S��Đ��r�I��Z�[y����`�+F#���g|�k�#�|��}�vG���;j����i8ٱ�@0S(�^!���Bkpi�L.���ș�%�����"cÓF&dM*z����:��\@��3C4�gGY�P4jW`+�u`�)�Q�����@�l�<ZHr��Q1�K
�2��:����]��ef���Ez҃#��<`�R1~ÓG%p�m�t�XV���,^vҏ�r��˖�{͎��������돿��<-楥�h���4�%&`�E�%,�J��ψd�,V0�;i��+��n�"5�Rۤ��V=�$������my^�F�@$B� ��"��J"[G��<�~Ò���    IDATE�F�άD�!E!��XT_���ĩ�dщ��˔��K��%��$���D��$V
��T>GcԔ�p�KuG�~��� �6�o��}���������E�t�H~�w��L6q����r� #/I��J˒ˀdگ�i��Y��0����HaHJ���0�����;���E��D"F"Le2�f�l���s�=��,�@��D�#%"(��#�z�*
���U�v��':+�2��ef�>��d#03E�MM�H�sȉƝPV�]��·����w|�u�e�E�[o�������㥺�g!]1�(Q�d�:��%�<��\�������<�,�P�@����d��j�d���E�@��H�T�YU��:�H���e1W���U/hϠ�Ԝ�|��h��wĉ���:��Y�~�K��=�o�6���Jl���h�
9 Y�Ÿ+!��G
qǒ�/�r��n+�~��G���g$���/99�0��(7���(t�y]����b�ƒ����7"g��F�3��t��Y]��}@�ըO�"���<�f|�'+`�!.�ߘD;�u�Q���:�r�3�YC��yl�yi��D�NTYs�e{�a��n,=#yl��EUM���4�� ����!*�%�v��<�k+���ۅ�s^w��~C�������{���ڃ��^F����V1��0:� 2`hAh�S�%�R��3	�b����G�ar�H%	P��N)�K�"����˜�E��0F2�-�)F�m ��U,���|uƏ��d~�?��'�]']���\f���7`X�������0D� �nу�z����������o`F7��f�c�^���q~�K�t��%>)��0gK�G��f��q��&4�#~?#�?1��?���#l�h{�Ep`;7�
�g���^��fX����A�Lg�M�����>��rj��rYR�r_4W@R8ɂ�f
V%>����fy�K��{��XtH	*l1]|ďO:�j�}�gn�y��x���g|׳ת��z��!Vٮ��I!

���]e�F �r ϡ�Ae]]~;�	�t�D�]�<ک���{&Y|�:����*7�+Luq����Yd�x�|$#�z��@��ؙ���i��Q=?�P�܀�0�d����r<
dl�����5����\��mg�/,~WjN���ŭ�_=�m�1޵6��ňL�]dI�9o�R2�*3��~�9�� X9�;Ѝv)��t�m�l�Yfg
Z|��8C�+ ������
�" �I�?��@o�{saAcy���r�#'�3���qH�x�s0L��X���%b��P዇�yޥK�������x��������j�k�;%�@23Pe4�L&�7��L�u���t�#�}��3]Ϻ$?_��۴��H<���|�d�g��X�&�b�G���t�E��d9<_�ꋷZp�N����m8+	�aZ�ꚯ�H}�H�<��
F��`|�;;�ܯV�t��zc��Љ���e����?0����KU�A�%ɷb��U4Y�.�8�"y�ʸ��S��6N��J�9���"k�@��^���{CA۷eQ���T�0��Ž&��A����������Scs3�I~�!I7���cIa�24�1�Aa$²�Y��SF�N�J�/{�9W�Xw�c¼u������[���G�=u��	��U;�J���l@/%s��+��V^��$@��!W��Kr�(��u���8�%�~U1�َ&��~z&�`c��*��L�6����R=��N��,:m�W�����mR���'�L�t�μ3�t�謾��1D����ws��\}�̥倩2&5w}�z�#w~6��P��˞�5�2U�9W_QZ�%)����lv9`���%���9���R����(��l(�$
:>���=�k5��?��L�/�IVn��^P^��Al0�OT��t�E�m�����`�R�l����U']{�;�yh����İx񷑗��󉩎ߒ��i<	E�2h�"yO�-���ǻ�X��_k��s�+��K��4{�_2 �?�	���nq�>�6$���'����+�tC��@A�^3;5*pD�����6�E��"����vѭ���oן}鬇00`��[~wiS߳�|����=+)�&'���hG����)V�+Z���"ٔ>��1O�Ʀ��XA��T\2}���o���'�BM�A�X0�! ��L����71Ɔ�2��x�a�pe����[��y��3߽i��r@Uۑ�Y��Ο\bP�khD�&h�~NX�������ƣ�3WML��[%��d3x�HS�]��=m>L�Ŧ�y���C�!�|�Y�pU95%C ���^��W֒�O=gA0!�����	�C��7�M-?��u'��_�O�̌Z�^�P��1���������W8�+®���;�ԙD7l1�Jv�l�X�A��I��O��~��MSb]�~�ej�o��;	���(����k�z�z��x�_ʎRǧ-�Cl��g(�O�G*�d	جǈy�v��[��G�c׿n�����,0���o���V���"ٱcÎ���sah:,���|��@���T'2�L�ﭛ�b
$�/��N�� �_����D&�p>K0�cX��|;>]�}���H��0מ��&7�`��H�@J��󉚍�NY��s���L���Խ�֛�}�Ɩlx�+��=/]�M��g�(&\�CWv4���B�N��3'm��-Ϋ��X->�����z-`�c���H^��G�?�)P�0�~4m6s��7�P�q�yIE�O�\�����������<#�J��;b/���y�/���..���(Z�eF##Ȟ��X*D&1fc��/�p7�~���� [�t�t�^5�rz��t`��2�¡��ۮ��8�o/K3�w�\i*�Y��� È��sՙ����M�vs�i���{��
i��	�(��(���D�h3[C&E���/��H,)�:�h�������K���^|��s�M�z@��GIMGd !�.:7�SKbi��-~��h���xNĀۦ6��v����PŊ�h��A�1Cn��n��T���G͉5	�Ê�2�dx�/1��
=���V�4=7��LM��>{�'o�Q�S�| O�Y�g�������m>�wڋ������~�q�H.J���%��F�g�a�J\�y�9�^d�Ը�˫>���Jg�I>h�PS�_�_�����'{O+��x�N��"r�S�4
U*I�X�OJ�4�dn�QVXSR4}�<>��>�v�h��Rƥ��-�cK��� ����ħ�� ��n�. �d |�%e�=I#��0��!��1�;��nXz�ſ+;r���[����ؘ�ｾat��;#�k����"��$�LaM�J3�3y�46J��J:ˍe��}��"�6���,OE�ڴ���g���N� �$��+��`�m��_�$&�ό6>=]��X&K�R��DQ'#|H�d�Jn1g�rrD��2�
.L��	�q���Q3���=xع~q��W�	Eb&�����هϙhy�J-;�4�ea� g��6��n΁G(0�'!���)4�WB�v>1ȍQ͟X0�6(ͫQ��()��9ұ~[�χf���M�H�f�&IaDq�~c�R���.=d�$��$pM���0�L>$[�R5S���q�M��IY�e����q�h��S�s�N�o_�~�)�Q��v�Pw����Z���l9>!�"�|� �M���E�Bu;r���3E�uDQ
2a�:͂��_�%E�L��a�e�<S�m�l�����X�?~k:04��-���d4�y%���$��#b8���Y��eJH��T��g�eA�
"$
����W-F��D�èI��8�g�'����?��S0��>{[�K���Zk��\�,(� :ua�B�a���B��k��fMe m
=)��ϋ*ZB0�R�v�U�-�*u��ұ�Is�*��	c���!J�TF0��*O=G�\[Β��Z�oZ���hy#�<{fQ�d�I��Jɪ��$I�@�zȦ.J�h�y@F�u&���Yɤ����b���Ǟ����}z_6�>K�`�?����O��aalaa�Da��X��ő����=YCt'����k�)(��)LD�T�p<�N6���fgӇ�V�^r�B	VX�%��2{�K�S'�i2�r�q�B�a{gW�y5�I����-#yd�9�f�>��$���lb+y��IJƆ��a���Q-�j��+2J$;W��f"&�=^��9�� E`�9d�s�L�0���������g��Y8��Y��g`Z���a;7����Ӫ�VX&"!ˆh��(Cd�91ɜ���6K+�=R��w��V�s��j��oG�[��&F���񡣽|z>�t�k��'S"yVL��HH5�I��f��n'�#���1��K�}��k��9��0Ĝsr��%b`�լe#����#��Ñ�Z��S/�$J��1;=�$=��v13|d\p�� UVX�5�7z��y���ȦEd�qG�Y�p��|��_��q�?��}�"�=�m�������DCU��؁���;<HԨ:�i�qX��ԚQ�6D��i�cv/8�S��T	}�j��;���p,3�[ce'Vxfj��Y��P���8!Ѷu�FDT�yꞃ�K�3`h�����>�p<� Ĭy"����9R��*�Jq�%��Ɋ���>ů���U�Y<ֽ}y�����Co�VM\��xh\N>f�S,Xixy�d9��KY|�����7�Z7�G�0�ol��ؽ�|驳VV�jq܆�"�fY�]�4x�F&�f����ak���ӛ�e3���h����D�h,���'Ɩ{�T�h�㖫�X����!�L5uE�(����$�61k4-�y�e9N2g;�.�'�j��D�c5ڵX��+˙Ҽ��K.�?��G��ټm�x��K��к�m4K�� v� 13���";�a$ˍG��=z�G��=�=��5�̖�\y����*N�-[XE���A��#��5e�'<���HN,�k�µ7,]y�����~#����w^�Fs��s��95S��4c�eGmӈ���&5���QJ�+��(����*�0ji�tHIX�������y]?c�]Ϟ{���{l�n{�Q3yn�1�D�&QT��r�У�4�0:�`L(�Z�����<��Gg�:��oK��?��ݙ�'�sG�ʊ).�CVy[�,��LYw��P�|��՗W����cΓWw�r�Ǥ48^ �X�w��{qg���l��]��&����&����s����`��K�\C�=j8W� ��Ar12��p��W�}��ˏ~׌�ͳ�/<~ۍ�:��_Us"!��� KQT�j�0i�`�����'�wY���/?џ�c���fs������N)�HD��S�,�!����3�N�j\��K._�:}���a��>uG��������o*WEʰɜ�t=]�!KD�����E[��}ݒKJ7	���L��*��׷����x�k��q�;�D3�5�M�0�L������Ol�	6��Rf��3�T<����SGv^�X,��N�D�s�G'm���΂��?[p�y7�~l��f<.��������N�K��;��x��\�(@��|��+>���^s~�~I��){���p��^Z�"�(����tLL:�p&����;�+M��ug?��x�5��ۇ�~��o)��Sti@��E^�cȍb�)|�����h��n'�>�14��?�xq���/�����bz��I�ch�DN(z�l���i<����?3f�����|ߋ���U��A,\�"r#�˟=꽗|��m�����}��'�^,��֔�0�)�c ��V���EG�uM���y�;೹��[�v��և�˛�~LB2�
!�a!�jO/��>����<UF����Υ'��z��oIS%�LLf���ƣN�NӪ�~�8����f!�h�f��R���W�x��Q1&M:�l�^���{jŹ������gzݳ6�t⍿�fE���7xc{�ZZ�ɢg`8#c�o9���?S��k����U��H��_��o�߮-4��G�@.�b��&���/zׇ?[uĻ;gz��̋����oۣ_mR���\I+�r�Uw��^^��]�3��7�qO|�����/�o�񕶊t2�![�^{���x���KΛ�ò�	���͡�M��c�#ߌz#�4]��l��,���θU��٣8�L�>�k������w}��'/���0Ҷ7h�ϭ8���j�~߃�����ý�����u�������;�ye�*�?V�x����ѭ3����1��C�^�m�}ח���m�f^�]���}�|��3v�im����۞�:�� g���nlX��GM���qOo5p<o�ܹm׻�n~�1[*$r�^Tr˒��tEI�kO[:`���ݽ��|f���a奂��J�k6ΛE;�[���7����KX&�j�VR��%��?(T���o�%���Ծkl����EOP�/]*?�zx+�1�����l��Ap��U=�VP^�񲪵O��Q����e�rf�L6��z��+˗��C�����F~a�c4=�ZTR�����[f�!����v�0�ߓ����r9'�|�0>�������2�����r����͆�_��ZKYq�Euu������30��ñ��OF�l.oD±TWV���x�>3�g{�o�㻺^�?42z�i��t]o)-.����%���Z���������/��ɏ�|>*�Y]M�w��C*����޹`hd�V�0�u�����?jk�7���_m���r93������[�x͌���^�����݋�n1-s���]�%����Ztל�� �|>o��ߔ���2V��C8���?��ٿc�� Se�4M�-.-�Dm�Bf��Yޯ ����i�>��e�p(~sY}��ˣ�3&���Q?�5�󰑁�?0���}��f�_������f��\����[^Z����y���F]��\Ww��ÇG��`��R]�K��?Q]�D�̊����|�=14��t.���0�b4�sYi�5��u}����ڱ��{V���2�E��%J?U[��/�@�tg��g`FGG���e������ﮪ�����j������G0�#��7s	ILQ�����ŷ	�@O#��k���8f|r�l6y�a�C�p��ꪚ+
+_sf����Mz`G��#FGG~g\�%
�/k�]L�w����m�0���S��5�i�����U�՗��WS�(����I�� 344���0�%`�H$�@5�j���7�P��ew���zdx�w��T�Pa�����E��)0����S�ɫM3&UVYQyyqq�������߽vxh跦i,fƿ���aV��}Ve$1���E����h��޲���JKKi�����CCC�	�I��z������řLꋆ�E���J�//++;�㘁棆~c2w94�((�|C��?�-0��K�'��7�zA�ஒ��+�ȿg`������v]w��j0�S3���Lf�������;j��>�U�5���f(QXD�����8f`` �L��[6��B.��ⱂ��UW!v�'1������c;�5M,L��f�-s�0���E���������P[�x�j��m�����[��w��v�%���&J/k�]Hq����<�;�ښ��dz�L6�D��k���LOO�ʾ���ڶM�_����yu�(�U��>�˞׮����7��Z:�
0�_�:�%f����n氐�+��Lâ�g*q�q�����7���z:�E��[6�]}�W0����t���ƶ���),*���n�s���N�ƾ�JO0nj������-���z��׾����7�c�i��D��3����z�{���)1��;69�u�1�H�-���^�O`�wt��Z���vz�\�1<�We��_c���j����Pgɐ�t���H+T5�UXX�����ΩĴv�z����W`���]�O�i_���~a��h�Eş�_���9�]ok3�O�\�OU�w�{{�u�t�: &QX􉦆ŏ�50�'?��G(�	���4�]w�{eLgO�M� �P�Jd  IDAT������M��@bB�h�֦y�������.��%`���0`Z;��r&���b�U44\}���C-M]�]7��t�(,�DSC�\�2Okk�u�xr���X,Vpgռ�/T����=�{:�oi��*�E�%��s���s��ã�e��H4~Oue啇:�op������W�����M$�?��4��r��Ԏ��3G��m��H8z_Mu��JK�r#�fc�_���_6��{fs:v"�����������"b��V�~����w��V:~p�k~k��_2���>�9Mɨm]{N�n���#��k�(.��ѳ��J`L���������_���$J/_и����~ILg�S�G�k���H$�pYM�g���i���P낖��_����S���s�]V;;��><2�=&�o(�+�lUa�!M�n]����S��ʮhjZt�5.y��tt��}d��{��+�Dc�U�V^^Y9��.��?/�b��%�\U0=���e�����#[���,������}����t|�pۢ�ֶ�3�	���0s�QF�ֶ礱��2`��U�U������)�oQ`��(Q�����s�Q�y����r��hߏ3_�Ğ����Lyy]�[i�g{/��m�Z���8,H�\�4��1�%�I���G����0r5�h|SMe��ee�-������CC��:��8�1���|��q1����G#��ێ�������Fc�5�uW��Nt��ji��e;'��:���\3>cb�M����lY50��+���Ƣ�ǫ*�>w�������ͭ�7ؖ}����D����-�Y�Y�rٟ S��kY9���K���E#�G��j�<ԍ?����G�圤(�D����M��$���rf����Ζ�Cý����h4�pUE�uwyh��������,������ll,�� T�ռ2O��lY98L���F�U�U~�P0`L�&�I�|{����%0RWW�����_Z�Q�F�,���?��n�hn����')��,L}g��ҟ
BYz&*�@Pd����U�����|U${�����C�Ɛ�t������)��L�|����s	���׺������eTFñ��j�9Խ2r�;[Z�g��:EQ&���75��v.�Q��������i��c����U���|��aO[�wl�>�SX���yK~?����׺v��秦�/�E�)/��֡nc����[Z��bZ�9��N&J�<�2�(��8��TWW�����o�V�2��\UQqcyy�!=k 5Pֽ���M��UU'���45Fe��.�?<T��E�H�    IEND�B`�PK   ĺ�Xm.���  ?�  /   images/b2b92e47-5c05-492f-ba01-c47f59068786.png q@���PNG

   IHDR  
   �   Ks3�   sRGB ���    IDATx^�i�d�uvޖ{fU���t�Lς!A���hRR���e���-�vPG��I)¦�e��EKa��-��	P�pؒi9H�d�� ���p�Y���R�T�^k�/�{��;����]���%wFtWU������|g��<|=���3�p>`��3�p�����x4C?8g@��E�p����C���)zx��x8���x8g�g�!P|�=<��<���@�p<���3��3�(>p��p��C��YEQAx�(�H��!��{|_DB����q��vcc#8|8+D��w�w��a;�}�֭�(
{O�(
#��<WQ9>��x�0�z�^�h�H���>�*�a��z���{"{�Z��·߳,�j�Zj����<�y`0=��؅��	��y�&�#��˙w߶��'�c�����wܘ�y�q6������-��(
,h'��H5��V�sr��(����jL��aV	�,.�8�,��:��0��<� �yNᎢ(�?��d�,��q<��N��QQ�y�$�<S��0���,�"�x�$�2@���y����eE�E�e
PI��</B�5���E�a����4M� Ȣ(�E>��"AD��E�GE!�8��AM�	q����"�� "�$	Q�0�<O1�Y�i�<c#�7Y'q�e��<�L&��,��H*A��8�p/"�L&��8��<�'Y���Fc�X] tpLZ�ׁ]�~����@��>O����8����1�� EQ�����^�E��x<�FQ\�4
�0�̂�VH\�YQ�����V��l/N
��L�EQT�8�I^�&y��g�V���0�</�X�y^ < �d��A ��&/ĭ���!�V$��<�"�3hj��(˲��18�'I�i:��Ss�iJ6�L&z�XǑ�y!Y6��$���0��5�d� �G�8�̄AH�!��q�q��(�R��@*��gyF�d��ؓ~�($�T*�c�f�d�U�$��"�nR�V�,�ܒ� ��(����g�#�9���d�v+�dP�L�(���aQ�0�q� i��a��$�GQ��1�@⢣j���ߋ� � 5�8�1q�"���Hݽ�E����E��q��X ��$IҬ����5����lY���Ȫ���lH����%��^ь�J=��V���,�VF���<���lE$O�<���OӴ�eYUr���)��$���72a�I��q\����,�dYAP ���I�;�������Q�ӂ� ��I3��Z��wը!�c  x�����?/��k�8���?�H�$�9m�8/~�q�o��,;����#=�������j5�m4�x<�wn��$ɾ{�{����1\��C�%�tAEdgʔ�b<�&����D�DqZ�E.Q@T�"0�0��x�� �ʋ �e�� ����B�<!��w�8�.�b��DqЏ�x7�q�$J��0LSe7E��0�ð^�Y6�V� �q�e�t.�,���`��';�W��� (���N'ҕ�2K��SAQ)��d��+ �4M��tT/&YuRL�4E��d2T�>Is
b�V�(J�Z�K�ѐj���A���n�e���-~r�0��m@��h!d�)p� ,�&�a�î�\<��������PA��̀�d�a f׶�!;I� �;,�6����}p���y�q�w	D�γ\�þ������(���{<>���k�߱1H��v�9V���I�3���n2s�$�T*�3�2`�`�'�Q��8��A;�t���v'��(�F�V�=�Z�ZR��Q��y��a8
�`��R� Xƣv{����`�;z� �(n޼	&��5�:����{�|�p8<1��tԚ���H����d�1�k��%�D�8)ta��
\I\���EI��4�-i�ZR�5x�=^��F�0�m���R��cNk��}�	�����	$>3���� ��	�1�ϘM^�|�a��b r���^E�������@��@��ӿ/���@��������׶95���v~G��(`b���@����gN�\���r�|������>�3\www���~�U�O$����I��A�nRM֢0�Eю�͢w� ؉��T*��Zms���	�@'���G��766�<?�K{Om�l��[��g{g�ذ?��1�����; 	#I�P�@�N:)%��ք1��V���URo�dyiU��"�f[Z� @�b�Ŧ	�Lpn,j=�δ҄ ݗ",��A�csf�-0\�^>P(h)�����Υ ����R��9� |��� ����Rg2_#����#_��0 �� րǄ�L����(j���vov�f��0V���s��
f���k%x��qL�3�p3�l|>��������]�7���5���K�$Y�$�8�YQ���H� U�x�R�_k��_K*��U��|�^��n�7�(M�?t��s������G��v�k�������;��mmm5���z}���jFP�ҪU	p&QHM0��K!aJ�¨7Ro��
���ȡ�G���G�ӞW{���MS��$Qe���f�iV[&J}Acuq�@��_� ��b碶ϕ]�w��o3%|��kU ŬoC��~ӈ
BЪ���O�fL��o:������ݻ��|�7k"ع�^!��L�{w��	�{�}:�4S)�Y�>�0�{)��)c>�: ��l�{!*h�����I!��P�N9�y
�!w�ܑ�~���1@�ұ�yM�X2�XB�U�D�8**q���o�k�sqR�b%I^J��ۇۇo�Q��?4����ܹsGww�>�����;��ߵ�����M��ٔa ��m���I (�[M��k�\�!1�D�K>�$�\�$�\T�c��;iw:Rm4%�Td~aYN=��9|��
�&P�Y��3uV�V�
�e�*���4�>�T{N��% ��Ms�v�[!�@��0Ơ�Q��i�7�0𳅦c �PǦo6� B@J-�9z}!���m��1c,������ϙ]���U)�3�d{4-���gK���uD����_\ާ��.�S���玿gR�a��<���E�דq65C�u���>'����Ql�b��qT�J�h�o�Z�8���f�s��C�X�?�@X����|c�������^o����vcwoOv�{���-{�ۜ���lmnʠ�G�XY���\G:m��� jW�]T+���$��~�@���I{�#�FS*ժ4����#����N��Ҳ�q�@Q�J*��K�f�ʀc
"&����[����Ej����.ܐc���`c���6\ �Y����q��h)�aA���^���΋Qj�,�Dar�Z��Q���,�>��(����7��̬�Ҟe��8��>�of��ó3s����|:6�,MKAg2GQ�x���H���pn��������e4�l<�x��ԫ5 ����/.-v��V�������m� ��{�=�����w������L
�^�'{���`#AB�d4�[7����&}`�jUZ��Ԫ�41a�`�+u�C�c��|��VGZs�QTk�]\���Uy������cR���P{��@a�ΔjO���f�S2@�ى/��
�/_8L��(��0=f}:>���@���<WV1;V΋�V�5?�A/f��Y�)� >ڽ��=�8�}����珟���58?5\ ��`��YX@��y�ݦ/�4��HF����ڒ��-I��
u�IP�wl� $��w1`�k0����ޖ��M2�F��7���j����j=w���;`�2
�<Ϟ=�m�/_�Ϯl����px$MG���o<�0Id��:͆d���]8/�.�Ѫפ���T�XZ��ԓXb87��dAH�d�V[Z��4:s�h�dq���u���G����RotJ�0A��O �v0ScV�����;׬?{8}����׼��]�g>�{_h ,��А�/3I�1��p���5�f�,H�ޗ	�]��W(k�P� s��M�:�I�����= �����j@-��p��ADm��:0i�sۮ5��ڵk���.�t,sss���"�nWj��
��l�9-��Ϝ��1N��$.]�$���4�MYZZR�?[�6��t^�����幅/,,,l�`�"gϞ}���������W�\'aww[�w�@Ɠ�Tk�̵[�8ߕ�/o�����֛2���B�-$I!I RO*�ۤըq�yQ2�4Ϥ�lIg~A���0/��%YY]�'�C�I��r�A#�&>�
�����������و/���s
<��� ԃ�����UhF��/�����e/�;(�1��s2k� `@1{o&���YFQ��9/����,S2�2�W���e�K��m��g��8�t Bp��2�	����v�
�F��3�Ao(W7�	X�G���B�c 4K�s��;����,�������[oqlG����^�ٸ�l���������x:8�vʇ��Ѐ��8�ȍ�?t�ʕ�Gq���	CA.�J,i�J�Y#P̵ڲ�yG^y�����oH6I��R�@J4��q"�J,m B�#�I&��H�z�T�-��ve~iI��ќ�գG�ȱGP�$��R�\�Ʃ��ܼF �i@��z��q��?�8�;>e>�NK��:0� �j_��3u���ՙfd������
_�M���0Ytܦ�}�?��ٵ���iEa/���@��Y����v]�/;��*��`-߃��3ӲL�7g+�/�·p7��~�ˍ���������dn��N�(*}�K/�ec�q��������^z�%y�7h� ��|�I*;������o,t���ӏ=�އ��v>���={�s���?s�ʥ����=	g�zv��,X�@,�B�J,�z�~�J��[7��/UΟ}O*Q(�JUBh�I*IJ��Ea�&~0��^�яz�#��9EgqQͶ,>"��+���"���p�����2�}�g?��D�&H)�n���Χ�4=�~M���jz;�&(X��]��o2�s0`M�(xM�{��,x)�R�c(}���wV�}�ʀٿoc�&��^?tm�dsa>�A��}g(���	���<���<	��� 	z&�8ll���U~oyuE�S� �Tk��)�u�E��_��A���W�&^~�e��׿������G>�2��Y�qT�څ����Y92�k��><ŇgΜ}f���߼v�����US�I�У�̵ZE���S�+��(��~U�|��~i��Y��l"A"U̐����6����A_ñd�H�ޔVW��5ߕF�C���!Y=|T:s��A�V�B�R����f̀�4�-t_��
�F���L����s|�9"�'L���Q��U�,d���{��e�}��g�����v~��,��	
�n��}Vu��s|�&�?~?PXF�3a���G�?�3�Ef/X�����ۣ����䥕e��	�y��a��K��Tvn���`28�?��x�"}��G�X�g��
,դ6i4��?v��_{��co~��CagϞ�ll���W�������#���lԴcX�@��Zo`�䨀�J�5�_�"o����XߐXri�
 |�(*��L�j�!͹9�[T��������
��t�鐢Ať��@��G���%��~Sd��5�`g������^}�=�� �guP��2�+)���t~�����5�����<�	�?'�,�X��,�*� U6+�Q	^��A�����XnJ�j�/����ܸuG.\� W�\��+�V�G�CGK�Vg-��d��1��5߈]߷p:��ښ|�_���yꩧdqe�̽��"�j������X����S�Nm}`q��׾v��+��[����'�:��A��B��ZM�&*1j�IGٸrE��ƛrs㚄�DZ��Ă�@jq"�XCE�fSCFA���p��$($�֤�nKgaQ�s�Ҟ�'P DZE�1i�6�2����?f�w����^w{�mVs�><^#��	������a��>����㧩7�ie����>��@���Z��Y��K�2g�]`�V�,��Y�c/3�!�D�;�oe
�����(,L\�ÅELx�n�(p.8��)��}�ڼ���B�z�}	G��2,k]
�6��d��q��a��6�pM��/}�?af?�����X|��7��]�*��:����>�я�����_|��?�~u���v�@�73r�Z��
%�:D�K$ÏF:�ɍ�y����ڕ�2�e�=G���T����F�Ƈf���P��c��KҜ�Hwa���G��(�3�( H�9�@R�ݴ]i�,P�jǃ@�#.�i��A@1���k�7�4ZS~N�ֲv=n6/�nh�@:禍o
���t���ܻ؆39|��ǳ�y�sɀ����nsF`wEu�)��� 
���.�h}�+P2��3�(�26���)'^w2m9`�Y:v�@vvv��ٳ�/(j͆�>}Z#w�jYO��+/�љ���B��³�>{�+P�+�x㍵����ҵ��cw�ߵ"��d�)ցE���E�/�f- �<˝�7����ʕ�d�ە��<� $q��Q�J��t)��&��"�vS:�e�G�P�ʡ#���Ą,ƴce���1Ӽt�9!�Ot4�OԞ���DBu_�t������j֩�4{�t�iV/oB��Y�9}�1��?��k4g��,�Ͳ]�z��3@Qv�������s�M ,�9r	4S�(>ϼ��Y���a:��2
M�6�����\�z��Z��Q������vL5�R��xf�Y��9�nMb�H�����^#%��<��h�H&s���L�V��k��_���_�0̏�
gΜ;q����������`8F�"���~�'#�'�( �.Z{<��'ٺ}�@qu�"��U�d@����F�.���r��#d��c��W�t5���\
�����>"���jiҌ=CsAὃ�b��8����_`������w�E��h����w�Tm
�
|����7P�4���3>����E9g( �� ��k=���g����^��dl����AJ�!SӒ� ��̴�ŝ;�e"��P�D@t�OTӊe�y0CC�mD1��ѐN��^����ԩS
�id��,����$��͵������o<�̵{=�?���(���W�]�x�����w"��IP0M6G��D���c��P�Y&wnߔs�-�/I:�K%���iz4Ҭ7�дf��e8N%-�I���):��Stey��L�qV�h%���hm��J��Ͱ�(f�bV��R���"�S�Ժc��AO�	��9 
&�>���n\� 1kJT=�ߣ�*��rZ���\n�}�j3�g��)�z��}�l8&��Q���B���HC�8�H���rog���k7��>83��W��p�;�2� =0�oǣ����X}=X��OR:H_|�%y�wH�{�1FTMq�S:�$�0(�N������_��O|��)�P\�p���g��;ۿP�	tN���Y�2P�1�p�D!�L�L�F�����ݷ�bx�H-�=e�" �D�7" $la����ǒ"Y`�l(��l�$��������Lsh��В�P��pF�ʰ��|����J��l��1��X�/ld>hZ��s��,Lt}��-X�0��,`�}96.�Wc����� ���d��g12 �?���?���x���%�M���^@���y8�@�5��em�t��Q\�v�aL3��8�,�wU�H�Q_�R�a���ٮ��9�&`]��&/����u����������
*�BWaoo�Z��V��啅�����o�A�ý�w߀�7��wy���nm����x�<�h*b�F0 , ���+�h�˗l"7�m��������L�F���Wh0������*
�S���d�,�(&c@����ai/�K�=G��.,1��h�V@Y��`jІw�Z�N\���'1c#[���@�ʉ��0f�paz�A|`� ���N��Mp�������i�F����qn�I�F�� ������A�m�������~7'�1�YF�o��E��    IDAT�%��}���i���t��16cxϜ����Q�0F��ˍ7iv�t�b~n�IQ`0U���ĭ/3ApnF/�=�e�n͑P�  }����� {~�'e��j��ث$���P���V�W~�{?�X�x���W޿|�/߼��_���6J�y�5y5� S@�D !̣(�Tnn\���g���u�@���'����	S�^H|�]WI�L��/�.k5���t�e~iA��p|��n,q�7��d>
K��|��LW�y�V���k�w���ʹ�A@q� ;���AAw7K� ���f��`᳀���A���A�K�&�3�?f���̨��1k��ٴ91ǆf��]��=� ���N4����.�ꃓ� �����' ���tf޸q��[Z\��Ph�
�MPp�����;ח�
�(��E9���<��'��'�"$ �[��עQ���������O|�~�r��K��~���+?}����d<W!�� �U����Q�q&�
�-c�ґ�X�&�.�c�`o�@Qeg#g����V�I$���n��I8�F�I� Pt��(�K2���X����|�U�����ȱ�0y�K_��<ܯ��WC�\~�Wgژ��_�i���wf���k���ɽ^ը��c����Y����Aa�,jtO��d��N�i��>�R�o���(����.D
n�2��p-x]�{=��s�d�?�|���[��ׯ_��9�z�>
 ���6>P{��P��˰lM���_y�%���g��/XY1{�*�5�wWV�Y_��!��_}��S.\�{7o���I���f�e�SD���&�Y,si�E:��k�r��E����EL?7@���(
�3�FP��"@�̀ٱ��fW������JM��&����pe��&Ȁb�&�@���n�0��@�:�1k,>(���˗뱡@�?Wï�8��(5�)г@��h�A � �,H�;�3g�RQ(�!��z>����V�B�x�((�Τ�yP���6�Ɖ���>P�<y�E\zܔQ���o�m݀V��٩V���x��V�Q ���l��T1�Z�vnu��_Ym�?����&�o@��+�<u�¥O޹��=�@�X3��^
D�5��S�Ҭ��K����U����dGM4�u���ǯT��n(������^�BW�5��j�|wQ�an L� �pnvK� ���8�QX��,P�Ty�Ga>��?��4�~A��T� p/@8HC�;���o��,ׯp-)���q�i���>��3g�i`c0�}�������~p޼�L����z��\�#6~מ�L���Yc�'���]6N(��`0*� ���@���ͨL|͜O�8A��Mc�'�}���0!l�=�
®/���|���x��'hր���>�؊H�Z�xx��O<v��g�9����������w�]��+�;{�FpݑY�A�I�&�.��K�c�Uc6��b��-I�=���L&,(d�@�d�m��qqU�5�4벰�,K�W��MF�������k%�0�ia6
c����{..�sA�,(L+�������|a�e��f/��cQ���l�;L�	�����դ� Ϛ#�B]��T3)�>��w���$8>/�j(�1	��et��pXgs��ǰ�����y�<� ���|��L���:P � 		W �[�n�<�ˬ5�(��@�3��L6�Ȋ��m�cNz8H_z�ey��O}�i:��X�+��J'h�R�������;�ϞZ^޽O���7���W���/�]���n���
�Q<��1�"A+��v���oc����;'[�nK1И�Rcc�jU:͖�0�#�2��D�FR�23�Q�Ç�57�Tn�*������CQ����k�I�@ �������&���Q!�N���b�����Ĭ`u��#qM�{���[&NͶ��V������c��Y����{~���g���f:f����-�}G�}��3�1�e�l͙i�`*�S�6�C.�E=`vP������L
�G͙�·���5�m�V��^HM�}�������/=�jR���0=aq�q�n��%�ί�,.����+����μ/@��Ͽ��r��?���=q7P �a"Y���Z=�V��$� G�rD3B���Kr����u� �)f��2	�@�V+��Z"�H��g_�{x�whI6��$�v�я�y�w�5����msg��5.0�o�}V�/~��-�w���B�5�b3-�(��I��g����Z��SD�͝���\�G�M��\��}�b���g:�Ε>�]yи�P�]�}0��
ʟ��Y��Ӏ���{B��{~߈�h\�(p�z�QP�Es�����)�q��H(Y�r_&�\_�����/Y�ߺI�x��g	V0�y?��ͅ��$�������N�?�>v���(Ξ=[��q��._�����NiHKf�@6 &b��x�d+�p�q{ajN���W�����Q�G�E	æp9!+��L����CP��( @�N[���e�    �ݙ�O�;85�X�ա*`�?Q���lڀ��i�?�pSF��k@|��e��� n������4@7_�����.pj��G�ìF>�f��,��e�INe��1�+���_�a�c}�cU���vO'C�������<�'�/�Q���3�h�`/gV������+����.�X�Ǐ=¨�Ǯ���"0�aR/�{|n �5���G���_�^x�`�Z�O���E�f#~��W'�Q�V�,w�?w�����������}a�_�ּ��{����q�?f����U4Y�hR���*r!b�� ���XꕪLґ��ؐ�ߗ���$�K�!R4�a��PY£q%a��>�X�&�pj�;-&]�'�ΑՉM��y������im�m�k�Y��ll��W�^@1>����m} �c�Ţ�1J�m�(]ޕ����S�{�Q�@p/�*�Q������Z�k]g״�l��<���ij ����S��Y|�[9D�L����Z�2��C�
4�°ޱzqQ��`;K
�����&.{>1��	�����ߒ�|�+��N��?�q��G:�~���v@�����'VN������1�s��ͽs��������tՀy����u�lĄ �� P �d��@�M���s�3�j��� �\
�)
��?��ժ�`z�z��bau����f�M_Eg{~�k����@�3
<0[`���2!M0�2bG����b��&v> �i�{�0&�����Y��O�s�  lK ��p��gE���M/��25�]�3՟�]�;˹�oL�� ���/|;!q�-G�|&��$�	�P'��g�)2۩��Z4G����V�� 	��g��&2o(p<�(P���-|n��LZc6~ ~��'��:q���[4= F��|��;��X�n����9��������;v��/?~��3�//\|띿t�����'KF�-^���^� �[�"I*���Q�4=PÑ��(��҅�r��Mɐiɢ�@B��� @��M�8�H'n 4@��8"�讬Hwy�m��C�=ߕ���u�(�D�J�@�G?��p��W��������05,�o`�@).��
Ӏ~
�	�	�><?6��Vr��ךK��/3�,����o��{�6/��mn7O&�>P�{%s���mn|BE�� e�m(J�����~�T�[( 8�ݬ���i�����B��x������G��X�� P �� <
���BM�x�5k�ͳ1FM����(��_S>���(�?r�	Wh���cN�ũ�jۋ݅��Щ_|�����x����ο�Wׯ]���(���U��E�L����v��6��Ѭ�`�X�\P�X�*�/��;�(jIE�x�D�t̽'��� 33�f@IE��h�7K�T��mW��G��.H���G1��j�usd�v� )eW�l�(l���΄�Eg����iӒ���[�>Pئ�& >���`��Y��G��oދ�(��L��cKF�f�7f����Q� 2 �����7�J��� {�7O�́g�S��ހ��qn�h B���<W��C0g�m�c��#�4�ND
��ٌf�p�ZD98"Ph`$\3���(�ӕ�[	����}�7�s�����P�;��l����˨�j���������S��k��}�Q��ڻGϝ{���]����9[�X�;���HG�N�2)�F�!{P���	؜	W��_�[�|_@��T�<g^ �f�x&�*D��h�(:��p	W��,,,�Q������a(�(e���@���>:g�5��;�|Va	�n�
��nZ��4�7ma�7A6�`�L3`|�H�$�>��@�rO\��,����4�o:��鵢�ǜ���^��9�3� �@��f��7��??6����yl�F >�軻eJ����V�dz�H���f�U�Z�1�
�a ��NW��i}#����^�/��^O�LK0�(@AF��[�/|�@q��#�uA�B��k�g�
�j���|�W9y��:qb��c��r��ŋg���[����(�r�B��P�~0=2�)r�
��Y� ��x�ܺ�@Q�©�����Il�jR�ץ�����5�c��.���d	W 
�(��6��8�-��<
�UT��hǬ�4&�kU��'��]��{ڟLW�$�������0�ڧ�v�;&w��8t�Ge�5L�NK�E2�'�E"�Ŭ�A�v����?��@�t���مL6��bs��LF?�	�2�l�ג�A���( � 

>M���2?�
���yp�n���
(��1 ��Pw��i �	W�G��䪛1K��%�Y��u��n>u�h"�3o���?/.��*�۾��diy���� ^c����§�����=���(~���x��������o<���zQR c��x�M (@��D[�իh��h�(�>���7$ذ&O'/��1���Aa¦��r5B�'lL�AP���n�A��t��nIl$�C�r PP ,,:Ӽ�
�����0�5o<������5�i�l��]5��hm1�Sf`���y�)<��c&	~��(�V���3c�Պh"��m�j(|����/�@�����B�-i\�	F~c\c,�f��E�ٵ!�"5����`��
3�A�޴mׁ�K��GYPmK�S�S��g��ҍ��}�X�N ��f��[�´{c��l'Tp�so����17�y�ݳ���/�-�����}��a&�/�.
*����:v|��<� �s/�z����~ikk��t�V���6��[��~��G���?ӕ����'6��d���d0b�U�iw <8�rBkv�bG-,9��r��E:3�\�cяN[�5��&��Դ���'���[4�_�|�����\8SM3�6vȯ�Y��&�^�}Ŵh�p�v�e�=���\�m�T�@ �hڸ͇�Vc�	j� ���\�L/���fw� 5W61�H�L���Hs�u���o@s�j/C�郠￱jfY���12��L�谖�u� �c��1�����#o�8r���[�>v~A���7)�K�L�Fx�6%��k�@�"4(o�ml@!�����K_������
 ٙ #����k�Dqoqa�W�:�sO>�����_�s����?�iL� @��(�� �]��U5!�;3r{}]�^8'��]��ףɁ��2��6$w��V$��e"����{?��ԫ�^\��e
�O4[mv瞛_ �лm�:X6���\Zl�]�񧦄���wY�P�.u�7M�&1�A�^s�y���C0.pv�*PX~*\N�	�
0��9�aSܲ�G"
����0�^�̀B�jb ��}�i&)^6�~�l	�n�%Q+�v�fzhB�4a̮G���Uf�����
d�ZH����k���<�ObU,�Z������y�I1���#f�;�k�3��a�0M�M��X������Cs�{���Ñ�h0֕��
5�-/-���N��w�>��ܧ�}qf���מ~��s�����nh(�pE��Q��q	a�K�Z�j-f�Q Ũ�'P\a�պvwDF��1�.�I��N6�\��F�>r)0����t�����$��y�U��
��,P��XF���rN��Y�Uj�S��~���6�]�ϡ��@�2��e
����rMrՙ��C����Qc3}
�D3 ��VS�P64��G�I.���f�>Gs`��	;�-�7�8�HA�:�Y⓵~PH�޾�Ƣ|0���-�@Yդjf�_��z�Ib�( �pe�E�=f�|��,\߀��VQ�bc0ӵ�1k�F������c����9gse���f�).�̢E�-yo�y�����1o쓁bl<|*��ߝ_��G����(�{�o�������.h([�LT����E�淮�#BO�D*�D��`?���p(��m��������ܒ	���_��"��W��`2K%�0��	��Md�_�H{qI�WѬfI؂գ����9k@����t.���tӀ�Y���)�����Pp� ��G��:1�C�(10��s(>NC3ʺ����X�9�"�ͤ3Mu��d(��` ��D��Y��;��:��70�	P(��­��Pf`��O�O�@�s��b@��G�+��J�`nm3c��X�ۢlFk�1('�V��"t���F!�Vu�Q��������( H�����U�l��Nn3;p^��Źٱͅr�r4���ƛg�P�GƂǱ��+Y�:�??7��G���o�����L�<܏�}��>v���O�l�|��SP�v1G�4c3�G��l�H�V�F%���nܐ����q��l޺%��]�H��c�Q����E�:�g)���B���,��23��Ҭ�]?�
4����$� ��&J��X���}2T+����*P(t�>9��0u��be�T۬�Mn~���n�S�u�8�ٹX��z��4��[�pZR�mG�H�U�z[��^�&O�tW+*��.�!��D���4�LstRHf�� 
����x�w��3��˜4Mml�s��1�`pf�}WD��� n��h���������O'�>z�\�&��780�Ga�kJ�"n}9 ����݉Χd��k�c���]��|���Q8K�8����IR��p�iw��cG~������Ϯ]��ɝݝ�(J���G�E!�̱�05h_�ِF�&�J�\��;w��ښ\>��vw��G�&	��'�5�1
 Ec�+��E�B�9���ך��,�5���K�ݛ�؅H�sf;�! �4�	�l�~hPx����)��2�H=��zXw�J	 ���Z�9�������>�ͦ$�����W��,O@Ao<�"�]�5j���(,��"��@��A�FdpT���f�z�v��=Q���^�6P��P��7P5�)�*���,O�ܘ�s�v7?������U�Sߐ�$���|�*��]?��|I�јU� 
n)���Z ��-��:�c P0�9Q6���K�a��s�α(vq]T���P|��Xn�b��vڭ����#?��c�]�$��q_�g>��w]\��ɝ�ݏB@TcdJ�4ڑ��a�2�*	��(D]E���m�y�\|�=��c{[��X�4��a�wE�����:GG���BC%��έ��Q4Z`�S�	��\�ihS�汙ˌ�-߰��EM��q2��zU�&��Z�[��n1P#0�[O��3U�vB��DhV��49�O��N�@H��V*��Yܾ��6N"�߰�?�훆��40�G������6�qє2����I1N��S��4Tk��B�iKc`Z�8�4L����vt-��F6�����۹0�`�(8��}�9+}�ޫ$jf�AXnRlQ|�滈z ,��@�Q��gGf���G�l���m�i�#���a;�/~����}���駟f;�V�-s�]$#���v��.=�ן}��7��?q���O���>�����£Ԛ qz|�    IDAT�܄!8:�*�4Z�R4*UV��vw�����K���b� 1@ο�4r*���D��s{t ���`Wb��E{i�졎M��qP�C�f��`�U��Q�m�⨦��=<5tC>�1|�w�s�iUDS�=z���� �7��(�!��i_4�1?�<k��.}��:r^s���P�jB|:d>�U��4�5����&���74��)�	fa���K���Pr�Kq��L �67�0PE�9`�e��O��A�����((�eW��΄4vb ��d+
3W���=+�>}U����΍=+��`��Q��9��\��|��2J;?~�[N�sǵ���]wy�5���g�+/��y�3@��5�l1�PPP�����o=u�'���G�8F���[���+���' l�X��-����~-� �Σ�H�U�j%�N��vx��m�zᢜ�&_��v����?a$�*���	����X4lUI�%0�XY�a!���	w��n1�BY��T 5��v�N8ԕ�I�Ӵ� ���٘�(�~j�'\��C�+Rox��QС��l�k�3��u��i!����s&`Q�).mס����ǫ&�C�w
������s�?�:4��!ޯ�aU�؃�1L��UFa~��ZRل��+�A:���������zߵ��d����GC��X��h0d%��l\G�	k�΍g�� �>�0����2�4�Pf�HO;u�~ `fJ ���J��N���sԜ���ŋ��ӟ����Wyn���]\�����9p��w:����C?񱧟������ۿ�o�]��ˣ��1d:�t��bf6���H�գ
�^�Hju,�:v9b;<0lP��7ަ�1��1�[���
DKH�Q\�Q�0)�l�4��X=:�]�J9�Vh�04��VzU0�;�D��c��3�`D��Nd>�Rܓ-R�H�XG�ѥ˙�31���R8 �V�7j�:e�r���/���h ��i��J@^���j�Y�� � ��O�����(��=�1@�P(�М��$P`[ Fd ���|5��4�F{,�K}����J�]	xS)�P(�Q4����2�&��s�0�p@���ܹS�QAT��8��MRe!G�_�?�)�e$e8���� �dT^����P�5%8N��k4�ݐȅ�����
�7"*�|`�;<8S�v��q���͓G��{�ԃEQ���O���_���pxR�qa��>�
�S�� 
Gs]xt�ݐ�N�����]nP��7�!W���/�y�Z�1
�'�gL���I�-�C����������5�?����D��:�2���FELs�e�i��ZG�[Nj�v�½���"\�v�[8p��v��q��:5��)TkM7sf�ŭ=$\�G�()������}��%�KB�(�T�5���q@a���(`VN#A�� P�=֨N�۰�~Bs"ⳁ3錉���aĽS���v������9+`��M�XwS��o��@�|��ԎUf�Y���ဉ�C�L�v�Տ � T����s\����6f2�:s�*�E.qU����������c�N��XXZ�P���G�i���ͣ�N�����Jrn����]�����B4�A\h��r&1)��� Z�n֥�jJ5a,�~On�o(.^8'�.I�4�\A�Z�x6Mdʹ�iȤ� �H�ZY\^����8:1����0a����ڎ.
��@�u��\�.�Yh����P�ؾ)��[];r!�^�� �׎.ת@,R�h�셚�L�r���vۿ5�ۺ�4Ì��I�&Ȯn�P�3�k�W�ԞW�`��������B�x�T������	Ts�v���	R����P����ޟx�6/���44�j5n� `{ 0���M�W�a��AY8�"z���=Fq���]F����v�NYr@⟏�]��[:Puջe$�
|@q��:^(�(�2�
��-�p&�z�7��.�W����+�4�]���/]^����! �4I� a�á�V���_hXc1$��h5�҅�{��c�u���3r���r��j��@�7:[���dQ��d�H� �-�"1��bO�#�Npsb
PiM�҅�l��0a>
\�Zх-�Wl�B���	���>�n��=���� 4|Z����4&�..��I��v��^U�.��qޝ�Ø����.e~�$.	3�>�'`粄&�
6CߘQ�ъm��/��4�E��7�L���B���J��a~
033el��\�P�LV�G�/�`Á���m�=�	��!Ϣh�'`�o��y1v�ޘ`��qi�R��y=��������L��o��2\��[�DAٺF���n޼-��������ٜ8~R�qVBc��o�YV�Tgu���w<u��Q<��;��_}��.]��[��h15t��,3�nD+�P9�b�Pci��iԫ�E"T��&57���ٷ�!Ͻ���&Za�lUI�)��җ�6�U�-V�v��+�����5�JY�c��edZ�	��O�t�N7ۓt%-M)�]�Ù*K��4m5�g���=��u1�q`_F��9�q�_�F	L#�v�P��\5$mǤ�L.P׊�L��6����Zp���9, 
uRQ�0���1��L�5�5Ѓ���4 .��ܦi�^�
IS��4���,��rp��>C�8'���~�%���q�=��)�XK�?��Z������ ������Hm��9S�&g����&�������+���_{��y��)&t��|X�`�)8��ǎ���(ξ�Ə^<��l2'��2v�±��&��i�sIlTKbi5��\UL&�Eq��YٸrYv6���眛kjw�<�� �<�U:��m���V����V�d (3��ů�>��]9���2	�3���=l�rL�]�氳Jɒj��+ن����'ʆ\�������f�*M&9y��T�n�r:�9�b#�PؽhX�$�]&(���79���sE���|�l�;e����۬Q!�a)��&*8������V��Tv�Q�k��DhG75�����t����%Ѽ�-(���*3u���Z�8*{S�]M�SƬټ(dļ���֯������(L���uy(�m�:�y]��K�o��.�����D�h�k���N�i����9q���=p��o����7���s���'Yс��R��ׇ̐%ʍv,��F�	��|i�݈t��x,7�_��Kkr�"�Q��07ߦ�!D-�u 1�BKR���\W�]�t��6��{crA���ӈit/�B�� TUb�>/��@���Pk2A$���N��yǦWQJAp���<�8H�/0�]�e�ގ��<��2���`J��C	0�/�{��i�G5�����x4����^���5J��A�E��#�<��Wn& ��T�c\��u97���g"2,3u�"o�P;K�����P��WWMk�jv`�� ��.23��U�b��Cj�/R��C�47�Y�*v)�0��ɛ�40�֜TQ�&�j7Ċ$�`��_�I��cO�"�r|���|�>��֮Й�0)|k(X@�����֓Y�uZs�9u������W��r��ş��q�G�I�\Aq���E�4_Pz�3ʟ��v�Tc�Z�H�vv���lm˭[7d{�C�Ӥ�ެQÇ 
<dך�����&K>Bc�.44ԅJQu��� ����Mq\ڮ�Y�q���̵)���:�Tk�w���1Õ8�3��v�v�଺�L��I�({2/ĺ�	4�X��W��B3��@����iT [�2g,R�k�.�S�i�If9��.69�h��o�(��)�`|�FCF�@��>� �ɜ�?7��``��=��|��1�xee�=8�g�\�XXƙ�<a����*\�U#u\�ˁA�L��ؚ� a�`�"���{<�ם
��w�|<�V�	r򨢬����jR�EtRk��fW*   �ߵ6�<�UbM1iP�(�дwkg��8ϯ]�˗�r�!Z>��
Y�x����ϝ8v�G8F�/�p�����������h<��&7�hB�W�Td '�	aף�EH!6Y��������Ζ�>XK�nv
����$�B&�9�,E����H�B0L�ij�UC�����ۘI�lu<P,f,ƽ�niWk~Ø>ێ���:�����Qn1��f����!�x�����2�
6��	6�e�\�6 u��	�;1V0>���φ`�����Z2� 5���[K̵FDM4\���!^{(P�I�7�� �hu.���Ew��d�eڨu A-���n@C�D�f�����{a�����5�g�*D�,�kQ2QY�X���z������3^�_��k�{�Y81�C+p���6j2��+1 W��E�,oaO�����X�ze��>:�2$�6	�򦻠e�f��9���AK����쉵���������4��@Q�k�+'�/Co	��4�'��y*{;�2j�9�9f9+K�m�9T�֬J���+e�i�j,\fN( 4�����H'hC�"�0% %�Mqf�$Bs�'  �Tq<<�q�������PC�"���櫀&`��-\����m��AC!�ʯ��4�g%R��b�X�$F��X�� ,z���z�s�4*�7s(�.�,Z�����Ҕ�m�DqE���h�3jyL����a�\tA9Fhp�  ��'�>��K�29'��턅/�D��L9X3�1(����p����f*��Ӑ+�����_������9RQ����ڏug�~��7s����ș�\l�vD�p�;[[�ǉ��V�"K%P������j���Gy��o|�O��s���vw�L:�Ѐ0=�na
$oؤ�p�9z�8�v7e<P�0<Ӏv�D���p�š���Df�eW�xF�5<�
�����J�(LG
���kB �{c8�Qja�N�р��(�-L
�h�'>�ɴ9��/��@)�@��k*2#k�o��f�C�UX�2�ҋ2mm��N}��1��/J�����r�!��+�a/�P�l���F�&5���,f,p�9�ر��\5<���[��Q��T�P���qD�>j#(�(�
��/	���_����X� d�>X�	�n��ﳚ�s>���A�������� tD�Թ�ͭa�`�DM�i�IjL�%��g�m �u�BSa�ɐ�2A��~4�й󄕌�
��̱P�
ߛ�N���ܹ~�&MDV [X���qZ4
1˲I������������sϝz����᭭�g�e!NEPi��Ja�@���fC;2�A.�ޮ��>x�fihK�]!M�D�Y� ��=d�M�ZBG(��MD���k)(@�2�9R:�ߍ)`�Ц�j֞�?�a��/�p3d�CT������Q���l����'0����X�h�
�0'jR�5
\����Ԇ5M��lQ;z�����>N�R�paN�oĞ��sAq���x�d��48f��q�(�%��֍B�M��z/D�!�p}P��&�a�? ڸ�' f4�b�'-��:E��D@����>��ld�� =�> -���U"'�����u]{y��{:L5J����f&�1Y�9i�,��`����ZV�	f�MQG1�O�f���5.���,DG��
cksGnݹ�Κ�z��|F.�O�&�j��KG����x��=��-��-��(�|�_����}A�;'P8�C�N����A�PCpTƅ�v7Iu����v�$���`�� �)��5��ٝp�`BU�k�nب�,\�f�#��Ij�̍v��4����F鸢��c��)X��EI5�l�����**mA�Ԏ�ڛ�3vA�%GF�P�%���ԫ45j`I49����`shj�$]�Le. �
��aD�R&db�o�z��#�G/�����&��@璟�>��ό�c��9]��Fʻ����,�l�P}��:E+��@�Gl�Ϻ�1S�1cL�f��Fe��t]�pfZ�sׇ"��a�df*�:��e�Ztǒ�pP
J� ~}
����v8'2L88�%V1��=W���U��.e��mxl@`:%��t� @1��ޞlo�1�\	L��z�ˡ��jRiiy�ǿ�c{�[F��2P��o��cg�~�S�{�?�q����T��E�K�#��D�p ���m��we{sSz��Dj�]93���D:�/��)�7�`�?L#��FM˺M Y߁�7d����b�ZקFqU�(�P��w�!��l�٤S��Jj&o�M��'�I�1�}q��waY�Iu0��ΰm�Q�f��l����$�����^�a*��nK�ӕa:d'���6�H�#��0���r��,�b/�A�ХaL	�[6#���ѡ�v�2�%|)�k�H \pm�~DTj4��p�5.��j��Z ���DpV�s���r�i�aI3?�ܛ��1i:7�r�\J8MI�$ԁ�ϟ5�^9j����t�{� �����	�/���}0j�J��٪91��3�Qx���D�<4�]sc��!�@��4=8K]q�:h�L�ZS��O�7����w����u�����2P����'�9{�WF��ߪT*:����6d�ud��q,{��Jl��]3y�uw10m���0Pƍ>�.����54�I�$��.�EA`�0�|J:��#��T��4�~𶵃w�����3Ԛ ގ��8���]�������c�uںZ��Dm��Ԅ�I;�����.hל��@c�rX���{<��;���p�����L#0�����g.,#wab,ȭ;[���yз�H���f�s��M��N2�]w:s_����x&0,<�2��P�����R���0����9�]}��h�,���`�xj����±�}�}�sP�� fU�(L�g?C�&Y�قp7�
��,z��F�M���,4�y����8ƃ9�u�ɀ�/s2����S���<�A�ڗ�;�����A�Z���:ݕ��h���ةS[�,�P��W7�rs{�{� �aXX!#�s��D��} hf�._Yc��֝M
 ���%^�j�Ea�o@x�
�;�u� 4tZ%5��hO6ͭ��X�
Y�$-44^@t����p��8f@�BY�љ����E�k��8?ƄE��%�c��� �u�KX����+�h�:(a��*v7C���M�q]|w���L&���ޗӝ�pO,C�p���P������b2؄��}Z�d�d�i����v�=�E��}�� ��ݜ�Ϙ�̦�3�قs`� ���;G��=���а����p|S��M��V���n���0,��/� _I�@�|��p.�LX�-�'�J�5H�4L)�dzhe��s��w�VÈ��g�0�֜�� �CX��a|`�ŉ2
n�P�^�Gņ|�������sm6�����?Y�t^\��_?~���v���o(��o���k����[�n��\�HM�
5�!#b�lC�ﰇ�����?P��ՙ}�1�c�4�u.u@AP�a�D�vu�&t�H�c1�5�^q~,V,HDG��+�:<���Ts��~����F?���9�I]�8G1�ZB�1�{Cz�Q��s�{tb��F�}�� ��{��;�9�۷7y�j�^� �jRU��@Ӑ��&Ǎ�U�����K7h9"�p9
��qN�����!c� 54G���ɢ
�< J�B����3�I33R���p���_�йp!y�x�	�Ox�P �<����[��݈����q>�fp.2�r&�n�̛O����a�i=�!��PG�%�1���F1�h�V�j��%zA�R��螧���
~h����m����|~�fK��nv̼�\�:0^M��0�Be��*��:���j&/t����P����ɍ? N|�]����?��������[��7˲�H�m:�����MF7���Z�񳡌G
t�:p2M
����fC&Bi�
��8yYz-����|� ���Ή�(��"Д[�Er�������i    IDATƻk.Cą�m��r�L���e����2���-e\Z��K[�Y�+E>�'4��)�)�$��5��p���Q�9������[i����q6O�X�s�E��/��ugy+�À�����;��s��/��1	hn���i�=��1s�j�����`L����q~2/Σ�k��#���x�gf�����!j煂Cۘ���uq�J��`d�27�bc�|Oh���������<Me��E��G�������O�F~�+*���"�2L^G��@��`
y��(�j®o\c�̗��ó���ӂB�b.Q�vn�+��۵j�������u���fs����hV��z}K����l���7n�����c�#L��U�Ɂe�"G�,9p�0� ���A3 U�@�`a����eP'��ϡkW����G�v��NX��E���
�&�` <X,Ko�CC:5�`cQ��
�"8�2*�(�Ę� �kF�5�,^��nqr&dԦ0�\�I�V��6)lF��M��N��������e�sԶ;M������S��V	�����d@gJs�@Y?r���E8?����o&����cse�RgFZZ��	�ӓ�æG�������4��U,�9��.��r��g
��iL$s9.��9$p�P ���m`d̏�m��* ��^]^��md���S����P��Մ	�{�Z�* �{=m��&W�i�2��d��.��4�۰�)�Y%W�(y�լ�o'V�|��g��� �(���#�/_��+׮����ݏ��0!p#Vd��᠐�Zo@_ �=f3�j*��r�r����lgؤ���� �dΡ`\0��:� �==L\�%��k��D�q�6���58���D�	��P�T���A�z{{�dŢ �MPS�=��> �5�����V�@a�������hd} X��� he�lw�<�L?��Vo>ܿ��C28X��;�}8[.�����ۡ@���9�?����S����L�͘g����Q�	�������1&�&[���kA)�Z�LƌJp0���N,	�S��\��w��Ӂ�/��󛠣���g�f���<th��2�1��D��߄�{ah�uJ-5+���<�����,�F�c���;�2��D�����μvq��8�>�e��`E�nf�����-&��;=#n�!��dZw�I��|w����=����`���3gδnݺu��ի?p��忸��s�?V01�T���j���k���^NM����w�y�X X��-l��ʠ5NM��+�2�!�}>�F\��i;��F��4|L*��|��@a&�i�Z�m�F �
���F=(�e��ڷ��֨ �կ�f�ua��,�y�ʦ������mx�����NƔ����#�����	�x��V�F-d�b	D��[BFڎ/A���
4��oQ_͉\[ �9��S�Fg��q>�
BC��� �����gL 	��R�m�AT�Ri��Q�.��`����*��ni�D���M!�rs�����(�,hԨ���cA\�ń s<��M߂K�um�5�#ڂ���Lt����!�������k�M��<�s��}4Ҍ�}_lI�e[�e'v$�!�8?��Z %��@m�аJYH=,�á�
I 	�8���ڭ}_F�F3�}�{?��̌s�zG���M._��O���w��r?�c���f�ǽ�s��8G^>�"�⌈�/�Q 
���bO.��#ZJIJ\��\�h��{K�J>׶��Ƀ
���g[@q�������k���n[^^n�x<%��zqp�R��Q�\��>z Ȋ��-M_ �@������0���DS$Ɵ�Q#P��"0�<b���e!�����fzq�4&�����գ"%+Z襄Y�&�Ɍ�1���RӋ�k��&�0U#J4�v 
�����dT>��#�K����H���f2�pNA�LFX/�%@'�0*`�K��.�"�L���$bPPG��$RoR_�N­A�b8� b)����Z��^XTJJU+��A����:%��-���b�($�KpVDXa�pKlЄȢ�B���t$vr��7�@&�V��{�����$�&QE�d*�Z4>8.,Z8�wD�	�'7���t���B> �h�#g�-tPu:
P����9���*V�$�Y7��A "�� (8L�$�}�X2~��;SUVr�[����/�
er����t8眯r.;�ZZZ:��x����/0���|����h���p�]X"V&�h۲�<Yإ��H$�@��$�H$�M9]�s��Ƈ�d��ﱳ�./�~H�k�"-u�����
i.(A���E��d�`���T���N�����{�	�(pY7v-�B)������	�b�D#e|h���ƂL[dE�f��E,$�Q�@5"����k�K _J�@"%�I,,~!( ���d��t$ԭE`�3�J�#uA��s�4�u	+"�	+�RȒ��n[2�I�'�(�&�B��m�Y�P/�p�ŇJ�+X����s<J	H�KnP���ի��������&ˎٙ�Em�@�1@iM�)��T�D�z<���O�fI�k^�[%5����:��[ Լ��F15�� �-R٠`|!@$U�Y߄\��W��D�2XΜa�E���ܼ�j�*>�ӧ/�؝1P<����ǧ����z���5���[a�%�GRy^�[(,���BH6���J�HY[�|w�BT ��IB}�D�r\E�� ��ԑȔu�����C���r���9|\,X���nX��&L`��,%ב���	�Ȟ�"�"�pJ%RGwXK���e�,��e#J-J�ޥhq!>���[Wt�ta���R�՘��`��KHcA��$�s 𘐽c�4�r>����Iiq�O�B���O�3�g�����@I���̐�4�Ő�ܫ���/�& ]*�,R�󉠺�?jq�
^$�#�����HN�]K�.ŮP��0�n�oh#��D�wi�EK�+b��a�:�<�x1�	�	��1�BkF��w�A/�1�M��*!a]���B`c(�3�� @"w�H�5eg+�Y����c��0R\Xrg[c����;�K|2����⾾��LOO߱���� Y\#�@D�1h��'�0>3)Q�X���/�I~�$����+K����6O
ق�l�+�Y2�Y*�(v�WS�	�V%8�^%X������-Y������B��<��;xv\��#`0F��E�ui�P�J2��eC*�^"șQIxZ{Bb�a�V	)9���,'�J��G��
�d@(_�t,�H�>�z�|(&��@�慌Ν�zE����!�#�3��H��_��)Bgp,�ǁh)�G��܍�������{����S�BK���Kp��;r�H�KX0DȳZ(��in�m(�Y�	�P�9��T��z�@V�ۄަN'��9O��".�Ѐ �6' ��O�-R�����l��5IA���U��P[�+I�s���$�F��cF�7?����Ϟjow��@��#��mm����Rm���u LE�H�K��I��0���@�RO�%�@M@![ı�4,
����.��h�L�߬j,+-e1��ҟ��`
5h��T��~2�W �x��R������P
�дP�U|H_r�C,,�S��BJԉY�@b�cE��I�����M�,�jP��n�D4��濘j�r�	^4�4(��́D<��4:��}̄O��J�@X�l���dB�P�.��M�K�>Ǳ���Ȩp�*��FA�I�$#C'�Zg$#��X���H.@t�I��6�%-
.�:7���'�cH֭�҄+"�/���b��s#sA�I���I N��)� ���}TЎ2�(�$	�'�.�0���b3#��J��(�h��Y�%�!��K�"�^��9ϕW������^@9��щ[&&ƿ����x1�^P��)I5��#�. H'`bmX K�S��n$�����e'aj���O,.�Q��^	����I P���v��>���.`�"-^x`�Ү�=*��,@�� 
,8���&��������{b,� ,iJ���e��TZ9�G��~�k�1¯MP��Y<�pRގIih�� ��;�wq%�Ol�q�;74�]Z
�0��KOz8� J��C}	тPX|)*vʢD�/����R�N$#A�-
�E�w�A�CE�-�p �Os�%��D�7Y��T�<����t2*���k%}~��c����G�Z͂���/�W�����ڱe�`�$<�� �Kmx��%5Wa�Pߕd�V�xp�G�x\���*���D�B$>�I
���^�y�y�mo�{�t]�����e]d:��;99ug0 Z �`�+��$v��n�(ǎ#��9Df<h������K%%Ǥ=J.;g��$�c�� wdL8��]�9���<�;�_�E��H\U,p:����h���9�a�u	T��ŕe��3[
2���� b��S֘��A�|vi��T2h)�BZ"H��ye�aA  ���;�1 ���"aVIT�u�-]\�KA����Eʹa޾(h��q��Jն"9�\C"�,�e�%���5��2����QQ��;�����kCϋ�@4DV�׻E�2�����!��@�D�����3	R2�@@�4� �)���S�.X�Hc���P��/�pƽ��)�iI0�Z�襘�Yi#���E9�!I�NSq~Q�-�R�HN�mӞ����O=��;�c�=[<>�w����;�Ѩ�'�t ��`��?��b�$��}���RgP�Tز@��w!zI���J�'���_ è���>�
<�|��� ��/����C	k�d�I�O����pXԷ2$(�d�Z����u��
�AJP6�<zj�X�ٯ��F'g)z.�#���n)��>"z�>�#�D.6a�� �K��I@(mצ!���؁�J�҇��t�	-,�0�� �������!��L{
\�G�e�X��,;Jh�)�{��j�q��ủ���t99�o� R�X�8:^�Gv1��%��V���A& �u'�Wj�HKcO�%́l8E�@�G?�d�h��QXVP9�X Ԥ����N4ub���%�����Ú�?��a��Iw��Vj��Ǥx���G�95��������V~�S�^2NqY��g?�u��D��KKK��0e�NRl[��Iu��n��~,�y�LN6�|R���wlQ�X���1T���j�ll#t�O&@��DP�w_
&!� �^&�Zs_������d��ԑ�z ]A�R>��R���T�� Ar�Ʌ��ˋl^^�p�I����v=8�C&+/�m㒱��/+uD��rRM+���^�����,
�=�]�3�)�;$�m(&�s���ba���F@#-;�bR؜�h���:ᵘ|v
������QZ`A)��`cQ���(R�X��(dL��}��aJh��m�T:#�oq}*�B�E�\l BdA�
'��Q�@A���v�	(��1P�W.�o���J:9g����C�d'�/ទ�z,XZV���j�?zө�h^(Μ9�300�ƙ����
.~��QM�7@^�C��˄�2�� �"�E��|�Ң/���s �G�@�AMPPЇ�c�o��9��d��ًd!�%%��@#&�^M��F;pA��G�R�l`�lJ�2P���ϔ�K7�c�WN�t)()���n�
�D͋��8#�4	�wځif��#t<REk´�}9(�(,
���y|�܏BlcT{$wxQ��`�����_lj�i���&,�9M��k����� �뉭*���l1���^��N�VP,F%�(D��s�D��`A�$�u����h��,��wp��n��H�,i&������,��S���Q���V%�iӼ�*O"�+���b�9���k?)�H�����	�%w3⫬������p������,P$	�w��k&&���x�XЅ|��ͤ�#���Z)ӛ&��)7�o�'Rj7�`�V�sV�a �AAz,�T"U�~�?��~2��1&�X����왉4΃.��nb��L����ْM�*�"���A�A�7�[��Ơ��b��Y��%�K��A�]��b��N%�H,Pv�dI���\<<dp°#q�#Z�rg��B��`%����q*`�Yn-(D�Im[�]2�(�7|��]��x�Mo,��h�8�����҆"J	P�A��ԡD�X�Hm�lH��4����	@Z��hA�y⿔���(�Y�IR�E#&��u�AJljd�������ng��ɪ"D�wB*
j$I(�-A�heV��HKb���;�GW�**���l�7O�>��"7�
\���������/��o�.
#�D?77���7�hϓN)Fh)˞�HI/�w~�y!C���;�8�@�5�/a*�@�,�}ZX Z�"�	 @P@A���Ҫ ĕ1 ��_�1�@a���솝�-$�Is�������B[
ٟ�	��"ԝt	@B��\3Z4�%�~0,L��\p�f�0�I���\�s`w������ɪ��@!���)�֤h~ڽR�	�I@��Ѹ��h��7� "���3ɹs-�(a��Y7�z�դ	�l��@�p���G,F�;PH�].hVv��-G�9#%�v]�Q�rD�9�wT�I͓ ���n�����":!#�k,}���F�9�fB ��j�q����=eyyϞ>}Z,����(����ه�G����@��d���&��"˂�$=���R��|	l6qT��/f��v�a
��)+��E�Ԗ���B��M' �Gf��I/,��º����{v��tOrASg4�dz��j�o��A^/�*��2t$^��� �s�F��(bE�� �IK�_`�&�9/�W�Ks�!�'T�i�w��ݏ'�{�����c��I�B!��;	�,�|����Ks8�+B���V2�ʩ�����'�\�˂5����%�,J�^��E!F�nc�E�ݺ8²  ��㹸����BJ��c�cGŚ�ƭ���=�Zҋ�j��@1@S���$�/eA��(j��@pҪ��B��l;������w�	���� �)���b��¼�V�T~���|��K��������{�g�ΙOz����|�&7L?6��T�_x�0`e��,,a2r�o'/�~�Xp2�λM�e����E!N!�ՉX<n�@ດ��.��$s,�<7,$���eZ���&��Қ��AG�l���'��5�%��J����".�3�z\�!�"v�na��#~�j��y���(�AZj�=u4�.0��Et�U� ����t�;�d����I@��3��;
rɪ�_�s`Nh�e�W>�� 4+Ȣ��Q�+$MYiͥ�Tx���EU)7��e����z P��x|E��J��a�%�X���Z�ؘ��i�%�4T����bVɞ!"8����Pp&�7�z����c�%���>}Z)��'c�x����'��V>���aQ�e�'&SwɝY�0P	35+N�F�|�R������E;���4}���/	�WI� ���c��]��a����Y{�ep�vE�҈;��H��Dz�fN�%_��R�LѼP�(]z饢4$��G�[�̩4X�y9-&Әp�,���D�_<��KW-��@��lH f���c��4�����k�0�/2E��	�Kr=R.H*�"�����"x�n/jW�
~ �W�R% ��h�˙_.�4To��}T��r���,s��{v)�/<�㸑Ȁ��)E��t#A�&7K�Wy��¤1�Jc!�������4K.m��A���PF�g�����sPŌ��(��Xg�9�J�˾{�+^�����H����������[�~߇��h���7�d����`'>����ş:VT~e��'�Y�\p    IDATO�$������#Us��X:P�#S��--0 ���@�["������럊eu-ҨT��d$vM�eT]��� ��5����mpwww	n!���������0@�;�ν���=�]���ݫW7��Ҹ������):\�vԓQsL��&���4�e\l�4�9�T�-H�on'7q�͚�=��mi�z�ip�A�(S�\�2�����2��R2�ԁPS�:f�s:ZA&�a�h��S�ҮBuK�Q��*!�
�	d377G���_�)ܡ]�/�f���j޸Kǃ�;��������	O��4)P,X�qd�%��	4�l��Q9#��ZI%���-b�.�N,�%�p�q���e�5@��6��\�D�+o,�b$̉��p��|��=l��jr{᯺7wGF�8���[^|���r�����Y��8����CFrrNx5i��)��G�4=�#���l��ۍ��R��J�_�aN�
Ϯ�盍v~��'�N�y@E�8ߧ�u���]q�A�ś�U(����H�����
1	I�j��݊��L��D6H���~��ba%S���J���ߺJ����}>��A�¹BS�4�4��e�!r�/$㎰DhW\j}G�J��
t�r2q��ٹ��ߕR0(z�ư�Mٺj%f.���ZBVډ��!Zd=K��e�"���w��拏�cj.
�!o՚E����I-Wj���y�y�P:�+�ZS�[^��FE�l�y����j|K� ��������t)��G������N�x���&��-�+&u_�uO���ڪ���Ы�&A����2��c��[)#��pe6�+����������@^X(Dz"�4�F�y��:Wȟ�D8�x!��cV�RX��R���s_~�Da��3A!�a�o�ӯ�J�Z(�1��ƻ3�҆^���L��^��T�RR��@��������tz��.C9q]��K���5�/ :$UA�d��t��Yp%���y L���������<�I7�a�T�x=rb_9�5^�]��"�����7�qLh�S�i��5
�i���/u�K���!�|���p����j0VB�r�����5�NND��C�S�@�|%�F>�����k,������f�q�t1Q����z'�;�7�a���Lp\7��^�I~]6!�z(�?�~xe՛��U����W��i��m��ի�6>��p[�&y���k�$
�1�c����;p�4hU� �>+-_�����,��/O�M��Pj�ps����k$��H8��X��O"%C��X�$�̬wd0��,�����zȨ��f��p��\�'�JQ��>=�P����'�Z8T�^�Z� T}��7��l;�!�/f��G� i٬�`W8 ;0�<B��&RLDz��;-�Z��X�[yׅ�5t������J��b9%J�HyQ!��0�T�� ]�u����ʴ2�s�b(Սe�]bB�H�`�"�4S�*�P�r2%��H|��s�s��5l�Al[�7�Z��[�jP�_��
0F#֩)<�����j�_d�G�^2M-oKW�e�ް E4[��g���>+��ؾ�_4�g��Њ�a?������Xz"y���F3S���ʕ��Z<���yzR~/U��o=l��W�/U�b�&�m�W�-��nf-��IQ�.�e��W3EV?lȑ�S�*.�Yv�g�`Ri�5]��l���e�YZ-LB�17���w�K5?�|�.]����쪢������9
�O�`x����� �I%ѸIB��}��+U��Я
L���M���̯��@Ah�t}�fFH�C�ｾu�p���94��y &~�g�_�S�&��l�dU�oZA��Q�ݥ���E��~_�%^$�*G���tNe�F1�s��Y2����B#�WE��`e�Dx�� ѹs��~ /)��L�Q��	F�T�
��{&]�8Ƃ����L�����̢;%���{%x[<�&sryz��6z���A+/Ρwo���@%5���%;�b��<hU����Z,**ꜘ��`�����/�U5�جD����D�x�._��aG��Ϙ���7jce�4v?�p�
�-F�Hx%3)|ͤ��ܽ�U0�璀��ږ��jg׭��Q��,��Y.�Y�LS�2]�A׵�������]���������"0�
r6��);х�7��P�/^�8
��h�Ù:&("�=B{��N���_)�7#����^�N��wXxT����r�O�kk�r�M��cΗ
<9*�5=�?G�Ӝ1�Br�F�W·"~ڥ�K&��k��y$��1)�$V%3�t�U5�����^�[�vf	�e<�7��q�YFȤ��Ck'���\%���+,|��?�u�#.~ҳ�D?wOEu�s��zשּՃ�A0c1��ʪ�����ӱ��!V>���E45hԬAo3��DI��MG���g�Z����L�b9P�\w��}K+��d�$���'E��"w��T�&�-@<0~���]k�}t�;��@7-��s>���G
�bmt�ny�^����$JK�2�F�P�q6���\`Ь��M&Ճ	��S���R����~TΟA�����S!v۷�Q|�hjq�AE�a�љ��p����k@�گ��-��>���!!k���	���3���%��:������8��&�z�"�ԓ���*+WOm��h�	��h�?ٮ:�#<�j�}��e)u]50���
��)�yEzp��'�04�� Ț��z-I�ƜYBQG{��i�FcyqI��B���b��ԑ�cQ�Z1�ssssyKs3�y|������T��AM⏯��r�	,1��x� 2�وzi���l�t�v��:4�ࢗ��mO�^M� 7�;!�	�+� �� Lj^���i����q��.&@Nc����b��l�x&�I�h��I��/�$��I���4�L��(��Y�I8_c��c~c�t�~ru��TM$F)#t��'s���WDm���)KN��]��v n�Q$=¨W�  �U��S�W(�����;l ,T2l^Kdr����/B���:TLSy\�w�tG�����<y �x)���+�s^�-mĶ�cI�?�R���Z�@7�����@K��$=�A�}Ԙ#��5h>}�Q��b�-���V>Fo�~叜ęS��ט�����U$./S�WIz�������k�Bkk�K.�	ul^���?FJ�c��ʿ/�D�i��J�Jt�Tɩ�0�#��m�֌TC^����f�ASL�b�~qHJkby��|Y�S_�mll�9��k��TalX�P���^7��*�-V7b��{�30H�6���Ӆ�ey��R����˖��s�f��|7�{:��cd`�;�O�I$��]q%RM�������ĈK��"Uʾx;�g����:��i���H���^_(�kaGܐ���[Ĥ_�ȩZ�@�!�����qC8}�9�,�����Pr!�K��7�Y=�n�,�`��b� 9�?���$��?+�ࢦ�P����eD�Q'8�6bw7_�P��6�ar�g/�{����W�sZ�οŗ]�zѬx28=[�6��ݥLk]uJ-���"�V	#q��䗊@_y>�)�0�f).�@*�H�ob|yQ4�^@ ��ߐ|=��hPJ��0��X4�l;��������M�򡉉��n��{�_����u�qyy��M���]Y��b�T)l�o�p�v�����Q��C=��i��H�����S�"#SQ:��%�U��?;�NaP����G ��#����m�M��L�w;���NB��u�<���\�*�ۉ�703��(&�Q�Q��,��cą����+���<�������K\-� "b�v7ŰSb2 bK~�rb����g$�Ě���Z��	&EEu��3���ՏA�>����J|.&+�򔠨k�+A%�͝� ��ऌ�|#�+�'���`L�M.#�^�r�K�Q�y��}�Vߛ�u��������{��@%9Ɣ1�ϟ�gJ7��$�-�Ʈ�9=��"5走㆜w#��}U(q�_*��mx��2���*�uR��1���H��zҭ\F����s��	�$1v���"*+��jvѯ�Q��gD����?�NI�sx�>�����0#{��Y�S�iwc��ϝ��h`U�.e�#�Ӡ�A|F�ճ���J���g�Z�A��(������r#EY	�V�|$a!����HFtx���c�ۣ �Ns���~�g�O./�JA�PS$
��x��R�F��#\�x�?�v�ԡ
�(���)ic�~䠈��1�U�����+�K���?�l�#�ND����@ٓ*%�4��Z1��B!�`�ܓ�b=5S��o/�/+�Q�����֖�32Rk����P����1<���G�	\0ц�G!HJ����;����g�9H�ndLX+:���^{�z�.�62����l�-��,��&�Q[t �07T~�OK�#Ϙ;����Sc���^�}6Ϯ/� ����Cg1����;���<����T�:1r;%�$������5K� 	+�4]�.����?fOQ?�z}��`�x�t�]�њ.��y����g�N�	��T~?�6���ڞTBV�1t+x`�L��Ĉɶ75���	���m��\�{�jkkӺ	��(��"� Eb,�=3�Q�F���\�=˵��#�}JHL^��A���ؠ�U�q]E.]� �?E��b#��H�����i��0�����LǚD�����$J�o����)0܈�ƦI"�˚Y0�	3~O�L�݋�9��g����3p��\Ds��aMø� r�2)��?1 ޽�$#�}T��Y�A�
�,@qj���$�G[��|0�BD�"w���Plem����2�/�'(#3S���:1��}zߠ��S�2���0���� <G^y{i9�P��lɜ�э%N�W]!{f�{����Z�*�d���F�(I~�.ǼZf{fAN��d�Ahi.;`��A5,�m�654���) <V�ަ�U��K����x����`�VA��/Y頥R�+Ml�v��0B��'�8�3���zsm�������a�=unjZ�pf?PM�9����Cl��XߓG��>ro��a�r��0`����ub&��2qV�I��?��C���fLb"����,���"�+���
)�d|��H$~��.mB4߻i9����I��R)Q@U�vJ� WÏu2��-�V�&�g>v�Y7V�$�M=8���S��rh@fPo*<
��1�`�d�
#�SPԎ���#���h!����A���!N�Ur�K��a��*���J�-�r)SWw �,N������|	H�c�Q���J՞��f�)�i�{����R�3d���F��Q�t��\`
���*��><�|�0
�y�P�M�݉��qݟY�n#pg/���$����-���}x�+K���M���BѮ� �yuk+.����Ep�a Y���,�{����'����0�yd�%}Mʹ���p~�����<�>� ]��:*��~Y����J�,�;wj��4�@�%�-�;\o}�İ�r�������{�����	k���n������v_���|2+'gAt\4Hj��e?���a�8��kO�=Z��[e�R�����s�����3c'�ȡHO��~���}͑���%96.fo_c��x�S2��j��A$<VTDU�ܬ�v�0B����aA_O�(�F������^:m[p��4#9�5ſ4���r�$nΦ�q,3��D7TÝ��BJ�|7�J��-�B��rE�pը�D~���p5LB��GD������n���.����4Z�TL��B�Z:���h<����6Ҿ���E�֖�k�/�����1�iBe/+�K�HP�vHp��bHE3T̅�h�mY#����ljjr=Dh��;�a�mw����FFE�:��٬kl4!!"*�V���mZҫ ���o0��C[A���,3FGK{X]��ݝv������q{c�CBџ<"r�;�@�$���]�E/�b�ս���@��D]��uA06�������uw�?����̓>- %&%}�VZ} -����%~����g��5mg5�J�����m7B�����g*-QTV��seL����I�%=f�-���o�s~�u���"X�φ>�{�顑�kSeM���dHQ��������
sCg���]Ɩ����*�^�g�����w]dd�7�I�í��_��e�0I	�RU`"���s�#av�1:���K����bM�@���{�~&`��j�����Ch�<E]��d;�?�Tͮ�����Uge��+Zp�����������Ù��[��v��hG������S�fo���za��G���_��߻�I]IW�6m|}I�4�:����g��ó��U���&�?�m-W*2y\����
��@B�f�/�ͫ>�75Ř�D�,\�Ҡ�������O���������d�)ǒ
�+��������k��. �����9���b�h�'$$P��ݑjh�w�::����H��\\4;x>�/�_��(&Z�cD�)��N\,,�O����qt�����{O�9?�M�?�j`�����g*�«��6Պ��ؼ7�������������ƈ�"8�g7\�a�%�i��ӧ�V����F��gE�rc�4L�����>՗>$�����!�m��#��~o%$�Ow5����w�b�"^XB���MM�NVZ�!A{I�M---͂�喑�h�|�cU�mmm�EIO\���݇B^.VV�eUUjzO������d�����p 9HK�,=����Q9���H��A;�|������^�Ge���v>t#� ZZ%}�P������5�FYh�����Y�+��S4�CW�<�=�4J�*k�}�"G�"'B���k��op	m�S�Ϸ�H�+/��f�
�Kԗ��J_+++U7�%9����p�~Xu$s�8���6}'lՁ�T/��z}4�:qc�����l]�>d�6��d1!r�����g~<��|b���i��J7�Cx�����;�hr|
w��?����:�����ӭ8j<��HW���q��-�y�.m=���j�//�[}-�h�W`�b�|��c���&Q�i+�4�Jr�P���������i��/mJ��.�:�W\2l���?����c�_�^xfm]q�8YZ~m#60WS_�I��m���!ed�zN������w�	SK3t���ѱ+&f�����]������lA�x�;jB��1]E��z��^��n|;o[j�ogw7݇y�)��;�#mCb��b	n���Դ�6"��%LϞ`�sJik�Ք��հ�5�ҘN���rH</��A�����`�V�F��%.���1P���~r[�A��F(�������q3��~�2��2n�(_�?;�J��"4�@hY��ST|-[=]�����p����f��4e��*��[�67+�p�kSD���@@�K"�kJ��.��^���\�d��-jE���x'2E�sP�?�۴��ԉ0��+>���l�eBz8�d���_���N��陡�Z��?9$7<��}��C��w��r�6�48$ע��1����e�+�A����M����Iu������og�o�y��666���=���i�q$��sKj[������x�]�hE��۪m1�<R�c�	��*���{�h�K�F����Kk��OІ��` �N����
�,���E��񾍍���ɬ�&��Q:::����`bAǠz�{WW��(�{p�$o����|8pU�qd��O�kb�G�m<ƀ+E_OG�*��[�,���Եm:�+���P��.;�e�\��>w2���=\F���s'�!6����l��\y�HB;.<�+jg�ҧ������-�:"БH�V&��e;�y/8��k��?���
%xcu�m������Wfg���8��o �x˺\�s\�wL�/���>�Z�y�"������]������Nw�&�¦�[V���gum��|��M{?]$��ڣ,�\Ώ�OmPR~_�MA @^sSg��K�k�]�����[���椙���p���*���0��MJ^��$2c��}�{��gQU��yݷݪWU�p�aU8YX\|�n�����b�l=�a���,��WVV4����P��'@wȄ�#S������IY���((�8�q�h���^׿g���0UG�3��ſ������kg�9����blxy�����^�
�>rt�`�������K����S���v����6A��0y��璐����3�k��a���o-hRnf�$q�Z��٣��OYW����}�Ȩ���$��`�eJ��Q%��q��v��Z�~5�P�U�/���q�}�"8p�H���F�8�-xKG[{n��&�B�}�ut����65++fh�.'%E}��������v���?�gd�44�C�.�0�7IÛ>�1Q����Z�ٹ�s�h�_KAq�'��c�k��ogS�����/�P]�[^�5N��������(v}�<�?l�{xxH{xH-�������O��Ίȭ�������G��u��)��P|_������6g�wK0��h`��oB߹�+�* ���@D��r��^Y��m�u�2@�����3�Dˍo
p�<��}���r�ȢE��:�FNp����4a�S7	�+.��i�P�dN�u����h<�k�d�5@^��׏0�����|���vgC^����MdO",�������+�"A%�}rbB�'�x$�x�o�gv�����q���G\,�W:�1����ٞ��%%/��G�h�?^ 	8Q����?M����eM0{e��v�x��������I���J�N�<��͇
\�J{ylRbFb�,**��8���r��Sje�2�~�Qv�����n?!XU��f�j<����%�N��Ɗ��#�E��ZY��ʴ�u$�	�\ ,�`}s�s�S�&"X6淽j�YeddT"��1�\�3���*eee-L	��ߍ���}��Ny��o~}5g?�&��h�G_Y�9����b���Sc;��C?"�`W}�+��'B��Ƨ��`۰9����[Rk�h-T9i�ຍ��,^��םͤ�"A�~� �uqv{^�pz�m/���������&jy˄�����\�dgw�
����󐅖��8�4�N6W���Ֆ�f`�u��6Xi���;ᖡ��80P� A�].�o���N]��\m�� ���Z�s���X{�������\!f$2�PR�`@���������V��\��+!����.��Fj��n��V��#P~Á��
 Tx��Ӆ���à��9���� �(+��kb�O����Ĭ�P=��H�嬮��GSU�ARE�`X����8� d���fn�����W2&���1���w+*oO�b�4 �N�8k����1m �jdɗ48���.��ݠ� #�LL�*^�q�H^I���! �-ϳ����fs��k��#B�����b�.�L�@�E)J�ˑ�)o�9�G{�1�Y+Μ���LO���7a��y�����->m���M�F������%�/��e�"@5��k:��	�i�Ě&�2�zz򼪮��m�_�]|�^�����\�O!�����iʅ�:�`<<=W,�R5TU�1c��+pcc��n�����Ա��{8a]�BA�Rݲ�*�ݙO0l�T3g�]U��j�F������v_/�]9߷����+���`-T ���-��t�ь	�oc~�.�V�����P"�+��o����f���Y|���m�ӆ�]L�49A�V�;��X���f袾5�JC>.*�cy��6\�΢|}}���S pk�t�C5J��� �o`l�m�ho֏�������5���6�ͷ|Poh�9>~��5b�G�.a_�,e�ot�T��Wl�M�k]-7�ܧh	iAG�2(4b���#f�_\�����L$�J���U
D�-����޹:=;�qM_]D�:�ST�?])�;��x�wv4D��B��zV))�G��(;㷭O�����_�A�:��G�S�KQ"��B�tt�_�ݧ��W�'��<����F	v`�������=%���Q�������VC�l��g���cE��aT����͂�~�+C�*M�5�|��9Ͻ��>&T$$v�h(dy�_:���w$C���Z���e�`'K��z��|���fK}��7AAI��e՚FR���@#[W�I�u]��*�:X�ߧ���<v�����փI�j��.��ɓ�Ԍ�:��Z��f3%�p��m�����t�{W�*�ߴ��`��QȤ��G�� ��O�Q����Y	�U���<fc�2��/om���8���H*}��Һ�����x�Q��,/o�WY#�'��r������o�؅�dt��
���H��חǫ�9��b�䬷�������[ۛ;k�V�5� �����չ9Q^��ԟg��YFX̦����<Y�mS�YŬD��t~�R��~�=qs���P����'t4��N��7h����&?N��,1nlb��#��䏌��nn�tttXJ�X�����r�"#X�'�@p����I{{{�Bq3"3��ӥ��[��$a�SS[���:���X���LÉ�	�3.n򖺦&<l��8X%R������)�������Q[�4�=��QQ�,�.)��޴��/�hm��ơ������CWK�'d���S{�����ΗrSf��Zn��)��j�{�ա�B�;��(�x��/���Æ �`5.;׀gkt4�	'η���U�����|�`���5X3�4޵ytW/�����U `b*AP~,��dbh��S�V��$_�N)x:�F+Ȣ)�����\�����uv����P���hX5b��sb����]����n���I("{e��g[�R��&���v�
��#�{���^����yzD]�%gCh��3H3���iGK�����9��e*!�./���_5�`�jhh8��=���'��غj�L� _[[�A��n6յ-�u+�h����U�nkS�.ƿt��Wmd�><��@�aj��V���J�u���{.���Uȼ��������[sva��q{���ͯ�����j-k0|��}��AOx���*��	 �aa�+�x��l����>Ͽ?4E���$q� �:�����N^��d���K�o߾��3O?r��=o�u\�Ki(�Ў܋|6��JX;��m4suăp5�.�h���z�tힾ�6�'v���W��!!����J��3��(vuu��V_�%��00--���/P����ն���k�^�jA�v�u�i9�?A���>��)>����$�$�8�YX�ٹx^����-?/,���s���UV�-*u�6�Ѡ��{�����nq��Q`RR��N�������J[[ڬe�ql�#�������#�i�)-���P�
l-������볏���A��*����\2vu�@���S�Y9���a`g7�����o?�kfn^�mF��B{͆��
"��w�(t]��7����Q�� hna=:�yp��X�Xxc-��J�4�G��2c�����;��*v���{	��ń�{^i�9�:{]_�E��k���sH����o* ���Ѣ���вm[��l�뫯>��d`��TϺ��2�҄�-�O��
�[S�
2Q�^�	*^
4���h�Q��Oݐ�{ͳy�N7��?X����J�Rh9��g��+�@��]���GG^�\]����?xt���������e�@��5��%-�-.?.��Ɗ�:����7�j�pģ��|��������ʱE������2�%in�������􄷇����֖���#36ր��ե���/� !jl\�o�	k�S����l��wdu���y������Rqq�P� I�/�p�A�}�˦��a���j�9Ϊoܶf�� ������p������|�+^je�?���l���"�¿���Z�љ��ۋ���x3l�d�B���,/��5~e��˙0�J��f�÷s����Q_g��
]<wPyrv����pL$A��N"걠@r�����U��j��>���h��o�������|M��S�>y{Y5i���o: t������,QbcM
^ǁ#�QhC{�]�44tMVf��n���=Y�{W<}��Ǘ���������F�b��eg�z{:���Xd�N����;�<E��'�{����v*;0�O>�hgT���9O�|\���Eꙓ}<h)!�H��9EDG���XY�o3��[��q;��z�5�JMK�LFTlc%����T^E%��5�:�1�y�~�y=ǒx�}�X��y�EK��tS�w�ᎄ�ZA]������M�F2>9���O+��B�C����w��ÿ��s\ޠ:שh�$\���u<e9#^Lq���G�WG���#7�����k�Q��V��F$�3�o_se��H&���Wg�o�s�;�(���;ݝL@�!�!)}�m�e�#P��.�L����+EJ��)���)��2�QT*!��i�Ό��ˇ��~N9�����)V�m�+2:8mev���[kw�����\6��N�����y���C�F8앫�b������-��r�}%����o�\��Q~%6��~w�}	���̘3N�U"ll��[�dh����G�ݾǺe��-���ׯ�>������6���4���d%���4�J_z;�ll詰6h���l/�uu�͗�I�'�N*I�{<��՗��BC�fg�3y\��H~*G�Lᦎ7�n6(��D��%C/�����4>ϻ���0F'3�eR��6̪
�OM���8o�Vq����n"h&>s������zy�h*�󰊂�"� �`��x(��P-2[&7u���nmi����|I�濱�ϯ����o��`QK�Ι�q�X��t	���y��a�W׻�`����-�CX
�?�����ڽ�>�ۜ�?��T	��!�_�U@DB�ۮ�\ml�8�i�¼N%�N��&^��`i�:��OI�M�����)����"��t�C�s&��-��Ј�}�N]�1�@�O��S1�p��)�{_�P�$3^������&J��w��mն�j�p?/!"N>��0��R�y��~IĤ���kǅTS[ԉ�:���ꗕ;ٜ�W�ޤL���+�b�B�ϩ���,,����7�%�tQ+��5K���\��k�e�f^��x��;3;���o��V}���Q�]��{C5Tz��մ22t�U[�����=��-n����tK,<=�L��^���6�NOOYE�~�L�y=P5C����K�2q�H�Hx��'߭.`�:JLL�6wR6�}��YRB�WS���|�E���F�3q��$�1/(((�
�����$���e�����km)9��e�a.��O��@�V�326v��O��l{A}/�B�g����J��np�����)000$M��~�쉣�Ĥ���;�
{���?��yAG��./ή��Ҧ�e�v݉邃�B ��v�ѥ�����N4�F�tS���4��"�Ēv����qr�I���/-.҂k&Qn)tv~>���	L	3���P�!8��� �稹�n!C� ��M?Un�m��,Ĩ�Ԏz�f��E��x�h�g���d�����ܙ�u�cq����s(��v2qL�+8qa7�Mՠt�*ד��#;߼�WIo/��N=&�?�B�~I��w8�<(��/	����k���Zd}sX���D��������������֤�����+�g��j5�d����<dN��S0����n����ŀ� ���外�>���b$?���y�M]}��e�ܪ��r��+Ѻ.}���P�B\t�'���$d��WF��slA^^���|��Ä������4��.�g�%�/U5�K�����㮠��v���+Tfm<���uwr:��¡��T�o���#37�pZ�^��wjU(h^���f�wa���Z�˭|R�"����/�
e56�r�
�liY:t�(ӧ��2x8��
wh:�y�m>�JI1�R��:��_����Y���$�#!����3$^�� ���������$�_oZ^.�gl�� }��D]���^�̖��"ڹ{��T;�Yɡg��Y�C�(�n�I�Z"6&.v�������b���O�j�^r���u��l6������S��ɺ�$O��ǅ�ɬ���Ħ���ee����ʅ���Fu�d�c����{�չ�]s���yxYޚn""��U�~�Z\	�����M�N�:I@����6�v��E>�����慂
ZN� ���ˋU��PK   ĺ�Xq#Q��  Ț  /   images/bb187b5d-1fc4-4a4e-a882-8dc83b4f659e.png�zW%�u�[S��d۶9q�mc�o�m7�M�&�fs�]�߳ޯ��9��v���42""����
��p7�QΕ���p��v��@��C�ң�C@dy�J��y�w��ُ{k��	�n�ct�c��^�%�k��¡U���)%2Sࡥ�h����"�c�D�@$�)cR�lYؒa�CT�6�MW=ߟ��*}{+�ms�.�+�Tk4L��}�Z���U������+]�ע���f��a������J�q[*��N����8:�����Boq��_=y=_�_��ݟ�g/7�s�Ұ�B���ؔ������6��{�?��_��`�Q^<���4�6�(������7(��N���v�[�M�,��9��-y��}�|��I_��S�:�7�c�{�;>��rFV���g߾J

"�5H��]|�ɡ�gtQ���z8pG�����~Z�^�%��y�
}P%��9i����q�k��]s�|,�${����u?��%+Ξ�_sp�ޮ������mfp;;��!`�Ä��N���m�ʊ�<!��N�=H���^o�q��h���hm6��"�U����ãgY0{(�:��><:+��yq �	�_Tc��H��j��WQ�
�q�/���e�T��bf�7�����[����6�?O����P��:���w�O=؟v���p�%75���h�
�E(�?!`�բ�"}��S]w
9`��a0aL��ה?��0�w�����'� =�����(�1ꟜѬ��2�������xI	�J\'e$�"��#�C{�KJ[Cv
�=p�?�<E�)�`M���I��lʞ���zA������ߧ���Pg��ߨx�����׍���J`����� m!��O�e���� $������4V�pF���͇�zI~���b��<UU���G쾽���BT��}8$�~�{se�%�ۯK�T}�81�B�s;{�ݚ��#	Z��'����J�X�U>���pU���qd��`a���׶›��iw\;<j�j}}����Q��������M�#�������U�G-��|WC��%=�y|�#��g^��p ~*�.o^�jnЋ��"�|`p�ˉ?�	�0��jO�q��23		��?�sx:���I�Vϊr�_Ð��R���ؘ��+�V�T�`f��B�=J��l�.$u�&O�ё`�t��?��ɰ�zLYѴ������+�d���hn�f襣#fH�ZvL�����VN}yPnĊ/˅vx����a���v՞�o�O�<��� ��a�
ۥ����^p����x�=����d���ۗ����ba
�g?0`'ᳱ��I����2|�F9���1�䵣Z=�?U��+ݙ�\ 7�3���݇���߶
���Is�kS[���s-����ޫ�[��/����|��BRW4(]�t�,y]�e�rw�cɅ�;sq�hw�$��3�u&� �@PXX�����G�UoǪC�����J�c����uM�o'n�͝���^8����P
=ƍ{ۄ���k�&����w�*8?r�a{����t�Zi\E����Yy�]��z��7h](׌寃����1����G'r�!��-cXm�QAo�{��֭oM�Xsиx��O,�]{fd\�qSW>�79n�n$)��}�s:�2:�n�?�o�,�4�i�ٯ�-�퍍��;:P��ٱÚ�z���[��Ao̝�-1��ds�c�ұ�Ҭo�){ȡ�mw2���|c��̎�"�4�%��]��n��Ydp!/��J�Κi77�X� Y�KKw��6��7��"!6��|.<}�ӟ=��=Φ����W�)`P���)� �����$�yT��&��Kk��%KK98��3�6^'(���Q��]��KHjesv��x�,��͍�o��G�-"N���
b/�L&�V�P}����r~bM��V���N�$�[p�u�W�_T��:�ww��f6cS�G���������ݝ����?ꓟ�J�*3��|;'I��b�c���v��]��m��H"|���~K���8S�Q0��ɱ����~���8]�u������Ϥ����;���xkA:���:B�����K��O1X�÷��^	�a�t%����sn"a����i��f}�K8t�o��S��XhB�d�
Y5*����BB$�":��<8w��D�=O�2�yx\��G�I$����x�/ہD��I�7Z�Z��H��>�E�O[$-���3Na$�C���8����#(df��f�Y>�-`. 5���b�0�s���6o5~m��,\ay���2`�Bk��d��y4W��AܙX~�S��?[�2�{�tH}�e�l��Y�j1�`�������:��c��eh��R!iV��rB������MH����)}�ygo���~5}�0>>..�S2�I�M��`<9�i��s&/���������=w����>sN^^mkg˺^�~�z�w T����pN(L��DV�m+m���W&���_F�����VA>>���Ws�_�J���˭�'�}����������,*�����P�gؕxۄ��q���|]��i��j����w}�v���"�%'}�s�p��J~�||-r�?�1N�������q���I�%"	覸��}���뇦�B������-�3q=!5����/��_;�]�G!���v[���d��_����7�m��.V�H)A^����9'И)4�x��n���~5�u�a�ھO5�ݲ�i<�z��qix�vSRdf������8y�d.�X��E%~߁7���&�\^u�5������/�����u17W�-�jc�%���ˌR��8A�<��RYTΈս�͊�S�ݷk�,�ux��_�nH�'kVD{�̅��p/��8�.����+b�R|q��(ߋ�ȓ��8J�Y�ܰ�?κ���_|0��o}�h���7���ŕ����{�of��'�)�\5�\轸�dU�.�zǫ���ՍKK�Ԁ��Q���V0�xl�9�<�
aZh��!�Q`�G�P�@"6k�,��>� 
g�*�k��@�rm���7�֤��{z�O������~�2����͌|`�+I*�BL�|}\}��	�[�����,������&9���ه�5L��%����\���o"Mq�=�<U<�!�s�)�G�w�5
vX��ڵ�v#���M��#x	-�Dw�?'��D�(�8�C~+|���`n�ni�}����Ԙ��Q����p���n�D���V�p�
��xE���G��Tkk(�c�x�P5(���D����Wqt=.��������)th��8U�d�E-���a�'��l��-f�յ�F�)B~WJ��!B
��埥9ct :۝آh�e�nû[�
�b*M�\�a��P���n����������Zl�T{����f�DCB���}�����sՖ'�����l�H�����Tj�A%㱗H��f),k��))7[�Ҩǈ4Hz��>��a=,d<-TJ��ċ���/,�qli����� �+�պ̗M{���]���e`��K�Q�S��wY�Fܙ�W,��ʠ/�K�B�m;x:��+�?#N���i�\`6)5�~�����t��ě�n{��h"4kd���7���ɸ�)�������n�
:�T�2����^Q������8͎U�{H�մeifb��|��Tc�j������W�c��Ɠ�U��-��\���`��Ϗx�W��4�b{�A}�Zk���!
��g#�G|Qά.�?���;�:x}r	⺍�85�I�?Y�EN
�W��g!������WE��Y�1^3F�2�(/�(ф�,�w��7����SO?~��JFG�ڍR�@�����O�>p3��m�VO�}�x,@"�eT�e�H��s��+?E�Vo��u9��5�� LT^1
?3@���k�x���i��uj&�6_�x����$���NŬi���d���wO`���r"�v�(�p���H�����^QQqÎV̸A��8���q�9|	�]��>1���z��<���ub�}g�:r�s[�<Sh����j�������w�w~����l�&�Y��yz��{%v�m��,�pgZ���l�:(�|���yM���7t*%���0X�xE-�8^�� ��fc�z{��rIf���IrQ�xʶF)���ȣJS���9.2l���hߞ�?N��mo�D>
�t�����?��h�����A1�ZWg�M���BA,gps��DY%iȮk����GLCD���=.YY�
%޾E�N�3��a0Na]cjݳDcxe9��/��S��\��Ŵ���x����0�{P��XL_}9<���~�������u���<�v���pK}�99���M,��Nl�v^��2W[����D����q�
�E�2eC�~cR@/S�!���r5� K�!�toB�5�3��"G�h5�M�0eϛMK��+�G��<�l �g�ws�� �ꇶ�m���w�m1xw��W6��ezq6�-��0�sȳ�����'�ji�h��J�����J���ZA�N���>�%��E@�g�c��a��9��7���y�>=Vc6�����{{vE� �<�~G�>J�v�HOLLH�t�)-|�T���Ĺl�5��1��lgL���=�>O����|SO�+B�7������	���u�W�y'��إ�k�Zg:D�
�d�Df���B���Y��vM :0<B�4+�:�?�yZ�C�H���&ɀ*���?XU�\38t$�Y,���������և�-��4���Eu�����A�*���=�6|��sCD��%6�&��g���!�$��2*xEЎ�J���
������F��Q��������)m�X��*�e�?�s%!�טM��9e�jN��z��њ��hz"���]��ʏ,�ʢv�3��:r��7�f�##���g�N`���ý������A�T5�1�����+y~G��q�I������9y�\��"���purE��~��5F�l����o�r4�S9�u��p�^z/>ykM�.����snp�L�r�n���B��9�{yBR��c]���/��LF��	��~c����5�,F�y_H{m~dc1Ź�!�|Ԫ$�aW2��N�e/x�����MPx���)�>����U�c�ؘF�����ro��|�Gb)/�IT�mG�F;
y��sz���� ��zl��|�0���~)�u�&��}+D��ه�	pm��=3LlM|����ymF�+8/#�z����|��)��J~L,�@p�h���I̳-��`wQ�BT�*�[{����ڍ:���~�_v�av+?��53�-��\T����Ͳ|�<�*�~c�^��PxL��d'���o|s�a�H��0�*2���_��� �#�58
�{����a����S��R]^�L�fG�������M��W��5�*���z.�$r�޳�ì���bsoB�ہ2�E�v�(Rp�u�7��ǌ��?슇+e�
1Ow=��LA�����RGb�F"��Wq=�P��.��#���WCR�������e0��a�UƊ��i^����o�
[UŽC��H;���x_�&�*}��[ն��)���{]#�1S|�f[<�h"���S�.�F4怄���n0O�� T��L\��v���W��"{�Ա�I$����R�{�c�9�����N��x��)B�����}��b(@p�5Lװ���=����6�NƟ�38)q�� =W�煀iEhp���t�y�_�bLA�����~��ś%�Upm�o~kv���d�S ������
$���u��'?�����,2+h��o�a����j�M�O�B�e3=�_w\�C�l�s�����9�.9p���d����$x�eM90/&=:7{��oo�ڶ��>��.l�򂼫@{�۟s7����o��t�5��Y&	c;�Z�8&t)��W&[����&@�QI��?����;ƖR,�த���� q���q'}S9���ƂF����O!���͞�n�??[x�6�Xo��d�}���C�0<?z���S�|���6�q����`�:�w�UY���L_����I�&n�C����&Sp���|OG/�M�v��my<��#E����l��ڎ��׮�ĳv��&�|@��7Rg�i�}���N�3���r�B�j�U�"��b��7u�.���8��E?�h�x�.�E����l�f�y���q�����@: $�}-����М����B���:���C@�kd���˃QQW/����*כZ�@U��� 6�r��|YٰP��e �����U4�w�����m��c=W/z?~dѻ���L���We���6h��y ������ς��F\$�m�b��ġ*:�4�j�_�o��j�����u꾲�}�s���0���#'�Ӣ�1'���x�c�T�/��ń��x�@��� .a\Թ���)�G���@�Qg�����J��I]��*l��ezQ�8&�x4��<(����d�Ǹ#T��3_�V@և��8�♅n�ú�;��
Β�@�� ����?G���L,��T�ڜ�h�Y9\h��X�ѻv�w���v�"R�I��7__'d��A*i0�S���]����6}������P(����鱭�>��sǞ�pd^Ŵfa�8)�j@D?7�ey"��t(r�0P ��$��|�}�A:�ϡ	9����H�Z�B��n��j-���z����Ֆ`���0|#��*�)�������+|���A(U6~�-���h�~�����myP�םL0<mf�͹sF ��g���c@3�����J ݋H�����^ �x$�^6V�l��0g����<a�Yv��U�DN�a���9<��;����-e�j��g
82�f�������8��:��4Dm%�Y�wZv�>��y@?vNNzE��b�`��(rOwC����J����	9p$�io����}P�HK&�*l���<�����L=��Y)��� �d#/�����T S�3/�� ^�����߸��W3��Îf%oT!W���l	E��r�&Gh���9�f�ȟ6C�pg�
�v9��jn�x_��Q�������O�W�-�?�����Z�_bJ���*��+`d���7��H��I��;��,��*x=�w�%ԣ��<�<���f��=�������;��%y�[CU���{�R1���fy�j'N)B|"�]M���U\�+�dw��,x�;�5~�8����4
:)���2"o��H�po?qR�-5�f0fX�|���z�W�QD7B�`E����o�T�mux��H�bG��|Z�d�;����N�u��oawO�/,���Sƍ�%!�L
��0�%���n�8����i�Py���8Y���D�(ρ��	m�v\�1�|hM��U�Y+	F%�^��F�S/��)c�Sy�C��3�ix��eH&20i2 �Ę���h�`f5@�=�����BOd?Lm8��܃ml��G����-�܌�˸<A�>k���r�t�9���ʭ[P��=~�_e3�gBr�Ǜ�jNd=>#�e7��N
$�,B�n>S�-]���23k�OY;��X,�l�h�_�DB��������4d&j��&���^������j:d�g/�%K?�]�V���C&i;"�E"j3��X�AsPDʓK THtv���ձcf8�./�ٌ��)Qz^݋hVD�,Y������#m����5����7�5_)����vǃٞ�B�)g~�T>����w��e�fH����ĀbK7)��F�*M�B`R��x���Jթ����SK~^9	��,���>��h��FL�W�v�CaߦBл)�6g���3��Q[�QѼ��.(����V�BXe£��kt�Ϟ�g��ܷ�<&��h�c�&45�u�,8ʻ��p��9��GK����a�(��"M���{w�Qc��$��W�8u�HR�ʻ�r1fkTib��Fvm��k��G�z7;� F�x��D�=�V$R���zMx�&~��ՇU�q��,����l/�'sG���8۷[�w.�t"iԸ�Kn���rhѢ2�������ѹk�Ԓ�F
5����\��_d�wڬ_���+��� ��`�j	9o,TC��B�)�����x�XJ#N�["��l�|����d�f��1�5&��W�o7=n�ݒ�zdŷ��G���ء��ڐ��|��s�Ǩ��tܛ��mo��x�S�+oyg�30Y\�F^�wbRB:�w��o�D?����'��*O'��T(c\u�Ʋ^�Hz좐O4�f^���ڛ*g��Ӛ�<ug3u�q�MA��Y��
BR?��6�3o�W�c��e�K���d��p�|��<�Z
�B�9Ӎ�zuI)�[V0b+��b.8l�Z�������/��n;�u���*�$�	�q�ב*�ܿ��-{ׇ��v��+�l��-FXs�i���|_$w=���{7ʻ� �p��}������ǎ������qfY��L��UM˭�8������j�]}�Q;���Pޢ��W/
�y�>��Q�f��0�@�~*"8	5*~9<<VU��M�_}�Q2��-	]�;k0A�Bۢ�*W�p�Oy��(4գ��~m��ٵn�F��hp���N��D20����d1�h
]�hCB�k[J�l��]���k
G#B���tc����e�6=/���&�x��U���wV�Ǵ* ӭ�5�����ּ%y�C�`�������e'�g$�����HՆ���D!9g�?Q���D�o�	�3i��V]��fD���F�f��~�����kZ��*߂o4x¡�l?�U�l� uބZ��V<��	�^6BDq�����ُ3��GY���� Ee�6�mi��pP���.�
�6�0Cy0��LO�Iu��~%��R�&�f5�@e(�fc1��8#�7ɱ�~S��%�&� @�+���%��.�F��;�_�qC�_��g\a"�E&�È������2����S��x�k!�ݮ�����[w�x�ۈI듲���i֕3�_����-�r8��T>��AA���N�(���#H�F���:a��/4>�0�s���¶3&d蠽o��`���5,�F[>��$Z����Pt�3	�D�W���J�����F���_��e��P4�в��7���r��n�������و�;�ꝸr��b�d�t�3"ң�y4\�5����/���NN�R8��Xqm���LN�f^�rIʵ�5̸���"� H�gC�lwٿ�^��Al��N�z�D���9eM4�6lR�D*���ʝ>�](�8H*��� �~�����q^�9֜S�����*սC���$���7�%y���̼T�.�6�A<n�GR��w�ڙ7)�AA��ȳ��`L��S�J����������%��5d��֥��R3� �ML�#�ZG�a�7��vp���6�y]� ��!���9+�k.~���G��ˎ[B��£�43W�,����F��9Ԝ�ɭ7��1��Ɇ���OG��]��";���9�3B%g�m�q�-�Ϛ�o�ݱ�'r��v���ͨ��i��M��`���FVV�;aR���`?3e�
�#X

:G�B�����,|�QAO���{g��F[����Ҩ���Tf�0.Jn�B�M��E^�-��Ԅ�>"+/���?o��t3���]�3=�9����7�Z��}����k����
��ޝ���Y
\8v��%;�f�;���^�?�}�?��(Zβ�����q���Rl?c ��s�&h��N����%�aು�_]�h�u���l-K��F	���A�`�4u�����5N�4��b�����f�I���Wc���>��uQ��.`h!Q6��>��q���\��h�Mۤʛ�5A̄�*��s�k��ew^?���ө�Z��l8�R�C���e����g����4�s�q��j��2�V��"�iQH�(E�����Cl�c`��R���id�(ċ5ʩí$>�1j�R��z�QAmu^Vd�%�����F�8A<�$�zĝ{�����1s�~CR��-7g3�$0ʉ�<~�������0Ow��H�p	��b���!��V�P�q����\���ł��Ĉ�;9L[U	zg�jm ӱC��Un����mUחa�Z~?v�F�q
λ��������c?q��N�O<Ύ�����ޮ���t����`$?��R�_�	<M��=d�H��]S	n��V;D�bIH�|�&^Iܨ_��R�����k}Fbު�h����f�k58�h�\�Cz���ͨ����`�[n_����2f��?&o�z�Q���� o�����Q�qQ��Y�F��[n��# ��;�Gݔ�ɫ݃e�8���UZ�3ג��g/H�!�qTe��
��~4r�9���r�v�M�������y|����8�,pQ�_8����\�Ep$2���&v+��V٤!!�P��j�]E[
��
�����*I����,��ʪ����@q�|�H�b2f��+h0�lpE�q�̵����K�(�N< L��Y�C��]y46)�v�1]}�R�z*�)�2k���]�'=�w�T��c����_��-N�l��a�;[�+0L0�˞����	(�����L��rjZ%ksյ�PӛU�7_�m#���`�z{�~2�|�~0�߯����	�<<���T�#���qFX:JreU9}�h�~�}!pb@���G��g����
N�×�f��p��A�8yy��+l���ue��[w��[�2�rm�:�>Ɠ��9h.3qBo�%�В!��h7�/B�ػ��\���_���ݲ�p�U�kDՊR�^V����C�y��?d0�`9��Q�P�sH��� �4���H?����?�q��}-T4N�G�����}��ᛛ$�e�9���#���S<�f$)]�Z�� Œˇ�F�-�py%t�b���������p_+�L��L9^ܙ��!�岟ɹ���m�����5D�*�9i�š"���~��V���j���"��5f���hd���v�������@��9Y_�-�V��ů_�E)�4���uelc��q��Jw�x�r�� �0������C��� r�yt��C���x��Aζ����._.�� D5�w�[�Q�$X���`G�����yղ׺�p�U��d�P9Üąv4�v�)��4;���-*'?�r�n�Qf�ߥG���!^0�'�d5f. +"�h�+��ʊGj�bC��Y��Υ��Ի�fxs��Q�6�Zet ��(/���]|�#�c�"����z�F��4�-�4�~�_�"l; ��D��m�5�S$M��2Br�)�yk8&!e:�5���j7F�3C`�`�z���j�D�t{�#�h��Z�ۂ����?��,E�Ҧ��JlU������R�O��<��"'e՞t��h����'�5�ʻ'�Qw�ӜU0��=���6�m/��A��x�@B�/��䒶��)L�o����
T�jY���GV����w:�=]�`)�jy�*��ID���B1g�cS��!�72eO����<��v���X��P�&l�L�iݳO�����>/�P
r�+j)fܪ&����|�Y�:���"ߙ�]����g0BC�v����"��D���FVP�g$g�7z�� �Qͷ�30T&�9�495�K����ҫ�16y>�;�s�Q�l˨��HҎ��K�]����և6��>��g�&����a�B! %�y�]���B.�.����H�D���>������Cq0�M1�B�i�3a�a��?���'�^_��`�M���&�r�M�8)��')�P���E�/$�"����=���+�hB<躄5ξ��4�r����ow&��n�=��tEj/#*��e\J���/�M�LB����������Y&�������<��q=A�B��&��E���ي��8�@p�ZR��ˆ����3��'=�C^\[��0�U��ke�������2�=R���k݆i5��L7�lL��	��M�`����p04�Tf.\}�{:��7{L ��b���u3���IP��z����%�łɵ2������+����RH�Ӈ��KB7��Y"�L��.�.i�N�u��+��r3|�-5�Ȥ�$�½�^��#�p�r�k�~'}'j`ei\�4�O,�r� �d)��#ץ��	^1���F�?C��ͫq��������t�D���^wA�/ʙ91Y��{o�S��57��'V.�����.�n���$��Hu�%���V�8��o�|�;�ET����̪����x<Kuw��n�%&	�W�,��]��%��!���Kw���׺b���Q��Jx�D�'��%
}v�a���C��FP}6r2�L?F�u?��戂|�B�I��k�X24�)�`��D�[F=����vT{�'m��īU���)���#]�/�&��y]")d��M(������5�ٜe��[����~߸���'�q���d׋�&g�������J�v^�zD5�*|tV�Q̚sq���'U
�`���񘧲w�ͻU�T�4����]4�	�l���@�9-���/����2��r�*˾"*0ھq8�-f�8��Ϋ1�#����U|x�HY	����Ԭ�z�N/�8�1gd���Ŏ��=T�<:^�\���t��n$&jdD�r�@�[ҐG�}x=�'8�<,���~���"EPk`����<�R_�mF�������������d���Ժt��b��������nb���:?	@n.>O<{	T0�4e�ll�Bӏ>���GEq�Ė�z�̙-�xv���v�����&G9���`��8��=��bygd�?6��'�TMٝr �U��bv�z���}6��2e��|G��H�'�Y�i���Ȧ'���H�]gO
Ц.5Z��ӧ������L�؍z�������7F���:�����##(fk���8nl�c)��,[.�:�O�똋z!����P��dI�����~`��l����N��"��A`��'�d>�>���Ĭ¸�۷�g��{~�d����/MR�;�z��i ;Z�d^Z]����?���F��d#M���߀��iG`W}��@6�\�{�2����k�F�%/Kۯ�_g�{(Rt8� EUP_�x��0g�J��n��&�8�O)+��&Q@TRpH�����}�KbN]Vnq�e=��F"1�1�:�V~���6}Vέ]����٫EP:���c�$�/�E�)��:Q2�0M�V��`�qEn����3P�;j�
'�Ak��M��p���uYu3q�����D cN��N[�]�f\ a�ʊI�h��O��@k2��J/�����c��F�qLb?a��X>������-�
���Ն�<J��e����8#�q�X�Y~<���A2J�z/��f�U��b~�M/&�s�����}?�q���][;J+@��x���4ԛ�&�3����	:��(��W��*s���y���s�B%�8h�k2���b��~sL�~�Ɂ�-(�'��ң�?bw�}�'�p�m-_9N!�Vw,z9������bg��dQz�AZ��L�~�;�jQ��̬ʀ�]wG��O���+�y��{},LIR�d�M���콂���L���;b0�NAVNr����R�J�:-ֳF��]�9��)�;5��ކ*UH�1uڽfݭ~9d�D"�Z�'5��Y�&�63c�I#�"6&&%���L�"_߬��j�)�
��P<`�-pb���C,p6u���������i��):����eǗ�k���|���5S��A��{o2P�<_�q��ve�k`��?�����&^�sQ�<�����t`��m�r�2�剂�6g��#7[)�>b��k6�W��F��m5+*�؝s��s����s��)��$2"�K��a4�R�>��c�u��95&j�}�9����ju9H�kܘt��o{fci	�vN����Z����S��y�ҁ�NV��VY������$�DN�T��k��:5�`r���?�� �0A8�z���NF���͎[�ř�x��%�!ʜ��<k�S4�.$4]F����y��?�%3b��*�|� ��q[V"Z�.�^!�R~?��WN��Q��,B��c��b�t�7[�~i�������iN��L�l\���?��iD]�]��Tk8D����0�����=����/��4��r���d ����1:�X�[�������xm�C
8���PEB��o3�ͭ�Z�윘�7�+�api\�����+�f^�=+��HD:+$U�	J�GkI��H�P�'��=���S��ϣ����D5�w��!m�u��5c7O� ��z�9(�9��}Y:�t>���%:k.lE*�xY�8�y3��*�oz���S����4c��B�-��6(�t}�V<��Y/��9��9i�T��s���FB8L�V�8Ep���;E��{V��=��	��%��_:�tʺD�#Ky������.X4��p�xΨ��FX.�a��c+SW�
��#
�I�4�xlA��a��\[o	�S�s�X�����������u�"70�?�a�I�d;�g	� Vk"Wh�_�����B�>[%�{a۴�9$mM�"���7����v��̽�:��u^_�z�}s4ou��t$�]ʢ��^Fc�s$@aw�s���J����ΆrSߘx^�M�s+ݪ��j��1a��
�j�p��v�9���àt�j(H3��y��'��Y���,b+z���~�&ˎ7nfo��hz�%�#�xay]�6Ƨhz��Te}O"��(�<!?����H���n
�ɩ��|e�slz\ƍB/U�c�,(�
�C��/�?�}jLt2���i`��GE�Rڟ��0t�WD�ښ�wx#�Z]RVv��ߜ�����G�2����q��>5�(��&���A���N�#Ƿ���al��� �Z���)T�<9���PF��S��i�~CF��>̝ɝ��u�����K�+��r���x����T��
)�w�j`o��`9��
��f��h.�b���+��6��/.9 De!C7=����I���< �X��Ts�@�T؀ZI�)	VlaL_��s#R6�}�E`�0�XȔ�uۓ��h?���$�%��?�di�`���2\� �9<�	+%v7Dj5<GB�d�U���PN
��?zv�>W�\�FK)O�ac=+�?h���\6�qO[�1�
�������-:P��a1ޫ�ݿ�	�#����� {p���'�B��-�-Z�SG� 	55��Ԥ�+�q�2�	��N�d?�ei�������f�z~qcr�#�07���� �60a��s��`��l�VȀD���L��oV��X�.�rl#���۠�4,<q�NNr��|����aL��2�!C���/��ś��z~u���k5���KF�N���ِ��d^�Z����þG]g;,}�M�Ղ3i�D1����<��f��\� �_�l!�ș 8-���I���?�r��y=�W��%�,)�NY���?��@`�<w�������e�W�-k�����Z�gJ���3�b���x��/ѾA�4{vi�m�B-<x9���N�f�;��Q��8S��H,I�!�<b�awD� ���$9d��x.�w�o[@i���n������G8p�f��A�@�G<�\�;l-�Y=�y���T�BS�ĕ�u��L�tQ�4�x�Ŗ@�<VR��=r�m������'���ȃ�G#s/�l�W��W&OV]5�j�>�B(7)<ِ>�դ����L������ˀ�SO=�s��x�tQ`f�N�Y.j��J����X�q\tA�.��U,��G�h�H@Z�Gw8��'l���6�Z4�?0�M��gF�.����E!s��&�?���Qj�?�u�T9�{)m�q7�/Y2鱎RKYǙ�%�ė��6�[d1(��JP��WA$d��1�QFl�m/��f��xzõ^������i�y
���+]T@Ir��b�� %�<�U$����|!7|t��rK�@���H��N�z`��T&���/�Iw���NY1�����`NH�y�T}��v�*Zk�=�a?�|@}�c�+��1�=h|��6�X�e�gP���xni){�����~�*�7o�hQ�@Xd�K�հ(d������ @�H%�J�v�s�(��]�ĕ��v.d��r�ꪶro��[�]�s���,������p�K�跡�U�Ja�ϲ��_1$�4��TS�e� ���+��X���5⽩�t,��%���--K5ċ�������]�1RZ�`%�J�����%2���k+�-!��s� DS��m��?�g(��%�!�c�����-��]K���{wx�V� �>"��P+G���ו��z���s��}h�L������E1�c�~�q:3|#(�K�j!���!%�pI�����62��+1�Pj��L�l�ϤX%խ�u_<Tb>�Aι�N ;P�J ޶l>�1	��sc2�c���3@Ap[��;��ۮL~�+�!��!���<TT�Ѓ]�W���Sj���i���ɾ'�X4�8HX24'bv��+�:���e;JW�@�-HV��sSI�y3Q�%�J�7p"���i�5K�������� q'�e��j̪S��|�Ƅ�5� ���-p4l��R�h�<�3�����!��9�{�"�Q�I�ʽ:�D�����Z�-e,,���Q�"���M@�b�I� ����4��I-���T)���(�,nE0�]�)*B�p�4�O��=>qW�6��9VA��u2C$%�/n_L܂��Ń݉N�����]-Ռ1_�Y��?ĉ s���ٮy �W6��eEK���3&�=츸�
�(	U�DC��5	�-H��A�]�%��)w"�g`Vh��qi5엉=҆[�AC`{	��~�*�	?�&d�VH��՚�	�iܖ]Le����Q�|B�+��@'�0�&A�ry~�<B�J6"Ʋ�n�D�
��%����9!G�Ҋ���#9���a�D57��x� &W������o���F3މQh�s�J���7D���a7/B�sT�Rr�r�/�9p��������@_�P�%���#E�>JF7}	�7zq��a�!㹐��R�'��$��v,x������i�4���-Ϗ��5����6���V�SLdV�pf��7<nAP�U�b�s��BE�PW5b`��-��(ݴG�5�<��m<c��X�fCCpR4?W@
n��d�DV-һ�������M�5��i"�$��,�5�1e�F#a.AnAϘl��u��Ȳ ��K��!g��-��f�ڹ����~ �a3��,$��I�~/��,�&	�NK�G�ȍ
fޞ�^���d#{��a�G���|*��a1��d��W7����)�	E��ءTa)%��'ȩg�>CN��	w�eKH�_"��ۺ�߲{�k2 ݺ���$A'�@~��5���`�X���&H,M�y.�W����;q^��Y ������� 0�!�6M��@�+��r70%蘃�V%+�?�p����Vp�9�_���p�@}+��k��1������K�&��P&��DU�:����ŪXylPD7�M �?ۨ�.�gA��0J��DB*���!��r.f"I*w�Hi� �_���JZ���?/Vn9��Ĥl^��[�T6���I�d��eu��(� d�Pߎ�+�?`r��-�䈰��<����*WG��ebr�W��`R��ٚ����:�9�R�B<:X����՘�<f��RJJƈK��=�~C.�/�K�=v,�V���-E����
���lb9����*�Ƕ���nW�y�^p�j����3,�B��@]���IE���X�bE(��i�|�Q�%��B�0%�b�Y��,��.��L�=	�sI�m����М�(�+��G)L��TT, �
�B��g�	����I�� ��n��q��m�^<A|<��Fꮑ����0)�^���y��"s���pD�@a�==g���R�Ǐ=Ij*aaY]A�V��y�����)���"���-ܰY�9-�7
̅E�MV]]\�����Ǡ���1�ԛ��=�W���"X��
BO=��߻#�hV��r.��L\ii��C5��t����k����aR��1eB���M���vY�63k`^������lEsYʦ9���ca��
SEX�I���QT�|�������}u�&��99�F?���D�y�]P�
ώ� ���d������&>G�BkR����(E������fB��|!ދ1B���p]\J���k�>}��8����F^  �C�ˍ�춌L[�Z��E���� �:��e��N]�VV?w�㚶/�|^�2c3�`����ք�w�h��b1�!��[
:�|��*�?��?�Ms�
~jA���-�ў�����xI#��l:H -�̌.nn�3z�WLbZHvW�`�]����u%!(.NϒF�����i�6}uN|����ov�բE-�����ݻ��Νc6qV����S&%�,U+v�d�ȃ�n�k�l,J
��h(�.�w+Z�@�՜5�e�O
!Ø$��X��1�
�m�������]2��*�	aѢ��f�gh����e³*^����3�1��`� >9,�̴�����#�"u8fZ����n� �j�"A���\[C|�<�&g=�~���<;;K���\�"¸2rQ!aq.1B`���}\�-�� F��H���ɵ&x�H� �/L++h���iaSlb���jc��kt%GZ�$w�9�^�I �^9� �1����w{M�՝��I���}���w�y�o��ֹ�����n�-ip+��]?l���)�X�ЎNj��.��L��a?x�����#E�y�c$"Lzd�Ѐ%�'����A���n�|�2I�Q��#�0�mx�"W�
t�ك��?��df�{�]���_s�m�Z���K�#�ƸwA��� f���p����\�_hCxiE��%��	D��ta%/�@����Xۏ�i���}��۬�I"0!�n�ҍ�K��/�>}rʹ1x���q8ǂ�$;g���8??�>�H�6�i���x&�!�ِ�%!���z���Ǐ�Iŋ��[ T9sA�|���g�gݓ'O���A���)]��ӼW�$�d^�~8KTwC�u��܂�&8'�>�GNǊǯ�@7�o ����������R�?�����1�81�����<��%�嵫����|�����~��_=u��n��ع�ãН������n�R�;@ �շ��ۑ������=wzzJ�l��4&�,x���w=3ۖ�M~{v�$+�����%�z�dV`���k��0蘨�XX+F�4ځ��̈́���\�}�YP�,Z������=��w<�������	�/���K���x	���d@x�+����D��kY���"��C��s_�k�b�����TGZԮ=8�����	"��U��%A-cs ��H*H��kԟB���b��CG� �32������[̗��1~M!��_�g<;���������?F�X�'_9ڹT��<�R�׌���|��78���{w���l.�J���B��Bc^N�F�K� ��'�Jq7�����Q���ǡ��	f~�y����\��礜:+�A��?d!���Hؼ�$������t��Z]'"<��)�����!�������^�s��7�|�S��Ԃ�����*W�Tmi�@�]�5��d�ҡr4i�5��������9J��1_�z5	~�拽�������=z�wDj�%k�K_�?�/��|~LVLHxG0�g���ɬ-B�wb�wlvi��1�Ek�Z4q��F#K�W[f�_z�%>�	�X�*Xs�}��@��-��O��x��i�s@����Լ��%0�з���s?�s�*0�q�y�H-y>����K�M���cWL�����I¨� ����j�4)r" x*_J�]Q��1θ65�2恹m��o��j
$�K���*3��X��16����#E��8q���V�q$ ���=�,�z��T����@3�gװy3$W��զ��3a�vu~�&�ӧg|op�3G��|��o��Ί���ߊ=6��q;�J ��ݬ%��g5:A
��]�¿��6o�//�|}����?��/��W��y�����l9�רه��!��)9s��ɨ!���VXx'�.	�<�̄�\����R�2��sQJ6��D(5X����kK�rA����s����ֿ�c�x�|	.��Nb�.�Õ��Ъ��/\��X����½X��R��yѢ�^��@Vѩ�jy�<z�N��|ȓ���0+��ѓq�� s�ms���@(��?z�򕯸w�C|��ߗ�=�J��&�=�����/��3�S�7)����Ã���{J���Ï�o���م�Nȵ+�Ű�7mH��c�f�ީ��0�	Ǣ�W�|=z��h�N�V�Q�eJ���,v�&��!���%#i\��#�SӬ��m���\����s1	U�F�kv��_y�e�3�#�仄B��'�q$%	}����3g4N"�#)�Zb"C��_��	Q�l�IA�MM����[���{�٭*$��rj�`	�%�����W�T���z�?������������z��OUP����ޫ�~p�o���d�-H2�V4�����%-��n�"�O ���'�5c϶������D6U�B�[�-�d���`��g�M2������=�� ��~6��ÿUb�Hx����1� *1� ���v�����JK�᷸&�T��acBk�I�z���C�o5������1�%cpA]lU�㱀��űc,&+�Y���S��Gt;vu!U���\@�m�E�𛝚K@F���GZ?b�@�"�!p]�2����o�����.�����_%w({*��3&s��Eh����r�:���i�����~��iH��s4�P=9R��S���E���������?���ޭ�y����S4�.e���B��gx$�/U1lt���q�^�c��b�iO&�	]�Ww��+O=������o���_��ϝ�T��������o���ߧ��EN�%! ��4���j����=�
 ������.�V�C��(�Q ��{ɵ�yW�u*T��\�����"Z��p�H���?f����ثZ���s�[���j�*���N"��]Zt@;������r=*ފ�;_XnA�u4 8�kX�;�J:��	p]L��'ց�9��({@��'�?�14�"?�5Y��l�ތ��ia�������9�n�nX�K���u-����\3/�)�:����P��BX�m#�1Έ	@��%��?���k��0�f3�Ğ�:/�+X�zv�q?�*�ǈ�Ģ�Bqq���*	bo�1"���q�"���_F���������*���cx�v=�h�Z��=��#[��D`����J���&����~!t�;�^fD�q�$�����+�J6?d���t��N����^@l;D#�$��$������'��_:_�����~������}ba���|�;��JB��{��������o�wۙm`�("�M\@3
Q\¯E����	D	�9!Q��q�����n��� �a^ԕ��v�n�H��J��<�9G�-W��==;�H<f�!���Ic V�mZ�.�[amSI�OU��� �*�.�o޲�b��`0�Vc_y)(��}>���G���Waѻ�N5�P�'���q�"r<6��?���,��T������}�;,\�5�EF�ޤ�q���+�&h~ˀ��ؚ�❡���;'��UZA�t��l�B��~,��z���U�H4�"l!h�G\�b�/N%i@�V+�k:x�D�2~@l��g���/��!��Ya���㣻yY s!ݰk�����!����W�ʮ�$G�+��dCW$4ꕃ9�s��;�{O�*�<1x��0@�4���l@�QKBP�y�Q��H�~��G/�$��������_��_��uA���/���;����G��$e_��Z��\���z�q��X8t�� �H��n/\{�wX����`���[ ʌ,��H	K��:M��`)8�s�h��9n�w�� ����G��V������0T��Ru���@Ֆ5("V����sp/n�vŻSϘs��y�������ѩ�t��K�T��8].��EA)��=�ਞ,0�x�^@q=s�6�>�����Fb
Ȝ��"i�֠0�r���\��:qyy��\){e�(��v����]+���i`�T%�/Ũ��:νn����S)H��	�q�8zA�r��8��#@9[��-
�H&���2/�]�h�d��Rh=�Q0��x��f��`�����6�xW=�!ǣ�8��Q)eOO���f�AD �-���'�؍��L��BB��S3����X"ke��@<����Ǐ��Z����

�*'�������~��Ĝ_���� K��3�۪`c 1��ઌt��B�
`qyc@?+DSVi��;��.@����5 By�#���7g�7��;�& �T+���ث�C�t1$�s�eǨf�[З�.���f��p.Ȕ���C�(��%���M��Ԋ�b�lv2�,j�& �d��_���uL�Z��&��_�٢�]=���h�'q�I�LhQ�p�6=���Bȝp;���\���q��X��=J�l�ZY� ��ˢ��}�WU �r�&oӀ��Zܶ�Œc������GqAb���^�W����+jd��V��^^��킆���a�yd���Jρ�.u��x��%!�vHׁ���E	�%	&��HC�� �J\��ìW.��|B3�8�	F��4ϙ�%+PTlC���C�;�
+����/6*�4����Y��w��âH	e4 +�?���/���������������ӧO���W�=���fW������Mvv$  �x1�"���D�1��$!(7C��a��\aP�э��u1��J ��9�� Đ:�F��n8k���y�@�u�l�Hظ��Q_��x|�f��ژ�	\��J��$��&qrg���r
F�c)��_�R$��@�Zc��Y�H����Rk\Z�@������/��<��D�Xձ��Ӣ�q��!h���Ǩ��H�͕���]��21��r:#��X��T ��J$�lZ/�.�h�tC]͙qVq���!���R��/@y�^ꊦ0t(�ݿ�՞�����:AQ�\4=��e/H)���u����ߠqH<b'��B=x�jĢD)��i�}L�N�ŋ1NF`�K�G�c��/sy��]HG����m��¸�I&�P�gI�Ì�����Rvsm�{w�Xʴ��'�f~������w���/��/5�ZP�-�귾�����=��(T�oRS��B'Qy��u#���U�M>h�5��b&���v�������pYZ��U���3��^�g�y7h���
H�˷�2��rR`֙[�q�' ��"�&�;�3<�
M���5"Pσ���g�@�ެ�#(YkI���\���v��˷'���|�XX�m-Q�z��}�y�"�}A�<���(D�k:tZr��j�\.]��\�*����%����t�i��	���Э$-�b�ut|�J�Yy>#�g:��l���!&�>.䤂�!e��,�~���0��WmȲ�`��P�&%���fڍ =�*(*)��:!��R���a
�ʯU�~�i!ĳ��������w�u�&�y]�ۢ��`R�Q���Z"���K�@tKxɦIYI�^�Ŝ�2��i|�V�-�/�9�o?����>��S�>����?~�o�-uW`[��L�xR|U�,���%��ʾ1��%*,x���ZAZe�v� m��%0Y!�l�QLv�R2���-w��N���6��)	W,hj�oh	�N�ClZ���j�<Lv���1�.��2��� T��ki7���X�s� g="��۸�o,]KL~.��O���|1T��}J�o�
Vs��q���x��|���`��a�Z��5�1�y1�84�>�B]�����̄+�9U�(��
�����L7n�y;6_@*Kq�˓�1�;]̗4��Y�T���>��������u��4{'�P�F����ܞ��B�1Ac
=��R��`tÂ��B:؎2K��tW\�$U��+9�Rj����+�.�����*p�(���7R�G�*�Y��}�S���~{����௮�W?�?�*:3�����ф��=4Z�:�=���K"�،�!1��o��Ɗ)�u��6ь�1������')/�Ȼ��rա�L)�B�/i�����p)??l�+��e�Ba�5��܇�{��)�Υ��S��}2��*F��] � �k[捅'[��K*;�B 8�� ��QJ�I��O��`�a�������]!�pQjlJ�m٫^�x����Z��_���cuHQ�T'3�0�>$de^�r_�-,�z�켦:��~��}A��~�]�/�<`�x����P�9.sI+�sT�����kzT�c"�I)�"V�\Q'�yYy�PUA�?���6��V���}�x|��A<T\�(F�z��]�]�z�ir\�}������՗��w��o��7�z����Z�vۿ�4�QZ��BMP�d5��:��:?�s���(ۥI����"�e��Ί߈6��uV��Ќ<�4y�+�e���b��W�'IQX,�ƙ��� �EʅM!��.U�<l����.�9���'TAW�@*��DMKF�L�����
-�*U�^o��P�-�(��U�3����	�^��@P�֜S��b��u�D��9�ꂔ���S0�s\ժjJf�;}	�y��\��$��ݶHE�Y��R�'���I���������f�
jC�_y�Nv?�聢�e;��F����a�ЗJ�RE��"��躀:)��!�;7�<�E`�k\�\={x8Ƅ�gTT%a���9�X�W�o)��3a�A�NÐ�<�hˡ������Led�`��ܩ��_>~����3vz��8=�J29^nۦJZ��g4ᛐ2'9��`$���Tr�|m5�<O~>l�{A����Q�`�d�e�R3۟�X7h
ל�v��\i�Ka�᳝��t��CWo�jT�g�w%k�vt�xC��Sa�8j��pl�Fy��E1��)��i�ȓ.�Q�����
b�#�P3����&x[XbE�^EۿK�Sa�,�B�fG6�z�n;�ۘ+Zq��l�ll$���9}44$�7�/��~TTf��J�n�����E
^��Yu����5�͙aZ��3d��A@(���E�I0_��I`�����A�B^2J��=��pQ�3#�S�����.t�\�V�4�	�_l7THg��v�"5��\sR7��>+�c�dr��n�3���\AA�?��xB�l���i��Darރz=�*5�ڮQI�%;X n�y�c��-��T ƍ%�W_���	.-��lw�T�,����ITlV��TP8�O�6E�g�ڢb@�U5Ho۠�& ���B�&�ǂ@�P�,L9��YNA)d�����~C$��w����X����tk ������6�ObɇJuj��Q����8CN�T(��A�;��mMc�ַ�HD�L��G9SAaCr#�"jQ��;z��E�[��n�,�Zd�Ҽ�
Q�n�H��DI()�!�Y���;�RW~[K��V���L�ɥ�O��}b�;��Bv�������ṙ���� +�qx|�qG^�P!�T_u�&�B�, �IH��)�+(�ޭw���t�Z0�)��K]��Ն��ه�U��m<�J!I<� �ԭ̥_�.&�b�%~&(��)	�-(80>�4�1�N��M8(��V=��;"(�D��H-R"��gh��uIPX����������q�r��g��
�ڞ���n�� C��֕������m����<��*<S����^F,m��G�R/��PC�i�H���I�BP��WXА����������Y����D'2;$~)�}��X��Zj^p�`�5�G�,��B�cO�f���Ժ��� ,1Y!�!���Fd�ܔ�=L%o�@�����hj~)����Ȇ�"���^E�<����y�FM�aB���q.�{tpTvϒ����~����UU?�q�Esa��3a��2@����H�妃8�b)�ދ>myg����&�j�:ۖα;���3��P��'����s�Tp�^�X9���	֋�@+RqTa�-��I������A0� ������jz3g=�l%o��F�<?��I�=���k�5H��ݘ�b4��p�0�J1�<u	щ=��k�I�B'��d�&
��l�����UGJa8F�:��7j�E��j�� �&B��%/�])�j�%����f�n����P���mR2��9�ʉF��i�K�E�sݏI�Kf�3��	
_J�>�d\^q9���h��(D��n_A̰�IJ���;P�=�W�@J�����dV�M�Y<@�
ɚ�y�J���� �aym9q���)�5	�͓���(�B����!i�wh��
��2�"U�쾱�kؖ]��iհR^\j����#����`ȵ��G���ԌI�x�����U
~���R�{`�nߊ*D��&�ݰ%��@J"4��e�V�C�L�7'��	���xa/�f4���-�������^�-C�3a��L�a<��w.�߉_ᔛ�֞�֍����c2�M���|y�M�Lѥ�\��RT��C
{�|鳒g-������>E������鞫��a���e����GΝY���;<:J�&�X8x�:q5H�M�KZ �ْZ^(I�Ej����^N�qb@H���QLV��i��<K$'%��y�B�j�\><\̾���{F�DqE�<�n�6�	�
=�7YZk��fn�.�pXG�7K���i�T����~t�F`�潉H��b�>��iew&N��¦�*Z�q���%�L�
Q�� �zK��0�_��`~X( ���K��Ω��CA���p9��� ���?^#զ�
3?��6r�4��QCN􅡟�ס0B���Cz:�&���}M�d�u^�������rf$��lI��y�8������BYD�d!	���*I� A�bx! ��I�0�![�Вi$Qəyo���?U��s��:�CIV۩�h�y?�}�V�W�:�;.��#|e��ؒ����#�������|���y1B:a�XO"fZn{��ɬ�� �mf�K��[+J��Z#mci�]c�6z��s+��P�����$�P�<,�PC��S�wp�G��#[H���\aM�s#I�[�>����čr�}�!��$�}B�?P~�����a9��~ml-4�OmwNP�=��q5�'rtt����?��|��?{����t��D7���F�q��J��N-��T��.{*��]>,p�]�g�c������~?LR�~��&�?�!�Y�(4�	�P�q����]��)�������`��$�u���B�r�"��ċ#N��l=�ǰ�E"S��xkYaJ���kI�_p7��;�[�{9&�m�a�ud7׃�}c��q��V�0�/4&
���\�!F*�<"��:gS
Q�XJ��4��D�(_Ij���`-�\�4(xK�̏C��������q#DT�D q�6��2�}����Vju$�&tw�Ӎd0�w>�w�����u-D2Y=N�ӏ���v��k ���_�P�ߩ�ӗ�i��z����u��w���_�������Ct[���s�����Wy�wwb��=F��=c|�1~��y�����y5�v���jC:G��$���%����o J�R�|����s��$jK��O~p�`fs!�d�7]�mx�9��/ J�|�Q�?jLF���L��O���E���[��iD���WI�Vt�<���٠��N�tl;�4=��|�X�Z�1�$3�	'�!���v3\�X}�}�ِ�织{���Ҥ�ۆ�$t�7���bEb%�{�ti�^��9Rl�g�C�ȧ�ngh�Rs�7�޺��z���֦�>v����p��������֙��_Gc��lY�+��U���&_��=�O���+D����� �&�O|�ݗ��������W��?���~"�<����^n�?-�=ypv�U�<��,����(;r4����_����x|���3�we�>���t03l�nOo��!��C&�-�R;��'����3��-\�H�ס�3՚b�oͶ��{���m0x�'>��*1��8�K�ܮ�!1%�J�x����K�V�--~.���(���$�kiC��u��K�l����-%�����m;O�R �U+���|�llɈ(d�`A�ck;sEl��@��/�r�̋�B���ej��P�0ڧ��8i����<�m�2��F��~�:r�-��ykX��O���2'���]OV�w���7�W�~�o��/�@�'ң��'?���_�����w������By?Q�u$�A;.�w�?��DZ���t��I�D4N�L�ᦸ���� {)s��.Q��]�NƷ߃ږi�c��ALſ ���k� �H�B�ԫ�z��i��(�����b	����R��c�n�W���B�mс@���ud�I��%���`������fX�I����i�Y&p��Ќ�c��Ё�������/���Wƅ*�d���gŭܦ�6�.(a75B)!�J�t>e�Q��([r�%�w���ؠ�bE��2�L�XI�����'�o"�%�rs4��R�r�fǾv��y�B1�vs-ǟ�Z`G����sG���9*J�q!I��#�s��}U���J�e>M��vQ�u�ֵ����k���'V�"�x�3��̿�:��D�>�)G֘a�ې���H�Z��l/���)��,|�q��&�Ns[�`�E���";C���s]0����Yd�ꐃXF�D�)��*�u"&h;�&�!���tȂM��Ӻ�6}E����IO�7�X�O��Vð�[rH����[O~���o3vc��޳���v��O*�?avcC>�5\�
�:tu3�	Uۓ��)�.��!F#V$�f�VJ �ZA5���,�#�I�<��Lf�K4��gO�� f�烖�����9`��j!�#z`�CR���6�rJb�b0!_�� *�����߃���AG�y(GO��3�6tG�������EH�|^d�kU���I]�4��������WO�w�������O�ӿC�-z�}��B���]O�K`�0l9��\Vǵ����_C�B�ܞ����ِM�v�E&�|/ݟ���n�h���)�48[.�qj�ؿ�J^*\����A�Ai"+�d���2�j:S�	��,J�	"��)�'�-���i:�4��c���|(�I��ٕ��imp���B�u�qa��(�,�Ɩ�U�m�@�>�Y��� ����v��n�*�R8�~X����K�����{��`��kě�6������w�l԰9�}�"\6�V3��|+�Y��{�uk�4�cj:B-���K[v]�X�!{�P�4�,�FR�|�ւ|��k��y��r�U����{`C]R��3��ƶ�1[��N"S���\�'M��G+�m9ݖ�c.s��i\���y�8��8���s\e_�{�������wO��߱�����{����w�~��o���%"�ҍ�I�_��<����%�T,���*��Q�#��W�5�[m�^bc����m��q� Q[�ٖ.�o+�B�6�_T�Z!�����8LzP�2\b+��-*��i��L�5�n���5<����H\��e��'D�H�$�H,a'6��w�k���rpcwG�w��p:e�e���$�t?_�D�f�l!"W$DG���k6�v�`���$���`!�E`|;N@�� �
U�t� j�&�&R��d������X�D'��?Cc#Q�O%�'���}������)�� ֪��
Z_q��%���!���D��9\4V�p��#rŌ3�*�W�:����?]��B��ݏ~��O,�/�������/A���/~�?x�7~���7i����z����<K1�;�G�=��A���vk|QA�O�m�`�\�G�/�x2���h��Jb!S�+;'ş�CòM{�=�Tt�]��Ƀ�����LL��%/>�G��W���<�����ՙ��j���N^c����]���q���.��w���|��������$�ɽ����(1>M�?}e���	�x��>�Ey:Ty"V�$���y�@��Z���V�!�k�5=��*d��sY�?E%0*�V�	��H(y"~���9���C�ҝ�9�bX�n��Ɵv�!�s��a"E(>c55�c9�Q�zغ(�D0�M�ީ��+7o���鼺�37n�'�E�X���S�a��:��+4�����Ƴw�����|�Z,ϒYx�h�4�R�JY%8�jA�FIu���6,�����_�����q����b����)���bX��
c�q��轉�=���V*���}��Ҁy��58�r�
qU��EKb�t������b���;6��xQf��+;�`+]�=!�'!
�I�k��J���F^3$)5����d�|��6:�\�q0�N�_/�+���.����������ˋߩ!~!�E��ߧ��D��������y�)ǘ��/܃-��2m�JS�x�A"�ȵk�;��w2z�wqx��,,��zQ��ݪ,��f��G��W�}��w�ί��]=��Q�1"�7>��Ͻ�����Fs�ߟ��_��� M�w��rk�^_�戦BA�6�4�����C�E�q1��Gw�G]	�3!l��k�Cx]I���yٶ��_��%�`Ą�L�E��LO���SjL�k�_���hB� ��^;���B�PˤH�x0$j��4�XZr�>�.����u�u��ϕ���U[�I������80����i�)��3Ix>�)����얠w&?o���>�v���d2�s���Vp}Fȕ�D#N)&��Х�5��d0�3qy�ȸd|l-ៈ�����|�w'ճ���_���%�O�R�"uۣmv!�o�����")C/_��~����Γ�eV�ɲ�ϒK��'��E^�9K�O_x��9�?v�㳟��9}�=�I��Gt�*"��W��Ξ=�w�w}�m�+4�pS.�cg���pr��C=/�v��d��B0Ԙ��(Ϲ��.�b'���>��Kw//\�ٷ=�t����][R��Hwd�.\�,A�킒�	%�r}�]v�}��}���0�~��I9��.޷�1!Ջ�du�ǐx��o��͸���\�]��u|,hy/G����>�NH��߃�[fd���v���G�/�8���X��x�ؕ����+.R�;���mr��C��;IZ���G���+�K\ڸԭ�,9#��^Y�w�"�F��_��ߙO��:*�k,��þ���E���ދ/��5������]�X?X��~9{xr�����}M�=K7�܀c�8Ǵ+���m�i�H�N>(w�%�;�AR���_�@W����;��W��.:���'�?))���f폾�Dî�lRߛsb��Oi��˥�l��t��3�t����C�&����kz~nӔ5]G*f��>�C����8W��/1Op�<o��_LCm������s;�u(Ix�;@d�l
n�&��j��8{��+ǽ� ��F:��=X�a+r+��K{�|$/ �#��)'������A�	�5��L*W����X�cL����x�C�<��׳�|C�ΐ1��Y�7y�.�<?-���<+�$�|uRU_/��������r�.?����JT?)���EQ`���c ����o�������$����Nm_���d�X��b�y7Y����ih�׾�L?�IR��N�е�,:�Lg��%n����:��Fk����h�v|�@��m����T���Ś��󃕽�kw�굯]�z�ߑ�������;;_�ȲrI���5=�;O��֛q����r��b�����43d����f�z�z�)iR:r�,�0�]N�V�5�m��'����������&%�\;��p=�-�j2r�Ak��>z�$E���w���1�kL*�$B4�����8@'	t!aK"��"�|\��h33K�Z��m-Ww<�������V�j�#"�P{���J�E�Yj�V{�Qj+j׮U{S�������}����h6�\�˒�`5)�L`�T�{6�'��S�D^�Z��Bߐ�e*#�^���J�u�xdc�d��O����o��\߲?}Ru�Xm{\:��(������LNj2	�<�{ǮLeI��s����&���"k�?(J���]#�1y�Qb7bT/u��9��贁�������T(�^r��d�D@�$�.ۭXb�RL�K)\���#��$�4nX�z_�ݤ�]bٖ��\}���dAY1�AS����l��¯�����E+������?X���1����:n�'�Q�;����R�P��?�������`-'8�8<I` �|~g��~!��͕[E���K���P"O�������*���ƫD�gʷ�G57���m�?���mR����R�ws��<��Υ�TNά��/Vq�v�����Z��y*�t����&m���0	?k7���ǆzr���#��e��2w�☪�{��n�h��Mr�xM	�\����&4�k��,ϾW��dG��Ĥ�O��m[`V{���"N.�)��
�AE�Y�2=&�����Z(�B|I?����<)A҈$:���N�G�\�u�Iچa4�W��D�.�L������}���X+�(їՇ��@w_^�ʀY��r�-�\F��-+H(�-ToQ�a=j��*	>�����ӼK:�����8����[��>���4�;{��ΰ�|��OJ?�X��x��bD��-&�&/���W1A<�`��X/��7������6���n5R6�.��&y�g+�Y��ؖ*�h�y�v�ف�����u���~�2ށJ��j[�G/qk��m����ղ��(�X��_^�<i�#lZ�I��P�(w
�����F4}Ub�b}���F�x}*yc������H�;�q�Bс��R�>�$�*�K��.�ƫF�}��,g�0�<9#�|��q����0���ưąٺ�u����v��M2鰍K�Xu�����N�O(�c[/}�inth�e;�Z}�3��ۯ��xFZo.w�b-�<�.�M�y�ʹ�S��3䤆F��%����̯��v�~�}幕��{oNom��E
ր����e
C������I9������d�l��[��:��w��N<�zRJ�]���v�����[��.���Z�p��Z�2-�����o?���9���F}��c�r�`��D�~���q��heu��n��,7��"D;S6��Y�뤘n����l�~�$\~�k�}bt����v�.+�bɰM=�j��cy]ܪ�ԝ��~]-y}��]^�LZL�W��/���˧w^���Cd\�mJ�c��Es+�.����������ʒ�!5�J�/Y_W�W+_�]'��U3%Rσ
��4'�J���/6����R@B��r���fp����ʱ�kX�&W���!U�T�H�^��������y��?�0Sp�D4���gK�k��^P�_��t:K4>C$O�"/Ш��I�]�e�S�-ה.��Ɔ�����u�=c-RL���?��0 �A\-����y��X�`pr2�E	��ާ�I�
��;Z�4q�*F���"Q�����|�[�M/4Ʌ��	FBI�۵��x�_F���JjS�"$t�r]+.���;�J����B>�+Q/�ѧ��t����$S13�=�rӚЫ��*^�=y��=��t�6�рM�G>7�d�����Å3v�$mЈ�B@M#k�ȅV��i�c�������	���,�uǹ�_R��vk叿DRh�'�jeR�g&B��?���gT������F� G��H���H�J�K�n�?����
駽I�v���s�4vﾲ>;�.��9צ�KS�\�:]tG-�C�[�ck��!�Q��<<��6�fw�i�z��U���[���ٍ�d�,��?�4���F��mT5���א��\��l���k8�c(^��&XX,8��������n��Ti�3�>����K�J#��ݧ�m��Y^+�l�-6�,�/>_�m%x㘎W%v�P(n%��~J���b
2~��_g�H,$˲��8-��X5-쓘$,�e*���a������~����꧜�,� kA��R�%:4U_��/Ȥ��hH�S��{2�c><؎\!�7Q����eq�-8�,��$��1�F�>�sx��dN>J!����ڬ��N�[��[�"ʸ��p����a�����n��i�����\��`;�G5�]N���^߀- il�$^�Jm��"�I��?3�*�m��dfR5��|7�d�xmjJbm& ��Ӈ?!r�\�B�	���;9�|߅2FB���I���za*y�� ڋ9��͟�e�#	���b~S�q�a?��a�+u�Sj��b%*'�{�	���}���t! -�R.
"�ź�}~ndw ��������LJ� ��j���u�tYP�Fy�ھ�ە+7sBCH��|�蛊P�эƔ��򚪙\#�ȁn�����_�m�it���D� <�B_��؏�<�)��6f%�~����/+�I��]o��o὎t����0�Z�������|��0�m��f������(�����n,Lsn�Y`E�q�'�U&�:�'<�_�#�s��]�Q��z�El�m�Lmf
n����k+�݁�Y�D��;�%�������E�j�+��˝r7�v�?���;��^��,3���Z|��r�o��:����4��z��5G�f�N"0��.놘�fQ�����A=c�Q�p�'W�iT�X�uzt��Ը��I���o�N�s�r,%Ն6t1�������7���5����𲳮���[M�c�:�1�2�D/���ߺ��ZI��CymEMb�i�4��ݫ?)ݦ��~MB�:��霅W���E>$��`���j`�Võ�e�V��2Ne9gMz�S�!v�+��NlZ��>K��OK���U	�Eg[�����������!&ۃ�0��Z�S�mk6w�T��D����[�lU#5.���2���(�˫{��d�[RǬ���}�<��'k�H����#�|V��Ypu�Gz�_���W���)��x��+jg�`�|�0I��ok|�WhF�\?�����q�a���0�1�d%����5:�$K���A��?Qȃ���xZ�=�C/�[E}�AU��nP]Y ����8����QU@�o�~>4bԴd��H_����t��'�۸�+ǫ���,w!�L_�|Gko }Wx�	�j��ʊ�T)�e3�;����m��h�����Α����v�j�1Y�_+�~oWA���2�+�X�,K��.���b�l?Ǯa�q���Qx.z���������A܌]Q��~��6+U��j�&A���QI�ì���k����s��S.�]�*��������\��ٌ�AD������?e@�ik��܈�T��3�n��N�k�/���}s��;��?��{.2>lg�/W8i����vmt��EF��Sʨ��W��-V��H<6�l�$�b�
�d�/-R4A�l�O���������^�5��\��߲�_�o`�j�Y{�G�})+n���]�<ߩm
�����l���{Q�j�1I���wK� y�g\l1d��ͩn��>��AZ���'B��o����ɃR~�-������[���L��ļr4����ư�{��DpѺrA����}Մ��'e�'���c���r�"i.��D�@[V0�M�x8���q;��e6�9��#o�8�U�k�����:��F�.
�,��QW0ii4�O��5����|��Vz���t�+��V Q����Y,힟H��U?��n.�Uy�*ݣ��&���)�I���܁h���[�A��%���1��
�S�c	L&��B��st�@�͢	;�J�_�"}d���\Y��o���a.�Y�:���PϒHM���?�з��7d�hU��̇f��$Z9���w�Otc<�)�W̬�.}ՈF<��I)��@�����5���Q=Ca>�#�F�;-ڼ��$I�B3)_B?НFjV�\*4;[єvR㪓,�RY��r���e�z�ż��$�!L�	0u����<�p>dO�����y�W!d�oa6{�-H���4�B�x��8@ ɸ�^�X��������`2c��ܷf�i�XS����b���}�#c,�����ׂ�ak1\�)�N�%�zV��q���d�e���$�%�f�K$2�2)>�K\�(���2wB�#1���I���vU\�v/��~������>ar2h�L�c����;�nS�u]t��h��%�O��$'Ë�
����Լ��4b�a��3Azq��o�d,��,w��gk����l4!C���5X��Oq�l��K��\��Ԟ�L�4��z\�������ae���d�T������
]!W�x�,\Y�j��*�������L0v�S�=���|�1�E&!eNm�;	T؈���Х_�!���m���$�}����iԥ7��yީ��j^�� ��Te7k�w�l�A�wU��$�>bF���$7���z��'W�Z����A��	�3P��jV�P(BREGF>p�����RC��I_���4y�'�+�-hM��vi�tf]����&�	Z���jꆄ���{MSٍרܓD������Cq�ƞ�fN�o2�|z�J/�:戣���	�,��v��@���vw���dr����b9�Ъ�Q�u�Y�P�tU�?w&#��#eG&�����~q��YUJ�'�L�č[ی�T��:-(8�Y�0k�:S(���M�x�d�|�LlP�P?v�h�~MSl��tY�Tּ5z�[��(�
\%{��)����(VҰ-I}8*0�3��,�=��{���t�=-#����Nk��
�8�F}�a����d�>�9u��zz�=�g4�����N��}GAs�ڱ�T!��;�Nj��2o�_��*��Y<g�nx���<o���@����WRt�������r�� pL[w�Am ���tS�?ȯ�ȇ���7� h�&�����tc̃F·>�T@X��R R�meNz���z6r�v*��'�FV�1���K������֢��m�d#EB��>�'ț�Ҽ|�.�����W1b~
�B<�?����#�����y�&�����R����L��q㼅%
�ʝ��ڋI�?DH�LZȝI�N`ڒ5x�2
:.U�M���d"ߘJ���I�F�	�p����JD��X�� 2Yط<j@'���*�yv��6�_��r��}
}o�@����و��J����z�-��`v���)j����ԕ�LN
���[�Pݥ�ec�ɨ\��8��3��7\2�������|d�ܜ��he�U.�}�����HY�T2j�/��OD¿�
�7������K�t�;�N�˂�����cj��L���i=W�W���V�w��Jo�ye�RN����W0���x�@�����QȒ�>�n���Z�+�}	�{|�_�!�`�"o��1�������v��S#���:=Y�Ԝ��O?�`��2 �M�X	3�Y�n��7�G�)����g�A�#���0l;l�YɞH)*=ؤ�G[W{�=&U����ҥ�~�c���[�*���l���"���u�P��>Z&�����Ǻ���97�M�4�������!�b���D���A��yKH{� ]1�N�5b^�����w��א�#@�j���u'gF�q���"]���<Z� ����o���3x��!p碤����-肹Z
��<[�n����f�i� d1�<�?-��>�1����EE�}�A׹O���+@F-=Y�Ǉ��c�(��gQ\D�~<��E����j�H�)��(Kh��'}�-��N��;�e��TG�i���Be\��qi�2�"��A�<���WXOQ4[�a���q�����D�K����+E�_4D(�1n�V�og���̛�����ٿ��3�ݕ��n�*ӊ��]���Pg|���ǃl^kW��U������<�7Yn��D�+%���i� �8�*&n�$Ψ4�m����Of`��VM<���J_���e���+�`����~�;��I�|��M��t�5�V�\W��+W."qt�0Kf�e��4ӸrMx���m�/�+o�碸���H�	���0�F%��c�H��%�����:,Q)R�Tsq���W<�G��l�Ğ^5f^t;D�L*�Q'����i#�R�A�yk�3���Anqk�I:>� ���,�^&��V��������4�?��O�R$�V�w?t$E�;�Q.����]X_������"hץS�`__�:`�j��?a�����s��s}��>��''�W�4OĆ�x��ozj���-��H)�!\z9"��̌I���O��� _��HW���ʸշ�(-�e�؉:���g/�����ϹV��K`�ڨ�~jZʁ;�������=�J_g�G��Ǽ�HRy�l)�^�b%Z��u���^��3��ޙ��F9���_&���<��JF)�H���6o�1�����F��>J���\f�=:ǒ��H��5��ID6��@XY��,*;�����"��6.h���>K��p�T<���h*��M<��h��)��PK   �<�XF��-$  ($  /   images/d88a5b0e-66b3-4edb-b452-47f46dd40326.png($�ۉPNG

   IHDR   d   o   %e�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  #�IDATx��}y���/+�ξ�o��[-��I�,�as�k�k{b����Ĭ���X�ځ=�����zc<�'^cds�!�!	��VK�-�}TwuY���<��ZjI�T���̪���z�|��}��p�����>on���,?�aW���Gy瓜{��گg��ש}�w����7@�tvT��2 ]��|j룰dO�f�>�}[)uP)�{���B����ත����0ۂ���G"�[�UEoUѡ
:#N���@l��Ӵ?�(��d6��F"t�"W�� ��b�rR���.(@޼~��`BS��i��b-'N�$�^G���L�&�m#���X�%O;��e��"�>��$<��v']g��/9��ou���	S��;/��!~ d*0I42q�C1q�b)��Jb�:%&�2�J�#=�N )q�Ɖ���]H��U�Oeo}s�����؂�8�ca$2!�>tp� ��.6l�`d��i�,��b��L���dSv%���ޭ�<�[�ʲ��߲JBj
A����c���cy��<����f\C�`MC$&�SI�B�{M�W����}�o*�Q;�й\������u.\�3��f΀V�1?����rȆM>������� �K"��f�⿧8t�R�<[:��ZjtN�H�'�P�N�0�C(�A/��M�6u`�z<'��.jF��R�4R{��8"P���F*�h��R��w�]\G7AO+���rC$�r��;�)��� �q����wl 9���iʠ����0��ފޗ�";���N߃��/C��Q�(�-y/�N=��ڊ��6$��3�f�C_K5�,E��-��Ș�5I���������9C�5���
����)ddK��@(.0����bٗ��Cli=�<�i�������М�pB�B0��;g,��`dd���+uZE��Ɇ���/�=�܃E�!�a6��+���v�F�2�B� #�����l{�3�$�1嘪�H�QT��	WR�@���b��4h�-�|~�, c�0ad0��1Z�@J�Ĥ���0���*!�?���� d�-alղfԮhE�D���C�X\�ٜ0J*���͛��s�!�N��c�Nk�o��F|�K_B�|yfh>��v���}��R�����8Z?N�������]�1����%Ʒ�ёhFk��^W�� �B��r���e�H��5h�$���z�C����L��.�1��O����l`X���9��Ha�PV�ԡ"������J�q�X�|9�|�I������S�r�J|�+_��^t,
A�4y
���0=��a�X��oB*�'a3�t��4P�����XVَ%��D�S#"):�`��I��҇�e� ���J�W��0�8�@�����V"g�W�ƞ�c�=މ��0g���
��3����2X�]�yÕ����y���_��9o�<|�k_�O<����3$�s��8�&����Aqm��݋��QX��.���o܌�<�l���0�e��Oh�ê�K�&�X$��ּ���3�"1�\��LW����A	a�z�P���0�H(���z,�h�����L���Ǯ�Q��aE�*���8�2LDt���>�0�g����P�!444�z���6�7�,,��ߎ_��gȲe����^tQ����_��ub��M�/@�|Ri����`�s-@�D�$���~	��,����#U�0\�pU�H@��[]�� ��baK����*��h�8�f,�h�p�������J��a��}}"�?84g#������O�{<����a�?~����k��/��&&&�Fz�t�k��@����������x�w;j��9�(dl��>�6 �>3����+��v�HG��E_~��H! F�Ĝ�J��n$�¶> aEP�!��v2�`��h�J���wJ�(dD�B����1�t���+�������7����G��v�څC����ڵk=PX}%�I�T���wf�TWW�pVSo�����"��/~��5�nˡm�'ȵ-@0L�=u�`&�^]��hX�d�R~(��,�s���$!�խ�
�3�S���H�-3�� j �WJ@��Q�φ�*�(�l�W%����-�:v@���p
�<��	��_�Ǟ��z6��<ۍ�����7�)��}�Y���<�0����3�<#^ß|�OP���I^��y@��yCGC��5]������dq��h��9�
ny� ���X.(��*O	=�+�5�A0lU�����4r���*ɵ�Ӷ۰���3�o���s�{̠u�i*.{�������-ro�\��c����sp�+=#@�����Ν;1<<�U�yU��8�0����v�G�0�"0\�}y�"|�i�0�??�4��'0E�x�Q��#n�0��3�;��WB�I�FĴ��[1$O[�uqUǥU�yh���%6�>�cAàW��Gn�B�����<����cŊ�<�3d*�7Ŵ���6��a�Z�9W2�@ gmf��WaUr!�I=�D:X%�De�gC�*��|=9�E฀ؒ� ��{�dDD:t�W�ለ-㇤R��+m�`���7���d�\P�.���M0���w�?�B̆f�A_444$�s�Z�䟮��gUe���w����-ע�\���� �f0� J^�q���\Ȏl�-g�*͕���+�tn1+,@��QS}o����VH���/�'Ɵ�.�.����$��,N<�'N�Άf�}2��5���[��E� �i8@����^ppw��� �m�8��D�i�t��������F��)��OM��CgUE@��߆�ߪ�[9�������v���� ��:���C"�\N���Ff0=cw�T� ����~)���<
8�������L��x����'s��dLP�5A�-�XE��.�(�NݿxyF��P�,4�j2\��u܃�s��<9]�iX�������N���K���+�_���Ӌ��-ۀ��z�=�Z�[�RHQ�́���
�D̆l`���U%�����T�׫�*��w�GǞ�Q a���M�����~ؐ��贀�t��u�U��� ��au�6���;Z�̏a���ƀ0X��'q�3���4ޚ�tx�n����I�λOvn�	�
v	GZ�wL�汫uk����销0��k���4J�e�)�Nus
��s���'?}D���p��B#H,%�az�S���T�P��fP�w;���g�!L��`wJ:=�Ćͣh�cA:y��90�+f��k��3�@�QW+�pK�:D԰dL���'Ĉ�b&b5�^�Lh����)��H���[D}��80epD�jߠ��1�p�)�dF@�wmO���Y���p�aUuC�*��jě�S!@X�ݛ�(��խ�S9=KL�p�3��������o@���$}?�OG�5��{gd 1���r����{���K��I:a�����^�ǍX-�������I$;`��Oԯ�k��A��÷'�%>ܘ�Puι��thF@N�PPE���
V[qԺ�~�H����Xe��hy���d����M�s�-7�s�O�@q���5~�B�����`*	H�MKP������n�*k]�R�J�s����V�E93G2ܤ�jؠ4�kpϜk��]/�t��K��J���������= <�u�c���~�?�����X��K4an�A\���<P@�}/��ڙeڎ)i�o=�]�������t,z�l:h6r)V�3� p_B�ĕ߹��]GQ���~�ignY,W&/!�v��k�/&b���?���%CR���Y��tv5_��n��X��n�Q0P�����w]G ��M�������"Z�/Y2���p�y��%��jQ�����XSx���%C2ʦ�Q�TQ{������N�Ԑ��آ��!����}������0^��om@b2'�bZt-��b��C�6N�Z1�c�Q�3>�Ĥk34�����t~�q箆����>v@��cM��n%0���v#��
 �R�Ib��@y�1�:=���(fR"��E���g���n�F�{fM�Z��^��Fv�"E��
���3z�=�u�[yK6K�G�!���n����l�l&7%��b�%6��k��*��"NcЮ�[�w��;���'%��|F	)���S���]˲�.��M��ڽ�q�'P'��K��dGܱer(�0=bp���awK�"%<�rab.���U�SAi�<}|#�V�`�4���>k���=��rs�n�U�t2%ŒG֑[]�wh�îH.�މ�"%��(,WF,|����y/��������@Ϙ�{�"��0��e0J���H_2���&/�l�A�,1�'tM�3q�PH�"��5>@�b�iY�f0g���$t��q
r���w��/[�Շ��(ъm�q�C߸{jk]�M�y*��52u[�t�2�����!�2�̲%$�-6˫:	׽�Y�U��v��r�<��k]C�\pF��1�h�S�H�3����Ɇ���<�I���$�rVY��V$	����<n0�#Gx��L�,�i�`9�@�}�}VcI�!ܑՕ���&��d����I�%D�i��n�9E�R�fG���c; ܑ���T}{���>?��H��w	���"�0P߰��rg��ivda���-�sj�v����r6���i�Aol��Z���*�8�a��r@��G>6E������9R��&@��A�p�?��0E�e<Ό$��p��w�Wk2 �՚�a10�`��,!��l'���g��9sr�(8�܉G,5q5"�VV�;\l�ن4��9,φDH]��P�� �R��?-ϝa̳ȸ�����V��k���~�7�D��}�Ό��?�����߸�IX���VY	ob��gze��Rr`D�NC�����͏4�Z<�> �g�%Xe���`f���#�ʈ�)�c���&��ޔ�}Γ�z�j9�3-��pY4΍�y�E��ס�t��^RgVh�Q/G��F. ţ��Y똚��"����v��t��	.j�,.��%`)���p�p���ʲ�u�dyF�'[Q�}'J�ޥ�5!j\Qrc�K��v�����	�REj���i��H����G�eX΍���݁�3�/�T�:�r~�,�7��R���e��ȭ0��B7W���ኢx.o �n�^V���� ��<��Xٖ��p�p�$��e,�]^#�l�k���P ��UR�I�����(ә�W�v���6�$#���Cp�� QvS3	1A�/�
�rtfs9X?�+��Eq���rE��l���ha5|���6]�Nˎ�,����%C^�M���#;�E_uҫ�ڋ�}���[�~�>$�x�'�dGr���e��®�ŵU҅�r#8J��S;01��ծ��?1��!��PQ':���Dٰ�!KѺ���ftge^M�)�f���ߒ�'�*��{m
��o��Z���a�T5�L�'~��^9(��#Wx8ȳ��!��P[���C~5F1�E�h�6BRR[T팣��Q�
����Rrz�G��%�bi�x���t����i}�`���:5���w����q3�x{h
 r}G2)4U֗��,���I)Zg&5��؝�׮��%t�6����4�;Z��V�g#2u 'R�H�NO�ީ��H��N��WYv@�lH
�������>�p�ŨI�~q$H ;�&IIDbe)9�x�@QMaµ�Lt�e�=�p�@�^�h9sF��^�n��_p`���!Q�rL�|>XA�O*t�����q��R	�D"�T����w��JB�K��PW/����q��W|Ǟ��y���:����p��rQ�1�p�X/:�sexPYJJ�7������T�{o젷�� �����d�a@X�"Z�,��_���5��`N�OG*���;����RR����#'#΅xI��1���C��r8�2�@�� ��+�����<��U=���2���$E�EA	}���	�V7�#�Ĭb0�f�+.�̩�wG�I<�����pq�PH�A׀u��ֈ�*zy?�>����u㪦U�6����waE�b��#�DX��I���g���!��x�����*�����o{���-w���������Mc�
�߆�T`�<Vt��R�ވ�D�<2�!�H��C�V)9+��&	���j*:����ޑ'���Tr���P{C�CRk1Hُ}Gpe�j�{���$.l78���{^���HGXCj_/�~��?>�'w: t
/9�xo�m���(��06����X�Dn�E��g��@$��iU�:�]�~�(��I�izz��>ˊr����[lRާ��D鷺ؖ�ƫ�\U/�.FbV�7�s>�f����,cׅW<��`��ƹc�QpP.0ˊrL8�5���G0n��LYg�.�;(E*"�Ҟp?׹�V���l��m5.�9@H9������kv�W�������*���V�u)6ѳ�qr�h[	�'�_d�0מ���u�*Ĕ^�}GJ��v��Kwb���Zԥ��\r�urn7dcgE7v*��O�/������|��|��o��~��je��<����c�
�R�X�W#|j�������&����G1l�c�r�dO�RإjXټ�c
�6� 6�l3X:~?��&�K��E�ƌbݱᥥ� L<�Ū��7T���<�X��Y(=�'�˚�89��!; �PK`4Fj�-C{�s����;��dQ��s�I�\�]1���-�Z����~� phxpW�,aSB�9!y.���2?F��/ḋ�Ԝh��<��%c���T�Y�ʗ���F������bs
�>1�b��4�]x�C�R�R	���J$	����:V�,�������"��z	7�>�O�ْ��J�!���?oA�Ϸc�ųV��E�[����0�a�����;];��@���H!��*�.,�
���%sۻ�[��]�+��D'���xE�Q������f�^�~�֭�?����f��t.�-];��qړ-�~�T��6���;5��FI #䃡:j�������~~�yw���4s`� g}/��rlܸQL�U�n�m�oh.
ݠa�����\a`8���H������7v%Li3���������U����;gޝ�`A��͙37�|3��y�MN:��> C_t[W�,<r��o�#�,j�@[��p�Զ���x}��F��ؖ�'�llOJ���z`�:
��������/��b�1�k���^:(%�(�wމcǎ�Z�B��?:�Ј����)�l����C�rb��硱�N~��d���Y*x���C�0�O���P����@�v�0lKˑ����E���$�g�%�E�g�9p�@��Č*����C�g?�6o����G��fa�	̸b/�7�i͌a[�.�'j�����I�E6�5�d��uHx=�#c=΍�=ˊ����+q��a�������w��W��_����UW��===3��Lx5�Ç˪�.�|a։_��W�~�zlڴ	������o��1�@��+p<:�ɰ��-����C�aj#Hƫі����zĴ�S�����Z���¸>)����,�7��W��oƉ��,�}�7�ݐ����ר߶m��I���O?��~�e׶�Y��W��������b�вQ�=�W��1I?N�����p��ch��Ese�T%*��.�� r���J�\��A��g�>3��efs��UG�**$�E*�=jq+����3`��I�G^��W���{�`����jۧ�S��,!?��Op���˗���ª�*�	&9F�������W��^�G�i�r
`xe��ѓ�zeKN�05�*�Ǫ#�����a
�(�s�ŒM��Wd�,���[F�᪶j
M5؎�
q�c���yM=�h��g-��F�R��~YY" $}}}��������i������ǽ�ދ�˗#��ʧ^�����F������'7�t:���ڥ)�>��+@������K�;\j0A���iG� �t�	f�((�V�+8�3�lb��Z����.��9��lB@-y��h�0*��$��/��N^b���A�S�b����oK���m��fvww��'��m޼y"-�!^OZ:ɠfm7�EZ�c"=w���ʔg�����fn<����������?�U��^���x��=Ԁ+������.�6� ���=Ś��.E{����Jr�/u2�@ngE/�x���_X���[������d����3p`�l.�ܐ�@_u0�'�E�W'��5M�=��l#x���")��.Y�;{d�=b�b�0^ӂ��s��zժU��v��I�r*L���6���QV�e��Q(��7P��&_��&D9sp<�+S@��P�}E�_WeØ;��5���5X��VX�1��k�=:00�36g��=��r�#S���2z�\�qÆx���H\�zL�
GM\�A_2���8Y�FZɋ�/�2}��ſF������VU	�<$�k����?����9��ʍ���S�ܷ�����{F��݋�I��!gCw�u{�O��L���'�>�@:n�|�ʾ�n���^Gx�1կP�כb�Qϣ
�o�l0��C�dy�	�֦�h�n4�xV�������u�[R�(��y�Gp>�2b�h8]����孧���TkSs|4�ZL��% �Q[APt���=
˗�q f��	��+J'�M�mz[��V�ns���A0CF&�C$H���7� K!�k�b����O�'�qi�%dk�&����S�8 HP;�!���c�" �	�~-��Gҕ�����q��Fs�Y,p�G�&V1R�]�=|��Ge@7�☗l�D>�&�H�`�sK��� /v�W�^�0�� �}��*�q���$H/�������G� ��[w�������B����l �(�G�������&��@�b�    IEND�B`�PK   �<�X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   �<�X�J��$ ?& /   images/eea7d5df-ba1e-450a-9b5e-b26e568e86c8.png�{<��><���%��9lcKSrH�L�m�Er.EQ���m[Sȶ�Sf�4l�0�S�
#�P��0�� ��sf�O���<?���k�u���}]��z��17N�o�I�'����SB��@�����ƛ�������O� ~�p���G��3xB��߆�N����:f�e���E8�yA .�����.(�{:'p�$�_�c~;�Kn�v��P>:�r�q_YƯ;���Xߣ�1}x����^�w?��i8�T������Owl�?o}������c�ʟ<w$�˵�*Qb�6c�Zå�u�7K��g��}Ϧ�$��u)iNj�������ԯ��DDx��Lp9>   �K �{�_�Kl����ev��&�W]%���ꂗY�˿PI��L/]����Ew�Wwٿ�}ٝj��TRZ:Ƙ���m�r�g]������F�^�#��m���E�����Y̌���)�e���U�AUS�ݺV�C��� �����7w����T����0��*����"��Q`���^h���2999���%�:Pn����B��g�B����k�L���O�/��^E$"[��3b�7HG�j*�y2Шy�{��\�M�sss�����nhs��W&��Y�3�*��RϠ�7hi���yj����W�0�	`���5��U��ЍĄ�SIͲ�h�_�t�b�MmT�]�.a�ҥ���� y_�w_A�Qe�����`��C'�#����^�}ߴz���nt&+ZxCP8\�ݔ3��G,R�ݦ���,B��cm T������"�#�����M��+-m�a"��.g`hhH��1��҄1�	h�r�l�/:�{�:KĐ�:F��c�K�>�b�.�v�(H�!qV8���тسb4>3G5I�$�y�������h0����`��&�����<�r��!5��c�z�� "���n�����x�N���\z�_v~�O��5 ����+>m�%�̋6~r�Y]G����>8< ��'7^�ތ�� jt}(,,l&66�.Z8�����KL�&�k��I��,�m�֌g<��A��P###���a�j�c�+���9��� �f-z��b�(��6S5�A�D����@S#�q0��O"�?�,dŀ���v��>d�8�����<CW��� ��X	'�����R���,W?�KN�*���\���1a߾},�0�S�@�C�FeߙQ����J`Ae��w�5t)1ׅ��$�
X�~Y�w���m'C=�T����y���׋�j4u�x�.� �$ ��қ�d�,���ݏ#�O�w�x�`�d����x5+�͓�;���J=�p��1��ݗD��P�Q	���2d� ���\pǎ#D�v�"i��!�c������lة�	
h�ӧ^�(��5J��G��đ�>Ŷm6���Cݣ�\�Q��E!�nM1fU7 ��`���*Dt��p]�a���p�	:p{ٱ�FQ�������n�����{��)C�|l�����CS~� ���	0��Jj�Bz�PB��%x��ʕ �q����谻XЖ��Ȁ|�o���7��D�y7��`C�ކT�	c�
nilll�ӧO@�����*@\(D�Te���}���C��Ew��j�vOOOw����BŰb�M;(�>�0�������{ɏ17� �:��*�� 1�i�0��J�\X� �P7�}��Y4�5�8���P�,)�)�P�M
����peÕ��v���f��k� Gd����@����Q]��0j�@4>�-��Õ���3�n�L�"D�!1#�����Q8�<b�Aɍ��$N��r\Q�;�\��}5�Ѿkii:{�6��!_t����0a��t�,-mp O�E.��<��ɥ=�����;*q6�s��R�{���)��nE�����c����G���@v��Ge�ǭ-0nQf�.8:&K!gP=���:�x��M���	4M������H�°�rb�fƫK�u�>tb1����kVH.��Z�evF���ϭY��� �Gw�ե��;ׄZm���{��OZ��̤+yV嘊s0 ��\�Y� e"#��zI?����<+����L �`G�G���G|�UP�pΈëy7���n�:b���UR^R �B��;t/��@À��
��Pͱ�u�5��j-�A
'�Pn�2ɂY D��/~� i8XIj����6���I��1���_��V���h?#�~���c,V�~l@��9;�z����1Zfk%�{��V��ԯխ���%�_�_�����k��Q�]�v��%%����0 ���v	��}���{2ܽ4(�Rc�
1����#�8�mҧ�vy��^DH����,��R[���B5k��d�d'���@�����p>(q�XE#��!f�k�|v$Gz�2c�+�S�Y�v�� � �����PD�큯��62]���0��p��%����ry��8��6�AXeZ��ݔ95��YX��hP� 
Qb����y��`���iLK����T����\�ka�m���-�j|U���Ѻ�r����`Ư���a�5��O�����mim]l���rL��Q<0g�}�Kő-��頯*�++[>��<k�t̓�~~]�9n
_x�F�E{h�ݔBQ�(�:#ve�E_�~}�����:����WٵD��~�P�a���K�ӥv��Z-���
q�h�R�JS�Κ�|�8�9&ň����gc��q�q�w����b#	Lҵgt��(���P�UU�9�Q۹�&�)�YNQ`�82�&1Sbߙ�� �U>�S�����pvzfF7�8c ӏ��_<��ʸ�M[�F��a�?�+}��@���Z-����x���ú��"w�B�
�3#]>��:p�}�Dj_'O��qV��)	��9)��Yg4_#Ҭ�ǻ�ɰ�1+�4�Qdd��N�_t1��S���b�A�ARbbb8z���F�TPe#>����j"[#��	�%Ml�2y�g� N�@��|�]f�i����@�"��^��:�D�v,��p9���?�[�"|����gt�J����.+\g?�ӎ�]�n!|�(���SSS�aJ���E���V��Ӱpv�g֝j��O.w�1%p�����l��ҲN=�a���{λ��.��`�A��z�;��D�S䉖���¬8-~�����"�VJ����l��Ɵ���r���="��k��A��������]�PM"2��Z�ү"/��#�'�x�.�O��k��]d�]�]��J��_�
S�O�k��s_��f���\ŔX��u�!yb�ؙ�%�[K�2>e�R .Ub�2��S��?T�����z\�F�5/D��u��������%��_�U�w��+B���vv}r)��5\b� ��M9!	���՚4��ihJ! �������+J����!����+�sP_���eK�wO��lO�[�k[8��r���<n�v��3��7�"�d���-��%l�����pm�\7gpp0�Ir$	F=�r���̱�A��`�j���G�%fL�-D�|��|�WWWЌঅ���u/2�|޷��
�[Z��J=����x��
6���X��n2��A8e/~�-�mpn�7�|�������t��Q�ГQ p�3USm��oo2Bΐ�s�[�8)Ts14��C�aԹLx�"�\et{\����]�ò=p��&�=�Ĵ,4�lt�.w\������
d�@(:߮�����cWwX���:�=+]jg�1U�)]c���,�G���:#$��vu�����W����'T��lF.,,� �,��e>D�TOBP��9��Dr��������o\!�W^P��4���װSK�� �φ���f?��t�B�cp�/�0llV�f�DF>�m$)=�J^�y�2��i����Dk��������=ˋN<�|���17Om�{��}�N���x!R!_H�:6��1Gj t�_��s����;���E!BMt�x�T��������IW�\�����%NS��/(��ad�	c��G���5lZ�"n���_�:tAkz]M�1��7���O�����T��+������3�$��8���E����;�x�o���r_��Em>B��z�0$��:�vt�~��s{�s�����b-Q���Q���RG�<���ŏ�	73�~-��p�{�:����LO����������"~e��n����w���F���ݱ���B�����ۂ1i��kZ��_?XTF�/?�����w��\�d��u�(2+-ͯث���3jdt��=�jF������Dw�`Ѡ�YQ���g�ƭ�J:��u�;��_]h ����@����
0,g�Kx��s������аo�
> z�n-��B���8�@�/gã���0N���&�q�b�~�q��O_�bWL5�} ql��E��:�<���G�����{UT�p���t9�i~j�XG0kի����t]n!�Ϯ�\�%��>�sQ~�����c��z��v���*�a����K���K�T/��qX�u`�S|�:�!���E���Me۷��{Z��Ŏ�p���9[Zֻ����������u����kF�7߿_����t+�.�!�8 �M�|�U绌�'k�jk�6#�����Df�^rmtt���n�Sg�@�����p�AA�n���h��uJ��k��z����H���8��3Q㕮�_�9����!BM����a?�ň�?8C�_���F+y�?
1ս�w����}�������M>�1v�ʅ�h�F�}ʯ��z�2>T3�i��B�̇/�� w�Tj1�#Μ����~ݟR\��g���à<ɫ\jp�
�'�+H9�ʵL���)�X�M��.�5��������]��W���@��#�VW���ms��A|���7|@S�Ao������Fk{{)�t�J�Շ����%O�qF�-���������߭����Ѻ�n���:��ŋ���j Y��.��:T�m����Pͨ+�4aV�u�8����&��C����E����ϬW�)'���:��c�^��!RZW/8���>�����g�]�?*A�8y7%>)!aa'�i�{؛[|.�a����<�	1玪�� ����<5�vLLLt��LsvΜ(��vz�Q~����?����P��^�:��3�${�'%�����-���F2�\y{B���S��¿�!�}���{M�qg�86w;��0���r���lǸ��#��נz���v:I������k�Ijx]T �r�	ܯ���*�]˗րm( ,�{�P�&.�ur{!,!��Ξ�6��]uGSOOkGde#���|L����|�~B�@�XN����`I�L|\	�&����Y+�dߦ��p����9�l�t�{k��|���� �1؝ht����"�-90������oy��EԀ����9%��9���ލ�I(�A��^ �g�m۶I��zbXQ��@�Ҟ�-�BjpF���Hi��6�h�p�H�Ԡ��q��Z�.������9���B�0�,((��I��v �����vPbes��e4¡a�V$x��"��f�Z�ˠQ�u�����U@�\ID:��,�3w�T��Jg{£JD&�U$�
c������ӏR��	���pI�UE�t���%�M�`�G�0C����٩��h�ى���H��+�K&�*X��2�(Z�+��% S#�(�t6F��M�igv��Ay�{gY��A$s?l�������%����׺M͒��������fāљ|Ij���,b�܀�����2��+U��_�'~�DWLE=���o��g�t������U���88\~I ��X�N�ю�Ѕ-��׷�hID&FA�a`=?�]����7������z��=҄S��)�m��-m[�������s��P������_�u���⢮��Y*���E�$����\i��Kh�CCC��c�q�����+��`�o�+(��_ԒBF~�$fv(rV�-�;�$K;�������P:qpjĉEg���q���o�Q6�6[B�#r �����J�3L�fB�)^��v%]�ո���u2:��d$?Gtx}J���Qr�C��3ai��%��W'�xH�E|{_��7�c�[A��y��F.v��	,��A3��z�b��mfCu`����C�<cc��\?6���pf�\7�ci�o��� H�;��e!�O�Q�0�'Y�&"�\cWzL�;�r�̥���D}<�7*����f&�S�v%q�߫-Ζ��O�`�����^�4vj��Dw�v{�N��XS����G�Y��Vw�֑ Q�E�<�g���H>�4Z��$�$Q<%��q����;�C72a�̈�ɼd���97[&=�������!:�^A!���� &�w}"�S�H�(I�O��g�&>U+ˣ��}���Uj^=~z.��{PB[YN�C�+0��9Ċ��.r\p#��
X�'�[��~09�+��p�����#�T� \���k����Q���쒒�v�<x!�M� ���ќ��H�_���������k6t�v�˗/�T%"Se܆�A`q
�Wg��_M��0ڵL�Dr�uY3p~�J�u�Ś�Z�K�����vTw�Bte�.�bW�3P��j�UС���|�%x�"m�C��k!?N�	�300�� ظ�(_�5!��"��Ehv+�q9�P���fD���F������,bP60Ǐ��^����)��u��%�z�B9�����ߍ۷o����g����B�JokF�^]?��Q!��۵J{9}H���"�e��x�Z���y�.4���م�a��M>���(P�G��(�|4��@�ê�x��%�����9[]|�����hie5o ���;�!"����.;��<���c����͵��s��,�;��N!�fl���e�QP��oW������>��^@w��,]@�oM>Z�z�z�2��.݅�}�E4�2�{秆<�=�/T.�\�����O����+i�b^�+�����Ѻ[���gazDͣ�r���J�ğV��0e�-=p��nP�}z��J@��yt������O:�<��T�78�->,V{e��$��e�N��$fF���tb���X�����B���ï�3@�]W��V�
�a��V~����G��*����~�)�j�`�W�<O2��`��;P���nZS���<sƽK���*��\�M��!�꣎�P�`�/8[�n�䔔ج��������w�s!Ϡ�<��T��==��U��UvWsUB�Utue@��o�z��@��f�޺�nE��#EXn�m�ԍ�j��O�w����?,�(Nӽk4�\��:qv�Fmm��37�2�k�Q���{�d�@q�5����4�nj�emT�A0;�e��7��њk�*[`�O�2.N(4��P�c�l�o O]Q� O	�����(�d���ۖ�󚾤�$���U�7��o���=�kw:�}���A��ϙ�p��\1r<�)E��3&U;|ea��7s�㔟G�ߪ�ow-�qe{���r[k+�0V���:��*�A�P\RR�;�Z��4ו ��5 �dDA5���0*��mA"�U���T(F����W��t�z����Ȭxd���v�cii7�r�3b���uQ۷m߮+�� r��ں~ħ��zM�}�\<x�<}k��
��Ѣ����W�=s�^j㍴4Ô�o�x���Cײ�-)��D��B�_t+����S냉�Mp�!���*�`�� L�:A ;�ϧ�~h
>7����-� F�k�p��G|4�Tw�����JPu����w�W������t��*3���<#�02�n��~~�,5�H�I���?i����~�2`5~�y~]�c~�$�(S�<+N+�2\�K0�BJX�}����k����_���G��'N��xO��N�ŃAȨ@�+W��t�J��`0��\�3F�������/h��*��=7��m�y]#������j����jP�'�`,�u��Й�.~.��-��O�����^c�k�~󤆲�,5Z��X;?vr���fsKK�`S:��]� �ii<P�9:	p 7AJm}��;�dѻ87 �JB���4
�������֍%{����ձ���p�1s���_Ĥ��h�zJ��7W�X��C�U@I���r��	'����g
@`-�/:�w}��,��Y4�i+ ҿ+-�e͕�<LK��gU�����4�޸ꥒ@�~y�=ۋ�����q�1^��g���3AB���Җ��}*�g����@���n��uE/����7Kk���̰�,����P|�����kċ}�._����xO��}̶EYW7Is��7�E���;/ނ�C�d1(�x&G!�-�LMm����w?�.|���9��mڢ�Y��:��_�k�z�l��.b$��_�}��-p����#q[��c�M��+;ޕ�Rx���P��?zi��ba1z�@�PS�&hv��3l��x�XͿ)������mמ���w��	t��VjNq�
�z6�_�' ��n��8v
&F!�������޽˥�����j`Pu���{���Wd@�,���H=ǝ(	(�Y%�lh����DPH�Ｅ&&&
�����అ��#PH�n爫W�j�&o�H=Y��I�o��H����a,�u�+���xͮ���9��ST$���@	��IgzkܫЅ�ު�<��Gzb)H��=����p\��KR���_������r�GT�^��N�r��m#��p�0@;S��K�9'������������4E��B-+�{w5�<�lޅ��"�k���)#�f@��� �0���9�˗/��h���Ộ��ܠ���p��Ίr��42��67���J6�tZ�޻�)�5URA��3�"�A����n�Y���hDq2�p,�P��$r�.%&0�����T���Bk��j҅x�4;���J��1Q	'�y����+Wഎ����ǩ������)���k�ι�^̠K��d�N[�,��6���[q�����}�)�t�M��Ą���10䢫�>�D-�PGo�Rֆ�QF�b,���\{"?�g N���y����=����)�}H��c1E��#Ü���!3����$0$255���
H�Q��@��3�H�����U�}CY��c&y��f�g˂14\���-\�_/�B��1�Vږi>|���E`Bqj �"t)�V�~>��ԃ���l�/\T���cc.xiH�W�E�ͤ���1Ы�`K��
�W�����;q\���\����؈�_�[��1B����U�^��譌�'P!}��+�G��}@�<�T�?K�G�A�K��
���`W"�\�X��p�p�\�3���6$$$������u�Vq�1ZM�Ja�=&���ٶ�31�9}��;��F9�6��%��U�_r!��֦�.�(-�����bqCU��o���E��u5k�S��Q����
�"ϵ�9Ǵ�4��_��9 ���`mX����x��&�iS蹋AV�[#n3� 	G�7��𪕀�_)B��|�X�P@�Mѽ���A
k�1�2���w���&	���/k��C�|~���s���c`��4���Q(�v*5t�ݧ����=��p��,y�M�x�8�InEg����O���J��K��%�ʌ$�0`'6&d�#��7�>�kK�˯/�|Q�8e������{*n���&D �B��`#��i8* h�i�U����b����@8�A!"�r�8��jF�LAwG\��A�A�R��W[=G�:ĈHҸ���	�S�g�&���6��(�H��'�϶@C���Q�D�X\�,@*&�N�A��aU��w��`�Ft�*�HҼ�>���2�S�W�2�$��|2#q>��,(Ԡ�b��: ��K����4F�����5�!8odg����	��ˣy����o��4G��������M��G,�P%�����h��^��E!r��ı��:ʳ?AL"��$���DJYL���q���@/<>����i�jUg�2h78���[�A���b |l��@�Qh7�W�(�U���2xz����Gh=�m�NvY��*�`A�r�v�1����/M�%WU`:MO��3�Wƅi{�H��7��H����I��KM�_�o��k���)��/AkT��y�G���y�9ee�0����ۦ8�b�S�H��tK�J�
UƁ���D���E�0�(�SJ4��$AG�Ɩ��óB�h�	e�j�l�6����,6������8f+�l[@1�ev���3�?}����U4	¿�|��b���\�$����"�aQ>�%��ǫS4�Z���b|������@�җw �!-��bpfAY"�����PM����.��[T����4uOu��* �3��<�e���rejPh�
ToN#��"�}�l�~��B�\�n�ݣ�R����TbvKCTQ���?\�w������@Tqf�_À�$��7!�kL��|��g����B�\[�It�K'��D�zXŻ��,�����=?�m�C�|ExDy���5O��gP]F�A��T�K��``q�%_DQ*�ů�R/�e��l�i?�`���x5B_�
 |�Q���P�ŻP!��j1&E%��
(X�	��/,�����pq�}D?�"::�5+��.ԡ�u	#�P`%^V�^�W�8�)p��#��8�ٶ@�T��"|����o���tJ|AY������|\�P�L��sj��C�l>P[�,p�b����#����м�&Y	y�g�pλ!����ؾ�qT�`t��T�n�e܋JH�����T�q⢠�DyU��A	��:l�j"�W3СN�sōh�s�:�B3�!8֟$S ��4x��0�v�e9������c�����j����)RN�N����O'� �SVv�&�4Ա�u5�����%0�J8g�AbkrJz K\OQ"�GH1�j	w+���^;r�6�����UqB��$c�7��>��ু.�R����3���ۜ�m`�C�9����K�����}�&d�;*�G�o�eUDﳀcA�7��۷Ĕq�{���?&+�ǃ� �d1~��%�6<ie��O�p����x�.��Ç��rư6���\��\�h�|5t3���R���I�+:��A.5vA�v����� TkRk~�#�6^�f�f}R�[�{����nL�5A;�%���ni��=5!��@Ǎ��Q�S!��U����qR��, L�{�4\
�N�w��4w��L����<��x�f94� ��P�
;�J&���UpΗ�ح �P���N��B�5ފ�A]�tkn{{A�YjA��Z��������BLqM�nE
nW��0�pH"2�I 
�������Sx��ʾ���%���SX(.g�X�%!ԍ��P��EA��۳�18�!�0��Gx�C82�@d�p�k%�0z�3�@a��eY��]�ع���w�~&����Q��Ra��q;��O9{B2=��C~��!7Rm��P���\O��]�ba�(�n~�Rp�u�왘�O.���T��-���}O�CNPZ�}~�+��Pڿb���+m�������������C�S>t��pY�������b�h\8��K�#�%5��$|z� ?�kʭ������*؍�����q��MYE�L��=B����WC@�V�,?�ϑ/lL5��-_�o��&�������O�W��.�?;v����g��������U%t�15��^�n��+�Dax��OC�b̎� ��KYWW&99YYU�~�#��n9�Hf�a�-h��	�T���g�pk�Ί�{�&�&e<Xh�-�����@egX��cޓ�!��aDۓ��VUScĎ�tS�_�t^R7����^����q�~J}���`wn���|5����H��?������+�X�d�d<th�O��^`�o�55?�kA�eG&G��i$�O�����Q���q��h^�Mk�**沪d�qĥce{�Ul���o����V/)�?��$˱J�e�XYܸ�w�繶�<�2� ��>r/�x�֍7XAJ�1�M�j�n�ݎ���b���"�l_��:[�f�\�2`��F"o�u�4�=n���/(Pe�����vˢ��<����N��O> ����nA�E�Yb��^Kh�c������A�1
uQ�)$���G��������:{��Vzy�8�����6�h��^�Б�_�d'�ǖMR�@�x�qV�1������X1W�g8��i���X�T�h?��G�������F�y�:7Ԝ1${.0���,�r��q��sR� ��8�f�s��[���;d?��}��WA[[�T�n[.S��c�D@��N��2�6����FuVX8py�ʓu����f�J2֯`��^�%�>x��k��b�ѥs�{vY�j��H��?I����M����3�����|Ô�,���g <��^��3���ʭ�!����������R��d����#�L����앙��x�[�_Op+b���Ug�b*
���V�&�G�:�i�K���*�' GF�SN��i�h��54$(Ʃ^�B�}��$s�h���"�/b�ޱ��)+˲w�܉ʷ�o����β�]��^�)Fc�*�M����Qv>��Y !��x2�%9�ٻ��C��O�ӣ�2x<���q!���ƶ�j�[�(s���F���?ٯ<Ƿ��������h<�Zz�������"��cκ�rq+r<yj����|$��M�R���io��Ú�;^�x���m˓#� <�CuK���ڋ?�ڨ�4��]�{M.W�l�v2�iк�g��� +��~m���}"5��F�9)��\�25PVR��n�3� 2����ʎ��1���6�Y7pi��>y��K���I(ir����[�᦬����!)��d�����6G�Ea�;̾nX�K:��ç~�������}���,�i�y��E��E,�~.�<7f�>���'+sFU[{I�^3�N����r�
��,3�0ms������4�B�Ry�ԟI�{T$�W�a$o���o��e���f�{�FM&�4d����Q�ɻDځ�徙}o���{��*78�ǎ�u��1��H�mY��5�D]IЯ���b�U�<� \<nG�Q�W�	����R(���WO��i`�A���7�#���� �*�(��ulȲʹ�A�ܠ^�A��#���8�h)#��ߧ�r��yV��ސ&�ю�<Ǫ[��@N@K`�Y����Ȭ[��6QKKK�mm����i�+++ϝ?��^��|m�Wю�Ug������ť7ݕ��3��0������bً"-RHv�w�
�cܗ���(��JLLl��* @W���;h*Ř��Xd�wCS/Z��G|�J!�\�曳�W@4��Ԗc��,��V*������>WNc�`�b����V�����!{�	?.'{Ξq�3<�f��H8L���x�M���B���:>�Zj�/ۋ�L�Ir��fhh�VuOUk�`����f�g�:�ǅP�:-t ��f�7$Z�?�.Z|��<��ُ�t�o8V>>�ۦ-&�����
1c���2:�Q:�y���gRi&;�Mj8��(GK�8#�g��d\Z��8���$O�@�D����*
��)`��7�J�4�"	�+f�,U�@S��������9@Oi�<+�s[�>+�~��	���73n����XۭH*)�&�@�"��4$�GP�sU�<q w1,(ZW����J����T_��2E�tdTԊ-��B�Fz��R���Y�D�^T��`����4衮�����6����9LE��3�o�?[,�nK��	L�2��2�%,�t�����6i��M`�E-�	��M�S[7A�L�.�ܦ�zU�R��}[�	����Al��6�T�|�z�E��ʥkއ!<��m+�t'n��@[y��������JHD�k�x��a�z��Y��=�yV#�gϞ=j8��
n6&����'�ꬂcMH�l�3�-��iVe�.��n浍��GD��.p-A^2��p?-M��*�PCv���*H�v*�H�``1���텃~	P�&��=Փ2�qo���x��K�l & ((h9˝���z��,��J��P��ϟ17�o&ZZq_�M̲��6�m:8_8�?�7�ңN{�B6J�T��4&V`�ѦEɍl�{�]���tӶb����x�;��.�s�qS����x�b0%�=UE!.ta��pk��ϰ%���j���~Ao��3̋�8.�k" c5���D�,�0���˅�����^pp0;B�\W����^���P(�`<~y���j�f�/,�Le&��7"�?hr��d2�d{P=��o̹T7>D8�J�*���ܣŖ d��T�M�����ou��ǯ�����	��4�)�9�z���
�>H���:͘�`rfF��ݝ�zI����#޾};.!a��	�Q���vP�j����~Cd�|F>`GA5�'w��-�z��%�+uH�K���:�U�S�Q96�32���;�e,>H�:YH�%��/���H�������'�C�SXl�	��GκAL7P����t��ᗴ���O���4�b)P��6�qH�+�%/��z��$�3'pa�=���H��,�p?C���2h�ш�j�
�����th�x��C�����:�2�U�S�����t+@�xF6y���8�#�3������M|3�<ϼ<*�}��������e��I�����R�!��8V���:n��v�:D���ۡ�g�ZE��J�*���ߒѕ֏��uV�O�Mf@�Z9W�ߑ;�*�qEܗ��q��Cb��#Q�ӖP����UK��]yE���JPu/�G�q+�qOLJZ�O��&�>#��������/&t\̧���|���P3�5��/�;�@S����W�@���_�.Z�65}�^����A�/���]����	;"�TG__5������ UR(L���;X��3�v�'��� k1��/o)��]���NqZ�f`X���$A��;�G
�5	_��} Y5�
w#��qƜ-r�2'Ӌ��-��HB��y��S��A�����Vd��I�K��������_�Jl�}� u�����99T�jwQ��~��9����~r���G�[���v�^	k�g$ݍ��5HH��R u����b�� v8�����<i�aj��M��j&pg=�d乀8�����#�'����L�`�l��yC�F|�Lt�";�EP�r����]����Ѕ�c/D�Jg:�y���b�0�����1�,4~@X�);�E܄�Z�r��.e���|�Mf=0^?`$���e[r=�N-��&<��%o��.��\�B1/DW���a<�V�7sg���߶>��k�D�_��\N��Q� }[P��P=U�=��'�BSE!�F-��c%F[9���a ��yW�� ��<8)�샸g=�Q��6�b�N.}�l�7�n�I{璷�8	Dt0�Ol)����@p�[�|��v!�vz�U7�>����@���/��� #�{ڡ�ҟ���0p�wp���b���fR�Ȏ^^}{n��#�D�,ի���U�:��U��l �t��|�fH��Qӛ\ ҳ����)d%������q���yOj��~��ge@l��(�w���	6Ĕ(����N�qYh��+1����]eB��>�4�y@�pE�}��$!)�e`��(�*c�3�{�Y[��<�������˃O�������W��x�W/N��<�ۗ)�	�2hp���}F;��.?�<j%G(����:�������S�˯4i�t��/CY�um�M��8`r�C�'-�|��Ѵ��T3��p�>���\�U��6m�R�FF�K�AAe<Ѫ�EG��cR�N�'���f>��pi/�v�$��0ѯ���tX+�d
�˿M.��#�{����y������-�5y���=F�U����(ҭK4T!�����s�23V�R�?_ʙU��Ǧm�\v@�����C_^��oQV�U��6� K ȴ4������ؙ��E#L�.j9�:o����7���z�8���ò�jy/u���ʵk�� p�'Ki��lE�K"W����1�lv�pU�3Hm��8�a�~��ZX��j`��4���������܃~31�3I! �{q�-�����}V`H�"d�o����r���PE�>+�X��p�ր�g�B��E|�ݩ���w�*�i�y�r��Ï�	crSHw�vg�� ���e�b5�!����j}(͊���C��$�a�\����oP�up��ӻŶ��e��=���!ζ�%�ۛˀ�n��:877gA����qHw1�wփ�z�G�A���e��22~�����s�m�Τ/[�Q��(Z�K:�՛�&�g������w3�h\RBBxwww�ݻ{��ϖ�B�dy2����4�{�t>A�X�P���� �����6�<��흁$��A�0%���3���:�SZB��@ǅ����' �I7���Ėh��[�NK�f;�~�{���QR'@͘���J�î�X������y��@�+�
Z1�
�c�n��C�>2O��o\�]�Yӳ��l�5ޕ����l/yB�n��Eh���+m����x4��ѝ'{�<�2T���x?��r��e70�~P��]	���Ʌ��y��@��@q֤0L�y���/��˻ �[71c_����F�7�an��ڰ�1lNX�}��2⿼Zh�#���3�2�]e��������FM�c�q�1D�Ǘ�
܃�,F��"��jC�R�@�q*�)qJ��~��i�_aa�NN)��y�`1��0���"�vʛ�M.S��˥�,=L�	L�Åm��mw��̶����i*i��u'J�[��!�ycl�#W1�[�ܷ��rI��ԩ�Q��:�o���[)j�u�[
/�W$T=�p����2������;͵���6g�.<�9]�S��F�8V��I�~�| � =uU_.6�D���o���%o̻���Wݒ
���
ҵ�+>�m*jj�)P�m"�w]������^����
����wv�����������(�")y�(b����1�4t�=�>�4T>����:^Š����wZ�\�*a$j�HNN^U�R�ؼ�~�.3��Q���P4	eʬ4j���&y��t�|3U���3�Q@[xz߾G����!հ
d�����k�qн�6hs���,wC�G�DBZ��ȃ��+N�=+�i.�yک��W�i�O4����qA���������>tR�>���?��<�͉������=@����';�[N.x���<�~�?-� �����$�J&���͑1�R���b3H������ ��@�m0�V��'\�:���+�~��`�5��(O��Y�;���M�hկ�u��;����+	�Y/��i�{�����y���|4X����>|�W>�qyg�ab�A�af�����?B���T� W���'�$��l�q�q˳���aץ<��y�+�0�m��^�w��zq���ۃF6�e{�C���ئn������.�N�3�8��f��-BLE��w���&ӆ���#�Ł�������D���]��-�2�^�z��/�Ɏb&����#c��+C�W�J\ϝ�)��h��x���1���r���AY��+�����Z.I>�����OEV���k���O�%��Qt��]�'��xs?�|E��E-�Kש�'�n������ຩ�:J��/lɴ�M�/GB�Z����%oI���j���r�`ęn�N܋M,�*Ȍ�,�]�7O�z45ԲbɘS���4$@�mn���*n+]�*�6�BDWr�����5�?��qR�~ZZ��Ɣ�m۳�\��0��
���41~N]t�\���j�?��'�*ܩ$!i�a���]]�Ҽ�+�?L�c^]����X�y����L���|���ο|�a-���Т��i�N��%Wú�p+�kmn�`�!��i�ir�E����-5�}F�<W񌹢/���0?�>yU��_roGc0lyb�ѣG�_(L����,�QD{"ъWR����z���7�-��7p�Ulf�zX"�� "�#詳�
� Ȣ��R���y-��jx�0�#kx��sq��Ԡ
�Xi돵_U�����$�T sA����i�7�؟�F�tk���¯r�{�8V�c��C6�vo�!�g�GZ�|0C��z<� ���_w�:�ڨ�L�$$��k�L5"&	�o���
MB��)y��S�_�`���\g��Ҡ0��p'��'Ξg\5�}_R����β�+��f	��9�4�zz�
oPP�}�M�/�7���:J�;��#AL����7��×!JONN��nw�Zq��yϞ=3��@K�m9�U	f�xF'��v,���������+Q E��Ø�R7z������\��o�n�Y9�"w�"�y�3mMF�kOeUO���)�Y����u�mr�+q��g��D#(�Y��C�w�qC�o@�K���n��l�:�G#�d�|w*l�����l/	���S!Y��벫AA˪���漨�1��/͎�zL�K����q��qM_���^���4u�����+�a��E��bﰷ�JTF�
T(�5��!,��g�~{����|r>�y���~�9�s.�8��A�� �]�a7x��I�Ab6>y*s�I8{�/%���T��&�����eٜk[�-(�WI�F$Wc��|��?���+L
��2P�ҖD�pspx�1H��)'(�9K'�}U)���'��K]�27Y�-�ϻ:�2vX�6�ȃr����j��-�y��ڭ�t�_/��2CK��H��gU�� �)Aˈ�4BkUTT4o��ۣ������Oϋ7|�q5(�{�u��:��٥CW�B��	����A��@�FHۼ�ւ�7�>��B	Ö
0�)l���=�5b39����;�\����� .b�����̙�Wlj�1����p����Y�-�j9S%A�UMMYy��5D��␟��S7v�� h�ʀ~��R��w�x�i�?�0���S��sIʔtb��夈?���N���^��v�Öt�/)&�DOy7�$v��h�rc���!����E1QQ����=
�Ms�1_d�ԫQ���i���ߙ�/$
F��S}$i���^����y/���9�A[�� L��������� �4�w����9G���T&$'�,�MUs�\�=���,:a��2t�g���Z��o�GuۊǤA�ލ��4����D�u��B�DĢ���@�	��`f�bb�~�Ծ�@���9V��HD���o�1�?��3�t��ه��?oU�[���??��#��:�׬o���t�/��:##o�)�y`�.w��ѵ���Ɠ�;�������"̣�-'r�Fk@�Xz���*�aP5������LC�{i.GyYx�N=n�D��Z��w����B]��J$.7�:]'�!���ܒ`�p^p	O*�I�fXp������*kȕ�{�=���!عSS�
�2����b?.��.@/n?U+/��5J� �CV��8�ފ��,�v=�P��w��LS7#}�"���=�`�U�3�3��z<ۋ@G Va���U`��WWW��ݼϭ�&l��ݻwג�ɑ�j�HkRV�ކLp��Ä�Xݔ��B�X�ih������i�%wd��z���C_u�5�s`zz:0��MԺ�Z�-L��Ƥ2U(��xfW��3�xK�g���
HQ��[9:\)9A>���3����r�U��n���;���D].1K��q&����t�'VXq�Kh	D��UġM !���1��5;�q�n�o�L����������u�
��YKk1$$�}(,��z �\��A����ީ�|���#�%�ݦ/R(e���#oXXn�dW?=�v��E�eUP�R(8i��\�e�ב;�gz�8 �"�������lA���b�Ȅ8�f�"���Pk����Z2�w3K�x3d�r�=x<���:v9�|��\��u��w�$��Kul$4�q�b�4�ho��b���{��H�5��:�;�s�}��|��k�8�7x�:�]β�rB���Euļm&���h	��a�gI���.��K?ep[#�&BT���_���05C y�u�ݭ�G��*e���"U��K�N�\�P��Ʉ3��iyt��iŗ��/ɝ��DD���~&8�W�8+��F��Uh���.��JZ���vca..������s�4!xA�O��� B%kZm(!��^�g���9�X���>��(�G�f8 ��M%�^�<_Ta�*����q@���%?�'��2G�<�QUz���؆Q�O}�}F��.�2�� �F�������to-�σv��L��C���W����T�6�ؤH�
A�Τ���,�u9��b�A��(���~�����n��	��p9ï���*`�4�rq� �fU,��V���j!?��%f� Зb����ű2^����f.: m��X�oJPh*h�V��7y����`��:�d`��w���|Ɖ�'��6��2��p0���M�	ԇlfhn��>t�+gc"�9�J���}؄����0m��QЬv k����a��è�iy���}�k�׮]���~�p�j쌴[��K�@�@f$s,���D���5}����A�yxF�iP�b�e̛F�?��	���y�d*�s1ݱV:�ʿ3�6����6CN�}1�xh:���*E�����d��1b��(��.5hǎ!`R�'�MJ�$Մ�,;�J2�BH>���mf}݁�Q��Sނ�T�; Z/��8lf4:z4��~�yPE��9�����{�ͤqJ����O��'���\�:�G��ms�+�66�|:�Z<S���e��	��&)��'���4tJ�J� N;�A��x��Н+�@�S8�9��2I��^/�i���X�E�gssӂ��o�����s����y���M�[s"��w����m���{��C��m-r�y���t��ٻ���r���X�?��Ì��~���o�<9$�|��;�Ա4�5@�Ų�֜���A7���IID�����|�0z1�'ȏ>\���_��^���ZAbo��d�οgLg��a�\T�I_LJO���U���IN�\H�-��T�V��Y�H�[���!��iw�2RQQ�����0�İ��#���X-M!()�}�T����)O����X΃�~�{�j<�0�E�Р\ϐ�)���t�b��%i��|d	�T���lfP��z�b��q�܂bd��e~�ȣ���Z>Q��s��lf�"Aw��7��t|�:o-3Yx��扠��'J0�,J<a{�C"��dl�(��b�M���EJp:~�~��INP��>{ͽ*%c`V�(��0:����1ٕ?	��x@�gd՜<�ֹ� ����3�Ld�+�8q"����TI�P9Y��õBZ�:��S�����I��M4baj�@������LS�F��S�q^��	����,�%P6�?n�H'
�3�mC�AI
|�V��[i�m��*����Cޛ��1����!�R,��MNs�v��u�DH�_Q4������G���O�x`y�e�3�):S�h�sc���+����3�: ���d��}6��,dun"�1�=�F�P�c�ߠ]����0n���@G�N��攞���Dڕ��n3Խ��,p�;�h����"��Q�;�p�a �y�`�z���L��v�j����p�������-��N��T�>��,p�E�)V�G��I
w��d�w�9�'g�AL��,7��@�BEN���	����Oi��I��+�J|�V�Bՠ�'V� 2�t�5������F�k�c���pW~�X6L�$U�h\ccc�ޟ����cI�����=`��I+�^R���	r�HJ�x%kiT�ߛ'ԗ_��<��̘�l�ơ7�Q!���s�����,�Z�A�_�����]�$�O�0333�S����l1��_�؛�}b��\�ΎP_������]�\I�$���)e��F���o$]�R(���OI8�0P�!OOO/p�_�mc�upK��z������ �e��j�p�T��=����y?0a�G�DΒ_���3��}H__�i,+{`�>3�'b+I��2\����%;��@��E�3ՕJ�H��)//�P������{Á�@�4'�\~�k��d��3���d�"��x ��%������\u��siS��������`x�G� +��ԴZ#�I�\�c��PI��ނ#���%uD�xeWK�ll�<˰N0�v<��ū;����<��Ǐ��?~<�ɘ�yNj2�s�6�a�3�^�"��,x�Vi:�1}?�	����Ԥ��F���ϟ������GUD�ޕaaҘÌ��H^��A8ɬߌB�R"������ �U"}U)M�w��'��NC3�ǵ繶��B���m���&��3�����U�ڣ�pJ�c�t��骺�tá�Vq�<�MOO�jj"�MLT)\>6�&~*x������)�\�&�#߾.���D`��s���go�����u�`�wG��'�t��(ǲ�����ì��+m�$!���/�S�6����m�+;4O�Xz g?|u�.GH.��7����>��"�]�>l�VU?=�U5�*����yb�����n=s�>`���Ns���p��}}}SEEEm3���ֳ�|�A�j�|^��<姖8lnm�h�H#�����g���:�%�����[ߐ��A���G��`�s�����:�&j�	ƣ�1����r���/i��spo`�^�:v�&w�h���M�~�4�c�O��l!'X���U��P�_}�л"ܷNM�4$�W"����y��h�����U�������V�$!5i��2<<K@b�ӳ{���k{��
c5B��K�9\N�OY��^����7��"�$�E3��q�$�c��?/��$���1�s�wq�ɟS+�un1ke��al[c�N�"��I���b����㬿#�LF
o*3�?���x+��N�/.2$QD��@.�5��sӴ��H�6	$S�L7,�?6���{ 1�:��B��Y�>�R3P�)�6��'W���i�b�d4�P��T�5H*ޏ��g@�xNbo���&>�� ^w����./L#��Ǿ�GGn& ������@��I'��G	r�ltK_$��Ŏ_Xr��#��q��ٗ�F�4�Û� ;�@�&�l��Y�O<������1���S�C��#���u�82�d�	[�1i��_�bacSI&vX �������5 �2F�
�;ǧ�4��C��T�5o�O���":ܾj���(؎�/��j���R�ޮ��>��zu�3�Q4�O
]��"����Z�ڂ=)��Z��X����s�z�0�?��������A�@6���!W���,4�!�����Sy���RȃC��v�*��6(�"��1�?@�@4_�F%-�]��[t�׸\Js�Mk(�AlB.恳�[�d!$u�����l�I�����1���ӧ>Xt����P���������0�-��5$J&�m�k�����=g`�}�E��"$�ht����i���zX!�{��ƫ�n���on8���|Y�d&�������oj�SZ�r�!|�dd��g��h%Hb������+�/Zt�lC(�JAy���%0鰼4��Kb���<e�a��`yh����kx���#$+��|<Nl;�P�����`N�2��7Xޓd�M�x�[�@�%�Pk"\�!�!���ٍĩ��?XG+)@S�Aa�jo+�qT>��������d�&r�����A���a
� ���2gn���ˏ� ��'�a�t�Pa�TV��>Ķn  
�w���lq��Z��(�F3r[�
(���SQr������A�p,��ʰ�3�����)��oԑ_�ZS��@9rb��iC���{�@
�.ĩ4�����..�da���=��hk������oa�����{��Nx F����Yl�7Ў�=,mK�[k��/��)��eX����~��tGh�6��°�ϩ\�| r	]n)ʚ���Ѩ�l�3a��٪�]u�6���ܱ�u�3�g'������F��*R��ڎ~+���Y{#!��m"?%��@����A��w<��x��9�m��
3 V��	V`���X����/���Nϖ#��zo���ѫFn ����%	ǘ:����~Kb'û������B���Ǹ���U��6�������DC����l���]��mΏ�w�l����a�<a�E��<�p�R�0_�{���\�T9���m'j�	ٞ���J�8���'['ӯ�c�F��[��b=~E�GhI�R)~	6;��6
@��|���e��a��%�1�)����jo�Z������|L�����dk�D��v=�p�q�	�Qf��*EE�1�L=b�G�P[ج��H�06Ƅ�e�&X�S���g嗧��B�t9�)�2�m8hN� D{:O�$��$*�{x����eKX�C���0]��7()�b��<|�a�P������k��\����	��JQ��/���cn��
���	�!U�;�gfަW,���'�H`*'0BNvt?r2jil�a�^��z���9*7��9�^k��m�g����a��:�n�@o�p��u���|=X�)������hGD����Y�&gW;��س���Y?���z*}Jۧnb!N�.�_e����Gz����.<�"䡋4m[���=���ɩL��|j�4/�nE�k�`%�Lm�ܴy����Q$��0����-p� Y #�^�>�
ƌ�Nw0ET��������P��B_8�9�-�ڲ|�狏���,���D���p!�"�sX�_s�!ėv�/�.�I��x������Vj��%��I�fj!���f���A�ܰ��{���!F1�6��u��iKSZ�y1��g�.����Z#�5I<�t�������A^ff��"<��Z��|J�3�u$��KK��5Rm�º�������b�R�c|چ�H�k�#�e�^֋���y!A���i�~�~�G<%7m�s�e��L?#
�D,͝i�n�a�'�����:>.�^6�P݂�Ia����G��?w�Ί�6����s��k�����N�u����KA�>]^�)M��(L��:��wtTi^��q7wmQ�^��B��c�N�y��d���j���0i��ܑ��Vl]�ax���[*p��z#�s�!礥e���H�M%ݶgq�T�_�o(Mq���!����=l�Ý��5Xx�"kt��M͕Ǧݕ�:����$�9OvH�9����1��4�����I>�x+�a�_q@�0
,�j��`�ͳ���a�6��nJ�aMO�Q`c�2 ���$�O�E.��� 
wMBj�|��/n�¸&(���꒎�*<�TxɍN�g����.[�ϯt�3\>_u�G�
/Q��Wڟ7��*U'��3c�ܻ����L�b�=�>Z�
]{	|9�˿��g�*�ܣi�$��ܰ�ﮊ��\:�s��I�LA�<���,�s?
&���T�� $���[U�&�Ni�=��Y��RǷS��'��F�_�EK��nζz����!Q��V��˕��3h�_8���N�D�QӋ��\��V��s?�W�/��܊���H�ֻ�X��'{
���DY�B��Y<nP�);)�ܮ\�-=y=����P��sq}~���҈�#�CqBzL|fr��F)�� {��YE�_��R�r��v��"w�>�	1iP��J�@�cͨ|������]e��(W2A�Z�@��h64L��2��� %3�4Z�r��Ud���T?I�_�t5�b�/��t����0=׹�X�F�H��~��(��FN�j����������,�ж�~�U�e�G��1�-K�m��R�I�������'�J�)2�����m��mDC�Ë�"��B�8s+ʃ�B�a$G3����-�d�Ũ쯷@G}w}��;6�_x6-�(HU��������OU��#x>;(�:	��:ͥ����"����[�
5��2J��(�[�w&5�m6�[�ߚa�Np���b��>hjpK�'|*v���D�4W)�U�V[(No�fu�l$#-r�-$h*z��2�h,�-4�0`���=P��w�$��TVHE�5�nOe`O"��w�ڌ�j��JD�Q��e%e3/�Ƙn��^QA�Ő��߿��'���v����<q0���ϊ@�yu	�!�CI��³J�LC�F�c~��P%�֋-����k���_�����>\���&�e>����Fu�6�X���������|_�")wGv?v�O�-�I�"Ng�w����^��'�k/^����+ ny�sB���(_�Y\ QJ6n蠨^_Q>��:b^�J�v�z��d@k�%V�P�o�[)6�ͼD���s;�J@����;8`����4�ի9��e܆�4�p'�����<��Bm����m�c�Τm�g7�h%< w!V���z �Y�c�$���
C�B������ŏ�?�NWiB�C,�����m�Lx����gS��\x�E@�Kr�`�N
w�r�<��;({�1��Ǫ�����ER����R�*�r;��j�Y���(��%�� h�p2Nw��#��{,; ~���I'J��+>]��>�����B�+����{#p)��t��M����� ��]���t�;��?\Iv���[�|�>���'��uhQw���s�\�(e%X�7�?�v�FZ8����o��~�y;T��z�69b���,ͱi���=D��k.��De�+}Lj�	��`����oo��<VC��q��_���V/t�jG ��@�o�@Sh:���bm�-�5D��|m�������U���-�Ez�?")���yVg3���?��x���Q>K���WG��9Xw*�.b<F6o/�-נ��}��^mff�~��DCN�2���_��$��,��N�:Zs�WE�wun�s�JJ��-%���*t�����Cn���wCв�Ҁ]�
�^��>���OR[l�,ߕ�mΎӣ�j�wA83��ڮ� 1W͸����?�\]�W�lX���VZp����vJ���{?c��;_���f(�w\�G �������0=����Xl���.��%m_�����&O�f{�%M�]�b�g�%�l���:�����v,���r��M¨[]�4�s��!u��}=0���բБw�zѐ7c ]�*Š�D��o,t��ӳ��1�}�1�<������n[
�˚���/ʔ��F:�#{���_���u7Y���\n���>��m��E^���xs�����tONLu�--ץE;�Kdux�7�$Ӭ��!��@��{�ʯ�f��'�\c~_>�����1>/9��-�+�c��m��!\#
6�$�̈�lG^�@_���w��?� ]z��gg��=y��Z?sn�A��������7I5$�̏�mda���!��͸���/�^��3����	�X����Ol��������r��z��,��|�������_���<��+��_��|���I�4�O�?�i>���,�Yq*���.�x[��JTTT���f�'� �u��}߻�'��W�-��`�e
�a��L�!o���X/���s(+��㭎1��7(ad(ՁK^x""����Ar�%P"���O2�d� �������W;�x����Q���5�<?wRS���
@]�=3�&�`�	�������� ��jḦ&q�Ϗ����f�Y܈z�EԖ��{��fF`��dQr��j��	[������;7���n���"���������G�X���E���&�����}�
2���c�l�R��bj��VIr޼A�/��I���PC�g�z�t�mr�-8�Jrl�r�f�bN��3�:�pcؚ��%}4���+��L��:�f��̽dO��
ۦ���������?V<�
ѷ�R���l7�4�<����n�w�A��]F�����)Em���6(�(��W%Q���
j�c~��C�ķ�������r#ai��\��<Q�S@>]�]�l�ph��ß�
=^1�87vfy	��ˇ<w*�¢���O�څ'
�����ϠAYQ����u���D?!Êm��R?)�Z���j?s�9`�/������G�߉_%)��U"^�s��z����n�-u�R?�f��
�0E��t'�sQ�Й��#��<V�T9�+�u�n>���+���ۯ�g�g�u�j/i���,��4K������vOn/a�;��7~att��u8����� �uw��>�҂������]c�������O�c�l��π%T�*�/�p���)oзT�f"�4�Xj��iAZ�����'��f�_PR �!�9����WP���$��+���7G���Dѿ��pڵ,��6�WaZ�#]������j����	�2�>��d�݌�|�|r��s֘{~|�lI�X	�\�h�������.��;<'�����;��l���`�3g� Sk��S�Ț���X�:N%���:Ara���Kнy�JR��u��9_�Q�o%9_�y�{+�Wᕄ"�3�)e��y�����Z��Ь����'���;Yۮ
_�U�Te�r�/Z�6w42�L��e�V+I:8��?!��EM��;b4}?���#>x�������0��~�C�y���2�����"2����zF�:L����k =���Q��)5�Zre�/�c���ӂS��(,��s�����_c9�4�Sf��..��]����k��]B��2��s���x۞�l�d�bq+�G�9�Y"EK�`LG��?s@y�$nJ572��4F�v��/������{	19�?g��['�mR��2u�V�a9A�\�Z�O��oɄ��̍c�~��Z���#��zٙ�I�-'�)Pg������̜�� �'�YVV6��,4���6
��V��*|���}_HF$�I/�`��$A6��ٚ�+B�/V?���r�u���ȹZ����ɪ!���i��
��,���(���C6S;�qB��"�Ei%��lB�Vv�+�Q)��w�l����o��y��������eY}~I��t��*���<���Y	�W�3 	��\
ױ�bڼ6��,�װ��p?�_{���5A��=�!�em��6ѧt=�2� �s�r�w����S�VN�&qN���a��7�Q`�٭�v"��濅��t�b~6�������޳�`g0n���k�1�'GFJj����U�Y���Ɣ`=�&�gh�t4�K��Aa$�<�Çt'T@?;5�Qn����(�+�8��u"��SxH�qj�3o�Rw�-��.|����ңj+��-���vX�z��S�NtT��	D�G�����g/��e0d�۟^vTI(�)�!b�iv�W�о������h?�]���Hx�3 n�1��
���e1>@1���|��B��\if"�8�K��RQ�uD��S)�sܟ�K�VTR4���ue��ȟ�.������Ȋo�}E�n�܆���6v�x8!n�E������da2�q0z�MI�#����{D��[U}�)UU�<�2H��F��0ލ�I�&���R� �V��,�Nm�R��S`a�v�������J膴�}<5Q��-�P������v^,%�KRe}����T�q�	�c����3��
Pf����.��K�Vj��Z���5�%'��*xڝah�31�wt}��Ud2���%�L+��!��P7-'q1�U>S�kh�e���̌$��?���	g5bE�/rm�.)c��sg(Z��n�%�O��	���ճ�(i2�y��*x�5y�(�索���%�ُw��Ep��A��7� rI�^�?��#�)kiud"me&Mr�~�	�D�)0�
�o���/g9;,�:����O�&��;���"��gN�dI���x;۳��u�Z�O ´ ��zM5�$��p�5� �ԥ D�3i��|���w j���4�bA�i�ǉ�7��9�"TU��<�o�|�"���|��q�L�+�~�*|�LH�i��YZC�9��d!�YE���F�^���[��{q���B@t�sBYn�}ppYK+ؘ���wM��9�a�]�;�I��y3B��)�e0�R���ҋ�Kڑ��P��v����6X�"w���8 ��=e>X�)P���F-R�eL_`�5�����o����Z��m�n�y�H����$
6���v��(�����5�Ύ�N� �^��d���x���W�^�17)�HG
z�R����n�Xa��*?�m�f�/��&����yX��h��o?����n��}���o <��ka��+�0`��������s�u��`t-�hi�/B��vM��*Ri�)YYw�Q��}D���:ϟ1�EJ�!��#�L<ݷ4d�qś_l�8omԖq�#�	�輜:�\0��o#�J�����m#e������W�
S=��9A"Y8��`���;d\�hĊ4�5�k�X���K(w�ӧ��/F������o��J�1"���#�!��5|f� >�*q��ih6l����.��s��Iz)��Q��t�p~?������Ka����4tw��ag�� �f�>}.����ۻ�q܈�q��m555��G1f;�Ϻܳ[�ː9���$�Lt���;7&�:)$�����'���a��A����%�o$H%��g�`�Y�-|'������'�(Q���?�<:�,�� ,�I���_���N$�*f@��!���`����w�5փLr'ַ�<�n|\�S��o"�zOO���ð��j(�at�5E�kE�R��عSvk"����+ڴ���)mUb���Mٗ�99Z�o��&����	<�Ƃ�K���ح�kj������e��,�DÛ��7>|w+��4�a��<�������cJ���J!��1�n`����N�$A� HR���Ŝo�
�����ey�p�+����P�wi��`�����緖i��:���+����+�_�J󑊪����^��	UP�Ŷ�IV���
{��~@�:�_fv�:��F|,�-2�D�\e5���F(}��E!��.���Ls�����P#�#͙uI��O0	ؽ���f�IjK=Ԇ`��U����Й�{�]N��̩N�
R0������I���Ko��Hƶ80��v���N�ҕD�&+��b%~)V�d�_���'�7s��'/l˒��	��<3�!OʘWr�@���\b&\���d��,Ƈ��[�Ѽ�<�����ףQ����.k�VGkC��aL!���+dQh���*+�8��]p����b�V���0yc(y�)j<�!�E���ev���\a�G�m?}F$3����9l�_�U��1A�ΰY����JܒXe?�%�0i�w}�h|��z�*�H`(;���ŋ1p���V�[v;v**�ڷb�ۿ���D,).^^�]�7��YI�P�.H�	~Vn�t��P�8u"�͉cDu�K��5��>�4����2��:i����EMͅ�,�V<���c%�f�qf{m�܇�:\��6�o��"cbT�[كQ���;�BC+P��j��ߺ6��x�ɒ{Y�������s�G�z�*"�Ա�(� Q�i���A����<��į<[����{�m�|�5���黭��7mڄp�y�:('P?�*W6��r��x9W�d�����s=dn�Ռ���&f�-8c���ߧ����-���M.M�xڙ2�#�a�H���0gv����?q�Y[g��3��r�,꒞�*�1Q��r��O,)Q��;�����C�o
�/;�@'쓯���ξ�������+%
L�x��Wá}A2��I+��������~�rs��9Aa^^^Z#�����QCk@:\�f��]�90���g:�rR�a>�/�� ���)`�	 	Ώ����D���W�x�}{����Җ���4�%�G_��l����А��P,���5�9�X����@�0Y����^"=�Y�AB���=9��_W���1�̭ͦ�i��8U�@��0���=��������C�TF�$! �������/^��%ޅ��#�vU������w��8�0�1-b�A�
����M:ĕ�s�U>��7Z:�`/��l�!�w�s����@s��!��RR�2(���L;+d��`�b��3a�d���c:�56����q঩u�1u�ʭ���w�����d����vBY�$���x� ��]�l��
��H�Ǖ?�����@��m2ǔ��b^ ��7�'�(HR����������@ތ������CGRF�	�'E��Vf#�M�74#��'ؔ�O���i�5$U@:����L��-"��ߪ5)�����m:0�'S�9�,��u�-%Ϣ��ZV��>I۪te`m&j#�Ʉ��"#���n�$
1�\A��t�q��ڣV�@�F �y��c��xC�i�i���DSj�o��J�RSSe���R�n{	�MC���m�z�jL&N\d#�;��-�^�?��@������k�İ�V�F�y�^�/�B��K�,�J�f��--.����R2�o�S����^�O����娫�[ U5>F�ռ-o��g�6L���R����\k�6�S R*}H=3�kNS�*�;�ؤ�Կ6�� qF{�aN���;S�u�ؠ�?`^�!���ia�{OI�3�=l�`���陜a���빴a���ԋ���S=(��������A�"x��d�T���:~�3'�v��g�R����0��B�	�si��Y7�y���^�צz12Y�b�p����mGL���f.3g ��ӞnC�G�)��+_��I7��퐻���k�+4�h��b��d��{�ye�D�iX��w�s�|�gcB-��]#~�$��_�V���ˍ~f�IDEE�0!˽�㪸5�����;+֊^�ږ���w���ʣ����pa��/����lc����j�E+�L�3ڙL@v���.��|����/o�B�ҝa-}gjKѳ����`%��y�t���We=hn�s���更P=����bp�{y����5U�k-7�^��|).u�f�Ue֯_���U�?u��afZ�z�m� +��uU�c�P��MU�`��s��GM5�)�ni�%��35[���h<	���e|��^E�f^�)�PJ��0�1��t�sN��0�>�A���%c'ek���J{���i�(@C��#���!�S��9{��vŰ���L����*�~��&w������Z�x�v[�n
����~ox�T�Qa�x;�C=)Gz%�>E냾�����eRX'KW_2 m�ަi��b���M�\�r�ڍ�ʴ�����pm7�N���u�w�[	|Y���[�Z4�����A}^�v[5�v=/�����d�΁��sSG�i�-1w��g�/�ɡ�)�d��`ʊ����!y�U�����xu'��{/_S�z�ǘT�,��6��c��3JW���G��V��m $�'�t����A��`��9���/_ܽ�[������ >I���w�1-�.Jzf�3z��wW�2qz\�_��`V�9�ŉ~��j��}H[�j�H:�5����G����>��$__ҹ�'V�בm�!�VϦQ[�k�ϼԜ�a�RH��n_W4]���i������Ļ5��nm�aKՀqU���.7p��T��2$�2_��	i�!��O�`���*����'�h��y3�����H��� +U�kE��)&1�!��?�6���O�kSϫ�ǭ�Ĳ�V�t�QS���8GE?प ����KZ��wcC�P��3Ґ�C�&9�\3�i��эSm(T�Ǵ�'�D?t����o�_K�b��%�0��[ k����,<4�����n��-<5��W�FV�x�P�L<nլ�laiY|�UP�d���/_2�D8D��5k֘��´���΂>���|�r�nB�P��C�4+]}0 ��g����׋�]T ��t�3>|OH~C�� O���j=���lIW�%#J�1��)�λ� �D�z�����^�@���N8�f�J��L��[n{�h����|U���ܦ�G
��o�|D�(���8���P�D���0��A-�3;�ӉR�isNG���7�>��Z�G7x�x������#�}AMrh#�Q��D��'���Ԗ�鑏FQQQ���99��f��E�X���ꝥc�ߘL�����c�AG�AY��i�:Z�TT&���J� �?¤
�F�'����i5����[�9��JL�~%q�:Zڝ��UEwF��unڼ���g��\_�DZ�b�~������O&���K��z�	*����2��:�Y�����4�xz��8Rt:�`�"�ߘb�Lײ�E٪�,N���tR���|/�"�W"�wh:-�ʅ�6c�w�b䴴�YB�m9$����x�`f����8y�^s���z䁹�%�n�����&��\=��d4^y��9�^���(�-���'� ���6�B_��=@�fW��g�J���G׮V�uEB�)�&W��={v��f�ˊ���L_Ԑ��<�� l��s��ZQ&u2L6�^�b���R,��e�����aː��%K�Q���Auf�f��>{��S\��W��0b�,*͎���<����-%'0�����E_��M�ǁN�+�C���U��.^$x�=���xd����<��o�׉���
�E�w�"u���ݦZ��J�Y�Js�T�'$%-NڑLc�3��'n�vZ=\΁I�!��Q�3-=W]a\%
������4?WW(����2Р����c�
�?d��"Զjr777�"���o�V�h~d�$Wmh�U#��f����W�1F�����a&�F-	��G{}�0��9\:�ƆQ:DG�r �Z��s߻����c�mѵ� �����Z�'�0��u�)�Sb�ݜN�X8����s��l�����r����I�g4.4��,�n=<�I����W��S���5O���	~*q��	ĸ^�ĸ�,)(�'�0����:@A�����E駯^�=�>����Ī.0�:B�$���ʭ��K&}с��� \����_[����]��V��QUի�l��j�&�q*ns�6m:��j�F���1���da)l�(CN���lM�)`L?�n[4����'i?l5�̢�����݄Q>Y�GcLk=vn&'�����),��Ւ{�˺��8�}4�&�ݟ48(�{�@�����I>���X��=���-=�(]7)�������Y?�j(R[@��� u�g��G<"�Wm�|�"����������p^^^���'��g�^Kw����ߋRv��tb�+�á����' }C3�_�g^a��ݦ�+��T�;�a*d-=~�P6�ꜳ`&���@����UƄ���9�3`�g�K��a���j�Y'��Έس�HF�=���4_�̛�u���%���$�	��[ۇ6F���w��������Hy14iua��k8�zt�=��T{{{��5��B�~s�0m��{��vs�,+�u��h���o֣nn��RC��B�:V"ꕈ�0 ��g��8��*����묱������JӉ��Po����M�̠��1}?*h0�u�g�\�����"]>5��g�R�%�IaLzE�茝�6U����ٮ��#5V~�Ӵ�Z�dB�*ԁ����?N^9��+'h'��[K|�#��=t��(��ϴQ ��0ƀ5��G/TѶA�ž %�J��Y'���7������$�i���^O�d������� �(��Qþ!u�w������z^�{�%~����2�����y��T�v4��{~�5�C�����,�l���r)�}%�f"ԇ�#�5"�9f�nM�g���JJC�{ï��b�;�z<�G���D4[�kw:G|%6rd^������l�wQ�T�u�hW��ܢ"x���6L��.kV\��P���0�`h�"י}%&i�jdh�֠�Lmc,B]�օ(h-]T��yb��}�����Y�4Q�
pxf*��3����b�ߢֶ㩏�~��*[�A�
��A<n��E�SV����#	v8����q�)�F�8�Eﾼ�zz�Yn�`3Q0�j �& �6���㨁+���*;2�Q��Q����։u�T�sG���Q��Ժ˨�ɥi�ΉPWZ_�3�,uuuO;:>�]UEu�p/.�
��)����p<=�+���n�=��k2k��k �2�j��â0ϫ+u�"5D�#֘��i����gP5-�t�G���NjM?�>
��ܑ���>�h���-�d���c�f���s�\�hi�M0_UeN"�);�jj��q��h ټ{��m�#�C���-�"���¢"�%�E�2!�+�� � �S��GH4�,���#`a�Y��s�b��|0����ї��b�����/��f� �3unS<����v�a^����VǴ���\zT��7�Ǹܙv�1�{��v�B���U�ҫ/_��B���&����"�pkϽD��h�ݴ�^@��.���&�D�$lf3�2�(����ɍ_��:?=�臃�:�1��1iL�%�C��ͬ%x�fV��~VOV�b�:(�c����ZFZSE���="�n��o=����q��N \p����t�A ��~��BV)���yޣ�QRɛu{��g)�9��y�<4�t� ?y��*�	�L Sd�ؖ��@,�O?J��T�*11[����v7?:�?MN	\�<��='d��+!�Q}s�Q ��8'f���1}�Y_J%�'�k�*|c���G�R�z���!�\�u���;�m>S�F�3G�<�EU�!%-}�c�A� `��sOw^�=�Q�"Jʯ��v��Yҫ��s�/��\5�&���l?��N������|\�C�v���تΧO��*����q���/"ۿ
��w��D�.�H��͐�ʸf��^,'��v�ij
�III�xO�F�c�W���`0/��ڿ��n�.�b�sX6��^���[�m�5*M�d�`�$��z"*C{�u�a�:<��zU:_�0줼U^nZŀ�df�&�D^��{K�K��Af16_��	��t�z����gcB�:{��?X��w�y'�ETP hK:-K���+d~���-��N��~ǾH���sM¾�Y��Ѕ9���8�tP���>|��C���ˋ��7����KO�]fUr@]���jjN]�r'yW�������}�`}j�6S��5��BL�C�����T�f=n�>��H�)�ß��:N��-j�2�|.}'-X��Ø�ޜe��������{�X�as#M��ir�Z�.b���0�r�_�����Qa�RE[��E_�`�������8�uϾ�2�?+�HKe\��O'�1�
|��߈���phngo �ǐ�y��F��9�F�S}ۥ�ND��-|�8q�������?��=���{�sRJgQ*�l:(rl���S�U�1��ەj'���+�8�S%I�3(bbFL��~k���������}����ܻ���]�����Z�V;m޿�Z�{�p��w�����֞�$� ��{�_�z
G�E�����<���DnT{���@#C����\��񿙑ӳp�Z������x���CE�i�6�~�z^�f��z#��Q���N��'����R����{˿���omREo*��Z`}���]@_(�>�=햌�J��vb�!�_vwv�J�&%�7yN�|r�F�����ג����HW�t�j��^�����I��k���y���|́������A�E=E�KY�����!�ϟ7�<�[�?���#����-E�!�����]	���,���Ԫ�򢦀-�Dw��	�b�7�Eg����R֧��tI��q���"�����F�GN5��澇rX~=$��:Tl��B\�Q��W�<w0�;��s:������D�%zh4ptQͫ���j��A ����m��{�G{�]<{���	�U���A%�;j"���A�\�J8��^=ł�;,�����0���[NЇ�%Z����*H�f���>JetTt[�+�zį��021��R�*Ɍi���a<�Hd�Ї���0��[�s܂���	���K�+ċn��%U>�+�>A��@�|I8���Y}}J��o��}���������z�8�S�C��y�[r� )N?$�=���|��vU�=�-sU�B��IO?�߭��uU�^&v��|�tmKU��Xu͹#�g\,748d|�Asd}џfm4�u�����i�b�ֶ��[}g�*a�>~�mGO����x�L>�8:F*e�H��22c쑡������U�G7�S|��i���Z+۫�YK���i�/��Z,7J��wL��[)^S��[Z���<ڍ̕��3}c<`<U�pwS�@��K?����V-D�͑�Z�\��Sl�^�؋~�8�~3a�U�%J������ô!�k{��-~����x���m�N�ށ�{S��%J�##�p���T���H�ƠX_�0�Ic�J��SZC5���)#L��S�T�r�w�,�C�{{u/N�7�� ��R��^4�ׂ�u���ǵ-��uhJUt��O�m��%���S��� nƁ�Nq�J�	��?�]Bl���Yד���K�>�Wrݘy=(P�z����E�����3����F�B?����K���Y����Q�Q��P�.�"�̕�D��ݍE���J�7J�c6�D�@�U�\+L�����W�B\k�t~�@��O	˷]�쮵B�>P�Ɖ���*U���u�!^$-.��a[ҁ΢��?z�1�!���!�]���J���22�Mj+Dgp�s�3��+E�����G�=���O�a�l�{�9�X7����MAZ P���J�k��n�"l�u)*j�7ab%��2�~F�t2��uK`�d
�ĭ#e#�߹sg��5`_���4Ǣ�;ʋ�A��@�n�h�L|�qi$��!om�(��������c�}�n�/��U����μb��l��ӧ�z��@^���/i/�ۨ��9ĕ��N8�i�UĽk`VX������FX�y-����2Ư?��N��m����UD����k�?o�u�u��.�B/��Ϸ} Q�׶H��
��lK�\LθE������Vb�XD�R�2�����.�Xڿ5<m(w��н%�[VI�����N�ܣ�V��ǩ~�8�l��o�����%-�l�ӕMo��0�}ȿ���J��}|_���İ������gn�Tު����s�.�uDg�R߾	�jUc��F���D�y}<bbr��@���]�E�:-6��_	�f���su�6¾i	��Q	��u;.�kkA���N�����
�/~���yڋ�.�����%�p�9,in����U���T��=}���Z�o=
]��Ztl�pء��kס�X,�������2г��������Mj�܇����&G>��m�!)�5|d�Q)�S7�X��MQr��n|e��Xho��n�Y�%��3/�Zy�qgl(�;T��3|Ϡ(��{�L�q+{e���sO�1�����O+���G�x��@[�W����eZ�{��b���:>rq�4Y��A"%��z˫ws�/��ߩ�o�ا��[D��a%��+ʌ�=J*�i�Y���$v��Ú�?~���IG<y��RWλ��ALL���쇮��舷��A��x���h�*����,��ЧF�QI��ѵ4q�����lev�]�iR���Eе�3ĝ�s��t.��U*�%���t!��C�-���@N�1C9{ v���˗�/0�^�P~�;-�ll��"����V��e��Vܾ������ց��x�'~�5����U����<ߴ:-Mk䟒��=���i=ֳ��
��.ھL4+m۲�Wy�B��֔;�i[�GP�������/%�U�)���k)��:�����fQQ^��+�->V������ :�F����\�@]ےX�>��xvk�,��j�{]ۼTf��
��m��|G�7���m٬_!3f����>2�x�#�K{�X�;��CK���p�.�	����l �i>^Z$Y���;�jތ���A����u)�?]$�-Um�d�НW��*�k�����A0�I���X7-q����K��Z����󱗭����Qzc����H�F*@z����W��vikk���V�hO��I�o�K�CuJS�6�u�j~s��(�/`56��Ն��*B�Ӄ^}~~��xq�q�R�}������̗z?�����t�o��̀A��_���V:T���&q^��� ��x?�L�ŋ��G���2F�%%�֖�����}����o�'�*1,$��qP[ʰ'~���'2��XO����ʮ�A�;�7�~!��i��7B⹣s������m���k�.�6�/o�H��9�PǊ~��)��j�W{tQ�Ǐ��4"��:z� �����Ul��ږ��V���֓��i?mg.ۡ�P�H�� �v)�Lq�.��G��ZVɄvr�Yc�~��?�;���1�,�sшju3�����qT�%P���=8���Mߗ4{���G\�ð^��2À�����BmQ#��?��y��ޑ���mn�&W͍�S,�oV���9�}Cu����eu�-Ť���VP�\�raO0WM_V.���>���Aߩ~i�7�V3��%#�1�<0b�Lg���ǋ�w��m�(����V�C��OE$�Q]����U��[���V���_�8V���0OՕ'N�/=�NЈ+&:��o����T����J���*����ሎ\|�d���X���NՀN3���Uw&v1��W�£�w�p�����+��f��dQY��t��؝W�ꔕqdO�f��fv�τ8Cj;�#�Kʤm�ꪊSx���=���x� �׹�~o��xݸ^��뜪*b��?PA�(�T���G����C���^�&���rW���>m:I�a��<v�k�p��x�!�|��Њe��+)��@/�cm� �XA�E�1�k���	�Qz`y��G��x��ʹ�k���b~�4e坧�E�_���?�4H���?�p� ��MU�	.<��G��#�Z�H�׽5�U�$��^���'�1���_���ς���So��a�O�<�Ղ5v��?�[�·����U[��)o��̙�ټ'�9�R�:F���-��s�j\���T�Z)J����xQH��JR���=�:�&��D'&{���4�B�x<r��;�H��>}a3����o�0ͽi�aƸ������OD�-�_�U�2�L� �T��XL�$����?8S�!��狭���w�tC�y#+f���5N��L��I��xΘ�啄�1�%�"��d=����o��~��P��t��B����/�J~m��/n>)�X���L�h��1���[���Ӳ�'���Q��{FM�J���Zd��u���0�>�����}��Jc���x�1ۗM�"^����݃����-����2�\��� ��E�=`(
�����JO��Y����ݲ�����=ffv�9ҕ_�n�E�kaX�5�F<5y��Y�y��V���da�o�A�QĂԮo]e]���)�.]�g����Z�!c["`zZISS�=v�(���ca6�y{�&o:�؄!�$�E>��#F,P8�H�)�]A�P�@�������_t�=J��͕�ʎ��I����%7��b����J�]P
�o�-�Z̞h�l��diq
�{?+~�r('¶�Kw�OƋ";����pg<;��YZ����HYB�ׄ�f��!=��5���]�LH��QB��n����II�9��9s����Y�'��% b-c��l#��6��	,ǘ����:�N� ��_�D0It7��s�Z�+k	��T��6Gt��2
_�"�"��������
e�:l����P�p������A�9S�R���II-�:�p�F'�I��g�/�x��Bh��N�RjJ*�ZP? 
���n�?Y�S��<��&w�m�|���R�ާ��;4��R�H!���gvI�09D��G ��@���YB��M`�<O�ӂ�����㺧�&~6{������@��}��U��D �M�lZM�+ODMs����=���X!�骺9��F��eC]�A"D�{N��U��ϛIӉd۾)^�����t���E&��p�r*�3��?�4�n����P؀��(��xi���͛qMv�41)���U�Nȑ#�{W�:�p���s�ER�9pw��ݦ��]W�{���e��zn\���a=���`�Z��˺x�qI���C�==&N���<J�·������*�Z�8iBl�*g��K����򮒓x����c��H������3��i���v�&!oK��\4�÷��~U�����hbm�rC����c��[߾�
g|��g�NǤBn�s�C/�J500䆿��oyMxj�fdf���b<�O�x��004tAE�[��/���b��׮Hg�$jY��ϱ-:F*����ƽ�u��߈3��Hkqiz�q��czs�Á�
銏���on���5 e�m+3��oHa+�q��W)�&�9���wo�=�UR��]:@fj<�#ǻ���p]峛��I[�-�Y�^��Y��a�8��$&&�AWǧ;�D���
u<��9AZ��[��-Y���C��-���Ȭ� 3?a�����|�H��� �pf�)����!��J*z�s��lZp�Ƹ�$<���U�U��V��Q�Ǔœ�R��\ލ���Y��x��]x¨�k�%EA���wfg�v��Q2�����[�N��w�����`��D+}�2��@�MC����)�R�9���TՉ�,%�'LLЉ�^�+m��C-�T�;��C�8�	��ء͞�W���OM-{��߶�K7z*V$/1���{��Ѓb��̻�ۏ�ҭ�ׯu��_��w�Uk���ku&����-3����pcT4~4�&M͐���LU�9�Ľ��� �@�`��W���).c�ά,±���bt	��gđvzm#��n���SNWOGҠQ�X{�(X�S�����I�!T������7#6�C+zn�j��y���61PB�{d޿H�ƌ����N��j����o�Ȑ�^��v�ڨ��#&�ǳ\��<pK���8���E<z���"9�(-��3P
��X�[Nq�F���S���#eQ6�sp	������4�r��$j��Wm��X�!ǃ�G��,V��^k^�����d�wk8���� 	��7�������C�/P8�e_�(;4�w�grHQC$tq)!7<sfF��8:�n��-��*����E&\����9�3�U ��P�2��ۋ��@�HMK)�'���
F=���`�A�݅��7008�i��Z���	Tf���~�wUr�ԠִyӔ�Q �����!��j��-�\U���+8�2���\�C���NC�/y��Tv(�B�A�x�#�/`�"�[�M/��9��S�-���eN�ƽ���i�Zy�s!^��rӸ��N���4<f�"&��J��ޫre�l�C�}�6:5��>���T��%�=�[���aR��4�z��:T�88Z�$��=��[W�A���v����[w��B�����'�_ .��G�(����g���.�Z�����������(����D ���n�V�'C���肂���8�����7Dl�D�@�
���*��.��[γ^9(�S��ǜ`HFğG_0�bK5�h�!�=&؞:�c����'�z�F�@f��-�v���;w��ǥ�����⿓6�\�B�5@K�y�!>>���D���'�`�C�����ME�!B$�{��M������so4���3GxM{��Gaq����ޫ-�	5����BF__%�=w=�k0�@�v�h7@�>(�Yޚ��{��z�و[�{6ɀ�yȇS˖����NX�v�F��DyK��y��GL��Eo�wUNIQQW}�{�w�)�h Y\��n6bLz_!o��>f�����v�+�9��_�9�_l�������q
�2�!���-J�A_��ݗ(�Q[�}�'��}��Ko�=�MA-9@Q��.������FII���ƺr h���ɮ*t3��r���8$�,�*�*<� �PRJJ��?��	�H���-5��`�2��`d�q>��v�l*�:��RP͹0��dZu)���~��9�8MN2�pU�9��Az��6�0�8�#&%�r��6M�P�O)mm��|{�Ǟ��>�}6�˦���:D^��i�2��:>9]ǝ�i����!�E����g@u �����Y�z"G=�ȭ筹C� 3�yx�;��U��9����D��-�O�����q�LilIȏ���z��C<|��
������@�;�AjÃ�� ߣ7��IzE����K��<c�];!̀u1%5]4hi_��&6���J�y �h���?m�M�t�NY�#
��O4 H�$�q(Me�7�C4XQ��c9�r�P�P����X��
~�,���fL�������WG������xo��"��W~��~��,qt�-�;{�ȡ/�X�H�\��9���U�m1O�pvw'�\D�i�͏�	[(�=�OpE+ly��!A&�`|�'!]�rK�*9n��;��C�SR_J��&:Gr<��xCP�F�r���8��%�lz)/��� ����s?����`�|a±�ĉ���)	���8@Q`Q �#��ă�I�)��jϗA��x>@u�0���X���	p����L���ci^cHh�]M�ALLyy�QT��=^Mˏ�{@W��� L��ֺfb�.&b��R��C�v ��>�3���PN���n|��y�~6͈�����&���C���#3c--嫫��r�»vi#��K��{��YDҮ���r\쎙d�S����#��[�r�OB#���&���Fu�0j8��ꐦ@A	���zO���n�61ߑ�A'C�?���
��΁��~;�.Վ��L�m��U:x߾���)`�H�^5�Y���Q֗��A�'%���m��]׷��#m ����\�W����B�b�4��)����b�`<&�]�61T�5���8�ӓN��݀N���)K���������]sO)�({�d))�
��B����'����Y�h�bH���m$�\�+�O�����9h�9Q�w`f��|��h��
��!�������76�!&&J�@��i�*�ҡ�2��B�a@���TF�Jиm���N���x�]+n}h�|"��G�:	�I��_��

T�<؏�����e�����!���� qQ��<ol�#"~�v�t,��Utjg�[1�??�Xw��M�ϻ�9�켇^5W�����b��;2uH����K����q��m��d0Mx���,r�⠙1R�{��G!�ZnF�l�����NW���;sC�bbNe���@k�MõI���CQ�qk|�̐}�T���(��jV[���O-R�ׅ�K�,�"{7$�8�^�?��'�G��ʦ�{����B�Z~A��}x�"}��}m��S�_�OՀ♑Ac��k�r�l'V~����TO�<�Г��^�����mU�1�[�$���O;�����UgO��+��Z�Nb���H44��/���y�V��I�@������j����lxCG��%5Y]��4u��0�g}�;���Qu��!�L>\/ g�?���mAձ���R�>�6��X��)oD+ȍp�^8���ҕ��{f�2>쯳B�Sg[l�!�|����ϒ��PҚ����	�q����lK۹�����<���p\i�	/+�C?��\�e^���/�f:�H��f�GD|�Q��<�|�〚ı��E����Ծ��^v�eш��%����B9����5��f��Y,�lo��hϕ���ܻ���)@�G�%O?ʃAyf.���A��:��C�0O�!��$�	L��,�Y�hu&��¤���U����>��m�|�خ0U�r�G�ƄWzz{�ypQ��O��i�8�f����@Od�xF������?������+�6�}j!r���aR��n����` �i�8/6�e&&i���>�띬��,��
��G�L�Ad��{0(Z��)TR�nZV��V
尤a"o�h"�՟QM�Ro$ؚ���r���d���5�.�_�Af�6��A��Yzc`�9���B�L�����>�����M{D�P���K���Z%u�����|��f�h������S��$�o��_�,�uyf��'%�y�<6v%)�0���z���tl`07��gxu54Ed�u���J��Qev;oa�<��N��ic��7k���G[���ÄiY�g�(*��B��w�}�ԓ�<Gs'�=�;�g��A�Ӗ[O�dV��������(�\	������]�b9$[�?��}&�����|Aȗ^~��
#��<���НQ�e�?d枣�Dh#�8Ňs܉�i��{�=��P"���p��֏~_oX/�c�4���ǫ<�R����~c]W����cC=���s���4H,�S�LL8:��_t*��Ű��v���e���||��jb%�֠WtiPW�FI2ڏ>_c���լ�<��ZQ�Y=�*�h�7�� Y�xA����n
y"���LգL7�M~�Wղ�"�ξ�5�LZ�)�Qm��i�� ��+�"�r��ή��aC�=��#��M��x��Q�DD�DWX�(&�C8�y�;�v��{@�R��@�'uL�Z���ƫ����*�[_��i�6�kg]J
�:k�Ԃ��`/�ԛ�ޯ�c+���0Fa��*8���:��ߊ-K�=�P�{Ug�B�a3��S�Wcf`#�)r1�ɐ�*��_1:/Q矇��S<��R����OD���3�o{/���kq_�s��^&àe��v�i���8j���T�P���0��B��lz����ޫ�,�㙆i�$�y`ZZ^u��Q���)���ϰ�Wh���1��P�C�|�O8�!��+(��2�#�1VaM���[{��Yyvj\:��
��aZ5Lf�x�tV�\�~ٙ[hy��q'���W��>i9��{����0�PT4��G0�=�mX��x-����`xi�09�"�!�V���{-��G�h �h\R�=t�����a-��
�"�ן�w�#&���C���_pj�#����<�L�O;��>����հ�"e݇� 6���U��p��&�5��6��D˂=�ȭ�8�M�Z=�v�9D���PBT�ܱ0�6 q` ���f�n��[� Z�� �ͽ.T7�~��׈f�u���Q$��e�r��{�|c� �k������}^�[Z�����>�ڴ��~?�?{�X�)����dH�b���H����?���Q3|J�L���,�g2܁� z@x,�iE�`�w�y����J�P�/��lvU-k��9ڼ�Zɚ���_��6��p Iy�C#(%�����;�(L�M��%v�$��a�k�5T+�>y4/,(���=,N�%�{�X�Au������J`VH�hғ��S�9�Gu�K�q����z�d�8o�ؤ�$��������4<�=��!�k��,�(Y�	���[�ȸl����&�dF�]H�j� ���]%ڀ�^r��UD5c"�avX<�ch�o�0��8-�o�;i�"D�.4�PݨX�x0��ͩ��R����i�RWzK�@���X���T��O���4��<eP��ұ�)�?�E5�z�Җ����������Y-&������S�*b�]T����Z��;�^�;i@}�t�_�hW�%�/��axu��.π��e��`� �I} C}5d��ѭ�D��]̲kj|�S��/��T���B�.�1�c�x�8���
�3��Eo��)��I�M�Je~�0���
"BAbL5e��IK�]�u���U�[��.��{9D���6်�p �Y�U�J+nR�&��=�{o�+6{[���t���d?7"9��<[�v�׼���;"�B�k@y����ޛ���E�����b�����5+6��E���[~�wk�3{:�#.0#��}̦��n��ٓw���	�"vZ����';��/Z�����^��%�e��S�}�[8�����<����[�Ì��,�(�s?�z�}�A���۸q�^��D�G�f�[�[�Ы�ߋs��V��H�/6`�׍��Kv�B�H�X{���;Z���<�_ ����M���B���e6�z:���?9^�x�C��ó��3�����o�ψ?��$��VO���(r��_36@�{�昴�c����Z{'|�h��?�XO��P�L��9%rJ��)�S"�D�[�p�O8�#���O�E[�jVL`U��U˄g7�&���%^m�k��LF�v�V<Q�i�'�3{�D�E'�(�&��e�6֓l,�dƔ�)�S���^#�oG��B���U�����z��k�#�~�U�0W}���M���i��ٺ�5����(}��4!��z8q�f�n��肓�6��8%pJ���)�S�N	�8%pJ���������0~/���pve�[DE��?_��؟��6��cy��ek!�1s�N	�8%pJ���)�S�N	���޵��,k4�>�c�,,�t�8��`�ĝfi�	[a[NOR���@�L	�8%pJ���)���I7,�d�`���l��g�O�.;�sY^o�@H��r���fL	�8%pJ���)�S�N	�8%�_E`���4�� ����c��9��y��IuE��)
�ϑ�Fa���n��0_���buS��O	�8%pJ����o�z�Q��ʛ|[|��?����u�2k�s����n���^~�VɄ��,�����֗��y���f�f�����т�qEH�&��Uf�/dWORj��n��:p����E��ǰc��%4�� ����?jkOV���6�<l�+T.tи<��y{ҍ�t�(I�'=�D�5MaVl�G?�<::���d�����P��d��<�xƪ휚�g�<�>&�#�#��Y2�#�Z��a����j�����2K��bb�GcN�������hkv�Y��cDD�p���ž,���u۱�%c�~G�W��zFinp3`�Uu���tO�{ڤg�Oz|���I���I0<u�ԁ��\��#v�-�ώݨ��E�8���O�팬�п$�]�UjH'Ǯ�#z,9Y��0G�VC����L�o]�X?1;^y��R��B�M�fr��y�`�8���-�H!�����K���k}�O��(wqN�h�۶{�1&��;9O8s��}�4�Ӵ�a��Q`�����)��զD�6����&�������:���'�ycY����T,*r
�`t�����$iO��O��:Y)��s�[�ZZr87S"�S6���!3{�^}�Q�ݺ˿��?��*���V3��f!�P~zrt�jz9IA�ڗ3��l���)�c�����Ȯ��x�X:�\&+���-4D����'5n�V�W~��!)�}괜7}������;u�ԁ��*=?������^��ꬴ���P]wee��3z�*(gNe�Y(i��E��P V�۲u,H>�~oѿ�4u�ԁ��^���T6����n{V��J�e
Lɗ�$�>�`2_s�����J���h���IV]��D�u���\����i��ѷC'����F[]��q���]��'o-*����tJ?�q:y�h�_۷8ˈB�vv�8FZ�7�� ��J����n�K��2_�+�F'`���Ts{��ȹ�M���l3�r���)+$�ȯ���Q��Oj{�-�� !�������8ី���s�b5��b	���i��Wd��T7�H�N�a����7���ၤ��;�a:�~ޘ.b���O�{w.\���1��PE���ҜNV.�L�[��O��ɺLn�'i�p���'?TqJ��@��>��\鬖��m�����年��ń�?=������B���u������&��j��]>��M�y�|�ǹ�h�sΊ��
X�Yg�(V9d��J��>��Tz*��ɘ�(X���1�{����m�7%pJ���)�S�N	���$p�<��xv�kh���~7{��L�cϛt ��/eƔ�)�S�N	��/.p�W��ǧ�σ�e}ld�ݝ&Z���xb�����5B1�Dg�_�.7�;���{3�NE�4I�c��p�<II�œ�{2YK�I�O~��ѿi0蟽�7�dk���;����O܌�)ҟ`;fST�� Kd��w@�  �=��m���IEO�ȣ?٘��Jsl^���ֵ_z�`��m^c4%}���Y8mN}o�M�X[��`۶�/�rVE�'��Pл�nmZ�z'�Օ��Z������g�&��GQ�[�8�u�*��Μk!ܿ8��Zu�H�t�_��>EK�t��ҩV���v��w�v_`����-,XU}�!XjGQ���ZI돨��2
OF�e���O�qc�=d�&���]�TS�Dy����9��JN?��?-������7��W~�/���H��Q��	����te���M?F����;�aоh����uBt���7��,��~�nj��0x�,\�H�H��rX�f��HQZo>{���~�-�t�3�Ӻ�oH���o��'$�	���Å�i���Gb�o�{�}	�R�̽�J�)Je���M�`-��b~+���$�7r�#׎Q��щ�|�S�������-�e�Տ����k5�������O��;����G���e�GY�M���Q,Μ#X5�i�9V��Pa���a��]��Ƹ���J��zչ��'X4����m���΃ʆ�����g���[U�9/؂�>D�[���O�՚KjQ������f�"�t<�K�ܮ�-�bJ��,*�ߤ�װJ��j�7���+6f��]uL}�b1���Q�Ƹ�A3U�me==adx�镴��вjܢ[+Lo�*3�_g�̔hy�}W��M��S1g'��Z�d�=m-k����]�����^�_��K��zϥy�������Rx����^�c�JZZ�~mdg�����IO-�R��-8�#�H^e��Ơ�A2��!��<CJ�FbB|�ʫk>e�J��$���}�z�췠��g�W�}�.��igA-0?۾��nᢜ��/3哒���N��G��L8����?�T��y�fa�Ӑ�f�F��Q:sa^h�FwA�;�����~V��1̧҆r�3&x)O;��۳g54_���'Y���[�|Q��]�K�{?ƻ���_�vWf�*��%�<Ǐ��yu�o1�C��~~�@��n)R�v��ڼ����l�k�_���Q�X�"ȍ[�]�ٯ�h�z���k���~�r� nէ�}$$�v���Tf���~Z�X���i�NӃ�!�R�ຘ�O~���4H<��>���08�W�%&&:&&[�{!(�,͞���uN�6�m���6Ze�oi\-(��_�nΚ����j�z���$�L�J��Փ�Β��"�����|}�����ڼW�߾$+�+N��zut�=��a����t#<zPA7[��l�|���4ǨW�6lo?K�d�㒚�yL��i��_yd��l)���;��S�ʏ�+7Vnk�
9�������Y�z��U�B���B^��KL{��>�����
oP�F���T/�j'K��'3U�(l#�X���8�9���ڳ��DjyU` ��T�BI�+b� Q�^���8�j�='�%5v�8<���Æ�QA���AIt�Z�#�fc��m��I�ѭ��#~�&��6/��M��U�z_-�n�k�+�wXݪRN�t|��'ep�HW�j�p���<d���v�N�8ʹL�T��H��I�� HԻ,{u-����ǉ�
{0B!���H�W�=���;��2c�K��u��*{�#�C�,�a�*H��߻�?���. 9lV���lZ��!��Gub�/p���]�O���k�����a�AX%_9a���2��y�j��tnh���G1�{�X�bik�fj�Y����������)�â%���/����nT\�ȏ��\P�cZ��m^1�7�7)3�r���t�_,l�}��H"�κ"P�<�Y���C�m�K�\:�L�
��ԸY�W�ὐ�p䝒~O_�D"E�#Q/qI-]��l�Y84�I���ioG0��s&l�<)iHv�� � ����B�;w�����L������k"��
�J����صe[A��%5�Ű4�6N��"�����*vm/������l�i�߲��z��r����FY��!��P�9�6f��.�aM�$���f�`2END�l�|���6�
�̱��wژ-ѧh���#� �iz*2%'�#�{��}/h���q��R��iH�f��cbc[�gl��ؙ���;�s�O�=�_y�u��`F=�R�m$ Sn���	u�:�6��IE���8�Z�A�����(d=d4��	 eP���%�8 �Z�c\~0�|��Ȏ0(���D��Ӟ�8�.�Y��s����f���R���]����`��!zw ЍK)J:T��@~�ד�bZ�TJ}a��^�1a�����GM�JtAsxY�^?��nm0A�(�����M�mPI3P���|�Kjd��*>gb�>0HT�ː��V���V��7k�[T����T3��a�����!��K�u�jV4;9�%v�2��s!��4��+����q�ڵs��	ƪ�Bc��{���Z�*���Z��li;A�����0���	�����&�b���4��ő�����*��c��ql�`� �d�gɇL�	�7��@U���C��ByC�ʲG�+Щ��f�Ys���a���^"��~�{) ���̙���A`�n*��>?֍�|G���r�f	;-�ʿbc��\���s�k�T-f��^%��ZA;?�O�:\QHQ�
?��X�GR�p�_��{̵� S���^�޻�#a}La="�"��td���(�|Z�4��4�>�4����į�OO�@3cC��@��B��ի��V��V�1G�zx�q�����ʋ������Q?�8���As8n��0_l�	-�����Y��I!Gd@�g/)j|�pv����Q�����I������f�,��)� ���cuF:qTB���Q'�G�_��4���X������:�w�.kl��_Z��*�0��J�1��d=�Mӱ�>>�_��Bu�V�Dl%�|9���s]J~�X��X�5w�y�~�|kw�����J���ȵWǖu�� �� �Bn�4�M� W#�Z��	�<�K7���B3���e�����W��N��i��_5W�vU-�P��91�e�2��
���_�zkLL�q5�@���=b�Z�~ސ�مB�#�n����V�*��վK3`L�a�f����w�]���q�Akߡ>�X��s�v m:���ß��O��g�Y��*�+�≺�1Kd�]�QC:�'R����f�c	�$�'�&& !�k�gٷVF(X��}��Z`b�$r'��"�`'�G1B���_�;/�\t�]R�҇�1�ۉR����)2�ű]�j�� ��~11�mc޳ǿ�z���!�|��Y��@ �IE���|��D�لPoF ��#J��ڷ%���Z]U�b�(�r��q�"�ܡ�����;���1*u��(=`-�ŝq~V����p��9k���6�h۵�%t���԰�6걣5;�.;��f8|X�:S^q�<M� ڥd��I�v��?4 B��N#������k`R̅����
,��
8���mA521�\>���8
��g_R�#��~'/�Dq�.� fsߛ�3lE�u��]��l�!�g!�s{E �P���6p��_��^ݶ��;�002��� a�^�����gm��hU9�B��ZL&�o�y�(��9�0�&��B�	����@f�}��>n�|�HY��1344����6�뙘L��J��׀G�pv+�8��B�e "�=���D��LOG���4o�'��ʔ�1���Y�7���]��/��u���!�
��ak�.D睄��H���է�iJ9�w``j*B�~'h���-�]9>H���@r�M���m�wb���^�H��E*ʢu�Tk��S%6�}Ro��V�����&�q���^�ź`�s��G%M�!�sS���3���!c'9��3����հ������s\��E�qvj[<]st(�'ƌ�%�t�;�}=�R�M��@&�)�~���
oB��&<]@�s�$y�Ш��ȫ�1ߏ�~nA����"�}b��	���@�h�M�Ǒ�p(��Kx��r���>�	�}�6{{]�
ȍ{��/]����rlL�+�O�i�%�;����́vLQ����}��g�&����X�cst�_:)�	�k�����"	.��4g/�ـPQ�C���c��L��	����E]
���:�BZ�:��4SV�?���� ����ݶ���?�ڽ�`~�PL� vw~�T�Q���}�.�T&$W��d����!r�M��L�8R�;�}
9�"��^GL�
�c8x�8q��'{(J��c�ǿ����t wQ��ؓ}@76�2��$:���6��:󐠕������������' ሌک�#'�j&ˇw�&��
��DI���tU��b|�ƃm] �Rbb":v��,�-� 9)�)��B�0�$3I���X�D�����X6NH;T%��<�p���L��\�q�H��k@�*Q�y7��1>���.��V�>,*������X�Ȉd�:��t�±�iI�:p>2z�'��R�/T7���+**P���rD����b̘W����Q01�O*	寈ZO#E�A_(!5.�<�#W�$��P9��,�B��\��qz6������J�D` 8�Չ�"Hc��QLa��)���٤���]3��q��l��Ѝ���v~&��D����� yƋ&�[��&]cw�مu ͏������A�����)S^�kH�N�V�2����N~3��'��4����s>m����@�T/���X�Q���A�l� ���zԑ�#�	Z�tEs�"a��#_����jdo���fR�k>b���r���e��;�a�Z$����"$.�L�Âˡ�����)�&_9���7r}c/��Z���ZT�q'qP����K�~���C�B�B	�D��=��f}G���k4���a|N?8���EL�۱!��	� �^�:\u�Xt�h�4�B�`iA6�{������u����E��$%�W
��z=|rFJ�Wf��$��Úh�!Y!�^��`�W�f|r[�#`���YH��=��=�����?~:%n�v7�y����C��=���ah�u�L�X�R渉��x�Rpl��	�����Ly�z�4���Y����Вq�\�[�a3�>K�D��v���~\�GJս��ŭ���&&�������Ɨd�],���2�kV`�:_f�e����+���va|�����i�0MZP�/boF�:��]K��8�^u.{4���r�VC�m�¿��g	`�/��1,MjW.���Yxn�5���8n��Z���z^�aY;�?�N�$��,��}�c���N��u��F�?>�ݺ\�b��m���(&1�I�����`�Yx@CJ�[-�yX3:�6fcu��O���ʠ��C�T���,,g�;	n:���;������ ��ȯ@Cf��O�YU>�=�?�+u�W�G�<��.ܦh����89����2��=<�.`����*Vf���YKU�R{2���Ͻb�F��$X�3H��,}
F��>\${�.Ώ���r=�GB��^Nn*w���k�8���)�����[�?��~��t����D8Dũ:��bR)�g�<�v����7ć&$��ߘC�K٪�kBɘyJQA�����ZM��q�|\�|�]����,�����wzRA��-.><�ҴՇ�������(�)#nc����Bt�]��~���A�3���9;����'J���5��ݦ�vrk����n����m(�����<��}���é�v'��}z��p��LՅ�-[��䵤�<��^�cM�@[rbF7��>�M�i?�����DK�	��AH��'s�O���ѕe����1�4�'Wv�y��8��{wY���	aP��ܜ��U	���PvJ<>}� ����X�BJ�������)��9�W�='j��X��⯹|(n���/d=����F�!��sk̳p������Yhibx��~�-K�Oe��T!�HX�]������r�Z�Mc�Q7x[(?xl{pP��zi��Q��	�ߏ��b>;�o�y�U��+�a�`����k|ة�c��,~�o�YWO�|<�r4����l��z��3ت/���WR�2I�.Is�Ź�r�����"P��c���<C���ǿ��f�qL����,�`=���7�GaC�
;�W�K<l��a�f8v�@�s����FK�i�ˏ��D�v8?�۞t}C�9�%�E����B��cZ[�/�R�c�=
K��$�P�"��j��ڍ��"k�K29��ZE�EJ�v	);e�v�<a+�e2�	�s�P��Le�7@����z�SY���m�9Z�QV�8�޻r�y���S/��`X}$�8��u�:p�RA�ޑ\��#̞����Y|VV<X���g����h^�iT��&��{0��r�sS�5Z��Uڢ�T��0R�I�bGv�-��ߡE����:�zat6ّ-:g�?����	�qU�̗��),L����F�����$c�.>�xs���qL�|5vE�������|~һEto�l�3�4��Xy�l���U����H�-����O۱3��g��5���}�>f"��O\��� >��qЗ��!���j?�k̶jU�_�yX�k�7�������Bs��5J9G��vJE�����M�L��TQ҂���Bڷ��#&DmS�H�$mڞ�=ifr��~���]���u�:��?�{�_���T˵i��p�^^�~q�A���t�����C�M���*n������2�u�_@w?�oT�.��.�O�����tcB�8UP����=:��w�#~ ��
.��w&N��� Řx6�f������j�5?(��X�"�hd���#�	�pC�NiO�}�3&�Zy����9����;���2+��/��P�AJ�����̐��^��*��.;a�����vt,.:�t՟XVA��1�ߍ_���&~䊁-n�@�(oM<}��"Gבa�Q��Cda�O��G��0�f»�����m2�<����~v&�ڤW�F�C��&*��X,�ފi�$��X扑H���_�U���Y���P
{�QFV�) ����O�K'����.�m����84�E �!ov�2;�
'��|�B��*�z	��="�0k��b�Yn��r�����R��U�n��4�����gR�'p�
6�����>�Rڠ�|��j���{.ȹ��,��y��^��ڽR�6թ��C��pdQ~	Ne�[L�Ŭ�W����fJ�H�>#(���ޙ���6t6�nz�|Э��л]���kkk��$�^^�"Vt��^�=���~���@(((�'T<{{l6`9����08� �\`R �555�C����6]���L���њ_��D�+���&�D� ��j֣̏�-@�ȇ�'��|AU�� ~l�5Z'x��nJ��^��3b��썊e�}��q�<�T��r�@=:{����U��d����+��W��G�Ӏ�ҔWR:j��E f��TI+d�9�y�t���� ��"V&$1�>��^�R�q���H=�A��aj�iǬ+(�N�@is����Io��$��1�<'���]"�.Q��JeE��u]VH�l��.E/�N�5魵�]��#�{V��%D�?��*ʘ.�E�����OG<�Y5�EC����5����_{�Ne�D7��Y�M{q֜ʮ�*�%@��S����9@����;u�/�_]�����12@��2��rJ���]�c����v�/zIb��C��. �v2d���=D�E���U����qį�������M*k����Q�X��w��{|���7�DN��}nLռB^�5v=8T&(ʁm��qВo�X
[������7��ؖ��B��:�#���~0�l��D�g�;��H:o���������*�G�Y��V'o��L�=wn�v=�J���^�TjA���Jj���I.�H2��j��I��Y,g��CfR��$��:���mm�5�$��{�2��g�.6���=��,���J~�k�H�������X�n0�
%����/����Ί���$�X��a`q(����ΟU�`[����`݌:by^��+������R�o`/(�3+>a��C�m��ݵ����:%%�(,��SCF&�P��7��֯(��[�X�����+?����ß�C�Ę�eT ��5�Q��1/��'[���r�x�����w�)Dg�;V�
���7�v�Ã�%ɔFk�+�7�lA�z�NW���3WA���oe�ȿ��=��5B��n�n����)�o����t)��jz�[�7�7�ue%5 ���U�dP�MR������]p���җ���Y�O�x�j����|X����zU e�`FA,�7YYY�K��R͙�VB?O�x�aӁ�����V6�~҉�n�f�Of��������Q�{��g=�5.���`OU��p�|���Um
Ś"B�Xu�����wN���=C\�(�kv�B!�U��5���glG+�����`������Ip+ ������H����S�2h�l�F(���WB��K����B����ڋjD�#w���ځCZk#���O�bh���-N����0�����ߴB@�w�"v0�y;쨄��$�g-=��3�F�iJ�C� n?}%=���U���h<�հ�y���%B��l��&�lߛ���bTm��w���z2���z��Do��<R�~t�9����QİO)'j�x�m���^���/��UCsT7� ��9WU^^��**�h5}j�O�Z����d��В�+8���_�ͻ�)�� ;_�݁q"�90sڦ�vh>z��L�}���	�����!��]�螛/�l�o�Onpf�	E�&�M��G��wx�>M�g�4���6�`5G�Z}��}� �|�~e�f�e�XJ�6VY5���[��F��c�����7%*,�!����S'�P�i5˚�N��`��!����6��܄ ͆6@(uڏN,m��\������[���T�V�d��G��ۛ1v�t�2G�������˻B�t��6�^�����6�R7�@s\#�d�~�i44�˼�WGz�N�@W0������,�N���q�.����+"��+YI�tj[.duS��'����Y��󜀆	� ���&g�:��8t}0�v����2��4����
�a^q/`KϪ~�_��!}0�}��D�,\��WPncS
�k$q�Y��O��>r6���>����I��Y�l�PpN��(��'Y�����b:g�M!�G���@�6:g%	잵����z����T# ����J�R7�H�le��xi������ڊ�oF�����R �����G������"ۋ�iG@#o"���M�?�r/d�H�l��^�E�ǖ����2v;d��*~����w� .���)�ž�/�Vv��G���I	<�	��\
���u2��R��&w�3�%������ʑ��e`.[�kې>Lx			�)�Ucr�|5����ׯ0����(�O�~����*((���?c��R�l�t ���(%"�uݞH�1�i23,kO���U;g�	�u'\	@��g��	aF�ml������z7��GR�$���h���I����V*Wx8��)h&0
{d~4��3����,�>%<�!�v�.V���ե���q��hJ�lq�����	������ ¡F�Sƍ�6�b^��� 6�-`��a�����{�t\��`�#{js��}N o�H�;0���Q���������ޤ�m@��<�����<�5�KV��;0f��-8|D��b�ȥ1v{UF�ɞjP"�'�J��'�h@.�߭͂���R3�w�4;��Ƈ+���:7-���E=��W�U3Q����0���Ȏ��3���p:c[Kt|��]�O`�$ �\��Y��F�ظ��������ZsR�X����q�َ7ÿ.�5 ?{�%o�������$Ad���|u�7qe�TS����W����m�G�Ij;̟��j|+��L���������B�z�J-V�/�l܃R��$���b_���@��5��Yw��h���A��,�́��g�M蛔1�/z�.�|d�� 8x8��PVjv[�hK��_��[o��	�5Q�h����t�M.��|���\ԇ��]\��Z�ڈf71�����WPe�7XV
��Dύ��@�%��� c��.&��mf�$�E@�Y�l�K�`v�US�_j̈�c�eeBCT6 �e�=e�y�ǳj@Xhq�n�E�	)�%�]\��8}������d.��{��Ũt�m�g՟e��>w��4sՓ��4ܜmY{�rJ؍��~�`^��ڏ�����Q	
J�飍�	��r�q�]W�ێF)����Hyp�8�
z�.���A'�����x���}���QYv؍7�C 
�u��Xe�\��W����m��BS#��#f�+`�H��ʈ�l�VN�$���  ���p�Hdap�Xv[���ļ����iH/�/��Z���b��@o�f$0�Z�Q� ?�s����x� s�)�JR�f�� ��az��l| �n7��Sξ�=����F��1�m��:�x:/p硁��� �:�R �5$N�D����Q�pyR��9fIyF�)�N����O
����)'�K!J�?��/�u�(+�I�^����d'j.| ��M'Ń����'�b�wΗB�����RT׋��lI�+��k2<u�ǟ��W�B'GNOR'�^P������x��J����&a��x:�e���7N��ƯD�E��Ԉ�2 ��U��Y��J�����'ߌҏ�Xs}s�T��D�~�Ie-��屒`M���m������X�U�qc�es�w�'���/��AZ�Ix�<I�P0��<�bp������k:2�b{��YM��嬆9E5R�x���l�)ڱm��|������&�b��hO�P|#�B�>�#	:9�D�������C?���p���6�l��¿��v��Z�J�/~2�e%!cn&V���7t�9x����g�6���gD�*r���;g!
"$=�%Z��^�4�
t�DMvn�(��:�!�B�d�=��<筤�v�Cm]�;��[.w�FUwxf82>�t�Eԕv�3���QwO�R��������"�W��v���Xx�.��D���]�rRP�W���aр��h�i�RuV�+�gl(Vƪ��a��(`�t�������R�t,���9� LW*u�{�S#"N�lǊ�{Q(
�
� /��_��	��݋�K�<�P���/1�
�߲���օ\���=&�<]94�,Q��w�+"�KI���������-`Z�1�&|������/���+(B[\4�*��|��t��K@tm��D�T-���D_�JS"���yyy�<:1q}�[�����=)yE%�C#��ץ���D(Ɛ6G�*��NP�kM�>��/���&�^�:��?<�3z����`���/��w�^�z�2xz����f����65�|0��[�[��뎩��TY����9�%����R���f����;��@��>��#-D]���D<��{fpn��4�>��{q�N��gL �WBWh�����̙�-�=BҁQ$u��мl�mH�5���:�a�^^�_l�Y�r@Y3*����O��v�ܺ��U$G��E�	 H��ea
����W��R�/��Z�/�� �4%�H$P��O>=�)�ጎ��?�4 r�,<��/������5]jE���yDȗ����:v�D~�җ �&�lOwƚ�b��7C���8�v3kO���ҕ��l�#!�.�Cy=��0��͐�@(#��ۡ�Xr(4�}�� ����H���{�Vы��r8�A��H�㤨��;���C/$���<]��i�?�T���{�o�OM�\���򆸶������[�1������$�[�tn��/���_�Y�9���.q�Z�/�C���|����B�8�E5��j�=4���y[����8X��<ܥf��zm���ê��ǚJ=s��x:vO�?��&�IW�,�� {$�r�I�YΡL�_<��wLϊ��T�D,V���[.߰s���R�H}0�]��&�_�0���׶�9혙�x�U/�N"�C��hXn�y�R'jz�z�r)]��y�E�#dF�^���%�EƣWNO�?�ɬ*�z�xu �_������
��
��ᑈ�~B��4:�hnH�Ke�Q�G��IZ�B����}�ml�"��.����'E޳�)Goa��������[=����������I2�j��\);A�Y_4}�Fw��{OJ2
���V���5����M���u�K�$\�p�.&�$3Õ:��֕��\et�/�U�9�h���G�e�p�5�>��;�ݡ��%�)i5��˺�>�lue]�PhA�PǮ��9�`K2,���O"CX�27q�u���޺��\T@�>mt����AX��1~�۵S����%X*4kD'���<���Ћ����ަ&���E�N����M��ރ��y�N<Vz�a�����6&V��X|�|�n2��e>�60g~���?�)#���U?��~���cV��N�`�tR~z;�WF����-"�4�h�3I~4�;M��9b��D��&ωΖU���d�.�}Ɔ�j��AJ��薙h~Ibe��lJ;�fm������m����.BU0���p�3O ҈(�2�o���ډ��4eE�
7qe��s��ȉ�I�_��Ѩg��fo�e���m���9!��o��z��j�ȕ�dm�񯢆����˦�E7�f3� -��<�N�8��`B<�=>�4�g��e�;��Qb�%P�&��b#Lp�������D�~�.C㶡w�&�c��v����y>݋z=��HZ�&U�,l���آ9lIuM�۠�ARh^E� q'3��S����� w"� }��j��ԙ&�ئ
���hl�gi�)�V�39���	�o�� ���O�֑&�����������м��s(�5iw���^c�A�W��:344$�NL=p�[������)���wށ?��.D�%�q,!�Cw�4%6�h��`~0;�>�z1���9�`�bcY�nN� ��BJ�d���:J��b�K�A��h+Ml��� � ���R��?jl�Ԃ:FDٌz�t����Z��C�wc�V�o���fݪ����H�Gyn�[��궜m)�W�h�*L�v��?���=)=y��;��Ť�O��v���x0wͽ��0�(���՝F��0�=��'�p{����^1�[�$/"����6bKr�_��j�{u��7�$oI~���1�VD��Z����^���� ���{�m�(9,�*�C(Y�Q%�~�����^�嚠�z�!==�
/��dN<��4�"�@�6���UV���%������4�Y�vh��l��[L�\
ܣQ�#Hr�t��5'ূ~��_t��=�^�����gA���2��=:��K^o��#""�Ȅ�#{��Ouz�>�3�7�R��������-& ���5�ah����[���Q��}��3k���VN�$���J`$�Ff��k���s��������1WMU/�͑G(I.-/7�lrzm̺�{�>�
ɻ]ٺ �������� �^֣g���A`�BC�}�=� �\����ӟNs�c��%z�tz�3_��z�͐��N�V�8Xu��Y:55U���N?_UL'%�C\3��,�7�%�[畭	1c����yu�B�<b��%�7y�� ��@��2ŝ	fzy�2p��dz����jZ'c��݉��~��I�)�9��i����8"-s���U�Tg��ɥmmN�ɂ��Uu7�]��.��V��A��!��32-��>���U|��{���$q�'UЋ9	�G����*� s�WQڛؒ���Xد��W;g��
>��*Vl�C.{�ViO���Vl-V/	�Hr�Fq����Xr�ׯReͮBbW<z�v�|��-�J$�N���h�&ݩ:1�,@���T��{��ࢌE����Q/�* $�dGj�%s�M�ٌ>Pswm�����ƎJ�������Yп��J�SA+I�ΦNk�'}��&��u�������{�������{-�.��?�����!v/#��m��b9B�q����g:C>�@ҷ���\7��(�i<�ҵ�w� W=���?�Ϊ��w�dP��ޤ��X%��C_�ښ��` �?�*l�!�sPrVNT�?�ٝ3k�|���U3�߅��'xN{���ZTlmЄT%�Vt'��$�I_�Z�@ݴ���yyu̚G������2â̶�b���s#o5X�c���J.�4Cn`OB%Z��A(�1�<<��]��'��bj6S���=\�L��*)��;�$��o+���y�;�� �r�C�BrG�����x|�/�}��L�X$]�:�o�ӯ�
!O�K�vt���G/UHE�'w�2�k��W}�p��T�# s��(W�V��U��<^�)��ʡQ�9����^���)���[=+vZ�-9��������W�ȕy��i��?��ρ��'g��	!�?����]Z�'�U�9�!�EZd���݆�M���g��wr�85`b�����2�
������?�:��>yUe�	EI%X�ԉs�U�۵&�e[r��k� ����	u�/A
��$�|a]|zC�NX4��ch��9әQ��@7��%.�XP���"Ta$�d����|R��E�����$�^A��I��� 䟡w
U���K���YX�?�؅0�v�H��F��Bs�J+nd�[Dj�����maKz�엯�ʩ|�f�aWj. rlq����/f�� �@����1�y��!`� �P�Lnp4�PU�8���h{���������/��q�%��@K�:�"���+���Krvv^�c���:��?���[0k	���)�s�N���z3c =(v4�J�)����UV�v������qK�@�KݲN�- ��jW��ݮҎ�P@|�2{}�ݱ9��]�8!�t��^[��|��4�a�Uh ���p�@V�p�@����R7^*�>���et[�N�M���7��VyӺ�AbP�UK�(3+�7#á�_��A��p4f�6*Dq�U���	>IE��M<]S��F3�M��\��-I����bl'���X]"bN'	���e��i�\��%���F5�o8/H��]����b��Jo�ڹ��%��Gqjj��_�n�K95��oc��(�8^����i�J�����oN끯Ӊ�a�@ݹ�U�]�[u;�P�|ٍ��[�)�k(�]�0#P�+�? ����Le�h�׃�>.�6�nR�dm+'�
r�΄r�O�:�[��h��l�+~g3_�J~H8z�d�$�!����|���'yl���^�O�D��u�]�Þ]_�?�-����+� ����; � `��@���(p wS��~rm��V�[U�_�;[�D�+T-�K�������k~vO�O�;�z����^�k/��O]�+����G��{n��V)w�y�zX�J����羆~���);��<BY;'��#�9[����8Ղ�3���~��֪�=�=zCqB�>xlg�36�"�|>	��c�9�W*=�зf����7T���1�JZe��PҖQUnl)d��F�>5ơ��"��4�s����Y����]�Y����;F�e���
�ͬ���5�K���⡊S�Px��ʺ�(�u�������}q����(s�h8������c|K��w��hFՑ�n�`�������	Ӆ4���X�a�Ks׼l
��w@���׾c�]�Xc���z����8�����b�= ���ƾ��)c^)J����ƞr�ǎͳ#������A�q3�t�?`Oo��HoQ�h�U[ܨ����l�失@b�3ȭ��2�"�m:3�3�+&}����LO��3~��'�z���M'�z�L��9%rJ��)�S"�DN�����ώ��{���i��?�[�=�p<P��-a�M����ފ��i���a8��7��ڏ�Sǥ���2S�N	�8%pJ���)��������ĳ ��(,��]�b���P%�.���L�S�tG�.�ivד����>��+��s�6b}�r�=�F��e�x��[Ϭ�Hk9=��fr�v�p�r��
��~�1�՟�6t���>����4�vz��VV��=�'�����?��1�8��8�U����{a���v!������@����S�N	�8%pJ��K��6����*�/z�t�I��'�6��͚����ٵ���-5��̪��>X��k�M:/�<��?��&�Τ�2���T��X�����Y�x��ϐf����?\ztm����ճ�����aե�츅nK�����6)�[�j�a]�NM2+�~��.��t�ҩK�.�|�/��zw����27fܯr"օ����ݹb�}�_ƻc��ܧ�ݘ\�J���Ѝ9����c�+FMP�*�Q;��zm�e8�м8�q6��[�ǏuD+����x��rb�C��_��\���.���:0��2�[+M'�����x\��*+u�d�K9AͰ�%�S�6�BӉ1�^|��t�_D��-A��.3��>�х���H����(r����A
�ھ��;P�$��
$&�Wl��u�x��v�K���U0@oF+�����F%5J��u@��zQ��^ZK�e����X�;�������/����0s�⊬�}�E�Kdy�1�f��yi�>��fD�pp�4O�g�;��K��k����36'pj���`�z�Vr��׭��70��*���y�%gS�T�J��+�������D�gވ������s�<\�;�؏a���̶d�W�Y��f�n�~��ھcG��\\��'�Q�G"M������5�c����.[�#��k*����5o�~�'�����.�J��Ʋ��Rܔ(�ԔL�Ũ[4qݣ���K�)�3�\�M�{@m#3ch����}E�aI����ո�m�AM>���]r~�ڒ�,k���?�B�������=����U�Ĵ�?~Íكs�7�6G]U�u��s��ctxБk�����^��0���'O�H�0ҡ�@),��c{R/���o�ew�2��bi�wە��w&����"���޽��X֜3�΃b����Y��7.y kr�h0�o��KB�*�X���}�����>>�\�-�X�O[nTl�hL��[��:�/F�������;����ح3-33ӅL�9G�K���E�]*�B.\Cww�� �����0��n\�OG>�Y5^.�C�>}2����,�j��h[����)5%��M�#:�o�ᦩuΔxw�4]��w��;�,B5�y��<-#1q�N��˵Pτ��������ˑ�m��LB\�g�ܫ�"�CȬC_z}�v��Ms�*�ڡe�j[Jb����)
jrb�r#ch:p]4�=H�M�?;���x��pM;��a�h����w�b�����VtrrZ���B�y�߅�� �n7���~����g�_��}��琹9��ɡy;C�n���s�0sX��7̨����X��u3iއy+\8�,���r�a�#�C�?�$�S�Z�<�m�迌X�ʸ�"�6��y���U��v���+�-%~���(��ݘI�_N7w{�eg��K�6�ſ^���Wj���v��:�{��3�Նe���D�e,�t
(HL�7*�U<���J�h+~�3gΘ�������+�Џ[�5��7n��1�E?J�8�vx\��#�ؚ�$�Q6.Y��<��ْ�7OJԊ�/���R���|��@�P�����MݔU��]�A����JnѲ�+Z�%cԵ�M7h^�~��j�3 �4��ڐR�^HMkpZ�K�2_�y�f�"�����qI�	l���O��ŋ8&�Aʱ������{N�5���^#㺻i{;�7P�7̰_s���|<GO�2.1G�$��8�	���`u����z/�kxK��6�m��X>�pU]F"��Y��T��r����]������ʃ���2+��HC/�U�Չaz+�h�~�0�A��ޡ'��݆�J�wgs0l�ވغ��i���I��,����9:%p��BP�W|k�e+q�����B�tJ��q��h̖�����}q�0�n�䣧2`�ZKK�����r!A1z��DwEEEY���Q�Kl�Ce�ĹBv�㒡��8�p�aɿׯ_?��X�]�x;�m�Q�~	W��(r�G^]��=e���3*^��!x�'s0Tb����wu��ܘY[J���
U����jE�k�
�Ҹ��Dw4ѭ�ի8Ð������<����u�z+����0���e����Ú�=f��7TN���۷o�o/ũ�������t_H���AEh䍝����LBŖ2��P�Ӳ�:��f��fB�?�n�π&��Ӹ�>ڑ�Lj�_2�f���յ[@�}Ԍ���������J+���Rc�:z�(%�].^�RS����6|�y�MM͹/P6׉1:Q��ݚ��
y����i R㙆`er��:�4Hǝ^���4%ό��Q˻'�8�~J�1��[�-��3����d�t�4�gG�����Q�Q�����b�Jqts�,V�mԑ�ZR�?�y�ƍ� ��'�_$��d�ÒtUI��J<��v��p�g|@儡��R�1�{x��;?��bھ�H��w#G����ȶ4�6P�(���=�BR���O�<�su ���?��k��\}�����nW�����\�s5f��9�?@rv 9&߆F��K�Τ��m2,At�ݱ�����0)x�����_΍���u�B�^�kxNh�(�K����	��؞M�0�dpspf�(�oeŝ�/��uu}A=��K���
l��%[�UѼ����!�7�]���ux�n��&�H���T���BiW�.]��%W�j�A��D 6�s�ZF� X�W4#R���,��4,ﭽ�@i�cE}����Z��v�R�?����T1fP���ץ�D�<\�E�#tb����T�m��H�26L"Ib�G��wʅ�	��0j�;���>b���0��67fm�J�R7C?E���ز����jg��%un�G研�E�i��}�1�f�=��~6L�)�L��`6���d=��
՘$f����<�s�X
,�հ�8'�MA�R��#��'�ݒG5
�:�VH��ufff]hΆ���A)Af��!!!f6a&e��q1��#�V�H^�ѧ��5���ѓ��HZ�h�f�=���o�u�50I(���� �T:i����������P���a����W�j-	q�Q�;��
epN��uu�Y�&�ʍ�*���o���7�=�Ѵ��K����gϞUC;'ϵ�6��1�L���W�5M�<�N,K+��4�uӨd�z���9�&f��w�������&G��5w|��d H��"�����ٱk��Nb�n�aă��C�}��x����q3?##��B���p�۾��_B�U��tX[֪��+:o����a��ߠ���&��0''�O�S�!#�]�����*��ђ o�VO���K2pV���g��9�@t�wU��o:���2��2.i�]�]�ɝ9�������%�g��Ԫ)�~�����TK��z�������q? ����& E��M�wm�i�6+j��C��=�c������0�dY�"E���|��*��Pc���$��_�|1y��]{65� �K=�����3/n-�~u"p�h^F%���f]�3KB:u|�}�͈q�0����ܔ���V1�J.��P����h�ܺN;H%���VV`ڸ@��8HZ���"K�w�e��I{t&���.wMwF�t߆YԄ�
8�;b��%CAō�_rG�A�V���UV��=C��[�i��TT�ɰ�35N���<#�<�
{�W3*�@��OHi+��H���?I~�,.�a��i<�z�L,�d'�=j�ɇqT�ލ�D�)i����?�����J��`&V�:�^ b�m���ȉa+a����W��������O����y8�@��)��Z�[B��:Բ���e�+��
��� ����Bڗ�Hg�zt�@��fȁ-�K�C��ND�~�z���Z[�� ��Z���[�X���QZ瑧���:I���	�'�׷�ZA�Ǿ �5Vj҆�"��;�( I��?|�P���˥���p�@"W/���!A����E0��O<���#Z�t_۽��ɻ{�n��Q�!�eeC6��w����։���3m%0c2� |���
�02�� �#�h�%Ǐ�Nl�1���g:E5Y�@�t�KD����8��(�8��\���R���I�؅�vvE�td�rjCi*`��I��6PN4�s��w��t��XH*�g��$:���v�6��do��+v�J����F�s�/������& @y�� �����`O�����-�pďӏ�5���1S0��YC����4FP๏_�4���o��t��=����A���Pʇ�����;&�bb��n.�!��Dz�3o���}9ޚjtR��U]]�c���E�M����$ɐ�����ܼ��!d�/Ȥ�A��i8��˱����,�2��b��,L�b���Ө���F�ďt?y�dl5�͎ʮ���f��f��;v�������TU
@�veȋM�!�ե�;�\`w���x��~���j�%�ﻙ��P��xk��&��rAx*��5Ji:�FK3G]�`��� �Z�r-��M�`��%��``\&K��,N��n\«�):�������AV��b1F�����Kp]L�A(,��c<64�8l�&7PNՎ�Z�susph�c�jFA�LNM�['+���H�mX]'��ytEb�\�E��aJ��f�<��E]��*W�>h���� 8`��^?�@����Q��x䤂�Nf���\���<r�6��LA-x���5����2��nk�2O�ju�ߎoy�;�&���h�#7'�Y�
�nTX�1� ��zzz�i*x�$�S����KBJJ�:�UC�D�#�q	�����N���v�P���ǎ}����E� x��O��q`:־��9܀�N�i���熔5?njjB�S�DCm�W�{]��j�����J��ի���@�g��ǥ-I{���F��!P�?��4h�V��^0��0*�~�ֿ_�������qK �ۗ/Ź��:p�qO���+0F���D�|�k��b<�pUM��5���׽�V�H��c����?N�2_!����b���He�z@]��嚪�������{�����Z����+�s��hm��(1��'�T޼Z�z��L��U�'N�;>^�u�8;;��:E�ϜRo��[����,���0$��q,���=��Ī�:3�h�6��Ԅ#��)������0����7̈Y[Jz��òvh�A��4,����E}89v�qΦ����,���?-I�ˎ�^bTr���H�h��1��h��Y�&���P��K߿߃��Y-}��cJl�p��Hab*��~>�dEwm���O��@A��
Qlr p�BaK#����_#��+Ȇ��.--uA�Q���w&nC�����;!ò�.VR����@(������"x+xB���,����.�ƛ�'��߿�`��f##%B�i>�����G\�_����?���[�tZ۰���S�g^�;������O�EB<WKg?�<)�Z��z[LLL� v�4pjP���s�ghjjR6����FN�w�Q��G������}����G�T���'���It�,����0Y 0c����
�u����L�Z:>���p�+)�K�g^��X�>o�[]vKqA�Mr8s�#)!�o�ܘe�1LK�Ry7��R?ѿ�:�=����V��9?O�XMx�~�ʇ��9�=/q�h��(���z�}xxX	�PP��*7���G�X�5��|ƈ=��X���	fL��-�0f
�GNd��=\WWs���Doәx�e��9Y|%�c���h�~��ёQѴZ��?�(�jq�\J2���~� y�o]mV� �%T��%7 ~}���|�d����3�c�A���I��J"��=*?�H��+6}|��Xzz:y��_ Di;����*�4��_�6֙!�=�I�d�����mt�w���˝^-g�_{B��٭�@��������!���։aZq0K0ַ�Q��r��I'M�c���G�n��0��-����PTX���.�1,��]��N�ÿJrM��U���af?t��\���t����Ļ�=��������.�?��ᱎ�ߝk��a��μ�3V�D���<k��{��zO��d_H�s5�w<�7%pJ���)�S�N	�8%pJ���)�S��(0]Gg3�M�g��[;%pJ��3��n�C�&�_��cK�F�ڂNe�]e]�&�@Jڳ�:Ч!��? p�ה����R�t�Gԫ�!S\�w\J$9�LSŁ%�9j�b�����ō�OK��d0�V��g�N�<n�;{������X��!K0��b1�q03�!�)z� jjo[�5��?"X����w<�{�1�Ǐ�A����a��ޠc�����M�;��#�-�T���[�j"+�aU����P����!�ٻ����[�� ��+�ؖ�cX��cy�r�����W�;�M��ٯ](�^�)
\���0lQ�-�O���@;���=����qqqh����'�a���,޺�\��X�Ӳ���:M����W�L�~�ֿE��X��zRli�0�����O��gci��vQu��h��̉���i�m[v��a�PK   ���Xg�	�;  �;  /   images/fb3f2d9c-813f-448c-93d4-6d887e4d49e7.png�;"ĉPNG

   IHDR   f   �   ,M�{   	pHYs  �  ��+  ;�IDATx��}	���U޹����{�tO�>�F���%y`�8���U�@0UvA�	��(*�J��P)�
��TŐ ���M��$[��K�/=3���������ޜs��_���5�=Ӳ4}GO����������ׅ��9����9��A����v� tSݕ���!F�o(�h�8��(U��VO�z���G>����ru[�Vl�Z�|�pB�:�zK~.7���|b�op�\�n��}�n_5�M��t���XT'�֗��������j/���XZ��UY��͞D��(i��f+�C_ű@��@����Yw�\�b�W� ����R����ᯝ��v��Y���/��h��f��RR�8����S��pOuf�=aeiOZ+#W,���f^�0�Ab� B#=%��(Q��W-h�g
dT�F5��:���|�����g���=�=8:�ߵg~�Ï��u?p���ꟙ>����n[����������hR�� �s�>NpA(p]	AP@<"�"#.Ci���F� ���#E*��T� k��m�gv�܁P���K3��ї������>�_N��8�z��0�ܡ�ą�����Ͽf��;[so���N�Q'��\���x.��@R ��	H0���.�I`bI���F� ���H�$I �|�-*�+"�v���j'^<pl�����v����ϼ��=�z��a.<����yꮋ�N�b�����܈֋EB�# �{�a���7�HH$��N(� �-q�@�X������0<6F�A̓��<?Cj��T�Lu��N�w.//l�T�h.������/�y��C����f���JR�SO|z������O��jTz�ro.jB/rF	��D$�4�����[�$k�%8���$,�x(��H� ��s��'�C$�_�������{x6R��>�4��Ps���م�۪s�w���/�����͚�׍0��Q���z����G���pT/����/8	t��9�C��cT�(�H��W���<�	 ��gp��!��Lx>��N6��u�	�bO�ALP���!q鈞�L�jI��6}z������G���߻k⾏�q|���u!���_�{<p��'?]8�`W\&n����$�����
��p\&�t�Dс'�a$&��qʉ[�tq�`U���!�bb(y4�m��D�k�,�H�U/@ei�R^�q�]��/>�ѓx��r�6�0g��Sç���{f��h}���u���M!�\���H��ǟ27�\�P��M�F�0K��0Bj;�4��	�ӌ	�q�
�X���)Ii�;x|����ŠB�Pm��&��=R�o����6��.��|�?x��?��5Cm�J��o���o�&���/���]��
��"�'�E�k�=��y@���.1�		 鐎�ߤU�Ff��W,�H�1����?����A�&�;șD8:׀	� 	~�uKw����*���B���������L�Z�զf����<���>|�g�E�8yk�
�@��"Ί����	e>N�`�Wx�Kڢ���L�A=㢾p"0gi�C6� ҈2�-��4s���H�����xd�xL\d)�7�72Rk��ʝ�'~t�U�]8������O��|n�j�צ����>����:q�#�:Ӑ�B)�� ����<g�x��O �IK���PZ��	&V����Oe�@zE�"��Q��sF��$�n�M���t.�_�r`��B@Dt�y����ʃq=X�|�?�+����_����5'L��W��~�[?q?ܚ>w�0e @k��LP�
�r(�"�QXޓ��P��$yB3�L&�FbL0�w�ETtLj9����0 �o�#��G�ȣk���b���hC����M��F�����(N�M�xs�t�S��_���}���kN�������O��X<sp�kAŒ�J���c�����Z2I���~`'�Vp`ŕg�> C�(wc���c�9�!�F�8bπ�~4|��d's��#�[��'~�����=��)^����5S�9=� ���8�+��)���������!4lp\S�L~�<x�[_��x��=EՄDX|p��49)�+�s���l�8l�V�fŧ(��j#�����Bi��
,r3��F�2���M�^d�n�&���1��5X�I�(���;E�NK��	Ҵ{wOij��O��?�4�xa�sw�s�П�}�[_�׍ٙu���I���hl�����]�+��1�65�.mջ5atgW_N1怰�E�Z����hKxm�Y��]4�j�����ip����b4�q�c�V�,|�q�d��?�7�y��~wz#�wM�x���O}��'μ�ֽ@�k�'Y��M�k���!C^im��0 �§!����He�B �!4#��O�
aRm�tr-�:߸u����NVGj5��|-6w��x| U�?76¥����'����?����kB���̜~�C�2�ÃrH�Ns9Y_��9l�3K��.FPU[3��3��E�S[0�`�ȧY��eV}���`��_����5�s�1����lW	퀏��l�G!t�n)iWn��]������>�؋yd]!�N���>���S_���Թ��NQ���i� Z(^��)������
{���	dq���F��9:+��"�[�CL+�` o++&3���,��C�W��5t��H H�ѽ��ҁ�$~K4y��K;^ }v=�xU	C�����;������5�FA	o�gW��<��3�q�Hᬈ0����Hɂb��hW�9�^[�ɒH�>t<r�  ֠�tN����y)���k���t��p���C��w�UZ�wϞz��s��ou߇���Z����\�;�S����R҂B�V}b���D���e&Ա
׈Z�B�$��g�@G�n�CR�O�>�}�p;#���U�"���҂a"��} ��zTjU{�w�w�(\c��aL1�t�赖ʻ���x��a}��S�ᇓ���U#�~�9o�����ɷ��ZŘj�xÞ�K� l3��� �dq�\�r(X�/I9+��g��xU7�����|< @z�m���!f�F?D�$Xm�4�е!
y��p���0Ǧib��ɔ�Ayd�\t������ M��EA��ZKOyߩ{O��%/�.�Y���g�tN��:��9W.�)�	dI^�ƙH�6h�a+ �#AYߕ`ģ��g�n'���:h���'s�k��B�B�O�Nd����H���Р�Z�:,���?e V�ޭ�������$�~�-�`������׏=6#y$�t�4'G/?�@����FQ�!�B(r�;֊w������,iD�(Km\+2S��6ɂ��&>�:�'�[���]����1b��@F�[dŜ��3�˃	c�t�=P�R̝R	cWQt�@M�Ǧ�k���z��{���Sx�ܦF�;�{�;�|kX��n|���A`���p�t2��������b�I���[�aXl�za�G#�1$�h��d�Fksvʈ�6��DΦk|a��+��K�	,j3{�a�$���� |&�w+H���z|�giq��Z����&Luzr�2s��|n���d�B8�F����n�Ҋf+=�fe��ϋ9�����+���Eb�6P�����l��1��8a�3|k��q��v��ݖ0�ڼi@�
̖�2;^���$\rx���~�n�\8���_�뽍+����O�k�*�S7�r]\u�cn>A��\�<�8�VDQtkI~xZ������F�@ibC>+i��X�%D8R�81B�X%��R��N�Xɱ���Ҹ�H�z��j��N���O�̸:�,���ZW����"x!��(Up�&��k�Pr������s��O6�0p��]]�}�U]�I�0��Vw"L<]9d�$k=s���HS�g��L(�X�4$��Ajh#�b$y�(=�4�4�y9o �c�֥z"�(Fs8���x9z	��~S�ӑ8t��7ܱ�9�9����16x\\m� ���(�D��"�єS��k��#x�Ħfn|���44�}�
EN�*M�x�}�U�ae<�:K v00bBJO I6
��d�]Pi+�[l���L��!� }]�q�q5 <'!IXS���0����@���G������;F`�' �/�w��o��hEduҠ`��W�)	��F$3G��g��AqQX�����8u����a����Q�a�����j��n�����H��IGPBE��b��� �u��EE��ǢFWX~�8���0�W�.Ñ3e�]L`��� �?�y
�;5o�?��ta[	/��<�T�W.�g'��N��5i��,(8X��=7��-�]�G��m0y�W@
=s���g�L���Ak���1���r���Dg�B���{��؟���m�NO�����oە��EXߖ���I���q��J��"�21������tC�zA�l��!s�f������46�ϝ[���H\��"�A\�1r�2��9�rszs���7�g�ੳ.��]x|w���P)+8=P����B�+�������p��HM0��{3hRZC�eǀN�����ͪ�<�'�fH`c�����s���z��c�&ޒ�ti	���u�� ���=�N�Z
��	�`�����jp�,���}#���ؽ���s���9x�����&��j����#
��ug �z)�ƅ��1|{��K ��kp��E�d�m�e`�/F��eE�)�1ݱQm^D2bU��8�o'i>jׇgwh}���E�!I#_)��N[�|@V1q�b�9Cz,�س+&���S15�>�Q	���vQ&��!��@i;�p�̓p����ӛ��.���AWC����O��B�yA"0x��}�k�mU��b��N���&�+�� �(Fͬ8C���MPL^b�|�.R�ۥ�Ј�Z��m�%��C�S��M�Ə�o�ӆ�h��v�ܣ����mORN�e%i��J�o%LK��R���A���2�QQmݾ����Qq�$0�,@;N'x�����瑘%߃����E$���nn,�Ѕ7��oė�\����Go3]�\	�4C�W����Y���rvaj��6q��o�8_BzL����7���kJ���8���n�Gq��wv��WA3�c�ghM3�N��cdƈ틂jí#y؇H��8SS�U����&*E���(��g{����n�Q|߅� �j��2"���)`9��@�L@;Xy&X�4� 3xU�a Ftw<�2�%�%�K�x.��$׬���8
�5ƺ	��c��7&�d��S�7o�1&?{�W����Н�G6� �CD�@.�p|%��/jB�^o��ܲ&����\(��|%\��w�ax0�y	��"���+���AE`��Q��//W���l'���G�ۏ��vb0J�>e���/�q���8UJ�E&3����ğ�4NW%]�U�c��漯�c&w�����t�����9Y���X8iNgB�Ih���)6a"*�ʵ�2��p%�KC!!�B�:������Z���=��P���n�ʥ F�Z��(�=X.��p��4�D1��u��h�����d�^2Ѻ���Ў�+���g�D ?��!mk0�z���-;T`i��2���Y�~�^�iX 6Uho�T�����j�+�S���m� 6%�
1$$*y"�˖�b��B#��Ÿƪ	<3>G�C�-l�x�� �C����=d}��� !�;�O����y(@�p���"�$˼��8�V[�rJ��69P30��
ZLj�4)Qʆ
tVnh\M�%����
�F�T�����aùf�q˦Z啊��`�f��J�0O��/��f"�R�g*K׺�����q{�Ԓ�Ó8<т���Q����w�}}�K��8��-|�Dsb>�C�M�����;�m�X
�{�y�x�v�����W�����j{l�
&�ICd��Q��&�ȃ^a��MDR"F�Wd�p����h&4̉[�處!;&����HĈ�U�b�E9�hm����G���3����A��u�(�{pv�ס�넪Q��D���"*�gg���+�0�D)�Sޱ#�P{ z��W2�T�����;���m����Wd��a6C8�o�l�l؃ӧs��
ʞ6�ʪ��-�lo2Si"9����y�&���PdIt�˽]	V�����#�:ha͡ayd|	N ��o�$zp��~ؽg��\D�6��-�~s9/��RO���ED���G��^��Po��4�xOl�.�$\��y�hK�}9�4��4G�w`�.j�{.;&A�A,��H��5ƺ	�b��\V);"�Ũ����V��o��CpI,9J�J�!���LJ��h��b�96	e4"��PiF06S��G*�F�ޑ���~h$)�|bNM�Exs�a^�tAs*D��6EF���م�@�Ђ̒�M� M����BX�%&JN^O��U�����H�M|K3��>v���k���M�4/S�u|��V8}9%��[&�l	�2Y+ʪc�C0*K9�I1��ɔ��(��x�t^8o�~꣱���$��!��Н���C����
.��JH���<�M!2��H���zp���4�G�*�wV��rR�c�dz$s�giO��X=;&�C@d5��h�u#�s^3cf݄	�i��2~Y�"̦I):1{���6�5#�F�*j:�P�n ���6���ߦLH%PI5����B�h�Dh߸0SWPn��F���G5����d0��5��J�A���	wd�;��\��SM��*.�"Gm�*����8mf�0���L���d��S/�np	�}����Ū�^[��1�3KL�>+x�/YL6��5�	�o*z�Y��-�{`���F`_�)E �����H�"H/���7��=CЅ�+h����;D"�� ����D��j�Pp�u.��)����1��˄+�R�\�����Q�cML�q�[��鏂�0�NLiMD|&�#a|����T��W��}0Ο:^qe���Kx/	Wz����"��\Wo�e��L֢�2���s�SQ����)n��<��ua�V��xTm�c��"1���O}|5���J�zPx���=�K)mU�؏��7Z�Z��S8�5�/��-ׄqpR��&wr���\e��Ҧ���������N��I��W�+u-��k�3�.#{�����A�-�K��s8��9�Eq�Bj؛��k��H�!�1%x1N�buK%�f�BQԄT�����S�@�	8b������� �/�����v3j��� ��'HF�yN��& �G���Wp�N�Ao1@.t�B�I�"gc���u5?���=:1!� �|'�wy~=W��
��6P�z�p9N��߁�$)�/@��\[+itd�eޓ	'�tA��v��9��g/ ����8'0��(������5`���Rw����F�	��786�-˳p��4���<��?��]�(�lK����cu�#�t�+M�:U�*���H
�a�T,�W�|ENG)A�L餎_X��i��kK�Bow�	
���[:�K�6%�l��8�d����Ҭj��T�=Ca�B�����~
%R��EY u	����K��z(Þ��&N��xN	SdhZk4��l�ek�Z�&�(�')�ӗ(A��jsW�������2D�%	6#�:l��Y���-��60y�0����3DT���+K3B<r��2��i��ɴ�k��UJm�%��Ѹ�ہ�y��J��i<\���(;.�9P)���<���e7:n�X�Q�rޱ6e�8�8%�V��C.�c�Fɤ�]b�3��1�4��	�!������PrѦB3-E������d�Q8A��ϱ�V�Ԕ!�C1Y����A��|a`�3m�0]nT�y��t�g�vm�C��Z̯-�׫�2i��(pj)��h�j\VZP���&1�b���sh�����XLĦ�X�@�u�x�&ݥ�f�!,�R�gnUHQ��K)��Z��ws� �[����n�HȦ��/'�,T���\6��K!
�g�"�5�q�����ȡ���+�	�!�POɳ��7�K�hwܔh�z#�.��	��Dc�@sQ����8o�᎗���񡢲s������Z�C���p���}X���5��)�D��i� %�K˾�Z�������V��B�^g��?0sz"pi�2�''2W��h�3���}C#�����͆��z�z���31��#v�zBZ�VmC�W�"��,�Nr���	��2:�?I��:?ST����|m�b9q�����e���Q�+&�S5Xc"1��a�I4G4����4�0���Rќ�0'���(�X��u����2�E	�.{�CWܤa㙘������݆�{o�Q�̺t4h{xd�:S�#�w��(�v��T�5fYp]��,FȸS�~�׎�x��$�ë��";n��S�6KCX׻�p��V�@G]�� ���v�d��N"8#�y�ia 7K�Pi�7�K2IV< �QfZI��[H��f\�����\qߙ���g��v��L�\څ�HƈC�h$1#���"�_�L|������L�c��n�p�d8�Fn�C�¸K��&�#�i
gBUY�����$��,صJ�R���J.c�͡l~2UP��'S��B�Jї"�0ٰ��u8xnD���D�
�j��#����Ή?Y�4��:��O�5{N5+�\O�$Z��c�q
���#�.�D�ULB�"� ���S`��AeŅ.T��s��uIG��u�Y
.�ǽf�
ߣ�g�|B�=�t#��h�?Sn�;���!�Kƣ�����9lP��%�PX$&��Ƕ#u�v]8�ޝ7��=��K0h\�2�8R��>ۘ�����a{Fq'W��f�����f�=�skrK�)[A�H&�&� ;�r�Ä�~�ƀ�I޶���w8,�����.��H�
ٹ�`7�0�G��t��X�dE�\b�<w"��o�6�Et�x_
�� ����gGw�[S��B����Js`�ӳ��1�z����S�e��S��P�ְ�M��n��eb�r�H^g�d��bʘ���2�*l�����V�؉Ҷ�)?$W�(�L�[ƖYR�&�$5.Mu��l��11L��D��Ϧ𗂁������p{�	C���������r�h��j1��Q��l���Qsi:c�dRe��q�l���fu�`�j�#T\���p�]�
׺�{�1`2Z��s��-l�l#B3����R@֧��¤u'�g�J��=zn`�>�?ㅛQ
���(�Ln�w��F���I�Ѹj5�;w�./�v~�G�Q<P���#LJSǹ'l��˞�:����%l����lj`��DK��r��n�*��[��I
ÝY��.҃��8�WcJ�;_�BCm3*��m��q'B�p@�4y��f!H)�.�m��̞�w_�W�0⮟k���_>]�:}2m%����9.\5�v�4Y�M1�?׆�؞�U+��f�����F�i;ѩu��)tB�����V%�12�+aT��R�� �8Y����ur�W�~a��0m��I� v��Ş�=û�z�-{�TF���ڀ�޲4q��/�5���bJd`��K��$��g$EMA	�f�>+V����J�m���'��bz�ƃ�z%n})��� X���'XQ�q��f&#��^ �NZǈ���)Q[��S�t�ێ��v����qu{�l��)���E�����N2�<�L�f-tNf.M��%�*[#��:�P���ڢ�9N�7G�Eg���(+�SG*��Ji�{�1Ft��W��6�$n��J�{��]#����8��v�W�0{!�A����4[��r�!i�D2��U��%i���u�������؛)v�n��7V�\:����LWA��1�1�I����je��v������Δ=��|w���]{��C������%��]"U�S)N'"O_T��W�	���޸x�J2����.�Y�
@G��ÿ�`�W�l��	3��V�Y�:q�°�-�R�'��q��y$���N���_)��W��J����\���8��约���}�Ċ&e$[GIk��M�$]<����t��/bU�m�.%�X���y���_�x1��H�T���G���H4	�ㆱ�#8#D��s�]�oh���J���cЪ��괟�ʹ"�<�}�¾J��Z�t*�mYXX�z\Z~�m�s)��%�0���IG����W
0- \�Uڱ`e�`�d�R�-%�p���
�d��S����Ƽڸj��;���#O�
����"��Eh�� N��]�HN��/��L/k�i��ǭ^���
f:�Z�	\�fT��k]*�lQ�}/��8��D���{6Fd3��e��crf��ϵ�K;:���f���W���~���n)�����.ȹ��y4�y�#���mC�q\�WW���Z��}�Z� K)�����f@IَM��ҭpY�OfֱlrHV�M[�lG��)�O�{fdH.s��m%/J� 窧d	%�^]�x�{�/W�0'�zl�≗���Nҝ��B�+�F\�B��<�>��'��(�=6��N�.�2���iaVq�iN��n!�Cu'��f�^�%R�l�r:�h�$SТ���ۜO�g2p�#�u�s3"�Z�8�R؁R�<��YF�.�"r��2UP�5Z������ė�f^7_����g���iu�IcG�\�I�n¸�7�r����7e�P<ĕFz�ss���%��՘��R,��P����3��^�Ĕ�1f������rR2^��ٓ��5/��T�
)v�,����7��	�$I�dE%�oFe՜� YZ�b:cࣺqT�Q�@�4�>����b`R�c/��=KS>�ʷ���yW��(���c�b��X�
�:�J�P̟����3'���e��mڳ8G���2S���C`�IX��u^7Nl�W�{#JY�0�A"V�$E�# �U�0��h�ʛ�wR��F�L��}�l�5�e��K�
�7n�֧ν}a��g�
�-\u��5O�>{������}�v�Z��)�!�Hnq|��/@�W_�f���#1YK�"�5]�^FCN�|���b�.G i˒(��_ӫ��-E$�A(Nb�"�īLI��~�Z8J�[s&��.@�&��#�H�;H�q
�K��rh)3tN��D{9�L'���&[[�h��(�IK��n"�"A���U�k��ݛN���o���O�W{� �{
] AQp;�ز�/dsJ�u)��ʡs&�_������m�&�z�Imz��Y��o�/��٬�َ�{�4�s .PMQ�@�-�BY����)��P!8��9�
eӓ�W{NMT��Nr:Rݦ�>x7թ�@��Q���]����trȸ��nm˩���8TЫ�iZ89$T+o Z��_�p��+_:%���5��'̙3�.�>�a]_��ӛBO�C}B�81�JN�}Y�j+Uˡ<��/�����il��v�xf��;���L?S^�U�s���iXߩ���z��	�.�Qż�m�E�ET��������[+2<�&	��y���&�Q�1�,I�6���J�l�����ӲP<��{J3�Cݨ룮��xkua�G����tG����z��M>A�:���ř��oWG���|b��S���o
a�O|���?<�������N0���娛Rh�)�:�B\va���K��C]����o=5���_�G��啕ZC?����x���B8?��,_�7�w�v�S�4�v�x�
D�W:��T�(�4�l�g=a��JS41e�g�O�$D��2�n��9%�-�9o�~q�w�22�@󦏛���r��cG�GNT'�W��~$V��n���J�M�P��]�Ęj��4w`���w.�xh�״e�Ӝ_�͟}/4�G���Xм�n���Eꀻ��c���74�����o}�{O���xKu�euپ���.�?�byj��U���./��j���4�;�{�'Um��U�'M�huR��;Q��B�-���F)2o:�Rl�q�1�Ou��\�5\q���"g_���}�&�}����C�~z\�+��d<_�{����]�
I��G3��
)�[Y�14;v�����	�����?{r4^��y���.B���R��|mu����-�;����O�z�C'���5���p�Q1���¯��,�r���Z�b)����L���(,�(*$�i�c�� 8ti�V{�,��E�y�7Ώ�Üj���G�8O�}������{���yU�.��nW�?(@T�B�TD)�@�D Ԋ�N����K�:O�:��0z��?|���ve��ϫ��:t;�C4#� ���J�d�x���Y�[o=)ZQ.��kp�5}��G�n�8��="�&�Jx=�*��t!=?�7y��G7��ٸ���Q���w�����#��L����^���^�W���>�ڨ�����w�-�/��W�#Ӛ	S]^��*�=i�]j�c2[B*tE����ж3�n����C�vͶ�=�ȣ��mb#�D�֏�y��o��Lm��fkf(��"�2sO�oe��f��By��Rk)���X3aڵ�Cٹ�OR���[(��F�߅햆(������#������V6m����8��O������� �����b)�bw��-=�r��8�EK�_���L!C�b%��$B�3�S�����\A��N����w���(x����>Ь=����υ�F�s.��<Ӝ{-)M������5FŮB���'���>�-��9:�*�JZ������9�͞�Y�7��z�G�g��w�8�8�O�{�q�O���J�NL�Pǁ5�5&��ǎ�φJ�[�v��'b��B�6#�A���7|�g�=�p���{:s���T�8����Mꭢ��ܚc3k&LO4� 7�
���Fm�U�(����{˳Co��u�"�hC�{�<��'��*���$ʏR�4�%�@ \H/MM͵�1�����n��IT��e�*h���Sݷ������x���7�|�6�������.��uM�J2,���n�C�����?�W���¥�D�Ku��r�
�C{<�����P��q佃����~'�|O.w}��#
����`A�k�T޽}�b}~�����ĺ]D�X���GO��z׿ن8x0:���9�L/O-ܐ��f�$���y��k�b~]����bX��j�2���d�;p}#s};o�z~��M������7:�<�slj��ۣ\M��F�b�t�K]vW�r�uf׮�ZcO������ɤ��i���3�����[_#W�?ʛr�G+�m�_n���e��N
I,�ܒ?�oR�������Xw<�k�����^i����V���t��\ǣw/�+�]^��4NPp����m�WTۿz��0C�����o���C~����'[��&v}��׿t�˧F��������/�5�ݲ&�?�������_���NnٕR���w/\�y�n�8�/�,����3<8�w^QӅ�c�5��B.v��n�EΧ��[C�@'^���Lм̥�H��rx�`��0���uS��V�I���59y9�k�	üH!($B{�����>�M�R����\@1t�l+�D�k{y#�I(!�\�K!}���κ	�yM��w��}FA�J��·�ؔ�k
�ecc۔����1(F�j������ lme��Zk�V=su���[��5�a�HP�q�����l۳+�W�E*̎ДNI��=a����0�$��#��qbWP�u>D,m�,�t[�+�q�
S�P�f� ��eTRB"�S���y�Q�[	Qk	����G Pp��VA�AǪ~�������xl�0�n����ୖ���!Y�.�Rp�y��!%�3�yt�(�>��͵�� :��!pɩ^���~�ȶH��Zy����K�`Re}���!����[l��ɾw�"����o�!.#��.�A���AAC p�[cd���x��s�`l�c�O��L���!�兗:A6/ӹ�D��8iAo�a;�m"a��kP�����J�P�E�4'�&P��\�AvU�!"�)�-�h��ϵ=4�M&��p��c!M4oё��ށIC��C$�t��~�m�c���T�|�)�M:���0B�RI���$�^-�)e��ѲP���a��pM�?_�-J�u�vDeZKG2 �U��chx:�0@]P�z=����7[�e6T�jGxܠ��A�U:��	�m�xa69Q�a���$�&����Ҷ�4���� �yjزB%��F����t\-��*��C��a�T.��aV�Rg���a8d��tc=1y'k�*L�t��u� 	l����5�ɔ����g8�n���y��u�q��8�l���V�'L >�8D�CO�RśO�qЙ=F�-�٠�g��Z�R�}ph����	�eŬ+=�����>oչ�1H�H؝!8��֙o�1c��B=׆�uO���+���W��@�*���Kڃn��4m��mbD�ho��K�i4���ұ1î~�m���c���^��YG�on&�%	~Bl��.������2�ƨl{=�^E�f�*���y�J��-\�MD6#�����1�>=
��f*p�jj�׾'��{@��(d=�[�e0NLG:���&��Dk�Άc��n�B�d _��lh/:6�c�l;$���"�J�5#ۊ�&%ʦs�9։�ж�[�*=�Ӂ:�8fvS	��\��[ye��UY����U���J]ʆ��Eڸ��uDv7B)e��J�,��+3�jb��`cVk"����f��-;�dǂ	 �O���"K�u�����:�Ni�M"F
f��`h�\�1_m�a�������iTE�`�!J���r6�Mr�LL��v��`��&^�mi���9д[�<�K	Ds����?�)�i�e    IEND�B`�PK   %�X��%� V� /   images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngD�eL\��qw������;�ݵ��݋K��www��Nq�b�nv��Μd29�I���L2��r�H�H�
�Қ�{�^��<��9�]���r�53�g�
�ھ&����$�O[g�����]1			c	S����##��/��!Cj�pNȈ//��#PJ@B�qr�Lp��-~AJ��h��g��ֲ?���+��5���9:d9{��#��.�>j��&`�cbϩvac��]��o>+B�Վ���	C�0�����E0U	��1.*3��u/z�a ���ߪZC��{��c�/�C��/���U����,�x�.4V� �|��a��Hbd�|'G ^��*���w�~~5܏q^�7ޙ��uF���{z��Ls-�7��g�����n�5����M@�����ǥ�b|��N$+�MO�����7�ਓ�Cd�-ϐk&�{������D����AUBC)����7�&D5"��GeG�˖��O��W\�����e������1}���>L�v8G��([�D���(������#O�BZ�C0@��Cd�I�z&�je��q�/>��ە�[1�,��(��dxc���y�*b5{��8�:���)0�zGUj3N���yb��A6}�ϭ��&�Q��XveH����ʈ{��`h�(���c˸����e����Vg�wm�j9�E�����=�o0f��	-� ����~T�"���XӴM8&/��~���X�O��T꽴B��>�����<D�ՇS��K �������M��!x>����2�qb�2�;CD�=F���ڀ��įTr�����*F1�Z���͒f�?q:��kk!E���j#�>�x�Vmջ�f�%e:<PK����5�NsⲂ�Ж�t2�2߂8����D/��+�3��r?yE�� ��B6y�Ő{:߈������ ���X;��D]��\��,B�r�|н+�g�_��$z�'�*D�O]��9���a����83~�C� �j�j�;5���r�a��Ë��E��O�H,�2N��BF�x�B�0_!��_فU��7�����'0P<ɘ��1�J�&�>��A�X0_�9Fb��Z{H��c������a�����D`�i1�\����(������#+f�*L[��f�-��K;Ǘ�)���ys�	F�L��f�.�Hs���������f#"��fc�G���E����Avt_���;(�f�G�j�I7�*�E�՜��M>݀q�f��\8G�h�P2�(�Jr��nB�]ƐL3��Fuj�]�&b������P�t���+��R��Hu�?Q�UT̀6P�7���H�%�n�*�����9a|�%��
�h�WCI�#�5g��&�;R�a�$��*�؀FSSs����l֨�����TRR�]��������S���� d7�BVa�8�/�Q��ࢆ�!n �7rЙ��&��\V:i�E'g��:NΕ9�L��+w�0�j��@]9��|����Ka���A���+�&�P��S�h�3��*c]���ꊯ0�PR�Isר� �w(^u��ׂ�=���G�K*4I�\H�B3�o^r��)䦋	/	�}�/��7P�@�r3$�h�����g�TX��,L�׭.���rf��7@"'qa���-�B*y+�E��Of�Ks{�US9�xzG@2�Κ(<}���b���)��Fv*�^ w�eHyV�7
��)���h������_�cI�L���'8�g��8`k`��O�X��/kA�͌��fT1�o[}z������*�kE�/Z�����W���@�W1t9�5�s>m?~e'�U��n6�C�����I)��xN��1R,��Գp�����7�u᧰�{��y�������e� 'RC��)��F��]�sᄰ�����؜�؂i�Bb��FFѼӛ��厎�2�`T.g(\FR�#?UR�2"0�V,%��^���P�ZňNQ�0�ҿ�5��x�&�Z�1�1�_�N�X޿Q��5��E���f��ce�#�Ki!�~aW�tZ"���"��3���>ڡ�3��{�K�&WϨ��Ց*)�\=�?�;����:�=�� �[����v�
[� ����gfe�N���+q
	G�`�����n��]6�]�hCh�d{k���8Kp&?��m��*P���1�01e����xH��h�]ۤQ�	��x1mjoz�����)����:���W�J0�Z�^��h�ؑ��"�|� ���2xY��n�l>h?���!�d�=���B+l�i=��N�C�&��o��,����38W�-((���/��y�x�FP=�e")1J�~�/��>i�P�9�s9���z|.ypL�@=��܀1���( ���>ӏ*A�5�5�ogrQX/���>ܰl]#�aّ��<���̼DOG/6u���^�濜����̿���u8{�����\�o# 1-Am�',o��Ao�|��ifUX3���t�
󏼔�lL����\5�'dk̫�o���	�H[��btM���u"(���������W����QoF����>�D��GC�MJN��F�ki��+y��k��>@ڇ��~8|�gNʶ�r$�E[Y|d�2�P�2b2��b_��ԓr^8a�M��vchn���8ܼ"�á�_��{p�_\�\mwǻ���uqG�vƦ5j�=u����Wh��/UBL��ocE��N�������H��x�$>��tgñ��*طZ�_g��DA�4���}��t���gG2a|R��?����UB�eb�_�SB�f*�{��]-P�JÈ��e���y�|#]b���j��1F�b�,r��;Y.+ �#Yh����kH���{_:���F���.�"�Ɨ�иfӱ���o���QǑ>�w��bZ}�Kk�T�J2�l-��Y�����Uի�L��w]���s		��}+��ӓ�>��>zv��L9��Ug��V�*B���d	�+�ڂ�� �E��f~A�?�Z��"I���_�[0��GFk.����X��&��R��Ieƭ7�{��lI�F�ǜ�3LM�X�;�)�>���{�V�9ԓC��w�s��,��ڸ�]z�5TiaR�9�*�%�b� y�-��1r3�?�A�!$�jC!�����"�
�����m�ϋ���	��x˫~�5@��W>�P�꤅�Ռ�*�d�eW0Y@����`t��T���/=������|��u)���\��
cl���/�_�C)��y^~I)�:�\��>�f=q!@��O-
��*�/��PZ-�ݢ?T_j`�`�<�u���)�x����r±n��x��t}��{�c8]�9�2 ��c.S�S5 �ĨS�x��,��Q�΄��?���e~g|�<{�9��$4��/!��~�����������,��4��W�vh�hf4�Wb�8EO�1��<�������c�G���CHM%Vgrl�BQ��P��^}��WP�����Ы����`P+��~�r�ŐR
N���2�`]���@��B#O�Ex�*c�vv��#��a����=��/Nu�N|N�}�~^ �ԫ�qp�|�V�,<ĕC"��Y�|Æcv=\!,
�w�e�	n�����-�5B��8����5������C��*�!����ZZ����,����H3!�9X%�w��f<~���U��Ʀ��0h:����y��ף�s�"\2U�]��{zP?��#I*s��L<�̾T.�r�=܅8g3��E�����>�k�x=\v>�B�;S�3����q̵>M�]����X�>>>�#�9��1x��#�m<�!*i�j�/.�D�����B@�%	AM}V����1	vl읾X�E�
^^I3�<t��wN���JgR�1����Kb��0�^�ܠ��(=R�=���M@��wt�r��ʅ�Q;yd#(T&%��/������b�׈si��1495r�����I�_t���)M)O).U�,���k�A�� <�և��^��� ����C��#�L�[��f�+Ð�<��'c�7bڸ�&�^=99�����E���H=O͵�>���e\Q{u��l&f��Zwc0�an�&b�P��U�X.|F�"��'Qb	u�^Ԉ^�'<q������������J�?��ʗ�	�Ȁ��OlP�z��2��_��Iۀv˒��2"\��g��.�	K<KS�_�hG���wn9���y�������B�²�9����-��N��dR֘Mw���JR�`K)����K 1������}���9H�G=3�MzsT�U6S�_�h){�>��l��͋j��{�\Cv+vVA^�+n7���H� �#�t�h�������ŕ�2q�$�P2�h~~�\xZ�����p	��t	�(q��%�&��d�߻�iW�.x���^�<�V��2ֿ�8�`[���mc�3��e�e��o���⹾�#�v��"Nrjj���b��`� �� �q�2�+��F��1NNrk�L^��;v�@l��o�0��~Y�����96�2�B��������ﮬ��/$80r����-P���N0��\�큪���^�bM�T�P�﮻�yv^I���r��%-�}jj����.��`�Gx�@n�aM�зg8'�5����(L���࠸����?<[���
A�GCd���W�?�p7��X��T�`D�~�D5�#*3�������](Ϯ֑c�A6��]Sc�����W�������(Bÿ-ѧ��m55ˠ �<V�\2�^��+�����ڴ� �hZ�%�0�1����o�$=āҾ�yA��>c����K��9��۟q"�:�NZ����< B	�4n���Bػ�^��z?�Voj?K{CnoyU;���}�LJV��卒m�5Ӟ��	�-������J�z�G�,!-�����l�W�(~h��JO̭<�19�S���.Ȯb�6���Ijy��'�
�0�^N�"�䜖�إ)�IL4��`� q�D��[g���1��,���Q��	*�E2����������9�2�V���g�`��nn�c�R9q�ɦL���P��c�R���;RQ3mˆ�.��D��"gKd�F�>}�+��	}q������zf�]���@���GDR�̟}����Nf�,��vl|E�MS��U(��3���}���
�G�����f_�"�ʔ�h��>LM�����#�fNF�Hp_Yu"���<��2��`eU
�`c�&���584�Q<�\��N���heov(jR�L�B��@]�'�<SW#��7,�������n3��sJ5h
G�be6�����O��]�XJM�5j�	�hh��jeU�֫;��*@�9�ޕ@�I�e%̩E���i-U�N��XZ��򔯑��v��S􍄆Нi"Ź�0[q�VԅJ\���:�ߤ��*�PNV+�� �4�K38�!fJ��iI'�$I���D5
x�x��������;��@�ǌJ�N g6�f0UӮ��<�!��O��j)�[M
8yN/�ҋv���Jlm���_�9�� ���lg��A��������#�O�&?�I#Sl�� �.�_/�!l����|�LӴ��6�ֶ�e����^I5/./c=�~qr��(�o/֑�'��ɢ� ����?��h�㬈d�GTǝ�,�������M� ��['=���}p]H<H��'~L�{����U�_M|\����y�����>������L$�Y�����\������6��|���ꦒVi��� Geu���^�����jvmfjwV	���@�s��.y,HbE��[��K5���T�J��c�!�{=�=�G �c������@7��>g`�]�J;f��X��X5u{��Jd��jo�����VJ�!����)����]����G��b����Şq��yx��Ơ<k?�j�e��+���g?�\i>���e�X�m�O��y7��0�"��cFɨ��v^󰦜�r��a.Z�'bUYjSfP���.&�̢̲��r�`�O�Y��d�eY��V)�q�	S��}��Tkf�����wE��k�_�u��Da��=�v���Z��P�k�w��ޣ��nf�^��ز1*�dM��#ʃ�,X����WO�.�O��
�%�'d���kq}��Ԯ�,���kV�\��v��iN�
fE�ld�\0�gY��,JJC�t�U�����P�y�~�m3!�>!�N�j̬d��jH!*J��C$Y�Y�~ւ����=�,(ɡ;j8�z3�T���F�� �����ìKO�-Mb��L����w�+�-��L:�9E<2"賨��"�[���!v��@��,0�;D��d	(�3�qF���k%�7��8Lg���R0�HE���������a&�}66�a� �f��sq%tEϮ~�;�H��$�1��*��%�����i�k[P�� �:�ˢ��	�p�̟�<�]���ћ��F�R�#�,�!4��Ѕg#nکgB�Ǆ�1��6�k��JU��g��+P���6U��`#�& !�,'L���M(�H?�&y�o� �_��S�,�t�#�kJ9Ws�2a2J���ڵ�eE�igC=+`t̃�|���l��P����2��$c�9B������D��� ���j8EʽU�7��G� d�E�Ţ<�5��7��&Sb�^���y��9�V����˽��������Vx�'x�|\�߫h�����0�����෰L���*�?�~s}�}=�哽�|��E|E5�u,s�����-},��������kr�;�vT�h��(!=S-�>0��#�gll�沽�g֨$4B���9p���+�$<�n#��&@b�Cր�7��}nl�i���ML??[�`��5�{>��>�%�P�ƯԬ7/ ��ó��y8�,`�J!�'����lj\�c�����p�z���Kc�ˊ�LU� �S��}�l����9q7Y����I��i~'@�B*it�j�N`jÑ�;�}�7$Pѽۆ7I:���a6�e�g`C���Aqإw�!H���ƺ52~G.L;?�*
�m�v�
�1*�{}������HK¨���D$E��Ϸ�HB��̩IIH��%D��v ��.�iό�1#�9ڍ�)�h�r|�	��6��0��+��|#�o����"��}o�=��j��@Rs�T[Nm!�R(d�Ij3s���7�6أ�ekbB�'�d���pLJ��d���ϳ7���q 2?$��rx�+�f_b�ߔ��)���0c�w�Q�6s8�tOsj�Ec���Li�<9w�yf%���k"�C�[$����-)�rr���|����:��r> �{x�O��L����8�)�=�z4������l���݉�AOҢ��]eM�&ޏm|| �|���r�hj�r�?)0�NOn��G�
2���W�$���G�%Z����>cO�f�{t�.P�­�+����p4Ϙ=�� �ue����Ҍ������|�ɂn0mlO�}
�X�dx�%��9�,� �_ð��f��\R���lKl���dǑ��+n��L��x]�3�A�Jxr����@��BN����@B|wM^D�-����ѥk	JU���ؐ��<�ѳ�&��y�kp*��M�i���tt��T���M.����������i!` N
�tj��NP?ص�{��?/0��0�8�o�]��W˼��������'f":��/Q~u,��u�|"�s��8{��Pm�I2�w,��?��L/�p�����n$((b�]�޿��gLx����~�3y�ܠ?��A'�	'�7;�q9a�C쎉���kaÈW�9���-���z9A9���;�l��_aa�����t�� #p*0QS��*X���Fc� w��CJ&)
]���f�
���W9T���7G�K��7���G�/L�>?lU�|�<Y�[�a/eC�U2Y���D[�+�&t�O�r�/^�:�)��o����_9g��̆b���b�����������l�b�2 |�'����
��F�J�� �=��%3,*�������$��Y|�oҮ�n��[�D }��\��h��yC��և�IF�����{?�**Ȥک�M�o�"^�k8.3Ӗ~���`T��O�u;zGێ���?�0%����a�t��:�̜sp:��O�$��	���j��
��栌�T��3Œ�>�~���W~���n� 0����Z��Q)���ݣ-�rY�ɵfR���=����|��/��~r��<�S1��V`����r�����R@H�����vls<OB��Q�f*:JZ|m_��zo~��I5W�A��1kXm�M��W0m��M��Ps jB1Ϛ����O�Հ]J��_��uuS��)�Q�l)_4���ccj+%"nm��з���D72u�R����tol�RPBty8+�k����ā6�V0H][1�!����M��[�&��OD?o,Ǔ��	���cV���U�t�3㝼��Ҫ豙I'��U�^����6-;�S:�ݴ�n���g�ͽGN�,�C���(��>oUƲ�����eU�/�~8���<l�םVNl8�P�r��v�J�AY9C��NZ�m+�=0u�!�ɕ�zp��!*����mXh�*W{YB�م�k�#�;}�q����t�T�2ad���������'���Aݣ�Ĉ_[��S�y��+����ý�7���I���{Re8�s/�����,kq1�{�GO����pa�Rfq�����K}�^��4�Hu���r�qb	�o��#�c2&�_ç9����.�18���鈌��ʔ�X��0ڳ�u~8���i�5Ҽ�k�It�3¢�M�qJ]R�L�9��P饣������qE�Է��ӫ�q%!{]3[23�FB�F
�;<��	J�@��E�c�)�(�d߀b=�^�"e���QfX��j&���!S��ݾ:�\��|?Q���^�3�UhzIA+��3�1�9t���ϞǛ���p?��o�D�;�:�_	�.��記0���:���aeej���g���&F)���#��A[
J{m�	��]���I�e��b�45%=�|�	�<�?e>>�-	�V>>V%�L�
������9��A��~B�Ɛ�Ϣ]����3X@³�g�M���`#�*|�/[��c��pG��6�ϑQ^��������?h67�	[4M稢M/N��qgϮ$K�h���=�η���\��\���	�v�#|xݚcm�w�P��b�Ȫȃ�zS�3�NW��1�|����b����}�*�u�;����d��3��H�|�SD�j$&ng^t�5V=&Z�����0���1B��*'�S9)��AmF]�k�W0C�x�,�Bb�a	�e��U���F}~4ZFtQ�K�Q�Q���i'��"�T>o�3�m+k�=,UJ[f/Hz���W
��-M�����fA��K�Hiȱ"�i��`�>�qr��X;��Yː9W.�u�mA��7ޜ�%[��ዟ��қ<�/c��?�G�,���^T��&C��g���e��:�ݾu#�����ꅫ<Ui��,��'
�������
�%~��^�qM��v���cj�9lJ��,'t���d�N���U# >΋�p�p]Vk�Т�#;M?�b�OH4:�BM�X�T�\��S�ŞZ�;�51|D�_�L{B�\�tQ�K��������ڱ�K�1��Դ«�[*���e�f�����B_�����&L|�7���@���7`������FiD���~,Sd�L��@
J;�?U�q(w�V�G���q�-c[qlL!�jJ�17�3������019L(�^h@AXq<�%���$8O9�����>��1>����PE�1���	"���>��3��B�r���0*�ə�T3��a��(O
AƆ���Ba)l%�Z�Y���lp![�Y^T���:+Ꙙ��r�l"ٛ��Ԟ�,�uH�,�q��{+�����i�Kd�qBDU��.�k��- �"~�y�5����Sۇ��,]��(�����~H�l�}�M ����fB *6�#1)I�]�n��[��?�{kS�z;,���w����F�����5�ǹ2��\�XE�Z����j^��F�N�6^�d�����"L�r� S~���-F�kj�[��M� !�Ďr���߷�F�9�Q�+��-�hq�Q�u�8^#�zE������Vʜ�}@�cB���Lr���p8��a�(VIhV�#7�z���q���E�ۃ{��,���P���Q�T����K��e�A+��4��y�����B{�,l�S�7�����?ڰJ=��M�C^��f��ԙH���w�z��n�5TҾ���z!1?2N��?4ax�$�ə7`V���҇]��ȍ�8��"57(�%�CT�����L3yka��%�7p/�/JA�X?�}=$���H[y���9ƴbU�ۡ�§�RE,�y/~<���㔜j�����1�
��f%�C��*v�
[�$�j��>N]WGc�{�*���Z��c˕c
�3�K��j͒��=�l���M����x��f=2F�0�$w[<S��$��E�T�(t��X������f�"��a*��x������X���tK$n|�=��@<�.������l���q�|�W�;�)Js��:#ԅ��c��'�|���'&֎ am�-���@N�6s�IN��2�r\�i�T�A�lӜ�~�>U�A��)�����c61S��,��(��h�u�d駂�MY<A��\�9�R�
7s���F��x��M,���2.��Ur��x�.�5���w-3���8�ܿ�E�+$��e��q�c��F���2W�@�۷e��s��/Yq'�x�wq-�1��ҵĖ�����(e�|�έK��{uH��l�|(sQ�������k�΀
ve��=r[c[��A�5��#[]c',ׄ����qg����T)�3�f�t`Ѥ�ɝ����Bب#��zcٚ��дޕ�K"����Xɚ��@'���.��G�����0{DzI�����Q��TF����;��.���H2'~F��Ӷ�O���Ϛ��Hx����b�oOc�/��W����ӄ�fv/���ڨ8�\�X=/3�
ϵ<���&� ތ�:o����:�o6(H��=�(\�e�&��\GEb�Wݬ�ܯEg�+���?�����QP�����@��!��P��M��c��g��e����Q��y�*�
�S2�ր%)tT��ǔ+��J�����+2��4��م�q]X�0Z�ݿ�'�}�	��~��	*�`�x�4��W�o��~��+~�:Je���] ��i�:��*߃�Wܽ��L���1h��:osO�`����ʴ�T��;Qx��(�.d�W������6�P:��eWСν`ҏ�(L���#�8v �ˀ��`���{&�+���Z������ ������׏ذ��аu�R��U}���JD+7+w�@k�U#n�x�A��xL�;F�V�g!a��0��XWۻ۫�� �;}�|�	N��s<\����8�7�@UqP�_��H�]�g%���;^�)�3�����_����=���ٝ��Fh�3���|���2J�{Z��H^��0��^�o���H���S0��L�8����Љ(��ɲ��	���+��m5E!R�(�\�dp��'����t�)�4��H��v����G^{�x�㿭N�'1�i�����E��D��B�X�(�G�s�e��t�ԣ�*Mg$pL���N��۳JC��͛���ᤸ)�L�R	Q)��2��p+�<4{-�S�j�Ɐ2FN���^g��;���b$6�NO'�G�`E���Gth���ac6w�1\�\��5��ZY�S��y���r�o���G��*Ŵ�e��%�9 �W�:x�����vq������m:pwQ�=.�L;5��,��q�&%�?L��W�w<EL���'�$z���
��ԷS���O�S�nC)�:�Q�#mR�P���L�5z��Sn(u���o����5���>���<O���R���L;m�rt!~�c��Ś͏�4�7���S�;F���1f	M^��uw������(K-�������.���,Ew�YWY(�Ǣ�d�	oЃ�
��\%��z{�=^T괃{� �DƬn̪���n�?�ڀ7��c��{��"�p��J���O1Wf 1R8F
�m��9����Wp��\R�uJ����ӣ[�P�soh踠P
2�38ԗ�����(	���{5M�eK�O4�̟ņ���O�Cq�YԴ��SS!O�U)>6��l���O��rϝiR�-2$�*�p串0��a�za��{�wN�q���j�2��<���L�&�}z�`��>�}z>o�N��m?V���8��}?���`a�H�ɸo�|nxEN�������O)ge9)h����Ǽ��)�����͌ZR��g�o���K�k�P;�̸�$Ƅ�U��τ��8P�l�f�;�S�RV���]7��Tl���XZ8 �,}b�|��|��7�~�w����+�n��]���ˍ��W��=�U��Ǩ?$@\a��.��4��`K�Cl#�7a>��mn�<���r�j��A��ck@�������0OR���Y{A�xS3a4֮:,^�?i�3���.S�T��~��S����Z!��mB}lM��F҃���l��$8Pn���2�rQ�)�J:�ȯ�t�K�q�>g��)�)�(�|=7�Y��XExI��s�	C���J:B���a�>1N�P��d���}Q��s�(�i���Xˌ�4#���T�? c=�|��stǬ���}ڏ㮵Ӷ�o��Wɇ��I{�<��X'޽`Tׂ8Xӏ.�~��J]�����e�S��0�ۅZ�����E��w�k���&��m�&g� 6gr �zQ�y�\�L�3�Y� $iMo�,iP���
�������e�DgӨ=IX�8%�5T⢂�gП{�Pr4��T4bd�P-�}�Z_Z!�j��"���s��B���^�>=[�����hY�{f�̈�ĝ��W,�G`�������j�z�� ��=�'�����PR�������Z���S�8㫵;al����%�zJ,O�3v|w���du�M�M		-վF+��|��Av޴
���]��V*)��>n����l�Έ�/z'z_���z��.l��_j�wIp|9�|��B�F/���p�{�[���h�Ϊ�J|�/�� �����[B�Ed(���D��ߝQB��p�]��&�'̲Ѭ��*��C~Ǆzf���4ヱ�&̒z |��G�9�Oj?�^;��e%^�}o�[EE6ޅ��.������4r��h#��f��t~�n�}�|��;�"vq�w&�������ǜ�N�3�V��>�����F�L��<�n�|r.�7
��9^�8�S��^����ґ�O� �4�sO*PZ�2qA�lY~�߉�\���F�j�B�����D�ѷ�H.ʤ2�!��ųI�]/�9J'd�$�Gz�;�K�W$�KIj�ņ]ȝ���/��hH�P��x IF)�~���6~�6B)q�G�<��j����'%a��
͒���^��<�3��9%�]����S����%`�z*��Ӹ|9E�����Bk��YNJr��nu�7����|%~5�<	Nxâ\C� \em�rw&�g\'��$���-_<c�ωuA$���;�KƲ|��n�Jh�5����
��# T�i�#����>��l��/'K"�� �) (+R	5{ -l�#�[���}f�퉊^ <0>^/�[76s1p�=�j�9	)�-7��M*����+���?��-��%6�~E����o�F�}`��H�_�����~��N ���>�'6���itNI�KB6���3�<k>ʖ��/�1��R-ͯ�-���^L�ӎ���v��4����5;x���'FV�t�ySR��!e�"�5%����U�M�r�3��$�g��3Z�p񄿮('4[+����y�%ڞ������fv��_傭X���Ҹ9�Ӛ�����jE��a������8x���B|����n�O�Q���E� m�r��sc25���a� �d�	��@e@�
��D`R֖3�{�F�Q��@��3T��E�r]р2.���$���BX����9�еM��!�/4ƫ��I��#�IG�X�x-��H�0f��_J�K9���L�Fv�	e���#%v�ǹ%�������Sw�r_\z���g�EU"�EJA?�|Nx�s��qq��!m�������ϴ����=W������y�BR��ZG����196+���L�{kR��_��/！ίpW������o��ޏkI8aN$����i�f�#�Cت���𵄣3?�0h�%��Jq����5
]��0@Ɩc��(��}��%"E�o���&ι�D)�m���M��1q�[�A�Sl,��lݡ竵 \�:��p����C;�7�0�3;���F�o\���~I�����q��6�,����$��ٙ����흷���Z��~[gI�=�*fJ��� �"�J ��5a�rU�M>�ϗ�#����Ŕ��`~����og�~j-fg����)Yz��JϢ�2�=%���{�k��$�W:�4�f)V̫k�
1�Z��%ª��,xs�H�o#�qZc�G*#�z�~���*Bf�TZ�:��5����5I6�U�/�|
H�me�9і�G@��N�gџ�|+�7�}�&���C���<Ӿ3��*�yd2���lD8R,=6��Q+EM������q��=��a�b�MƊ��06@.C�o!��t�����N_v���Vs�#Vťw2	z' "�tꥏ}��%]}F� ������#��ڨW �*���
}%h&�JP���s��0I�Vtж��nKDjG�lc���x0麟��:4obd4|�L�;O��QG��*%S'o����Ǜ��e�+R~ ؏�8�=�|��6��5����ڝ��߬J�Q��R�� ['����p����G���E��a놢����Ze����l�~U,�f�3�P�|��3�F&�  ��9<��Oj��W�e?#��Ty�<�	�]���%�y^��pgc�U-LO2,M*�h����\{s���\G�]�����qٖi�����X����{S�"&�^�i�PNsIޛ� ��x^�@��k���[e�g9��I6��N��Wo��3N���_ⶢ��K��`U�$��TV�� �v[8^w�_8���u��F�rَ��~���6e��;,���nv��?��bFF�o���s����!��}��e������D|W�ӥ�m���d�Ad�d�p�L/:P�	I�_���vs>)���j�.�!��OX������,����g�ca|��ct��ac��%�|�K�&G�Wr>ߟ�+���`�8�H����j<�D0�ť��rq�7�O����v��4���(����u���9���ﲁ�~��kA�s�b@)�qE]:`�5��܎,�gDZ}�5����.Ѩm>;��,�G79�Qr6(O�fR��/Rp�_���r
�PC&�r��^P:F&*l��XF6����+�L,8F�G�>�"
SO�gw���7�[��
eFy�<�l^����>�3j(w�Y�x&���X�%���N�r�!!��6�"y̝���zt ���6{u�V���@�)�Y����;�z�b+�w��ͱj1O�ߘ��[�Κ�)5=~%��OJ7c��sE�l�>�j#���\Y��"�F�^K8�z3~S
~fnr�c��V��in��%B����m��{�M��cگ��֫��ߧ��}h��J�VO�!��ۗ��� ��Eְݵ�f9z��V�w7����"v��8V�������Tר�6�ϙ�%3<�>���Z]�O����B�h�_��\єm�.���|��<G��`�2��ő'q�,�d6z������FVo��UXc2���dۣe���IN�LK�V�ʹ�6إ����KU�xA�6J�m�CY&�|x��"������R�4�>4\��ԥ1�]�GVhhAo�Ԙ� �Af�T�6��c<����tU3����g�7��SQ��oF�&����PԵ��l��4���F2^G���g��K�Er�/z�a�u!q�M�"<��z)q}4�ť�Z+��37
qf	}��a��\��c��n��谨^��	�;�fu8��h�b�x�Rc�~��I�I��#�L�VX�g��m�p@����K4�MC��Eb���:�,@ӿ6�u� ���`Z�):������"�H݋���H^ 9q��Q�	&��`�5�bcc�{o�p}~���53�ݫv^�FA�o>���W����y�o)��r ��ǐ�|-�Ģn}�UZ���{xse�Z$'x��x��Zm���Z��	�i�ݳ)�p�����2�;e0V�F��.�d����.
f��㣉e+:Fj,e��eoIҳ�t�������=ɝNNt�N1U'S��9��>p��3<z���?����|�ҭ���}��?����p;�3�q{��"�����ȫ�p�晆F���A��շ���;Xi��w;8:ڋ��D��h_k{)�
��S�17$�1�3b.��r�0~K��J��<��|w�x���k��s��{�Ê�k����d���Jϖ��p�o$�P0�@��M�N��u�i�����%��e�P���JfW q���',�)6��V_�Yƿ��o�fg
��s�:A���*+� i�ű�]q\�JCͦeS�F�&�.��~�+��U�0�§l��%����	s�K�Aڐ�,:�� R$Cʜ��d�a�/�H!�6ġ2?3�R�E�[�?�N� O�^��?�����ߘ_d�1&Ƅe+)7@��ZM��P|w4Jc�͓#l���������_}�oߥO���}|������&��h�^�an��k7�ƭ;����Q�����ӏ����.^�����}���QES��HD}Cʽ�s<\��|��c6�1�L���/}��V�������x�⩈�H-��;2���M�#IQII�(���Y_��DM/��ɝ۷�0=/sh{G@��OޗyN�����7�ǾU�R�#�l��Mq"�9J�q.ݾ�\������4;����������O�;�P}�� ��L�lVAmJѱ��M�UQ�.b��1
)�W��Pc��p��%J�.��mafV@�^!CDF�E�et�뒖����"o{	��rIE��AP])���I�?�@��"�T��8��z���E�.�Y+��f%,SbG+6ݠ#^�D"�k�QmT11?-%v�����Y��&���q�3.�T���6�HS�/��3�	(k���HM��JEk�Y.H &+qcq��X�X����[�Q��|g�����Z��;�0�'��8j�#�?0hy!��x��]|ia��&�O���'x��!�J�f�)�d<�V��Y��;s�R�m��s���[R �'}���Яܑ�eٌ���ʓ7PxE~���� kTi巽�/[}�mnIYgbJ_�Ru����zUz�����V�O?�ç�0�8����x������|��w�x{���&���U��ʗ$=+��Ə |��Vg��������b�����/��`wGr����9j�^U
٨�s�5��7*�WD!)��b2�ڹ;��᱈�nݺ���x���BG���~�����%HF�c.u�b^������Ө�dcoWG|��¥]m.Eg�r7��{U�u�-A�)�D�
�Y�J�%�X#;��]���y�Xlt�[���>�v�1�w����n>�.�x�F�/�gLu-�g.H.�z��@���Ѫ��(T�X�3#��#Q��z،�]�8�B{����� ��Phl�z��M1�e#3�u�(���0��)��^�|�o�ۢe�f�1&��#���kbCQ�*W�B��R�s�
��a�`W@x��������krk�;����P��&*F�~��ﾆ�_�^�vY�����)���q����^��o��V&��9"��I��i9�8($�l{=}���S$A��K����+7o���ma,=����=��e��jbnv�SowDXEG�����4�,õ�=�v���'�$�s���"n^����i)k����ǟ}��}�ؙi��"�T�������"r�(������X������Ա���Wp��u���%b��'���h��4��� ;�ڝ�2�E+ eo�Bp1����iE���ʨ�a��s�ٝ�ݷb�0+=��73>)LA��c	¼�إ7s�E�wLU�X���2.�sG���*�d�9����/Q�")Z��Nҹ�V�./�u�:a�XJ*4r�9Yj%&�'�bn8ϥ.��ĴKa�{���X����,��W�yݯK����J��R�K��2��BO����Y���Q:���+����_�[�m�FA�{��ş<{�_��ޡ�>�KH�R�@h�Qb1�EX�����k��ʊ䋲�1�~~k��j���Q�F��EU�҃�eY���s�w����d�����l�|؅�r#�(a�y�(�/	̉��/��zc����_v���|�5����1,,-�Jz���(�
�5���q��S���Gx��48x�7p��=T�g��Ώ��G[/��;B?*�y������կ!sudai��@c"� |s�&�77������S��D&s�|p�Q�����"���0�i�]�:A��0�v����%gn߹��[74��>��O?�/>�f>�)˖���	��Q\nsǎWe�i�+����M�%">O�^�Ad1�(KC#⡂�*���� ���Q)�O#�F"t2H�1G�41��߸��}�_�\��t4ċ'�� �Za�N��"Q7ǎ`,��p��iI�P)�o��G�p�\)]��z���I��NGup���Y_�n�zP5M��$N�gFãL��)��(da>�����ƥMcbs�..��7���w^����w%��3<|���?�v~'���0GUk�1=>�v�^�.���xnǌH�E>�N��rw�,í[w�ͯ~�����o\���w�}���p0�ݗ�T�V~�/㛯��W�]���?}����\��wn��xCꚛT~e$z,wR��v������&>{�[g=T'�1=�,����n,ߔ���/�����|�����Ot����;�o���5TÊ�27yi�����:���c<�B��OO����5̎�HZa}}M�����H{B������,�Z W��]'�D��C)���x��)�x������������>~����?�Ѡ'�R�����ƨ��+K�R��*���>�'aJ��]E�Ϲ�K�7�'���Z|��wt��YO���F����t�ũ.�0�h��DU�.�K����.M"�n!�.��e�t�*�Q.�_>�B�#_�u���G���a��YJ�ؖ�cnn퉎�_F�q��TE@�u+��c��v�m��T���wc�%�R�{�s:\��>2�,��*��Ca8N�4�JDc�Ǉ���r���^�� ��ߙ��������?�y��&��ȉyʪ���&�6��=���������Ǉx��'8����̔�?�dG'YP�V�fi�A�/��i�ab���v��C6�Nz��
��b�@�>7�	���J[��h4[�+�n����_�\Uc������
)�8=>������_}k�{���#|����/}I@�Uq�;·�]�_{�ճbÀ�	A�Q*"�!u��Ғl�Ψ6�RV�'��	��u�y�c8�X�?�	=�\rzA�f�T�2��� 3�qܽuoܻ�z�"*c{'��@[��e��۷�`��u�[�{x��g�����vѥ��%dk��격�l���w���h��r��[��"�&���*�"���Ar����t���I���9�*ǖbh߉�F9t?�m��\�����rkY������;[�/o��cY�_���s~�s�ꜧ{�gv�R䊂iB�HÐ2$Ң(C@����+ئeS /ŰK���ι����bW�^��8����K�6�U��zu߽���s>'���&��.#zflP$�"��!�6�"�L��u��j�O�Kt&��h:��K�es�Z+�.-	+%I��<��ӧ�Q�͝��M �	���� R�r���E���¹�8s��{��O��l����U��'?Lgk����2��'�	Q2%���_n�Z���2�ss ;���<��s�"|���;s^���{;���WX;�A�Z�S�}!�WO�U�D9�ƣ�����������8���qD�d�r%�A��U9U$D���B�����&�w���t� �;��edd���'�����󧂌9-1�fx`gO����,N�$y�7V�ƽ������m��nbsw��2C�`};��X�i��c�^L�(dt=��BFA��Ē}[�&Q�����k���:59#�H,���[���-��P�dh�	�_��]3!M���m�7�AL]S��ߍ<ኚ�N�t�ku�M#���ʲ�+�aC
�QS�!Q�ϓ��0���lh���#���֎X�6~�JM���][;�7�OS�L���Ҩo�1+���zk�C!s�C���ֶ�w��E���y���8qb�DDA|������җ[$M:��:��Dc�Fԇ�'f��\w����+�0}�e�䒪�侪��W����&�jvwD���Ӊ���y�����Ww�_��k����j7]e��:���khu�s�.7E4���1=8�S���K��I���"�v��79wht��#
�%ȋώ�'a|,�v\�XkT�n��iw����3��o��EN9:5	�_ ,8�A��6X��_���I�t�B:�b��R���w;W�_�#��t��C实XX��'��"��m.�u.�2�[����������fL�*�4�ov�wֻ��<�	_X���R�wo�ŋg
�p�!&B�B��P�d���c(�f���A�`�$pSn5q�����8J�9Ұ��q`;}�;����+�V�bp�A��ӱ;Er�G����Bh�d���R�,x�2�0=���_K�df�y2Y�ƎٰO�3L� '�b��KZe�)]ˮ=:�`$!��\~��E1��������T�����"Ѱ��:�CG2�~켻�%1>:�X$����+j45]7jU�\��͇�����6窀;fD_P��B���qŊA�%a4j	��F���LV����!��N�<��'`��ID"9A���l��ǟ�X��F��� F��Ba��7٣$%c2���[�*��70`d/�Q�юɉi\9}W.��BO����s��m#K�%��M���Ϝ�;'Oc����#᧋pp���A�s�,�F�eցvC�8C�o8�9��͹�G�>NiҶ�h�#�皍���Óh����Wx����Y�#� �Ο8���Y��^��%���'$�$$V�ɖH�\�\�rUu��à�J�8���=,��� ã��#*М�ɂ����M�)�))Y!y�Huۇ��e������/���.���s]W p��r���D�{���ޚ�y��Lk¢D3$i�š�/i]B���? �\6+�U!�G&�F�J�AB�\��0Ƀ�Y_��u����;_Ci�q�=�"��ςd~h��A譜m��ș�e�,k�[3Cuh�T<ɴ�y#�]u�~�L��u�s��ldx}�=��'��8�/��p�AᗫW�����&q������R ̀�r���h�o�C㕴�i2���C��V����V˫+X��p cã2�3�3~����^��w������g~�Qs� �X�(~n��yh9�M5O�����$�F�џ��R�a��sl���C��͉�9N
"n��P��:8����ߓD"���E�[���%x��ۤY��M���M�i����&঱��`H���ju�k����1���o�!���b��ۇ@$��?�cs�H���/>C0���y���#�0��w����ldS(��"�IX&!$���a�}����9�E�^|x�
./,`,�@�p�����z��ƣ	��c~|3��z�����lEӮR����l���#<{�
�٬����D;�C�|p�_`��l{GP=�G��0���`�+���0e�*ʘ+82
I��Ml�Y��40+B�&=�����{�IL��oeKdf�h�l�	��.��q�ǯ��!�=��l�����g�H�>�����`�l;�rP7^��Q�4d�879���1M"�Bmժ���i
#�6궝�ϰ��N;��6*|J�.�~���L������Ôdv��_����~�I^������^�����66���F077���i�xѓA�}?2��_oয়�DIJ|Nȩ`H
�\ȝF<y?'���8b ���-�l���{ldO��Ջ��5�I���74)��M�4~����qe�$��QH�����{x[{k89?��ΟW&Q�.�������C�6�ҕ2�D�B!4�Ad�Մ����I�k�מ��ۚT�~���&��"񇥇���n�,����(I��a��}�u��&����T."�:���m&{�k0�s�͸��P�(b$�xz�
���B^v�l��>���C(���f;��Bٸ�p���O=�ܦ���F�b�\^(`�V�n�T���9��"������i��w�8���KX^^F�莟{Ә^�����[Y��&q�E�"kYzZ��l1����B�,�q>Z�o�WƮي'�&ӷ!h�N3	�D�>�&�k}pp��i�B�:��O�8���7�#�����sq�I�Vʨm	]%:����	8�HH�P���$�	��O�e5��dz���QN��:V�^ck�)b���ȟ��ƌ?��-�����ɻ�k�t#���{��'�%у�Z��y!xஶP�ˠ����8..�cvr�p �\�˯���9r�i��O�bz|B�vn�"��#u0��}�'���с�UC�^�$,Iu�F�e�	$}�A�٩�W3�mf��	��n�����XY]��������S�0����x��)H��o ��U{��t���?��X��g����9�gw�Ƴ�+X�$�",���6Yd ��b��&�^h��� �6�.>�t	�0�L"{��;wo�ٳ������1>0��pjz�������I��b��d�q����=<_]�Q�����}�ҟ*d�ŭ�����J��2��-i��lm,��h�lHÿM���ے�y�s�w��z݀�����z�r̴*I���룍�Q���#�C3iX���wg����ʼֹ�a���0��+��}eVW�����E���SSS�����+��!����4�Ƈuؒ_�]p��Ӫ��'>�o�ږ��N�����|A�Ʊyk5�b߯,�as{G��p�_'���: �.�;�4_�l������=C�*���!��"S�`}k_}���"����h��%�;1:������)�`! "Rn5`�zU��u�{]�����sp�8��Γ���w2i���r}�(>8wg�1C8����{7q���X{�����˗U���gS�<��ӻ���歋Z���l�<6'Z� Z6��8��$z��D-����'q��-��F�E����L��!%���{D�D���ޤ��T>��l�`�pDB�É5����{��Hd
S�؆�f���֚�W,`,��.�h��$w�$��s?;9��xRF���
}���Ѵ�P*DCl�X�Y���U�U��d�U���%ɈiWl�H d�4��y��Ǧ�>_73�9���'?�	n޼�X"�P$"�!:��$�,3����h2H���lk��oMÆt��,����4,5��G	�$_��=��V�nH��U��eul��8>J����X_ٌ�ę3�;�C"U�������U���l~]���J�g$B�5Wc[���g�j�ᇃj_4���=�	@�� �o>���kZG�Y�����=�o�\'���f���/~g9w��͚7G�Ntv��n�զ��M�d
���͟�œs87=�T��c��"�ص��9���̌���LV0;���A�%��MD�:Ъs\��S���6hdnP�V$'Bj�4��v�t�B���1���x��	�8F�Ş��j(�JXz��K	�P�q�"����:�(�g#�rav��B_߿��/�a�pu&��\�G�a��$�D��JeGeh�w��2��A\;y�9�ف>�l���;x��)\~�:װ/$����w0;2�����&%"D�~8|.��up�}�{�    IDAT(ʘ���k�ULLN�l�����1n?��[�+1�جi��̆�Fv1	
|�5�������єOPÇȰ���a��Ci˄���%1�tBS��H#LZq{��2�M��L����m����b$����~��������q��+'�m��&���Q�:���Y8&FF�)�V+��(�e3���D���}6zf�d�I�[��6��\_��bm}�;j����Յ������I ��(Ei��Ζ^�4D��{51u��n���"[�akg_|���,�n�X�V_@��;|f]�*��x�{x$�]�ْ�_*�G�����8�����_WN���.n=}��4��y��l�z�1|��%\���XO/Y��q�ܸ�6��qrfJ����B���<���6e<.�ЩZ��խ-l��b/W@��؈��N�>���q��,�,���GX|��}�$��&�QJ���E�ɏ�j�Fn��P ��"WW��qx���2���u-��������F���+��h!�W������u�=Ṣ尡Ԭ�P�
�f�8�cJ�(�@�P��ξ��'��Hz�v��6:l�>��Ľ59���DdDRe�8:��ޮ\�(��j�
�T*��C��v�
K&����#|��������3��(�F:�%I��_K,s3�����-�٘b߆����W��V�v���X��7֘&J(�����Y�0�~�3��*	���k�C}r8;J��!I��gV@�S�U;��NN��:��^������g��ܔ̍מ�M�\���-�$�+���������
V77�p�0:2������w��s.���(������;�����7ocG T��Fz��Pi��B#S@�P�ɉq|p��?��|�/��au�%��>JI�l�	Ny��p� �r��Z���D���H�#���h��M��:��n7�s�o0r	����	C�:����r�;�XZYų�/�G��A,���p��5u���O���a�3p�K�'����N�{�ȕr����ѯ��e�첣D�:3�U���ՀqHP1����lq��<��Ϟ��� R{[�{��>{"ؐ���7�]��3�G��Jl.�'H&���<���n{âps��&��14:�p$����<����a�\@�ӐIm
��ܖ���ʌ{sɦS:�nG�0�j�	_Qr��I:E�=�-�=mHF�.�F�I�v��0%YѦY�����F�;�FKE���$~��{2�	���g�H��$"�I�x?���A��LI��ɂ�!�ߏ��AL�%�pr/K�C3Mt�<R������X����s ��0N������HA�x�xB�C�3I^����{�jU����t����`o���y �b��2v�v�駟jj�K8=��7��gWr�c���#�bp`;[x���RAQ��BV����Q\?w������	y������%�ڐHW��.^���Y����u�n��
�k/prv�/��﹓T]���4LIht�Q�T�cWc�x��v��v�%19=��/bzv.�/V����GXz�LM��P��$���196#��p�/��O��u��\�� �"�v��~!"s����B6����Yl4c`�S,�X0�=8In��yҔC$<�M�q7u�k�B<>��Ԡ&���d���/-8W!|_�7�i��u��,2$���Y�K��Ѓ 
h�LBٳϱwt�ׯg��B��X,iB2><��x_P��'?�_}�b�p47�]3���DM����Q�f��G���5���o,)�9�=Z�5%[EX�im�ߵ�0�iC�f�y(E)eȔ���eQl�������~I%�T�~�ѝ����P��!G�����sC��J�"�bq�	^�|!�U���"�e��jM�	ዄ��olmaswG����؏G���/��s�����G�Ϟ?�'/�F�w�?��X Z0m�F���(!���kWqfa�\Nę�WK8::���R�G�u=K53g$���[�$���� �b���岌�q4��4��c�pfWLU9;�bg�f�6�+2��S�������\��&���M����M�x�.�������s��$�M������^�r��˶z�ʶ�v柒hd�o2���fː�0d[Y�v�!��U�����S���s�����ܻ�i�ߛ�� a�J'��0?>%�jfQo��i:�5�P���:���R��R�NΟ���(��R�n=���O�a��U^+�Q��b�!��6��5=8ڷ���,dS�[���V�,��?�C2;P�l�?o��v�F���%k2�ŀ���`,��!f&����D)և�cS���?�X$
w����Ed�S(V�Fl^���b�����%��u�X�����F���-nw�h7ʰs�ީˍL��lN�~�ƥ�[mJ%2�*�$f9�>ll����k������%���4]�ϟ��sg�JF$�dF����0�"��4����d�����O�Sk�Fc�&�9sJ����Ɔ�}o��GK+˸}��`�|��\���kbl�.���>����Ζ��$f�k�\v%����х+�0;��d�v�������`kw'f���3��w�]Ly�q�����q�S|�g�˸�dK[ȔF{p��i\��N�>-r%u�O�<�J��9����L���v�܋�I��S�t��6p\(��M��b����*�Ʀ�R�X[��������z�1D�>%Gѿ��?�=j�L�����u�<{�3�k����c ֣�.'a6{t�Q��$5�d8g����T����Tc�{��)Mx�a��<�e�C=k�Pv�Kś�!��C}CH��j�y_��/p��MaN�(� CC�OR���{{�U^���5Q,Cl�U~�`}����l��_U�ߞ�%%2�_�Φ�4�&�_&���Y���p1�O��'���O�ŷP�%��rjV�ŢS�9�s�����ava^H��۷��|Qk*!ᰮ5�
>�ܭ��H�?��
H�N	(���������Ͻ��_�n�/�����o4��,HJi���0�@��U�p��2��~������
�^.-by�!t�?���1|67
ق.2!5��z35�<n���'��&\�v�U˩�y�F j�� �ł�>��F��R��r�%;�T:�6�Ǒ8�C���L��X^]!��AxL
.�[�ھD��877��7�l%����s<�X����Ƞy�������e������I{�B�f�9�/���-��Í۷���C#0�p��[����	�ZTR�CG'�ب��DPnV��z+�;8�eQ��EV;s�;��������-ls��9�$�Jt{�n�.4���/�/����[�HN�v�|���7�td����<_��X�,o���ьx�K�a32������U;��F�}�09��~�=�&zhv������!2�,r�V�@�і�s�oP��I
��k6>6���D"Y�v[�kEc�kմv����@�Nc����Q������˕�7��-m��?�'�����ށ�#|B]����-@�Z�6>0���1�\�"����v�j�o���/������wo�������!�Fs%
������/�D��@�^G�P�nkhh����+V�N�?��s<_]Vf����~����b8W�ݻ�q��g079��'ψ��~�!~ 3�:��<������e<^z���jp�}"^�zUr)�)��/���x���"� ���0���a$�I��)��#�<W)�ZU�������+�tOr �O���Șo�jU���{��\�:=FOx&�X���|�7���N��k,�ϟ� ��A<;1������f���D ��{��'�l3i�$ucq�s2<8���ii�I����v��d�H6/wڌ��Y$b�ߏf<sj��͗����ۚ�XP�AŌ"e<^/k����5��_��T3X�[F�%Q����͎����{b�����l}=��K,q:����kptt�t6���u���z��Y���Þy�햌6����(�%� ��H$O�(���!l�7qm�5 ���������!�+y���~�C�E�$N����P��߿����G�G�n,��J.�[���/�"�8�f~�#�>����@_ ��x"La(�@&s��Ϟb��K�xvs�k�:r��n�T�BA�4|��z����r��$�C����QP�����0�/N�v7j�2ԡ�/-ߺ��+�]؝�g�4H L!�Ӈx$�K7�j���1��)q{�z�C=I������9D\>���7_ai{��c�m]T�v4��*"�H2AMRc;�M:��3m�+�7��kW��$<�ߧ"������Lĥ�k;TxǓ�ҟ���y��Ʃ��J��"�}0}��mH6q��Ua®��Cܸ{�<���j5�K]n��ňr��ED�R��`��q��p�Q�����wr�1��9�')����T+
MWѴ�>�)9VV4�K)�"��$[PZTi�}ft�|�L�{G���p�>�� ]����6�嚈V�N�VՃ�&����FF��ᠳQ��lE�8(��nWQ�=&_���嶡�"��*�8<~ll�J��i8�#���(�Սu�ri�)�	�&��̟w��3��*�n�"�FkF��R^r���/�w��6}���J�N.�Pq���C�r�K��/WW���&�������v�2.���߇T!����%��z���`8*�h�^�>=1��c�����je��bztT?=8���`x���� �G��٨�:x���ŕel�����H�Եk�p��E��o�ʺ�E8_������<��&�z	D���e�)�'"�
B?.�4	S�OM�Q&#k��g�bfrJ|��i=x��mBg���W$�WK��i��D�
���bT�X_�a>/�jafN�������
���G��e3r��^�֢����zi��F_O�ٴ)	Z6f�Y)8�Pq�%�J��*Y�$��P����/dB��b	�!UPo����)c�M��i3؆g��"jL��N���oEZ�ۅ�"|��!�$.��e�dV�`3e��<[Ԉ��*��oM�d~����%
�4&}ZhR2��a��&�+i�M)[���ZU�ao:&�8�#�
�*���+^��di�����.�����ɑ��<�?�������?\�����wVs��>hԂ��y��;b��^�"��@0��Ӄ��^���	������G�AH��D��q*�|� Ȁ</r�N�_#K��5,�h��B�a��N(͌Φ�>C��B��.ػ��j����:#.���e�`����y}��$z����P�Ţ"|��y������4���!L��|�ݾ���]��(2���5�dS�jNu**�y��c�(S3�.�����û��`$��7��!���"Ls���a�Ē8<���z�än�Q����,����:v��||�LN�#��`?��� ��ZI���ܝU	]Ɋ���dx�&Z3���.>�7���a$��{��Ƈ��?o��(43���X�t������Z#��)�~���j=� z�𽹓�k�g�Y��R�zIh��ڶ&t�����va�O;���!�%�#���<N���֑F�eX����@���_zw���wn���+&�;wp|Rnd+���T�!9D8���gu�q��%132��!��mM����BN���Ѿ�:$g�SGr�����DB�n�L6�o�0��,�/����E_��N���2}~�&�6V���l\6_$O^�]�I"
���ʟ<{��O�a�� cC�<����1$i+��XIb��I���6�����t�%�R���8��=�<N�8%�eusU:�G���=<w�,�G5;��È���Cއ�L�븘A�ZUZ���M짏�&q��E��=!|�Z*h5�� ��#Rb]^xY���њ�l]i��ż&�ͣ}s��j���<�&�U������sMY�^���=��t*�f�&��Y,,����FzdT�a&s��g�/�noc-S���d�H�-�r�χ�ׇF��b�(8<O��c�5��V�4r�����2eYK�,ãڒ'};�ϷIjշ��*�oO�1�*�Մl�߆��asʳ@pt./v4w�2	Qf���MDѤ�P���v�iD�f��i�A���#^F��!��P��z8!�C~��kM��Z�����WR2��k�zݲÁ�h3c�"��ϛ���������/����F5 BZ�+�"d��}��� �_�?��9 �N�ѽ�x����u@�͒�_S����A����1�RBH��6����J�4���{�<Fi��$v�>tG!w�Z�Z�jS�,u�1v��BpҎ�{z���1nt�r�Ih�T�E��|dbJ���7�\��?���2�HUJ�;-yG)W��C��nC;L���-Fk"�m�ۇ�����K����=>7���{�%��C��Ņ�S�!{/j�^(Y
@0�G�)-̎m7�����`��+4;N������?�����G�#�yx7Ʉ����>�?�ǩƄ����"QV�}�?���ɜ7!�4$�����݀��+v"&O������:kN�
<��c8�ڰS%�U�Bf��Ű$��O���D���l��O�c2E.T�9lnn`ms���ꠏ���K�{bG�*ƲQ�I�#C裵�����#H�$nd��t���Λ�o��p'�j�Q�6��t͚ҥ2�������� �}�jA��Ӆ�^6���zg&5����b89:���!�N����D�Mds9��~���-1g3�c��xo���B�d���N��BN�`w8G8�@"
_8�h"��d?�N��i���~�[G�ȓ��v���~���IYV�Gb��0f�������踈Y�Q<*_hR6��(&Z�<��*<Y~���{�����$1�7���q�G�++�߻wG׊�߅�Y��z�IEGf%�C
|�m��V[�dJ��޻$����*�g�N�MM�"�mȡ�$��X��	*��@.�����)}�a6-��y�i�[���C ��mKĂ�^����%٩҅�rBJ_tޑ?�A�c��,�bE���ǵ�0Y�<W���������mvD�I$�o(+����8��7��;Ϻ�I>��H���?[8��מ�N5��lM�yGlM��d����ǀ�͆̈́�y]eHM:�:3������m�χP$�t*��,�m�6�V�1o�	���!�V&(��X��A�?��9��'O5lp�~���1��<� ���S�f����X����=�ǏoU��?���?z�<;�����R�h�hb"�����IH� lscvp�p~n��
��ܺ�;�n�L�?94��gW�&{��5PoT��Ã�7�bn���ؼ��v>�V��3!R�y�-�N�z�AJ�BL�͗H$�`JJ0.Ȑ�Y`.�$/�7�VN��!�bzxc�/��,���}�3(4��,3��i>M�2ʙ��_�<b�*��{D�����xC��� �g��K&��n|�"L���y�V�����1�?*������Y㱳~��7�<«�רԻG�x��u�N� ���p���`3�C�e�m>�.��}�B��N�g�P�M�i�A(�+�n�G�)��oMhe��P��a�A��Ņ��܍����%��yO�}%�$H�}�K�eآ&�p}jc��v'��^�����g�8�F6_����P ,΁�h՚�u}4A	e��K!���|p�lm�ݔ��)��q`�O;�9�3��v�X�
aa�{�і�\�\�Z�9L$��E����F� !0:W�G� �J]V��6g�,�m�ۘ+݅H�r�K��>ؓN�Z,I'�{L��<d;]�P�E�{��]<���x�h�X5���.��>��|��SGx����Ҕ��4ߎ�׏���0:�~A�]��K�/�ʧ�1��w�P".���=�&�MN�V/L;��dK8��d��8��Fџ액NN�˯����C=�JI��p��$J�`L�J�(Ґ^?=߹.a�J{L�)R]�$L���N�]��9�PY��X�w    IDATe
�ˮ�+�D$
'�T���S�Tnl�^�T>�Uw���BVN��a~n (@׿�dGg�x��9�,>U3�g��ף��Z����ƁȊr�U�:�Jq�i��95��~a1aa�Z�k6�|�����W��9ck��oC<�T��*��8M[�Ħg;ˍ`,sj4s�TK�dA��$lV6y�LH��/[{�ad�s�.�\�X�˿�v��:�|Ǚ,�3]�-��9�}m$`��pre����F��+D<�X��qa1�$��Ŝ�R���g���,L/jE<Bp����݈���SM�J�͐��s��i�w�\��|S�~�۵W���������[-�m��Y���6��Lm���0�^Gb=��k873��d�l
����[7�ɥ��ux=�Vjڏ�qI'a���c�\��EǢ`���`'��V��q��fsz̬Hڳ�M�+��d>�n0��A?��z�t����FW��|$�����%�L��/����3)�ɝx���\���ǅ��pH����@�TA�����n$�e��PwH�Oǁ�'������S3�	zQ.�����D�	�H� �ϝ.�U�+�֦��s��7"�u��,����}d�U�f޻�Μ:���^T�e�����/�z�B���v5d�6y�9�	�X��d`�]���e2m���uho�C�74;GP�����4&֒��&Ꭾ	2*�V4�v��@�&P�#�`:փ�S'0� �t���)��ы'���\���T(j����!D�^E9_�^3�rc(�@2B�D$���lʫvR7ܨ
�Q��I6S�If�����P,W���\��Ad��s�N7��(�i�>�h��)������X;�:���LLa�!��n�����|���}�JIP1�D��Pw�!�]��g>Z�0��B�\B�������%�?�}Úy����.��2�*�ӂ���I|��u���J@	���Wx��6������c��xA�q�ȵ���>Q����6vw��I	��?u�N�Rq%q)�e�aoO�>��7�֎��"���ф�0�I��T��Kb�渎�M�P%7�s�SE�Ĭ�'Y�m������C�d9J�_��o0ɤ%��QJĴ�G�qI��fu���nY�Z-�?}gO���̂(n޽��o��Q>k�k�vI�t��0u�JW##������LS�}�3�{}�O<O*�l)�E�E�5��X�*ƙٛ��NXh�`d���0�6�L��T�kHy�}%Y��S�M=���aak�U��[;e� [�^����<�-��۟k��2@30��H�&&���L���l��߇hB����h/٬��s�FM�`A�����k*.H��s���'-b�d+V�|���ѾZ�R���c]�.?�G&~836�?~����C��"|��;������;��[.����CW�6�u�ޢ��HQ�����Q9֓D�Z���.��7�h�7���|������M眢�Uu��{+�o:H��Z�N�<d\r�2v�
wr����ś��D�n�D�X0,GBq:�Db���4��)��)á�:���nv�ÒӕK����/?�����j�x��z<����5�����ر�	Ӂ�%N�v橺���_�.�͡/�G9��N���(V+�$��ŉ�)�Ebހ�	��ʭ�ih�$L����k,2���(�
\n?>��Ν;���A��e�}|�ݹ�M��v����:�	���F����7�d<n�DMX�q�{q��
��e��4����O�I�>����u�V�P��3�j��f��,��dJ�,� �ͮv��'gD���9L��;�ȧS��_n� S)
�b�r�RG�f����͉�S���,�Q�7��2���0hA]71����Y��XX����(r*�J�:�����x����N�#��"����M� I4�y��EL�K���4&��亡CIDCƑΥ���c�p|��!¸:���V�(�#W=t�b�@�~>�	��`���3�|�
X:{���l`��I��ך�����)}(F��
^�z��+�d��K�c���pX��M"Bʀ5���:�QY6�$7ɺ�V��)�ӂţ��2�Y�X�5���_���f��A��'g1�7�kC���t;���m%��GOa�ze�P�U�/_��+�/��1f������v�l��L�x0�����`93JqhlT|50U-G�ITtq��y\8{ss�ܾs_޾�c|p�ⲩi���\�q*��S-,��΋�d q�ǐ��㺡]k�[vl�0�&�4%�x�����+�H��>����|��I`!!���lk0����)O;k�8���Gk�k�n���'�tɲ
.?�ϟVV�C�q&�ķ����l�m���V�ъtd���h��DX�G��YR��A67&���F�afq�5�>�ү3�Fk63��e�[,��\�L�^7��Qv��afd�?Ώ���`����w*¿�����^<����Rq.�� -�ݍF�-�W�������&��1�����&w�6�6k��?7{s��7>�܋��")X&C׃�4�խ�4�1庲�Z�c�{�3�~�E��6_0("�f��Y����t��ɋ:d��|�L��_����>�S<�XA�\B�;��XDi4�G6���x��
�G#����R��������~�+'N�/@!��g_}�[woiZ
z���%㜓���#��&7�	��8p��{|����39�J����裏ELB�^T���=l��ȵڡ�����qN���PTr�r��L�]�<E�^��E�xD�""�Y�#舐������v�FJY�41���!���f��|P�~v��azZ�����PW�f0��G��B�� �+�9�C�rtQ�]~9W�m%��*M3�94K%�I�k����m6���-���>\MJ4��Å�
��ˍV݆��kMEr��q�inS��/Cbp�^���`�-#�P>��L�b��$���c�o ~�!̗��a�e��,�������0��F�Eu��3��Ǝ�lF]��NE�-��`7�B�Y��=�i3�`��y>��r�^-ac+;�88N	a�5�'W?�j�Ұv���W�X]_ū�5I�Bv7����"���-�kj8H�a��4��6ﴔ�M�ǁ�a��.`jh����Ą2����cܼ{K�n�dG_�|M+N� ��>�.�K����|��Y�5�uDc=�����{�pU�g��z����O�N��N���+W�U/WQ-��(����V�^.��ƪ<����!���K�t�"�g�Q����R����z�[�
��1:9S�B��55R�$�rFo���,��l���Pn05��kp&&��"��Qa�M[+�x(��#
i��t���UEWiA��3`V~}+܁EXE���ZE���ZRC����M�o�`��͝�_G�=[��E����a�p�"��a���H٦/���A��"��D�:�ﳽ�Z�.K]�V&드 N���e�b�7���&ǅ���X�;�;L�,�e��0=8��������w��NE����_�ꓽ���.�N��**9%$���p����۰!�������	���5Az���4&3��T˿����C�_��{���MKH�Lh�oՍ9�p+�Q������o*�ӄC<^�������`W��Z�1#VōՄ])_`n�!�0� ����m���<{��t�m�^��IL��`btD;�j���lI:e�a���bm�3����ۿ�Kx��	�C�e�d���Ay�W�:v�I��:fd^��)aw�1!��˻���XB�c�/�'}�KW.�-&SʘfT���&�$�uZ�:3��N]�f�r2���]�w�����i��D�7!M*={	�ӭ��J���T�aa�zyĚ1�
I�d�Hq2<c	��U����AN���Cb�Ë�P�&�1��C��B��˯���>D���k����c�J%6l$2�)��
y4+e�p��%*Y��g^��%�9A�K[��H�ǖ�jN4���U#�����
L����� ڛD05���\�pG�\BYx��E�855+�O��K�ｉ 8l�U�X\z��8�t��By|z6Ԕ�e40�G��C�HĦ�Sa����������q|��{*�4�aC����r�
���g��<���1����v��$�{k�.�B4��KUI�����h$��*udD�lZv;�ՊtԴ�É�i���}&˝���ܾ�#�7�
��N��KWpn��
S(��
�|�k���.>��s�G�j��~|��G����ܹ\F�)?�����Z�eO/Ν:�3'O)�JhI����a��M��q��?y�LnYl�������2��ܼ<��?z���
}`��Uj�B�U��|mCҧ_���4Hh3&`��l�9����څ� S��p)�2�����O,�$�Y)b�|y��H��a��\j�=ɲ[P����5�J^h��&^Yd0�g{��ec�w뾵��U�4	�jMB���1y=���EC�R��5�0�y&�ĈB4v�W�|ތ���]�{�Bx�q�5�ҁj#����gW �����Y����Z` ���_F'~��h4��Ѡ|��{�������m�Ŏ��ڎfӰsw]Jb<_����.���8=9W���dy���҅��h�@�Y�˔ŏR��H��~���iɚ��b%,��];�t�}�:3ʝj4:7e1̓�r�Q 4�lxCқ�؃�#�J�5&г���X7��:�����?���{�6�8,�Q�^7Qv/j>�|N��X��?vy�"���EM�	�D�*}�)��sS0(%!��K�����a�|MCk ퟩ�#$���b+��A��|��P����\d;������8(�P��<J[Gp4�FX��0��Q�Ԓ���  �X�Vw�P����O�5����4 "�UH<�t�l`�0pU��c��Ώ�3�%�c�J["�R�i�я���T�H�|'q}��⽈�](��jm[rc3�ßMC�Bc|C��b��
=��T�Y�\v�aȤf����v�|n��i��F����>��:�tt$i���
�$�!�"�ܑ��M"��q�ݔ4�³�pz�i990������5��2�GGm$ݭ��@*���;r�fZx�X(��ĹPDE��� �f���ua��=�C���%ˡjucU��ԁ�����P,�c G�pe����]��m#ߪ(��Nf>���k,<��&#��\Q���H��{U�v�$����yL����p���`i�9��u��7u��N�����NϞ�=�:>���jT�Kv���%ܸsW�*0X,9	S��޵w�[�g�"�}�ӿ�ͧҪ<nɌ�7fx� �f[H�������6��VT�	��U='�.]����%U�A�����s��a�ATK� s2�	Ul4I65�s$��Ź��-w��/�{��IH���H ,8����%����Ȃ��x̵#������v��#����XE���3R�E�Z���#�v���lM�V���1���p��;��h6�f)S�Ôܩ8鲉��c�o8�ڠ8(�ɽL�2�+��|���LT""��|��aq��)�%4���*s���w6������z`hP��,ĩ�c����(׻�c�?:���������;ۿ�:��j�f�;TF��G�뀫�F����Sg�хK�8=!���S��rV���F[!�,�
q�/�
ܑ4�&����إ���b p"Q!6S8X�Œ3�3��Go�A`W�}a!������WU�s)��3"rm�Y�)��Cwpt���!S�i�\���q�,-f�٢$��m��b@����jf�%i�L��6�9�$|ea^E�\���/���|-b��X�0���u���K�&�xvd��u����vSY�+-�z�����ŋ�10<���~z��xtG܏:�:eX��$J<|mH�6�_��_KP''B\�ܻ��F]�C�,�<p�X�0���U�n\=���p�%��d6�?��k��_5X�>��\�Ȋ�5��1N���<&"I$�^�JE��-�5���`O����[�jؘ�C��;���1rGG����H{1�����E���aA���;J�IA31��a���a$��M��K:�L��IȺ7���>ɱx�0�!J��k�u�m��o��L)��K�G��l���>lPy��ǚ~���R����d2"+ٺ��&z1�;�O��@�?�a��
�Sک�>'s����Ѥ��4m!\����M�|v5�$.Ҥ�h��M3�d���q>W4�B^�" �ɯ����t5�3�3Ss�E�A��vv��=}��ɃM�S8�,�G&՜�����ޤ
&�S�<Ք�_<�����^���r1�Q����s�@/�#�^�,қ��f1|������%�}�H�q�#<SX��\���s:;��x�;�i�R_�4�T�'�KX��u�H�H@b�<Y�x�$T�2��|]\V(��Y7��}AT�5A4�%%�"�,��b%!}[�y�򹳊0��6S���`r8��(
b!��IR��"l�����k�'n��ZßM�-��3�����bN��J;b̽�x?"R��x��5�	5�n�Q���dR�H��x�2zac���q��.�u�s��ZC2?��h".N8&<q�Qȕ��􇃉�?|wd�[k��0�~�I�'�����[�|#w�n�Ӓ3TU:1c����~�D:N��p
�=��'O;]��V�>!�z��5�+P�VC�)���E�4Ӡ����C�alH��^4ª���Bl	��}o��J"����euy�E%[!{TZ���I����C���E�׋��1���
U���<X\_������J��kgG�)�{(2u9��X\�t��GV���pin�QƮ���W?ŗ7��*IXAB�}�����t&ep�>̈́j���n�erX�����]�����ǿ�ӧ΢o�{�����U��K�]v�����d!e��:`�S�3L�a�*�"�l0n<���;(v�.�Sz]�X�Z.��`:oq�ַ�0��$A��<GSJj(	!���7��֛m��-��q\[�T�I�UK�K`?�B�UW:���LCm��c��ݝj���Fl`�����
�R�J��&7vϼ�x�1Ӕ.qDX��jZ�Os"M(���Ԝ����G��ӭ�W�D� ��<x�hL)��zY;,�i�%�l�b}�.Pi9o��P;��e5q��CT��U��˘����ب]t��tJ����T�����`��s�����u�=��3ҁ�7�#�涺���[X�]G���z	�6�-Ʉܡ�n�����C!eLy����*ַ�`102��!��OM�`~t!;�J�8:>ĽG�p����i����?�~��pB�U�YA.��K� ��/����?�'@3�t��P�����<���Y�n}�
�>l��)����+X��Wc�=2ܚhKJ�BN�7���7�d�j��W�j/|jnA���Ǹu�.^������i�^��k�����#�����|ٍ�-Y�
����-�6��:Di�"�~��N5W�=��6�N�;bL��$�{�g%�o��b��$Zu��i2��-����A?�A����-k�2c\��.���F(���%��v�a�	S���HY$U�vt,�cG!�.8�ߢ��~Š�th`@M����.qL�$��V_ڽk�wkh�3ĉ�X���� s����r(U���w#��ui��N�_���|�to���gS�st���?m�Ȥ��%U"�o��8���	|x�<�=u
�j	�r�J^)Itw"���"lZJ�Fv'�$a�h��W%R��&���Mk˺�Ī־����n��@�!��t��%]���1�-��V�����PO�)�Suj��&#�D���Y9���9l�-Қp�W_���
��4��� u�M�I�G)! o���FWy�����f��Q-೯�/���|���8]�alY�(�JSx��Y�]+�/�4�r�"�rkÓ��G�����	o�ᳯ�"�[ʣ�.���[���CKRd�F�,��w�)��pic��<��yݜ$gթۣe%��1��Xl�h�9Y�4�l�_���Jx�p:�.��]x�%"ְ7��͟�
�*o    IDATL�_�'�f�jU2�6���`��$c�a��E�R#W@�({��b!�)���+���#�L	3t�����t�+�;i9I>#[��T�!���HD?�$&tgl5� �5��t����&E�"feCE�ו��ˍe�ln�(��M%s�iSɤ$��e��UQ�}YF8cҊ��&�*�I �ۏx(��� >~�}�d����ʨP�S��	�#�	��c:�֗�����\�O���x�i�5���K%d�%���q��3X�Tɸ��.�"#6��J`a|
'ǧp��9<���W���=5N^{_E�7��r�cL`ux�������cx#A�1�n���㓏>VLa.����
>��΀׏��5LOL���8���3�^��|���y�fÝ��q��#5*�rA����%���I��ݻ�bͤ5�.�&*��Z���0�@�O]A_���"��\�/y6Rnǟ��l^��ݨ�p���r�d@��Ģ��������Lm�i����pb�&׷W'��^���J��CW6���]��o���?��|+�ؘ����=_��������5X� q��c��谆�x"&��b�w�Np�ͦ�h���^C����gQ���F"2Ҹ�^�70��&#�.��2�ޱ�ٳݑ����!�����"���~#s�;~|�I���ዝ���9�^����E���eC�ޅ�넳֖����i|r�.,��V-���+��m*�ّ6��J��Z��cq���I��)�R�اƔ��;�F��ZS�6�ʕ\��0F�E��{�H�$Q�W(Q���UB>���,�ˬ��l!�(8p�~�����PmTD��!��q�h�v��|�j����vUx���g��]M'�o���I���;�MeUe�,�}w��ތ0 �K͒�\,�%�����}�.A�+�(B/z�YJ A� ��i�m��.o�\Vf���s~y{��^�0lDǠ��dݼ��}���i�W�w>�'��FgS=2�8�ݾ���/akkCl��C��in��%�Ѯ��$�G3Y�<�����Y�@4K���}#�=<�"��ނ��Y�u\�wk�$�t��^Q�p�^%�2%`.��/����fu�l`dʝ\<���)�#?��0��q$JX_G�*�\�02Ȃk�\ZS �,*V�����5t:#�3���Q��F����5AIɸ'罐,g�y�ǆ�M��$�<��_F2��B*��;�;"��@�`�w@>�DL���-���Zu8q��R$g�X��C�6P���:�y�4m�r���5� ��fe����bU^/vb	wv�uM���c�4��}���y�E#B#<Լ��
���6Ԉ�P�� tOc�}�뽴���%�l��.:kB���Y8)Qډ*'�Q}��+��F����&�6f�N�ɳ'X�XB}sBM-���ҽ����ڊ�Y �U~xh�C�i��ױ������S���`���{�w�V��"g������[k�8�� �ޏj��a��1����@_�����,�<}��/_���b)��s���O?����w�фɿ�rY��T"F�1&���ǘ���z�t�A��r� ~���h6����3���n����Ҍx�Y�?�65<�/�)p~��)˫�tG�k�k+~��7���no��O��<2�<d�Ƥ&	��#�����IU��j��L�Gb'�?Wc�c�Ĭ�������LϦК�p��cl�I\i*x���P��f�i`�wV����oѬ�$�Y������'��\Y	K���,-x�H��#@Cc�d���W&��;�2��Z��ZW������O���j��2��
	��.S2��"�#.1�nq;�4�W��o��s==߾N��U���b&>�,��DYĻ��_��HC[��_<|Gv�������x���槐/�e�(�V������� v�q��T@%/��&2���0��J�!��=����.C�1M�5�Z�BWO'����&�5sy�-1�N?�\����v�y�qh���+�]�'\D(X�d*��3S�g�H�XO�0��JlKE�@;~,��s��괹PH����}�!��Ewk3��$�޺��/)�	'JiF:{�V]�I��d�V2R%c�FI���*��$��A�k������������$|��m|y�:V�	�]� |�]7w���Я��T�������V�$��u�(��� u�pE꠆�PN�K[F��g��gқZPw�$��d���,Iif`S$��r�j����݇p�w�M�
�s) ���"rB3J�hd��p���T@�1�y��w��3s���)�S̢`sʤ!PU�F�R;>��B��$#���^�K�����9ְ!��mmi��يBlx��S��,R\����������m�[*�'��0^��ֺѾ�H&I	4�	�ֈ���"�c��C�
����6V_�j��ih��Ϋ`m���5�	m�c�g�=0�û�ʿ�Ex��ܾw�?Bm�mݝ��R�G�Sj��!{�6��LN�3��zxۛ��nDWk;B�������յ��-�����!���v]�v4��#ˠ�͠>X��()����􃞞�����N
�ĎX��!>�$L�d;�7o&��_��B������Fs�Z�u�0�Ю��ZF����	��?����s� ���c��A��'t����_he��Bcs��:��`�Y����|rf���%�r(��t�g���!��ʬl�Z���/N�SS3�wq��������
q��$�O�
���NZՂ���Z���ϭ�xX_˚�9	[֘�ױ>��ޑg�cQ��X;ʦ1��0Wz6�ET" �F��af����w��	v���ʋ�ë*�lny�)�02E>mEi|�".�e��$�o$�V����Q��{T�P�Xq��Bl����zo�g�D��������m���l������뿾�rm�/�"k�X�3("c�}u�t��ܰ�:=��7���á�!�q�x� �����M'ڄ	�pRp��R�P�ޔ��������	��/�;Im�m�$��P�u8Q��b�7�dJIv�݃��!��5c���8�r���h�����N.�9a�-��aڧ�����.�jMDp��=��c$�y���X�cɸ&q�l(��^ټ����N�c9��j�{~������%dp��������B}�hW/�j�h�W�X�2wMO2�(��Rī���oh��S8|�7i���:n޻�"���Q�^�E�Xj"�0��irJ�ǳ�K�P���V�06'j>[�G��ݾ�]�3&2D�A�'�r�t���������g[ŞE�X�~���|"�������>��wA@�zO�;f��4��Z�{���/�I)Pڸ��nC.�B>�BA�C�4x�l�mm���ַw�=Ї��N�ܷQ�K�biqQ��'���A��C�82�����5�1�0I��嵍'v0?�|a�4H��?������*�t�ٷG�^�mM�Kd�W'�*��I���-]�5�	����'�JX\X�y��Iaav��B�At�7��O�O�
��-\�qEZ����Z,rgvptT{���AyG�ݿ��7�bbn
�Z��w���f4u���fd����.M?k������9�C��^0P��@C�}��.|#����9�r����I�_KMH��ɍ8jk��hC�e��<{����DCk3�ڟSj������y�&�hb?��/�@���*^�����Cq��L�((Q����޺!k��yJ�_�����,�/�kmn66�Du\��Q%��YliC( �q��$	����z�Ɗ�f�$�Ɩ�3�w����炎��㝕l�FI�Йd2m���
�1��M�u�깤Y�e\Qi�Ɋ4��}_��3YN����� �߳ɔi�;�,�C�^�0U%JR�Pz_�0����!|���+���v`cc3s�X^^��м&;"[[���|��I�����`�_D��<��5
m T���Lź�&��A�*�RI.]���Y�U~@}cÕ���?�N���oRO���͊���������0Y;���H�"����9��n ����E��#GppxȦ�z|O����k�>��eH�h�i��<�+"e�@t��i�}*/��ܬ"��Q\��Ig�+�d"�n���;4��F��g�(z���<�b�RV_W�`u@�;��	�&�y
lgRX�Dp��S톺 ~�{���&���._��o^j:ɹl2�H1�d[W&<��t��E��
�b"O���ۻ��9߸sUE�7�5�ܗ�VQO�:����y9gqJ#��e�zWcq$��H;w5�Fp��1��Fxk7��¥;71� CV�s��0_�Յk�$�IC��b��I6!t�����e�W���,u���eqbQh��A�L�lZF�**L�!�~�2�0�8N�>����$�I$��tf�Q�;tGw�Q��ӗ海�_\@6_�ٳg1�;���F��{����9m��f�)����{��k\�{�H��C�5*�bN��TRi`/_����I�tu���C����Z�}��%1�z�=��_Q/ʟwl쉮'���aM�<�_����#y��KI�Ǳ��2�XZ��L����=�5�R�}�bȍ����T���-bmy�^�3ہ���~���jAl��ܐk����$/d�ٻN�Ɓ��j�޼�k7����Ե4�+A2[cKzG��>�$0a�a<܂�Ɲ�ρ&�(�0���OӤ��F,��Ҭ�0�#F�-�Σ��#�}�e�z��B�|*�<�)z�f�[Ե4cms��r�c�x���m��,�������0hˉ��eO_:��QW�D����MAx���ǃO�^��U��ӭ(���V�<3��LoiiBs�IIW|؈J%@�?��Jx=_;�}q`�&�7ߑ�7�J6�a��DKX�9�Q
)F*�˗��ڵkF#� ���'��J^�/�k2�"�ZE��U�M�66�V~gl8�n6��76�F�oκw��{9�jB*���]F�P�RI�<��Ta�GC���?��
����������4����s��]N�2��gC#�[;��֮a��$��,�o"Il"
��dTzH�Y�����Ư��Æٕe̬,bm{MM͗;:���;-�E�?|���re���׏f�L�h ܗP��/���E�9���?�����Q8���Wc�w�&ތ�Qɮ8T۬,͎�v]���-��ÈF��@�;}N{X>��}���>����d�0/�Nn�a�f"��a�o@T��eu�G����VW��� �A}CP����);�L�l���]C<�7S�*������wT�c�|��_`l�)ޮ, ﴡ�q#+b�u7f�B{M#0EEEXl_�v¿��G`��h� �����ʗ����*�-�Z�,�9]��$�9#D�z'��R$�7+��L���Y��	�;{{��b#��kwoૻ7��#��p��&a��<pޱ�y#��D��YYv�4��Ή���Մ�"?�0�y�r'Z�T��I^dYw57����L[�m,��be}M�?�6���M���c�˽~�Qc��39�����Gpj�4������꛷nau}U�O>������0�9%+�tO�@���b�_� �����FD��C�ȡ�z/���q��<:���y��=�3g��ȡChmn�K�$d>܃����ž�0f�,��k�n�Hq
c�������ך��C>�g�8��kx��^�v*.��������שqY�XG�,��,������TL���x���¿����wqm��a���,-�9⾔������߽��"xp��}Ϧ^���]�=X�l�d�|��|(�ɚ]�<h	�S�KXPNM+�jO�{�e�J��3
Y�]j��=A{�Y�-���[wY��,�1Mv���E4��bm{[E�D������3�����W�����O��ӻ���#����ӧh;�թ�Hl�m�\��8�M({�Bo���w<��/�f���WV���k�)���	o�g���&�F%��
Ɍ��	��!�ǲ7tQ*�f�C�VrXT.]���W��\�i�d:���9U��i@�,p���YŖ��w��~a5���sXE�TS���l��a�[E��iYlhc>���+s�����n,�F��F�p������3�����Uli�4;;�fju�!�fsJ�"B
5���C�����˗0�8�!���FA���U1f�����J�p(:m����m���~���oη��)J|������Ĭ���^�$�"L֦�y�Z��[��z�OE��8::
g>�������}�̾�^�����[���^�	I�b����ے.�݇�~�����z��5u�|C�$�q��ʦŪd���)�ɠ��I�e����p��)M�4`����B��rϢ��2���tYN�>B����!t���}�5u��#��?��O�0D��Y�ܱ���tv�n���h�b�fFoځ:��s����[Q.fT�/_�Z�!z��>�������o�о��8������ە5,mn#O���ԉ3�p���c�yS���U��XW�-8Zt
�S�>�?@�Xsh�Zf�_��~..*1?F�F���w{�&	6Y�w�b��R�B~�٬�3��1(�Nd[��҈�u�@��f�"t�Ke'����v����8�:��0��5ݻ���5�Q#�u���@��4��oU�31�zp6M��ܥ{w�卫��S2j8��0>8~�K΍[70��gg��=|��GO�a�V\�l6If��j,��Ng��"�.߽�l�(��ĉ����<}�B�luC�w�)a�F�6�f��ܧ��7;��ɤ~v>#,z�E�!���1<73���Z��Ceg��7;����!B�$}t���9*����7p��5��y���.�4�u0�ʇBI��V��� O�S��*��0��nG��^;���^x�.��Q�ќ��d������sT����
�.9ȕ2B(_>y�B�0�Am]�G�D�jo�ƹs�p��1�UT�'^����sl��ERTw��~�A��h�A�@&�֮1�u��6�;u�#��N����{hH����e���7!?���]`���l)����ѡ����&�I�/,(7ziuE׎�3md�>��0tSS˻"�B��W_�ʕ+j���-��U(�/���W���d2{�"gY�0W1�C��^�
���hm�������L����U�0�����X�9l����ȳ�?�-�t���h@�D���Z��F:gHb��i�&��#���=�KkH�˗/+&�r+"d"��7��*���*P���6����`��LH��󶣽��]���L���MQ�E�O_�����,����kg飒�qZ��lQi��9}8�?��O����! ��ċ�>���ya���=������]"//aB-ܵ�c����/e7�_�{����E�䏕��dV��7��� �̿��;u�؇��&����	kj�o۱muQ�(����]lk+��5)���I��g"�ƕ_���1L.��q*�r�r�"��a�I:�y����儇$�x�7~x��>����J��q�2.]����%�׸���7`\�<>Y��h�M8�����1����Vװ���H,��
'����s&�!UL�����1�i�h�|*�$�)Ɉ��^X�XA�"+�4,/4��&����I�D(hlA���M�<��Ł]{��S��(_u'��|8��o'�|�\�b$P�P�|�{�F�߯�-hzi��ܑ�p訂B^?��۷���3u�]"޵�Z1<0(a:jo+��`r��p*�Ć��7�����؊%���wX��˩����������##J�RCGS��!��#\m�����#���10�����'N
����i#I
�;*εȦA4� �M	_{&���ʊ:vA����
�
@novY��a���n�6>�H�*v��+��\��[#E8{���ŉ����S�߇c�|��i
�W�Đ���2��4��p:�a�or<���QSP��N��}]=r��c��4�d3i�Y���L�P����z�~z2�Rtg/_����"���	:�    IDATܸV�6�������=u'�FCm-�-LL��/��\��a�0�M��FƼƴ�d��fӈ� D@��*��[�f*��a��Z�C���R��}eu��&R�t����tV^��HT4clX����ʤ'���������c�/�o|ml��9���>�`2�Y�	E߼ySn|"R���6��pMƿg��ݚ���ʓ,�NH�&�o�U|�~�/�m����mlg��c�%"�Ju`^�
�<��@��庆��Z��Q�ْ�ΜDgw<^��.�6����ׇdW[)Q,�l����hm�R���;�n� Ygk�����PUS+�sW��{Ss�[Z�������֞��7l.�o��7�	���O�=/�xzc�c�M'�^����m��[2��J�x�0�3>,���'�0��!��}da�و���G$/v)�H�ry��Oeae�ʯ~�+1 �f9z��U�0�0/��$'h�@7�6��B:�����#���C8���/��X	���d��l�\u���uj�ƽ&��?���G[}��|}�<z�XK��m��.U�J�@�(�KM�ׂli���pUف\��sGa���l
Wo|���\��FX;�Pu5N�=���.4Q�O���,�M��r*f�'����6"q��=uF��辽�Ғ@�O�o��"L�'�0eg2�O��t�F^ci���f�-�Ĥ��׉�DN��]�5�)��Cسk�",�v���;����ثqL,�c#�c�O#��tŇ�t�v�w0���#�x�8z��0�d�n���5�k��f&�n��O�jkk3|U���`�afs�x8��3�"ۭ�oi?t��1\<A�fv���ܽ�ɉ7h��oatx�=��L\�k�"�Ѫ��a�߹U�K%0���{o_˻���ǙӧQ��J=1���}��pfmg��!���D*e`~:�2�����bi��p�Ю�b�ǆB0[��C���C�lʲ���y!�"R�a��h�I�2���>,��
�z�4#�@J�8ue%'��hnihe�C#��!�C��,���9m҆�f0mM͒��m�b��[�KE%��PNt�0�9�׉,H�J+���jyu+kX\Y����4斸��m�C���P�I���~��߫{mt�wb�޽��)��\ES�]�;���&m.�,����%llG�{q��q���`����&��$x��%�8dg��!��ؓ���UC�g������1E�M�@�Ը�$�^]M��4U��1���5d(c~cbEm�w��m���?�ZEٜ[�a�����tK2�#�\-�8���p��C������CYMV� ���7�M�^l�H04�m��&npx �u��n9ʏ�
izS�|�Ue3�u�������ud}�TM���
ei�YCFGGU���&�ʯ����9T˴������������OQ������'�s�qr}��wJE$Jyd���εÖc�!��M� �tt��#�e_�L/��	*d������V����G7G���@�l#c��KcC�ҼQ9	��z���s؈D���Юau@��yA���WI�N3��67�����Jxe�o�j�`A%bymi��/�I���Y�0&21@��>��4�"��杫����`T�ܚ�yM�f�H��ts�	ji[x�p.%�غ\8������A>����_a3������āÊ3�km��0o`�V.~/� ^NO���x>9���(�Ξ8�ChמQ�w���{��f%��b�������T�������Y�|mv�S�鋼@�!���勨a�����Ÿ3Ԃ�#�51��`��;���h&�7�s
��\^D4�R�eWt�W��ع��3��gƅ������g�p��5���aF8�,�]�Â��{;��E(Ԡ�0�H�0"t� �G/�c~cSz�h<���~�s�=�ɞ���7�x�x
���I���!�d�I���6j��#�@�	L�󳘋lb)��f:!���|_�/|�l\� #�v�ك��$
)�Dkx����g��/�XZ!��,���{�*+?:�����,�mL-2�|N��D�λ\�4�����^D��PW�Y6������A˙�2���g���W � �̜.�ux�~*�a�Vl���✰��>��<���k��_�����qqJgr2�߈�ى���W���E������EOG�����I���?��҂�ǎ:"�����<K2P��Y2"�q�T!��]��a�>t��m>�SoU<�5~�>{}�-2�ȧ��U?mQ������U�`��F��0av�v��u5uj���}[S����B<��U}_����(�40.�aB��=ճ^�|5�����ZM��C��D����������5 �\h�J���e��7y�1�4�6E5�D��s',0y4J���]�34�\�"��� �f(�%96��ť����^6�6�{��%�$��r�*��*'Ps]�L^�:̂�#�5�-�-m��������Q�o�������vc�wX��(�o��|��C����l�� FۻT���= Ǭ�gO���-,�� W������FOG��O^d^`�&��I��#{���������)L߻of�W������HtK�#@^���&5bB�#C�8z�jj"l-�̩@+�I3���'1ԼHx��
�`=���Rsح���#���#�LT��=�=N$JE��-��W�q��GX4������D5�)�c���]���ϱ���*��M�8�� ��z��ܦC��'!hn�([i*���<z���Laay�9q椙���ٍt>�n���;�_D���$bѦ����aȨ��$��	��Cb	��(f( �IX^�����X�m��[��ZW�\,���j�]C衵#�|N$��tR��)��a$��(� q��@�!�<��
L`�j��ǹ��q��1t�7`r�aNq��!Xx��(����Ѧ���)�#	Bl�b��EH<��"O{T�1�7��{HOK-9���[7���C,//���Jpd]u����#�GC�ΐ@�ەڥ�.�ى&���Mx��6��%�ƃ�{�[T2��c� �W�w�>x<~,����o�WK�V�H��H�:(��,�r�%Џ�aB�"Y!ꐌ�#2U�j/B�T�]���J�����p���O����p�{�2r�=���sC9��n
���s���2�������V,���L�N�S�	�ρ�`��P���m+W��U\v� ������;q�mE���SL����V>s�z;;�����~�˿�=&FFr/M�~>G���ic����{�`�Λ9ů�0���x6+)��ٯ��՛Wx;=�k@H�丵�����TȐ�l��HP3q�^���=b&s�e��N�ѡtdsV,}�]��Jƴ�욄)W$��������wE�E��6��"��l�}H�(�Ŧ���(�[0�!���m�D�v�֚�}��OM�"6a4�\޻��9X���"��	�2a.�y�P����EzP��u�6�`v��Bz�x��$ƨ�b*bi�E�U̡�R�7]��9]���

v���x�g�ݍ�P��]�m��ӎ����6�����͟~^�󩍕�zW���CG"���9��2BN/v�wⓣ'��TN�1���&ṙ)�s��^��5���W�� 	
�Wf���?�׫l̛�o`��b�(�*5Y�PU[�n�Kv?���x
�,E�)��N�����CsKH��m�D������Ң&�x>GU5���Ξ��������	��;�N�q���~t��&�g�,E���.FX�p�)�D�9	�%Թ����8sp?v�t�V���_�����zv[�$+����$�?$+���:�n	���^X_���"&f���)M���ELٻw�]����L��g�.��,�0��k-xɚ�Ⱦ���������Ʉ�(5aes��A������kT�}X�[c��������
�Pʉ�@8takM�Ӌ�X߉"C?�bI��E�6q|����m5��p�>8z��A�}9�[7�ʯ���.���]����{!@r�����$���v*&�#c�$��m���Á]�p��Y1��"�v�1�nz5�Uf�t���Z!�A�OG�<�
��/�];]�:��+�:| v?�8v��k�~$cQ<���d�T���z�u�V�]�(H^�t,h:]M�dcr4K�`LB��0�iK�X%[�k�V�aH%���:�2��l��W�Y
�I5�L�k$l˃Բ-�ME aA�c�:`X��&X�)�1Qr,">�GX�z�]���ڂ�S�q~�8��]��s�(����q��S���Vi�L�2�_\���
�k���S>{�z������7���/~���U]G�R�^q�a�͟Ŗ/�'[P���d3�A��d����CM�t�����3�n0b�?����5�'�UQ�-�7�8"܋
���hg�������4���Z&C�*�u^�S�v�Tlk�����7A#,�*z0E�@�f�7�͎�:��]�
yew�f/O�zSFޗ3�4M�I����w;��I�$�ɚ(w��0�%�IaN���4
a��p�}��G`�B��\�0��J226��̭"L�d��Ы��<#c+�n�٥�՜SP���9�K.hD��l>��5��i���O�����"��o���g��1���q�\�N9oRw�\�Þ/Ù����n����;�N��}�1�t�9ݻ�����2�z�����S�`˃�7z��Z�������a�<|�Ϟ�mgh��� 6�#Z��ͩ��UFJ�Ig��'u�yM-�=xh?z{���_ZX�Mh�"���EAM�	�x�I�!ɔ�[)������w�?xx�����"� w��Ln�@��o��é�JvѠd��Fw~��EM»��h6�"����X".ؑ;��`=��*�^M��x�r��UV��$��Lbyc��M��v�9~Ο3<�I�ڽ�`~1� b�^j�+9�d�Z0'wN�z@��\y`y8���i�u�8q����B���+/�|2���y�]3�����n�5�i��*�O+�tRrja��֕��Aw�|A��T��	���T�?<v���}�wn������H&�����	��=����+��H<����v��S9E���䤢��&�����v����]Ѝ[����C�}�Z�z�<h,������$x���r�v�0������3kh�/X��WMIG��-<�}_I-�*?N�?k���@��B���["����9/%q�3݆�&��]tb��vE߭ưM�ɬ�FؕL�=�yr��d�?��t�5w�p�쏮c�9;�*P<�,8R����1[�No�,R��E!�	9�S�*���i�XS%���,��b-���2�Ns&w�^t�d-�lŉ(�����Сk��4��r#�����
ghkiF"���So���_b���TF�+2������ڜ���ĕ[���!�>`�M&��=��.����jf�=��w1�l�cld-d��+W0��2�{�ŗ��7!J{PQ��RR�_&/i��e7��#d*{�|^g&�K�>��]���eɀ�"l�o�H���=洊�?��3��)�j���\.�N)a}���DkMgvas^�BBr��ʲ�.F"i|�}UպO
�R��̚��:P^���@Uu�dsl@3i���������0I���!*��1$2DJ��sJfT)�\��2�6/:�������;���"�W7r����"��;�������(��|�];a��6��;�E�ًB"���Oq����L��E8�؎��Fݐ\��-�}.�B�e"�pǘ���<~@r�"�GF૮Ѣ|ym�^X��=Ŷw���#Q�7�So�f������my����CA�י�99�PS�ڂ"��@����ى��?I%�I��û�y�6��y��Ӵ�E�D�U���C���� ����R!�������s�l<`�v�T2�)NwV��/M�:�Fh�@�E٫�sX���N�_8w^�p*�1�ʽ�x���d1�۫"N��Œ��R�lX�9!��Q�t�,�l���gَ}�C��7�j���M�hl�������)bVwW'Bu5�ȋ$��~>|������-�z�FA
of��������\����|��I���`v��޽-ol�GL�i5c�P�l�Ŵ�d׫��lS~�j\�$�Q�So���]��:�T�i�@�3٬�n]�[ڛ7�!��;�!���Ԡ��qfh�0�)T��Vj�g�M&��zޖf�kj$�9�� �}�lF���CLL�B���A�67*��!�ds����Y�i�b#�儔HI3KdB뙴$��}^xU2��5[a2��愬)��MŦ��DP,W yÂ��ŝ���<��	��!["�lvφ�c�étF�]	B�TR�KJ�b�&UX��Vc��Q1̹��A�I���k��7���̤Y�vPb��"�aJ�l�TFp9B��s�،}����3�D�jij��z�5~���a9�$ȝ�?�(d��:�����GJ��Ћ;<~1�H*��/��~�3�����2�+7�+�:_�km��#jX��ӳT`����n5��^����eFx�S��'��"gJ6Y���-��2ai�	�!B������4El&U�	&PQ�`����L����Ǭ�m�����[6�|���_ϸ2I���S�e`銓��
rc�d�=ͯA䍱�K+�������d\(w�%�O�1V�)$]&^DT������St�8F�5�{�㱸�|��#�9���üb6]F�a��BR|U �ߙ-�����pW��n��?	���OϽ\Y�˩��3	I�����C���]'\�"j�N�56�'����ǣ{�{wocq~V��e�`5v�J¢��ފݻw�#����@'���?�s/_��]I�/
'a^Tv5\�3R�E��<������zd�]W_+X"��ޤ��I6x$5����zt!����5}��o��D(�O��G��Q�̓��q��<�x��ێ��������l&�o¤]�f�k�N8VD��Q>{� F�:��&4	�կ5u��$�g�C8N�!&��@(�N,���KJ��Lf�ϟ:�I�6o�|J��wnbbeEE���+¼y�;уZ�ue�u�!͇�d�b��*��L^.L��ط_L���l����Ǖ\��]��}���Ӄ��l���#D6ԙ��܉�c����}�+�m�Ƣ(8\�0��@���Ȏ>q
���X��Q�~�lL�04<8����Vf�4���<j 9�ӷ���e\�{ӫa�ӈ�p���}���E�C�|�2�ܻ#^���!?z�v�Q�rz�'a.�<c�^%E,��fV��z�-f«�3���
���ᩳyk�؉bl�)<~�'���k��Cu���V�a2���=_V�+����̞e�TJ��	WךL�Ps�D��5&d'=x� �B��_Sl%ҒS�BH�v����-D77�O&u�Ry c�e#��
�u_fsy�3�����3�a+{l���/�jq��a&{�9�{qykE���L�ij77���.=�D�h�� ��-�$MF3h�El;�C����Ο��3g��X�x4�Wo_��?�bxI�2	֡�)$}�v����.�lǃ�P(���l�"��������a?&���JNe|�X$�Ӭ��Y��r��>�$�]N��s2%������6Cs��&��%i	[��}@Mkc�Vrʜ~��������a�-�˰���h��x?���H���+��w�s�o��ZP�;*�JV��7{�Jm�Y�77����4^�l�p�Ďfַ���a�Y,	��~׸�e��P=5Ȑ1�a�h�t����v!��w��0df��fP�}t��!^Iq�����$]�����?�����;�/����?��^;��YD����9	�p�����F|��\8|�dϟ<ă{w�^�S�� �;Yd��	�Ji7<00����v�\V�'-N��5ී�zhH��UWIwL(�Ł�Ir��'�'��n��o$:k�5���sBBө$�v�{{����~\X\���jiş�����n�&�ѓǸz�:��G�e�0�K�a�KJ3�T¤bM�%Ih�D�e�>�p��;;�����k_��_K*����0����ѮQzW�u¨��    IDAT$�0H!���S7����E�7^\<y�Ξ����(�s����y�<4�Y8]-��i�gcE�o%T���(u���t���pܛ5x8�� ����d4��%R[Qd&��7:e�r��>H/a ��`;���ך�T�ZZ����x�������9]ȱc/�D <u� ><u��i\���{7q��5=0�������?"����4٧
��Ц�{�go�����ѽ�����"�|}��޿+^��}{qx�>����F�`�_�N�s�h�L
�TJ��s�K�\]�Ld.��u�(׷���T
o&���gx1�K�M2�hj@SW;��Q{�/�����Xd[��0k¶�����֊��VIo�������V�`F|G��U��6@��(Õ,���N��C�k�1y�D?�H,���E���H�,�:.x��K���x��9pMM�: g�sx��%r�2�^�X�K�a!$Z��XDKc�B8³�}9���(рr�S~Ylڋ������h� �bb�������ʢ��E�-h#B�ޮ��&�3�HmĐ�Č����?����N,�gϜס�t�%�޺���x6]I��RԺ���e�#}z2-r�f�9�}���>��),$��
j��H�}f�4�H���I�M��$P�tF�ZX5�2	�BW��Y��B�~�>F�Ε��!��	�Rl-=0���[���ኑ��8%�P��O+X�c�^�Y�lxiV��2��aB��D}�~8��Y0+`��I�Ne�$Fv�e{)�2�+Zf*{�w�bNh��5'fʣؼ2Տ�8%����˃]]�����o���W���K�9�8�r@!��x`���*���(;��Ј�9��E��ŋ'����==D�	WUaqi����H)omm���d���it��d׼�����5�������;�N��H@��ɥi�7K"�@uM��@+P�J����Y���s���$�ˍ��z%Z�1�����ֆ?�W�=݂��=0E���]vdx3x�(p���XE�0�e��"�i�/�W��|��'�c���DT����5��bg_H�p�e�?:�[$���u���y�����a�7n��L�\Ю�ܙS2*aD�Ͽ���"�4x�ގ2'�]��Z{6*�Ɇ��(R�	��.�m��8}�:j���`{uMc�"��*�j���10Їֶ&�3)D�;��)ѿٯɍ8w@��r�
��)���+�2����p���55`ei7n_ǥ�W�1��0�Q��5 E�H0?\�S.k|hY�ޒ����q���Q�6:����D�$�pxW�_�N��zǎݻDګ&���Pf��hv��l
�b����x�8����:�p��I�L|�[^)�Տ޾B�1��֐���>�MbHr�~�ˈ�@�h�j��x�[Z���ݍ����%�[�����9��ő�CT,򊾔�SJ�*��wN��t`W�<r���16*D�����[��3[��e�l�T�s%�4qz=�� N<,8�d��o�x�9\�>�kHr��ē:��]W[���ҟ���xp㶚^��`�~ʡ({���EA�\y�Ķ�v�~��ϰ��h��ː+RGOBm�פ|���l-� ��͂�_>@,r6�����Q9i��<{5���ob���D�4�|nleVK�Eͪ��LV1�t6��ˁD{nJ��$��"y����c�!��J�Y�YE�9�4�7j}�B��"\��,��j�̴k$F�^�2ڰ��ռZE�fDYK�l�Sd>����B�F�h	
eyR���H��j�@m@�?�E���	[p4/��>���pT��VW�!Ǿ��٘(����B�s��˝:v^G!EJ�*�Jl�:"�!�1D��	9G̿����`uu�\�M_vw���g��߾Y�_|���//�x*�~:��.�c:b_�����W�p=>�p���ݍ�E��QBD��VL+h�@��߉E�H E��,�l�ɸ�C6����2��hf`�wt�P�v\�ë� ��whO�ݯ����4�1 IP�iBF����������M6wcO�+�hl|E���I8S!f��b��q�y�(尣��by>\8qg����A�	ܺuWn\�o�t2-���`�6��c��4���o��YXT�- �N"�����8s�ܯ����[��������u�����ܤ
4H��(��.pZ%ZIJ����$\������H{'F;{0�ցB4��u�����*)!iim�����G�UScP�o4Ss����9�~���d�I���4n=}�gӓ��&<��./��هs'N����+K��]���������'80�W�Ry��/8=&H�{0���ڒQ˃�/0����:m��Hp4�Y��M���/�ե��^��G�{dXE���Ȧ���E>��
��3�1I�\�Y�E�Jj��o#�͡��߿��kC��|-n����K\��Ȣ�������ܑ�S�w �)�i{c�<�rPb�4}pɱ���0>Mc�i�b�`�NEX��l�X"w�HX��鐮|�[jù�;e���3��p)�G��憊0����>���]�7�^�������ʇ�Ls���>���g�T��T���|��;�4qz��?�B�a�Gl�TŦ��ӈ67������~��?��������&4������≔y�˫��m ���M#O���P.�l�����}_��	�����%��ڂ��^x^CӥS���1"Q$2匧�b-5��1w¥\��FS���	u!!��;坔X�|?ؤXE�d�А�3ް���_5b.�Zf��
xPz�9O5�W^��Ѵ�Ϻ_*llM���Ng���y��ׁ�4�{�m+P0}�-�&گr������q��g��ou�P!Bʔsq]�b��o��ѫ���m<W�|�VL����ϐ��k�&���9�<�.L
��@WO�|ݩ_�x9�`m�/�;z�����_��'��|��N>[^��ɍ�w�f'�Ҙt;Kv�sExv��e�@�����s8u�(�����s�Xʼ(��X��&��DM���M����<[S�m���$����	��D��Q��u��&muq+ka}.��#�!k����]˥��f�`�i�0j@��:�\Q�?S sﮮn����+��yܻSټO^���"-i�et�"�R���$Ex�Y���l+YDΝ<���w�\����k�v�
���C�7����t�Q�iT��D4k�������"2X2����N��A2�Qƭ7���+�ZY�������_�a���A��́�+j\	��!dT"wN��-��-��m��ӇV��
HD"2E���"��G&w����^��]ax��
���wL,���"�����>~��/_`�&���)�q��\8u
�!�����ۊ�#<G���=ؤ�<r�k"���i�u��e\�K�����a|fZ�q._��Ƒ=������v���|��)6����ߋPC�r���T�QΑ��5֒"��$���Ƈ��g�����a�^ۨ"�Y�$����&�Ø�Z���El�2H��HR�������Gqs��5D�7�����pC#��Bb�S�G���$zy)�~��O[I�(C8�I��3&���&dh�H�b�V.''4�ˣ�,��$;ҳ�����<��:���K�1��EF�R���UN7���ؾ��58�d�������눗r�
5���M�%y��.b���c����$R���U,Nϡ�ʣ��_+*�O�8�ǎH��f���4~��/0���	�������kK&�t0T>���D$�B<g��:5zz��ɛUӣ���G����! O^<���w%w����vz}�(�@�hU��G�UI0?'3�'Z��L�(�>3�E�����<����9�L�ϕ�^xߑx�g�8�DZ���4�����"lHa��F�mp]	}���:�Wh{�kU�+5 Yk��?g<��ͦ�Q���ڊP$���|��w�A��X�u���k�H�#'��vtYtre�{�e�d,�,���V�Wx���0͊өk�3��2�g8�ҷ]�"�j26.p���Ő�����@�?��v�٧�m|�E���c��?~����N��4����c�L�F� W�W� _�.��'����#���x�Ϟ<VYdhR���7hmC<�*�3�5� �QrY����®�ף9Ԡ�-�Laiф@���ͭ�X2�h���bjwm���b�$�/� lzCt(QII,��
�
���T���,��?�$l�4aZ��P�.$琣���2��pÝ*�gs����8{����	��_����������ޡ�����䋗�R�Ix����� ��	�!���_^�'���GU�i2��w��M|}�2f�����1��Y��h#H�''d�����0���\^Ը��	����C-m��؝���XZXD4������E׍�Ԕ�q�ǉtieI>��TB�:�0���9gM��T��>{"3�|���hCU-N:,N�ˋ����&a������k뀷���U�e+��I�$v-�0X��y��U���S+�x;?']kk�YS�����e��8� �,ڧ�w���.Oݱ����v�8����4B��n>�a�cy��௯G�m�b"���Zu����,p]^[���2��I���X�$���x���6�3E�b��0����"��w�����]��9��1��+*в��$�9u(���U�7v��TX�b�����,O�|�|�`e!�o�Mr��T6�NYa����˙)̭�be;�C�p���C�݁]�8�� ���a�~�6V�[@���.��kM����%5c�6'�R��anr�X
�U5A+�Z�q��a�>ym--�1s�'_�+[:؛�;D
��ƹ��{)c\o�TH�;��kkj��K<WZϿO?����'z�<{�k�n�I/Y�)���e�ݰ͹[�����ޝ
Fv�$�BX(�UX������钉���������m���F��IP*�n�be0�3S��p�o��)éSA����W_�:YN��	�aZ�Yk���`�J��g��Z�'���誙�}�7����0�����[L�Z]5CA�M�U`�պVD]��՚z����!�i7*ZT�k3�Ͱ�]��<Wˀ�>�&2��l6�U#/������c���WÈlms"���P���G�l~�E������+���������I��@�xz�"����ޢC�,?l�W���9�=~T��ZxY��AH���g��<�����Z���Nq�ABC.��5ux;�U~�ѓ�fw �JH�`+�n����y,��1�?{���a�dS�?ӛ�E� oB�*^������������ |~�B���?Q"��g���)�P!'{6$��4�?d��bc@�R�ݔ]� �9v珝���{`+eq��u\��?�N����ݧ����w�2�7Y]}����RQ�����$L]�����ԙ�8r��`�[�o)���f_�i2
��nN�=ѭlzfF6�4e��:X��˫Ԣ������A�����5�B��f�9=0^WZ��3mn���Kk+rBc<d:�ԡ�i�gx���������x�j\��LAE���g�é����+L����|���,��������87<�8���y���+��l͝��][JI5�,����;��p��ܿ�ETW�1�ׇ�{�H���F.��^��6��~*��/_h¶W�li��&���0�c;h
��Ӌ�9B��Ǜ�����B|�[�v��
���#O+�`{eM�!`�hy�t��cxh@0t=a;5�f/G�)1W+�O�R�I��\��ؤB�l%��L@�"n+�oC��]�Ȝn�i�@�a6�g�S��4(�]]���[%�-�����C֯M֭��G�Z��*����k���%�*�S=zw�BϮ!�l��)�"D�qyIG�H1�`CG]�\ks����+�ܩ3hj�G�֡3��/~�D>���:{{���N���ѝ�H8����fd�uWK�,<_=}���w�ݏ>�G~�"���c\�}/&_��fCϳEV���8*�e%�q�d���X�"QWDM��E;���p��H��Q�,�-"�Շˣ��l,K�Y`�P�Cu��BHdRȽ��Ҙ�XEXT%t��O�7�r�����+�W�AŠ�EX���>I�V�0��	�����~�1�M)w��ц3�b�&�02?��"��$s���@���8|���@/i����KgRx��&''uO�֯���ԕo�zQæ�k~�@�/%�T�-5%U�\gzA�@xo�.-�������w��lt4����饡�jy�(��ܫ�V�7�Q?�9M-͸x�4�;{��,5��$���,\����fZ�9�FW�P � ��'���N�X��[fxٌ�>�Yc"�tf?҄@��re��ԍ�r�r��g1��>�|�7~��������D� ����ܾ����)��]��ȶ8i�)�L��2y��|�m��\�=~��ޭ��ֵ����W�C�����BC�-�'&Q���ݭ���Z~Չt��Z�5���ؑ؝7֡�Gp��	���gܼs��^����,
����{�ؕ�Wb����9�Yd1gv�n�;��W��a0l��<h��_��o���7�X,�4��G���f��3+�㩓��ֿ7�#��.��������[�
�����X��;:U�g��p�M[��=ɋ�����]��&`W:���6�'�q:���(H��.=yّ����uDKg�v�k��[\P���Ɔآ��vw!�ڂ���x93��3��U(�7E���]��&&�ceiO_<ŗ���Ozw7w���]��<����҇��i��0|��<�;;�ux���EM/����Ə>��P@��_��w�>���"�	=��g1���ө�Og$$6ylΨ%�ZYF������x9;�l���d#~�G�����W�&����kL�/���(�� 
�2N�22�(g�jB����֌��l�cW0`&)�ek�"L��u���F��E�M�Z��Kl\������2EV<�'Y�lb���2�`�H�2�W��+��7/el���+Y�|ܐÍCg��B6u���)����q�K+������]C�p�8arm),׌���Y���k�đ�����,��)ܾr���'�2dc�������+����Ds38\� JN Ms�bA+	jp����\dD��%d��������mܺyS���1�<}���9I2�@KS�TcqCZc���1-FvѤ��'C�m=.�M^י���3� �!�M]ɗq����T
�hܘ��|*���U����i�(*I8]r���[b���k%��n>�4L�2�Qئ ��T������[[j<X���"�D��'Zm�3�$ˉ�Œ����:a�U-��PNʴ	=7j�1|\YlZ����r�&�4O������//��(�/���	s�bɄQ.r5@B�K1��)����c,ml���8�}����Կ�OΝ;����������ѿV�Ȕ�D��YwR,�ܑt46�0����:��T�B���t��^Hn&t{ក�{��*���m�#k�%�K���Z��q��$���NM�k½�)�M��>vU���{�9;C�"�J�gj=��qӿs��-�1���o�>��ׯt�V�C��e�&I��<��=�*�1��KYC����uܸx燇E����]|��/%�hmk�~z���I��Ʀ�C�u@[���Q��'�H��+�q��+�/�֭[�t�"�������+,n����9�&2Yz;NLb��f�L&��20�T�X��}���D��#��7W�G/�=�Ծek���y�pY�@6���7w�hǲ��cX���gf1��ۇ���Hv����^��`lnN�v�qw���!��;׮!�aqiϞ=�����T(֡y�oX�p/��3�;������9,/,cue�B	��m8�f���l��?��4�������������\]A,҄fh�g�(~��nfj
飔i=nL..biw��fDP�yu�0��?��O���"��7/���#�Z��92rd�8�^d�4�Ul!�Y�A���i"oki��5�6�/�    IDATƼBdcG��eާ,X\eЬ��3v��%�W�K�a�^��FI�3+M�:�h�X�.�׃�J���>�drs���=.r
�}��g����/���x�Wp��WIaGF�ʘ (@׿����G��{3t�
znJ"��O(��1Sfj�Cg�9�J���s�������m����,�xIMR���;����ג�P�Sw�ԄhcR\Ƃf���8#�-f�g�P��p}8��S����׮\�ّ�bOON���ӧx���I����Tc{i�Nu�J>G-*M:8��=c�Z����Ζ<�9rG�b�B9������r�����g���f����`¬j��.s�hj��֔� Kl3���� �� ���k�]��)�\b�����/{*VP�`���;�OH&c�c���?�Ή#DH�g�qEHF�zl8�&j�k��q�m���O~"R$������rq�S�h�	ܐ�"������ǐ{�ۣ�P�o� b��6͆=ӫ�o.�:�;9�k+x��o0��w�5��߿y�~��7���-��o���I�7 w9n��A����H�������>��w�Zu2��á�Txjؤ1#�D����At�C�|��7��b��]ݏ�՛ǡ���]";�
;h��I{դw� ��މh��UQ��Af7kUgސ�X鷻st���,,-�F)+�<	��~U7��0NP{�e��c��}�n^�"B�_y����'���d˄���u5�'i��%�}�LB>����P��ffG����+�s�6.������op1���z����:e�z�i���*��~&-���o.v�-��j�BW�^�I�ӈW�����ԇ�B1����9u�|�Y��b�$��7$%E`xF�T�!������A��r��F<x�K��^^��Y1W���AoS>�qw�]7ExaO�<��_�"��;��#8���J���5�<ډ�w������:��Puz�7<��ǇÓ���Y�G����JLZ]_�w�ػ7ؠ�q!��.`C�N�X�E�����%T�.L//cyu����(��o=�5fg'~�'?U���ӗ/p��}<{g8�t.�/�a������������N���G�i!Ad�VʺΉ�0zj�azixTL�v*�U�3�Q�edh��|5����v�5��$�
�7�ߒ��+W����"���t���]X�l'E����ɽ��]=�:2���gP+�87�Ͼ�{;"�9B~1��D��@�ʓZM�59%��]s �tk@� g�� �3��8��c"p�51򹣞]^�(�r��8<���a5Q���F�L�>[��0�$)K���w��M�"+�O���G����S�Ex���w�G�|�������}8'F:�)`fc�p(����uMlI�DN��r������x,� 2�iw��_ �&჏)Jt���ơ��;M�>��X��1���-Q��
��Y��I�Jh2��ba)Tj��rQ����B�"�3���~�l)��,�$@�
�jYX���?��8;:��&}����ff�ͥ�8lNTT9�U��B"Ԓ��� �sp(.
L�~l�Y��Y˯ҼV2�miԍ�-L.����"e�������ůc'���y5��?L�,��	C��/�(X����HE���Zs��H;:�_?@�%*�*%Dw	�Pv-Vj�,�a\��w�Q;� R�I	Pԕ�o��'w�"�Ԍ)/j٫��>�jAʢ�[N=|�Yl��$�m���c�`��<��r�rSSl���=vE��X|�F&c�;`�c��ګ�]*��+Kx;F	̊
%�7�+�p��yM6�ܻ��~��U�#5�X���}��F2N�P\��J��� ���l�`�d5��ś���܇]9#y���߈y�"|X.��v O�K�������~6�,Sp���ђl���&���$�Ɲ��O���	y2+��7��R򴾾�"�)���Y���¼� �d���h�삷.��=��a�4e�e�B]�:��2˯�@] ���9<~����R!����_f�a_g7�Z[��ݲ�0����5lm�bmmC�3�����k����A�l�~�?�;��������ԛWҜ��������*�蒤D;���GO������%�o�'�d�ut�'��7U�=�`�/|����W�$�Ǩ�|p��x���EH(��GwW��X�Ȱ�*?ɉ$��S����
w�4�Q�N8�|���C����eCfVCN��&��\��rA7$F�J�P��\�k����M(���يh�*<H��^�� 1���\��)���ζ���k�4H	 	��s
�֘�0�E�!� %^|��KS��Z�F�љ�@51��H�i�r�}}&_@U���R���&��X���4ծ D6r0���!5(U�{I6�4b��n�>|�g/�J�S_�@oO~��Ǹxn�r�"�WRz������^��7�w�������G�7��X�X�y�s�L�r��|<����?���c8b�(�����
Z��4Y���&a�i}������z�
���Fey�����xlx�Hs�g&r�����|lonij�'p�|�E�S.Qe���������������)T��3s�	M�|+Q�"%�qgN�kw�,n��D@=yl�u䘴��S�h��.5�\��"�*�#4�Y�����y���9���_�����/�]z���?�/�L8�TWn���&���e�)�2	xd�ν!�"�������):��8��H�}&�W}4�������/�J��bF;Aj�����|L��՛�EX �L�x"�6���;.+�]�v�4����2���^O&E���M�+E�]n-��]�(ז����sr/Lw�|��<��+UL�L���g���c���֩��폔������_����bgG�a/��x�X���rA��\�?قI(��<I6Ų�y�^>?�k�.���K(�ڿ��.^-���p7����+�t�pIY�����.�2|${�èK$�[� ��Ó-�}���$��=�20�S����R$��Q
kۛbV���D{gfHD��Vǻ��&�^�Ѐ`��L
o�~|�=�^�:5M�j������7o!��annZ~�_{�<]�<�d��h
��W*)��tJ��rف��Il��{` �PP��=z,g�����[���P(����K�{���q�lobxp?��S�w��ZSGǂ�Mx6�Oލ��1�(���ܼLIz�:�?�M�|�:����o�ᠴ��	�^��*���7ݻ\���7��#_�q��h����ZA�퓯5�=�C� 
����7�Q�}�B���uŰ�H��m&a�9�A;^S2r�C��$&R�HJB��T���ɩi,�.+G;g6
�.�9�O._�پS�<2� ���l�h�Sq�4+a�Q�b�D�t�0;8��t}PRƵ5�<�8��S�+�ij�pH���!]-(%��H=y�����vB�E^N�,�z��K�J%�x��}��&�	�����k0�8�_�$�T*-���z>Z��w��K�c�f�vb\����x�*..���hT��z�����3���?��\�h��7���f&�&op��lC�6b�^����!x/o��K��]��d&٠~�C纃2*����$ςȉ�!;D8�ز��YId���G���|�v� �ݩ�~�������[�Z�����ذ�y���X4	U�n�3i�̽0��T�Ј�����T��N� �ld~u2i��O�s,��j�ȗ��88���������������K�����^�.�O������p���wӕ��{�-*=�F���5Z��a;?�V�!o�0w��l����2�:3N�071a����S\�s��2^Bvʁ��}��G��ܵ���nE�}�A��B�e^��k}���F����d;������وq����xW�ɚ])'>���E<y��>�N���G�n���[�t�<��#=��'���-���<x]&B���o�B�/c�.���y��̡��A"��*���x��}}/fg��QxPP�'��ok�]�L�S&�	)ҘD4Q'x�!o��:��r�|��,�q��0Nw������`@QbL����������zA�5�D�P='��wS)��2����!��
eM@���m�������ɍ�����ܻO����&���D��xvԄ��jH6$�H�E �n�1ь����1bu8)��Iaum]7%ؿ�[?F���6����=y���$�b���ę�a�ҁS����k���A�����ށ/E �q1��O�!�+f�'?�M�������_����_������ '�aE���b��:��Ԉ��Q����DLV������Y.+�룦��B�XTҋ��5K�
~��Ѱ�:jz�e�(�kg����AO���H�G�?fs�k�\�f����+,���)�9��*pa�4n�^���A$}Ax5's���{��V�V�n�?6��6���!,����ӱy>�|2���)�ϰ����*�F�)i7�(��u.󗔮D$��ɟa\{���S�_>�W_�����1�Ώ�E{S��s�K.YD_N�SJP�O$E��%b�l��`f~�++:�t�L"w���ɺ:$�q�h���>���Klo�2�-A��b3Y��c�����C��=�b��-�v4HO~�umM���[�,Ҝ^�|�xs���.Ml������c��dz�ϓ�$�̒��,�j�Ô#��d�?��KW����M� t����I��Mf>#߷��F�[��ʅ�ۿ�;������=��:�*c@�v((�u��li�:�S���2�:�f������[��f���G/������3ã�8w�������.2�#��+��	/v��~ͮ�:C������Q�~�7��B�,��(��c,�D�	�˩��Y��/.��dEs�L�w��GF�B�ө�"L��.Sb���4Ic*�V���:P�P`�2���s��t��%+�U�T~�����a��j�M������C��E	�xSܠ���+�|��=�g�+!O/�B��\���.��%��L�+�p��`"�HơĊN,<%	9(�4����{��<|�F&����U%�UCu�$�:fN�*�ᎆkI�AJ$��:��C�,L�J��Σ��`sz[��F&�7�'�y����K�snhH2M�V�d�Bx��>_����R�X<�E�ZF��;�E5�p���\��O��D2���2�=���}���#Ч��k�%�5�C�����2֗�T��O�@�]^E����4�OR�H�s�~�?Q` ���_~�Ǐ`nj��z4�r�I�b:�JL3*��><>F]}��v�N�����*䱸���s�XMuȇ{����V��4�Ѱ��X�Y�|��h�o@?m^��0�
%6P%M\����	j�]d�ל�	'�Q5��y�o��bmw[;a'5�t"��)�C�k�=>˘�a^��4�b���G,�T%��9�E��7���B�''T�e�Hß4	Gnv���鳸6z�@P�/��E�--�0-;���J)��>�\ˌՐ��#�C���<g*����*����2�}��ـ9-Jjh��I8Er����0/τrM;o�*X.R�VRQ�.��/_���_���FC"���j�j%_����u	�CE�Ɋ�O&B���j�����r�Ҍ��V���)}�уﰻ�o���;=&�Jf1��1֛J���>��R�,�g�5�|`���_��!���`�[��s�/�K��?��qiK!O~���9qV><Й���n�dI2�����&1��F�I�.Y��X�v�&���Sm<NIS���&밗��������|~!f[͂�Rx���'��ެ�pw�PCE"���=]�/�_��`�����O��������7�����{�#�/`��Y6t����槑#����9:�P��=��'?�j���E��C�P69�nȰf�t��TS�F��Ho�
���4v��s��N��r����A̴�b�l���w��d~�ߖ�%�f]p�_��,��[z8���%����!�t"rr���B�|�.��� ���!����W���7X#����+�p��%�xa���N��%3�%�.�T�I�{�(;68
'��4lS�����$%��~��Q���gO�v�Qq��!����B;f��9�[�ڐ�X �xD��(��9]��^�S�Y�"Ru�>1��=ݤ�U�K�����ކ��aߘ�K?ev�iN����������}�dOdTA6#}����!ݕh��^�oܸ��hD�ݗ�^೻�&��uu�������A�k���WJJ����ց��vh��݃�ww���!�5�u����}�V~�K9s��Uߐ����o5֑F�B�N�J)O	0�������U֓�o侯�����*�4b��5�1�jWGy^�^/��:�i>�Ќ��$�D٬V���M�\�jc�A�<#�h�AS�&�D�d]\;;� 0�{��d%;����|�|��ъa������6N&#�5��{=5��}�k��C:!�]�
Q����&����E�da�i
%���נ|��;�+�{!�$p���9�4Ҝ���s��E�PC���r ���8��keT<�gT��U�������F�����18Ѳ�}��Ξh')BU:��Y�e���ЬF�X,K�����n~v|/��`�$�`sg[�1���7� q�ǂu������[�똛��F�`�P�_4S�b���b��K��f��|�`cO�z-�,h��Ōc�����+���,ȿldP2#����5^rg��b��cw���َ�e*m&�"ɱt¢�C ���9��9�R�����?�M���I4f$���8��B8(�0��,3>o7 �O�8����σb�$n �'N���<N/����������1	�՛��y7�'뻻gΌ����i��8վz��}���m3NR�6DͰ }N��J��`����N������S/�P1I:�]4���mb�����z�C����P�([sog_$$y,�õ<���b&�ޜ$0�NP�U�ν�%	JD�LF=;d^$bZ;$^�f���Ȭ��м��فI.2�ښ[$�~����յ5M:���F�O춮]���-�=���`�O�����K�iX�Msai8����f*M��������e���bbzJA�Ufor���b�_$O4K<.��6egڲ�>~ޙ��K?J��[}"��8�hЁ������Nt�4��q S.c�����3'���û�	,omamy�U��p��C7W��\EOc;>�v?�����^�|!v�����0ї��^���"D��;�"<�{K`�����W��o�#���.����������~�c�$��������o�ݣXYY�!��>R�R��]�!b��v�^��̞�}���m�l��|��bzq1N����M�2�#{9��w�L�PE����N�+JKI�[:hQڗ/�%:�k�\ N{JS*�#-%)�a!�mr���ڡl��}̤.�4)Qf#��H�`H(�H ��'�w��<��n&,�+c�D��JM�NN�t�FS�Ijkh���:N�r���ߋH2�Xs�ѐ�T��UP*���h�^#��ȗPe�{6�ƈ2 �	�1T��}�7�f(�P}��P���oK�rުCʏ*}��6��O��ZQ1��o�'ĂaE�� ��K�/$󷬘��ѱL8I�eO-+}�noIA��G$
~�Y(�hѢ��ś��R��C�X�����|f�U�Ȧ��mm�
!SѨ���E���`!l4>�-Y�I$3ot؍�M�V��^��8A5r�Y���6�u-�˒8�e�����g&�X[ش�6�J�.H���7�����Q��H��ω���H,�X2!�#o�/�H$�D,��#�9�]|�<k��{������ZM;���ɗwƧ��dko���������.U<�_�l	E�Pc����N��8	�\���gF���}cC�O
i3�����*V*?��u�L�D��^ڷYF�>��������/��`���4�T�C.��ô���oB��`���b����Ύ�C�D��߳ ����
$�ǋ/����Ds�{T��    IDAT���$�ˉ�T�L������Fn}co�����w8Jg�'0z�΍�V0<*%��Zic��OȈ����[bxj�m�Lh^��`�$�]p �66�@:�V��I��C�������P2��k�'�z21��&o0`s�� �{�8�����	Z�T��1]��0��$����.�\@�R���1v�5	3�����������'v��cr�)��V���N|z�~x��b쮯�������ϴ[��A������A��FC����Pʞ�Za����"&����ǰ�>���.	I�Ώ��D�����/~��ϟaai^�u_O/ΝFc<� 6J�hB������ߓm�F�DE��vḔ����Db���L�R���/�$.«��}�zN������Ü�����\M��9�2ycѩ�kY�w�<|���0"�{���oe�*Mˊ�NԎ��"�qи܅C�h��9e���������(�Ed���#�����
V�װ����Ў�䞘ϓͅ��$O��46�����:��ܿ���."F�ea���'Y�N�?J��32-e�R�H���C�W�.�Dk��2}���LmK'�)�T�i��EO��M�f�7��/ٷ�d�*���0�U�2!�\��H��q@Ř����AM5r��d�{r"�7�#j�����HN���z��/��g>^����JQ��a�Cـ�r�JŖ�Ѳt����MN��8ĜQՠn����
�]tMR��nd�Q3|��Ҷ�Թ@�����6�3�>��;\p "�i������q����J�,M��:Vf��iu�� t��n�	�c�43������s�5���/�� eb&�;2�0mH���s�������_��>��鹥?���=30t�Ϟ�`g/�"޼y�������4��P��
x�!YM����P�`������PW�����+�'[*�����A8�ĺ���"LX"��zs��ꄑ\��')������qZ��I�F�ds�2���.�^���W�j]}��*A*%�H�/��B��<��I���О�\�";򊚉e� Cx�?��嫸s��/(ğ����O�g<���d���<\9�0N�$/����K�|�90��l'}���%=�\�"c��N��`���Z�X�ign;�9�UK�$�󂿋�Rk���L'�y��-����v��OF�嚊`S]������hko���L�tJ��,<��]Z��o1�0��׫Ʉ,zu�̡�9�Yߊ��_Ǐ��Bk<���-�}�?��ϰ���t6��a��Op1M1��poD���b�	�!�Ig�x��_f�lNE�l� ~��m4�b8����{_���[���~3����[O[�^��\1�s�frQ):9B@���` �jYьl:��VDN�]ʓ9]�H�f1��ZS���PzS�dQ+�;ɢ�Pu�<�H�$�9oE\ ���'��E��;QbB��0.�����mHtG{�@H{lMƉ��&Ѥ����"��{��H�ڭY�ME&����2h��3��B��捫��p�GM��ن�h��B�!��8AE���M\��T�\U�f�0���>�;�p�q��fe,<�;�UUv��� \_gt܉�8��p��i�_%�����Q��h-bO|<DV�}Coh�)C򷦞�n�9�r�&��d.~���."6���JES��Ȃӽ�eY�	�f�Ntr=��'�Ֆɥ�\4��f�s{g��v҂������X�/���E����H��s��~���}�b2��Ĝ��(98Y��z?)M�UEHc�u��H�:��PH:�Ӷ��������<y�k�Ow���ɍ�=	�������ƣF�IU�k��w!�����I�����ٸI�b|k���ۺ������{��U~��v�q��[S��vsggd`hD����^ŷ�������biy^�v��O�����`T�Wt���hE;]�8%��"ȗx�U������}$�v��ڪ���u����A$M�X;����*v��t��a�I���сn6��O;:B�;�d� �DN+b=���
��E3���:2�ޓ�|n1�d�kU@��y�$�L�Lk?�u{7��*�$����IG84|W�^Eoo�Il*�����INR�Q6-a?���!�{?OjB��#� 3����,�v^������)j�g1�����W��EJ�JƊ�a^�j��B�����^ռQ���xwv����Ε�;!aj�>^�pI��L�b��F�И <5��I�&qx\H��X^]�ӗ�057��!B�$� �\(��c�����p{}��=�{�
?��ϰ��&8��j����o甔>Ih�VD!���R:�;C�@�0܁ �vw���,o�ݹ��?���=|�͗�����޾���'���@"���l��j���t C�wN�/��D��'qD#~���Z�zx�KE��q��,r&#1L"�� p��(��4�f�O�:�&���&�"��޹,�ۣv_Zb�K�2_3��PA��d�]�-_�`Zy�ވ���H��'tNv���A�{�J�eA.B�Ti��uc����#q$Hأ�܆���i3[��o��H�־n����)G%�a��f����W9����N6wQI��@rI��@�y��e3�t���͍��#�z�~Er��8*����d�ZX��R����=Q��&��&�*v���(NVt����hOˈ��sk�,�
�<�Xȍ����d�rz��[��b�/6������ЈL*m��3q�4FD��\/��Y�W���;�bf�mˊ��w�Zw}�#��Q-�a+���f�ƖgZ�W�K��W�����W~�4�Z�mkR���6a���;>���B�ͭ$����S=7i�ɻ���Jy�$3���u���5�I{���	�����$�H�A�N՚�IyO������*����D_�w�������_�{�"�W�޻�va����?�;0�ё�8��-S��������d�@t��]f\����ӣ��2���=��k0�h��Je���=8��e(B�>��XX^��N���d67�����r^��ڎ)�z��d/Hhv|⍼��!�/+�o�.e����w6aq��+f�`ѢN�<��듍"���Κ��01	X~����6D�1cX,�|���Wx��!2�._��"L�:ulS�x��9������z-܍:D�8]7����=�X<y�����$SXD���!�V6]��r��L9�m=Ȁ�$���cJxp�<��ʖ��?�U���DV3B}��++x��ӧ���b�o���ql��I�q��%�S#���ku�(��i�s����4ӇύL.���-�|�+��888T�J_�L�2������z\9�ܺ���vlo���'�{��.'��,ǃ��.iػ<,�8*y9N*�(��� �֊*c�|A
EɎ���ik�+W�����}�w�o��h����� B�^�ɹ^%ZQ�
��$�_, �#L9Q8���o^<�	���ZTH`�5���6��2FIFh|V���{��Ϣ������T��m�_x��[@/B�u��&u>WNQ)F]z}�Ɉ4�!r�I�T��x�������0�$�Uae�����E\	FL$��{h�K���ȉI�����/0:ͯ�h%Q`����i�Y���2-H�5��)�k8aE��+����xx��A
��m�sey�K*zZk� �N@�Z��hlo�~�S0w´���MT�����+(+,���S�,�c�Y��KdNqS̽m&F��y}��@6��(��3�T��!P�V�sD��O��{Xޫ�������S��UD�N��T�/d��'k�\аA�$vӤ�{c�϶��-oҹB���������K�f�%����Aq��l��mb��v�&�lO�f�����s��"��Y�0��3����!�#Y�R�ޜ�����w� �\�?~�>��t�M�:��|�S�Ǩ0Q)_Թ�)��7�����/Ow����:����.�-������hW?Ν�HW�����gF��4#:���C�č�71pj�\�L��0�ۃ�d�XTP�:�bIF�ǺQiI�ԅ../`v~k��s�?�>р��p�ŋ� �́�/(�M�i���������*[�Ei3&{G����� )!jjk1i>��J��!���irrRP5/��9���r��4������}i����@���.��?FkK��"���\9�k׮���QR�t�G�{��,�ܯ�@.��[*�;6��5	�O�E/d3���R�W�����I�Ɲ��<���c˦��4b'���KR��=���H	[�9�s���zF'.��*K�tm�*�o��cG}�ЙӒ<���R�Ģz�Q�!�q)c���������nʉ�
�\�.� O���h~p�
>�s�-M�������w�����]��gH6e���r?JȾB�a���!Ӥ���8!�p�����������@��B�x��/cva{���}v�����qFꑠV(�0���<�S�H�f��h���1^�L!G���k&�U���d����)�@��ɒ�դ�%]��T,�4J���2M4}���b��*#� �AI��4"�%�}����Gv���s9�t�k����8Y��K)N����� 1?sN�ԀsR�#:=^���$�)WTX%�c��r W��|��ˊ�dQΔ
���,��Z	�4t�!�� �xE�/�$�eCJ�OB����S8^߆'_F��Jޠ(rݣ	��Og��ނ��445jM�B����L�dF3�xp���e�2YpO�8��n�i�Y1�RM��Y�ݮ�Y;�0a%�o,�D�XXK3~PyOr7.n�=��)�||}6�艜h�[S��؆�M���ey�K��(f�t�;����4���ő�L�\:3�g@�"�5��ưw����Qq�'k[JR����Q�<�l~�D!�w8$�(��:�Ɨ�k&�[-�(�+"�,�)J�4����C$�U��[�A5#8ia�ح"L�=O�ni~��7~y�����������ͅ�S�������gό�lO?��^�|���caqFTq��I ����퇣iR;;t�-�H�c�g�tw|b���N�Z�prЧ"L����4V�����#;ƈ?���Ɔ�t�LɠKU�ִE�#�_~�<�L��.�>�$x�t&�����S�$i��?���eO����>�:uJp�4w�t�j�0��vvΉ$�d�*A����M|��^�}��j��E|��GhkiU<����=y�I���+hiiB���vujzB1u�B�\��EM�,��<@SCښ�������,�����A��lj�k�z5� �;���"j�\�܉�a:w}u��s%��"0�I�zbL�9ʱF�G�O��aic��ں;����^Y'=���ĮJN!�]䌯,����f��)Qc�/�}�v�Ƶ���t47 ���٩1|��]LMM`�###�~�&FN��Z��4�⠗:ꪢ�8����X���]|Riٜv6���i��!���1�N����
2������vt5����gN2:���0��W�V�^&-w���,nl`ugN
< �J��})[a�=���aw}/���J.1^��J.'��B �f
㵡ݤ�%/]�K��kN1��4�75!M��BH�����0��3y ���bEBɋ�ߜ���J�Ƃ1)cb�K%@���@ �hL�?�1M�0n\������F�RT����,���{HMc�"�)�pt}gm͚�K���E�jZ���*�q�7�˫[�*�Q�P֤,/wB���ɓBN�]�zE��a�	��ϩ[��@�;��R�;��3�W�&ZU4S�m[�B/��=	��m�RY�$�$ه���E���ʇ����Φ7?����'JM���E�r���4˄�m�^��%�"���X,�\iq����ks^v�:���q+4���忳�`��x~Y���mhZ\����4mM�Ĺ.㺲d�EI�#;�+�P �(I�!�-lΉ����9Fb���e�JN��ݨ�nUN�
Z�r��7�x�����Xd�P���\ׂ˃�����m����:��{t���٩?]�ٻ�yꔊ��SC��L&�n�{PNçNK�wy����L�=�����DSC��(�[�{��?�^,N[�����R��҂
����V7��t�_d&>C�i��ɛ?�����o|�/�r�v�:��$G'i47�"���u�Ԏ]�zE����.�s#geIȩ���ʊ �H4����F��1�䬍��z�F;Cބ9�}����Y�߾~��zx7o]Gkk3�v����k<|t_Vn��4�]����Ύ����S��\�X�uwu��E�
'���=]���{�.Xp�1�wir��L�~��J/�x<*��ql����ur��/j�m�=��ۇ�|ZI7�={���y�9�s�Ϣ��];U�}�Y$����H! L�#'x�(�8o iv���>��/bll\{vBњ9V�h���+������nmF1s���)|��g{�ZA.\��[wpzhX7�C< #� 
�2�!cyT)a����V�v$�b��?��ۈ�V{'�|���y9�I"��hFiҒ�!�	�� ��\jO]�>>����I��<�d��(L��-���>E{�Q�A�oRG�c�mNݹ"�Gvt�$nF���<�}4c�H�a�(�Z<�i�Rߨi5�i��k��R��.'$)R�����`�a�6l�vwT����s��i���Ʀ�cQ�77#���^��[0P=B���H',�
`mGҭ��ul����>��Ϊc�mͨ�h5�v��a�)t��"�-!D9_����%��Y
�G�jѩ��:�%����c�Y8������I��<p6>$a�J4
0�}r�Ss�Bl�����r�"\�A����n�ڃ����,C�lN�&޷$։�a���GV4eK���Yp�Z��֟��.���O�k��X�j�X�h{��n��Ւo�&��?^�,��b�x�qn֋6����������j ��0�9�>[�d���д�K�i?o��4݄�e)��e��}D ���{AE��0�~7�=�u4"ܘ�I5o�0�U�Y�����k8����F�,ǹ�p{}×�m]�k)���ޥ7����w�p4e5�*��������w2�Pr:��8���G�OJBD��x$����C���.r����=�bq4�����͐8�E3NMarl�����"q��t��=j����M�!H䃮�v�?~�P����]8�?$�����S8�~��w�81vf�����M��@�f��Ό��\I̊�T|	���?��q�)n{S�}��\�&�RWG'v�����E������G�T������cܿ�5�ǩ�(��C��8�޸��/�:8�Y���}]�x=�Z�����Q��1L�%���gR�դPkʋ�7*'�S}�r4���VV�lv�.�O��E-���>4ExzjgϏ*6���;�Mj�I/�?a)�[�3�[0:%"E�sr�b���
:���2&'�������a1�����틗��۷��Ձ�I
��*c�pr�A?�^��"L��lN?�0^0B���.'v�y���`���ۻ�Eb�m��a\F���R�S��n��$����|�ɖ,��HQ{M����#��v{]H
X�ٔ3�u�m[="�L��R�L�Xu� ,�r�ˊIkL.r��*I�d5���;�(�g�"o�9}x(*Q ��i_J4��5�|,��V9KL��kcaJ�M���̞��P�csu���ƶaI�)��!�ԠX���&��t&"I�>�%�[�&��x�EӠ�����,V����F='����&Է��8ړ� S���Q�=���&<,�$8�&e�W[��	xpx-�m�����M�7��XԸ�"Fw?���Ei�U���V�䈐�)NڗѲX���)n�,�=d3�9Mʷ�L�B�,0[֔�4f���຀�9%Nl�������)6�t�c�dg��3��f&nQi�|��u����u����c�f�t�i�E\��Y�-/i�O�.�|�����&{Jf����Œ 	�!:d��������7��f}�bA�j0hiK���4śשF��P$f��B�E��	E`    IDAT��z�Ӎ��%������&�ev����f����/8�GS�*&��6���=z}����W��_�����޻�jz��Vv������+��c����C�L��H�8���։��3�j���I��(� -@ҿ��i�S�����!rJ]S#�O!ZW'8�y���Sx��-֗�t��5��%&}��\*�����Q�����A��������[᳣�h�w��sZ_����2���084$r�h�Pç12tZ-�����s᎕PV&s"��7jli�{�RHx��A:���QZͅ�p��Miei/���k<�}��p�������L����x����XF�tGjllE4V���^�wu�3�d���t��J��f5�~���4���!��v�P�%&w�=]��Q�{I����m=�\ 4���͕+W�=���5�g38Ȝ`veE����6n޼)�<����2�wЉ�r�"�OrP��WV�PΕx-d���tN�c�ǘ�����$�66���ԓ�p��e|��G��@�� �����ݻX��Uf1 O���E>�~Jr�j�耟��N`���,]�*%gr�m���e� q���9L�L�ū�x���Ѱ
f"QC��?����}��S�R��I�(�a�#�|G���'3�4�u	$�!��S�Ā�
�a��3d��C	yr�`�G&�|*-�4%54���I{e�r�lV�d-u��X=��ܨ�_K+��Xk�H�N�����=<|KE���X3��E�ϋ�)�y�d�7�4��T��^~�,�r�Q%Y�ij�`�m,�B�E���f1ɨ��-1Q�)���f$Y�i�i�Ś�TIj")*���+]@~�'˛`A���j���?w�d%90<��x�Z$-Ky��V��=�_����,���Hy3
Z�e�N�~���D9�h9jY���U��>�R/bF�a/[���az���*��M>�	�9�\r��_��_��0��ڃZ�!k55�lh[�dO�r2s��l�zn��S�!��M��:l"�c��EA���KKI��X��r�ˆt�"̿�jQ�y|	��)cqK"��p���B���C��@}_'�}m�6D��u�"̮H,p	�)�t�}�9�{��.(�.��%�_��v�������.�����������~����[�|�SoQ��$�h�o�P�0:�;��Ҧ}�DՄ�j� r*bܗ�����E�I/��_����v�F誳�����i�ќ�$������D.}bE�uI~�������+�ya�9{���*&;��Z�%Wb���T�澗���ޞ��\��3g�h��̄������I�0IF�`mgOE��F88<������o`�o G�x��%={��S=�y���ڱ�0�ׯ����o�Q�&��Ճ��A4�4�!��P�S&���W:���t�LL����tQQfG�M����8���S�Z'���|>�s�#�v}c�8�8'G���e�/����5���iϻ�Ej���+h��0�JE6���4�n�p��hFS��_�T����7�h�K��VVְ�L��*��v��q��%|r�&�:ڐ?:���8��w�3bԓ���7��A��X ��prx���!tvw!�!�r`�����>vK���CwK'�t��G�^1������3LNO���$\��S��d�P����n�N������&���=�{�D��K��~�G+�x0�D8�x ����M�-D�J&[��/�&�?j��Z*)��
���&goG�����T�5��c�$G[Q���i��IJHmdY�	�ӈ��m&g����a  ;?��R'GZ�:����(��soG�qK{�vĜ4x8�!Ɏ�i��$���BW,�|(y��V/lmbfm�;pFC��4 �� x?S)��0�1,&
Q62��"�Zބ;WB�hz�"��0�b�]:w���!����+C[$���">^��*���[
S�x�Y�.����=���ԣ�U^󖇾�V���ӆ���ELa���\(�g:c��1�؁&aH��,Δ~�@��Bݹ��}�~��q��b���<5������Ţj+$� sW�=6'�v����of��wr*��P<y����W�Җ#I�|��ߖ@);�<���9��T���i��csXd��a7��q��`K=�mI8�Ȼ�(��ɠ�3��I��6;����"L� S�x�9h�'��$���\��~�N���ğ���j��YܗZExz�L&:[�0�s
�}��jL4���h�OtI������a
�޾�-�a\�zݽ=""���bsu�h�7vL��-��`�\�JAa�4��P�b,�_�f6�ٳ�p��9�݃C��j�(4�E��/��g�������;w�4�a������E�+p�9V&MH��?�w�"Q�nqwL[��#畒42xG��x��<|���~\�y�������������?W&%%�$kjlFo� z��u���_��ي~Ɲ--��V�<#��޼$b<�9�K8�?����v��F� sr"�����D�
���&f&d*B���ʲn�Ʀf�|���t0
������b�xPܸuK�$��<��D+j�]&�C{O�����h$a�e5��B�����$�D�������wcX���A{��yܹr����X^���$f���/�$�q��p{��5,�G���DK[������z���`�v�p"
���CE��а���r���x;�
�K�Cn�����B�[��Ox}����8ȥ���[$�E����Ǉ0X�AD��$�\��T������*)�,yz�uX2�TDJ�� ��,��"\��]�͂~��O���׃��6�g�4���Ʌ����4%�/i�F���\^j3� ��HPb��$"���9��9�7��`X&�*���O*?��:>_��f3¯���#�y�A������d?����
^�� ���*�� GЇT1��ם�G���	��Ȃ�I�rY�0q����ו�Md��/'B2�y�R�H�X�qܣ��i�B�4�4�
�
 ��*��NSV����@������h�]�(�f����|~�,₣?9�u���'�ł�_��ω�E��y�D*N���!϶�|��R��<!�!�N\D�8�(1`�\�b��>ɶ�鵠mU�x�:�=l�'|�l��Ž�=m�\!۞υ�W8���I]f/V#`� fd\$�)���4 2ɟ�ǲ]ɢg���
~��"�&� r�����Ei�U����p����B��BK,z�+^��)���˯&��luw4��"��š��K�3x��!&߾Rf>���l�BC�a�X|��$���vaso+�;x>����r,���(g�l���m�-/aiv�Ô�ԭ�l��"	���	�MM�g�P!�����)/@�.]AgW�)��ct䚞�D(CcS����g039�s��	�li�c'pd�l3�������ޑ|�$�`,��8��vgt)�p�>�u[�	=H9a�p���On���+����۷H��$��ȽK<V����ho��ޚ�!�=__��/_����7lGo��N����$�r�0==+�p{k���6���l_�>^��&�W�^����"i���FE���蒼�TA�ZV��<tnݹ�+�.K�q@�)-3��w�{d��R�HC�����UCt1{#�qDNU�[_Y���*�6�dzn` �=]��֗����o���+E�q���ݭϑ����u���h�^���h^���:��n�=nl�2���slJ6�tG/.�9��b;X�X���8&��tpW�ܮ@�9]u�*�_�n�㼞V���\�0��"��j�w���&���)3��*�f�01ϖY���0�er���q�)�6�|�I�ah���DB���v�w�����H�p�{,�o���8^��D�l�r�;I�>5AƓ����~��-�&�
����3f	n��^ēI����g�g�Ƹ�&�(Q����>���9f{G�%�\�B�
X����Ζ�z�d\�'l�)���V�|&ސ��,�H��=���
�'"���C��L�ܝ�7p���*|VX�>���=SH���t�q���U�C>��:���*xOª*-L{UKw/(�֝N�y��?�A���5�lwmj��qﴜ��Z3��"Rytk�H��1r@��eA&���ME�E��4����e3��b�=QL�%���ޛ��G��ʚ>}~�>�"�dmsӰ�-5��of���>������gaN�D")��ޚDTj�y�XZ`��V��D��~����-�cJ���>'iZ�)�I	_���j��,���r~
��"JQrn�!�"�!G�����j�������WĈ�{
!/�>�ےl�����ǫ��*����J;����+�'��tm��}>������y�{�c��k'�"|��4%�e��u錈��	�?[��*¯������C�֝���F4�,�Lc��;LOLc���]>Y�-�2��EBF/�}���}>}H,v�����c�͋��B{�jEE�;,^0�nWr���ԇ��E`ymU���G)��0����l�锜�X����'L�Y�}���n��`_?����;|��>�{q���ho�����^����gG����444�.ـ��f��Q�?H�����S�]�������ҔN؟d�����Exwka�/�.,/.!���p��(��u���L�9	��������� �g�Q6�T��������yD�as�}0o&�,�,�r�"ϔ/MB�|1�tG	��#�Q�ɀ�yEř�L�.?�?�Q������mAO[3j��V��Sc��ڕ��WؘQ�{|�����u�����|p2@� ������fu+^�^��cOyʡj��+ofᅧ�U�z1#{fe׌��w|m_]��RKԁM��9g���|߃��$�(6������y�����P�����I���٤O�R����Ţq�tf����;�}P�U��¬��x���)UIy�-y*?��>�q�ͅ�.j}w����¬*Mkr��1�T�Kj��+I�ԕ���GͿڒ�d �Q�!&$%Q|	1��LQn6<��+%7f0�#պ�IG�P��̱cf�����Y9�-���rfN�''�lfNK�ht����&�Lp:,5I$�L���=y4�)��h~s�uT0H�4�V��I�����)�5b��-�k��g��2l�\|#�we�eT�E�^�hvg][��R1��J�ݶ߅M�6fB�A��1������9e�a�a6�F��$|���u�u#_���g~ڇ���+ޙB�*W��H�j�{Z��w��C�I��o��қ�v�.>�R@�BJI���k��m��iIU$�FX�ts#8��o�]	�0O�;�J��#ސ�9��7�ȉ�d��1q��b��C��L�ތ{��rnl��M&S�י�y}$Rn.��o�\�h��x�)�L�,��܀�9e�ߋ��L���Iq�t;�]�f�0�ɡ��bn� ����dU��+���!@�m�_����ão�X��^���#a��n�w;�s&'�yjN�B����Hļ��t�#�������/?�v������u�{pPׯ]ӹ��5=�B�n�G������Sg���mO8,)����Jfȋ��nn���d���J���L�\*����=kk��7/
�b~��Ψ+�J��"���4�dHb�c��ۯ�qYi��d����F��A_ʍH�cxi��ʊ�g�zM�g�����ukgυ���O�=���V��T.���s��[o����u�����{?uRo���&Ɖ�[ѷw��G��Pk>{�F���BJB�]6o��I���W.[�EA~��;L>���ޞ౉�:����={aC�y5��{��o���#�n�0���1�{��)������n,p"���49;���A�:w�$��t�t��5x,"�Ż�Dt"���fKl�Rls:4	�2�_x,�0�@sL�ݙ�����?���VV׃$�����EK�o4;0�=��.��+8����[oj����
���z����7��9�Oͼ��涚�e�q]=}�S�$��W�je��=&B&zB*�ʇ�R��]5���}�`@��n� L�V;�z�R9 ��h%o�Q�n8y�V>���Ο8�s�z��̠���w6����g�����f���T�����:�P�h�L�% ʞ����U��Q$�)	����}��	���:���
2F
<�����u|���뛛Z�\�V�l��xL�\V
qWF�TB͚�*{�k5�Y+i��0瀢��uBG@Z���-���dS�	�	�N�"��$t��y�}�Ξ8��L��4ﳢ��WY���	�}0�5�uC�ryu)�\�F��杽}�����N��Т��?��u�A�x�ϮTpk6-���R� ����6�*�{
����l:�"�/�R,r�?yd]�/��O�]:�,nz��0�I���`�ơ�!|��~�@� ��֜�W������@��������Y��%KPu�@��)�|�����a�%ց�^� $)��}�S�:oh6��{�����4[��NBje▩��`]��"�;�Y_�}|�[^��� �>�/��h���_������0	������W$JxoBf�z�5;f=�|��>�DO�S,����"@?��4��#[8��0�:���O,�r����-�l+���?��wj�����7_~����J�/�|������D���d�{|v��q�07��{��\���tT���}�L����B�-�"Y�t�]łS�p¢�{����Q��(ڷ�l|�HE`��y-��U_�K7��������U�O>�Lc���	���hskUw�|�_~��,-p��NI�s�������N�0��y��i��PW.�O������:~�68W���w����MrA����絻��SgOy�!���+--/k�Z$Dm��Z�� ��2e����5��ę��N�j��RX�J#�vt�m.]����� ~��{�fArHY���G��4P.�
������V�4F��8!�Xx���t9$x�pez
���i��i�	�j��aw�ӣ�~�M3�hz~F�^�,h�BS�[�����>�LLʥlPQiմ�����e<�qH��嚶���j�����M�g����6�@*C�%��$�@ZV.WT� )�ҩ�o��-&U�4�Ng������JH��6���fϿ��MKw��]�y�IE�� ��p�ZǊ�(�hĆ8�C�;�t6erEx��1u���liuwWS�nn��%m�l��%"u���q���^�k��L��q�!�lZ�Bg]�|�nӅ�ʞ�`w��U˞��-0�ᕗ3�s�6���h��ճ�ލ�t�w�.�+�ы}E��sav�m3�9��Z�{)mm���/Ι���<�^�{�;��uja��C����ޒ?b�q3~	�������A|���tZ��>P_O�'B����-ܔ�O�����,������Sk�m@#鄛O���7i6h�{��X����k���;l�)�1'ja ��Ղ��C�N��a�K���!{�P�.@�{W�N���#:���=�ł���\S�� �v����V� 9g(�L�9�����5���/4����LDʧ,���A��I�8o9g�F���Wq��9,����r��?10���,Ĭ����o���73+�W�.¯��d��ɗO����1;a�|8�����w��-��{�{H,��"��!/����Qm�[�D������Ą!���W��n߾e}!�&đ-�N�@붵�J�XHG���_�4���f2���z=ة��1�P�)d8`9��Cχ�
���B����pzt��q�=���"7���Z������>x�-���M�t������ǎ2<::n��ѱ#A���>��C�,/��m&�egΎ�N�fV��Þ�Ϝ<eO����2�[�0�xK�;vn2R��2�V*&y�=�f�t�v�ӯ^��ύ=��=O8��`��?|D����ʾHu�)쎶Cʀ�G&R&tϬ](*c|���r�    IDAT2�v�y/@,� �"�
V�!��_���C�@��ޮ��_~���U��9d�2�N4�	8��Z6ץc�Nh��1E�)'(�+5�/��/Wй��z���n.k���N>׷�51r:���s�g� Ԁ6��1� g6�v�F>�7��  �t"�m�C��MFv�P�����Zq`<z�0�'��zS��y�������^U`չ��yEK����s:�_͖ʭ�Ӝ����
9̚u��֐�b�p WV�`��0�x��@����U� ��Jɤ*�J�[��M���{��i�fyc��,Z�H*�|k���LC���/2C�&�!1�F��nԵT�1�L�:E�C��Z��.�nj��+��c�f��:P� �t+�7�_��o�Й��� ��.���n�3Y�4�;���Ƚ�L���f���QЦ�ʥ]�nnx�\��P������4�@�L��	�n�~�={�/'�RsqE�<3�2���x^�l�3�׋�)��@��,���t�ۻ�d'ܕuscr �0����N�)E:�P_W�FF�}ZY^����?��u2��&N�Iޥv,S�Ʊ�Lx�3^(>��(�|p5�%f|r��#F�c��ɇ׍i��49�WV�}]���ĭ���>�㜱�h��\�yC��^-����[_j����DX���n\�[-w`���W�����I8W&SZ!�g�{�{������3�(�͝�.�{��߼ZZq�v���AS�s�t��o�ͭ/�����U2W:���:��vVμ' �Yҫ�yͭ�*�ݣ2iF-��.b3���܌>��}u�k�>��Qw�3s�
D=�T+{
GT)��I!a�'0�F�Kn�:�}���\��@β�6�r�e�s84��P�Siǰ���v+ѕv�8�f4�@/HM((ཱུMқ�����@޳���`�O?�Lc'-Q::vD��|��~���I�IDS� ��ӊ�c����q�"�,ө�'t��qO��~s�$����!�
,W�}>��g1��K�c!����W��2I�/=��ԫ�9O(K�~��ι���=j�04:Oj,�|>�aGNp�xCw�4�.�ن���,�B���a)�5+k5$�E�Ц�@c��4�-	� <cyQw���g�/��F�m<��N���)����[�����S?y»���5���6�5�7��g.���ok�حrs_�=��|�;��s!O�}rtB��V0��\�Z��E�f����������Y�6} X��E0UT�%KX�P�a��l�c���7��4�hl�OG��4:��Fmؽ��,hiv^k+�����B�a���.E)L�D�F��)�LCe��X8��K�FF��L�=7���|�39K�q�d��(ՕS���ؿ��7q�p((�)�-�4�\;l+�Ʉ���R�=�:�$�\F����ǖw���4\#���(Zj�<��ꆖ_L+\�aR��VD�FX7.\����a�p����f���:b4�ɔr�`o��l��˴W������� I'&&���֗����fi�|&l806��8��0CQ78gн�c~���f��ٗ_�;��0��M$,;Z�b�쳗/��C
v��CM�ΘD	zǤ�����=���%E�)aH�Já��$�����B<P��H��F�47���h4���Ͼ�A]"����(Fcb��t&(��.��"�:��v�`$��Ҹ2F�`�CFc
��� ݯ��������c��t������Q7)�7<7��w>�����Z)��wni����H[�l0p4E��N������m�E��� �B$a�����pbp��o_o�ON���[�r����jq�rW_�]���M�v]K�szp��[��e_(j)��c'�&����"�4 �V��=~�R�dJ��\���?йsgm�����O?��~�����b��1�ϫ��Z�QQ�������w�>~ҍ:6~�M�_���σC�8o*\?�G;{��]��L�Ň��v}G��3��=0�z����G�e���U��\�9������Kk+z��~������ѱa�n�蛻_��_�º\v��rC��*�f�7+-��G�F�-�/�?V��O�S��/�����+w��9;p�!�� ����2���L3 �
��P<���}~�Yߵ���Ke�,/;F��b`xXgO����$�`M���v' ��0���	,
*)��pL�AM��_����T��64��G��T<b[A�W���T�Z��"�Ӡ�KA1���]4�fXO���P�6�17�d��n���w._���yGC����*���=}���>$i`Y�u�	鄶'�ֿB����t,=@.ܯ�{w���#R+H����<:~�!��.���[
�+
ժ�\�HT��.?�Ѿ�ND��L2+s�\[7�]L�:i3�A"nb�QwpE��K�83(�r��!����ףQȓ٠A�U	Sh�����Q.�"<xtT��C���R��Ǝ�VW��KLX����;F2V��0;ڐtO�(慬�=EO�[��wE��F%`�c|adS{�Zx>e�!�h�*�0M�q�7.\�o����g�S@��������^���T������/P7�l������DhqzZ+�s���Z�n��>���M)İ(H@Ս>�g����$�.�_߾�$6t�>S!�K��ď��Pw�f��Z��@Buc����夝ǐ|�D�'�f�G���xn3	��i�Ȩ�<d����=�
�$+�����ps�b�Iӂ��[o�冔�t�իW^=J�(����g
�^�t28�0�$���=A�|�, �r�(n����s��d8o8�v��922������v�Q+y'��n��
Lt�!�S�5E�Y�I��mCT!u��T����ha��3	��۟^����^\�T��wWtpP��̔�|��j�J�5�5�ѱ�q��h{�D��x�hP�q��E�ƭ+%��/��/tbb\����o߹�{h{�`υ3�(���:�3EY{�����t�6��K�����������~���#Q��?뼙��Y��Z�{U�S�@���H"��5:0�j��'�
�9dӅB:��$��6:��~�;�=��7���#��\��o��/���A��U*5CVhJ+��JX���ݫT:��hH�į��ޟ|�\��ZZY�t�G����R|�0�1�o5mx�ɍJ1O@�ù(���0!�W/����?q�M?(�h����|a��|P؟|}:m��t4�l,���kS ` K�Ч���;t��т�gf� �*�vN ��jے���ϞjqiY���FG�[5+��٘�7x�@���@&R���wT�.���q�{����f��{���[_���\�h���i��kuw��%e���{�dʓ,�9�Y�_+OK����A�d뻃C�Z�	2�Y_Q�YV�ZU��PO"���]=wFC=����AC�3Z��5<
�S]:k�{_���jM���ql�TY��bq�q}�V!�1�`��I�@_�z���MaNS�����KUO��V���w��	�����]t@z�&���7z�G;5
�-F��/�o�ؕ�� ���|e���Y��]}��ȿ:EZP���7�hv�4k���c*��m��,�p��UZ��3�s���MP*0�q��@fv�H#��ɉq��2z�⹦�>�;z⤛�|h���j����PA:����546�d���W��ͷ��oy�D��=�H�d���;y���8�������B&����\���W��&0�m�@��/��@3����N�O�=��|���ڕ+N���75�B�S/����:��P�	y������~Y/^<��;ap��&M�w���J�z�)#��lh
?�p�XPO�ǲ�/��b�Y�@��=h�	���67\�9GG�G\�3��ڏ���4���m�鉰-kA�@?8_�02�{��~��J.�T>��l6������o��O�������O��/S�K�u�u���y��BMM>�>������V���ѩ	�1�1"���ۖ&�ե������\��w��|���J�ǎjd`H{;�&���\S�N�"N'�D+VWع�U�onn2����F|�Z��C��i���1l�l9P��n��8t�A��70dx3],(�M���W��7 �3'4R��;m������-/���g���ub��{���j��������b��ۭՕ5��<��cZe܈8Ds�9j�򅜻�C�	t��<�ߑ��g��d �Jӓ\����h��M�
ˬ�6,�|����Z��>Ϟ=k��}P_Ө 4���D�.Q(8;�T{�v�œ�G"<k(�L
��kGJ3@!�=	��T��)�N�\H��f��&E�.�`@]�EDLV�J��Y��ĕ!Sx���z@>g1��}��7�[�S�����������~�i,�0��^sOB4a��y���"���
bX����)��-۲5@m�f�F"�e�;�^w~nV�uEu�J%��5���0zTg�G̈́N'qM�jvzJ˳3����29�RI7��XB;�������,t+��+�J����m;���NG���Lv\�T6m�T�?������JZA�ҕW�+�D��l_��ł!n��/-�y�U=�ƀU��DL�B�C5��d�V6�DwAIHZ���jf6�خ�������K��t�tU�Z� A2���Ķ��W�J�RM������\��ǹ�?��?W��[��_qQ���X[�d��8�9|�˛[�x�Ό�k��G��f�����S�d�2~��0M?����J>wےG��щ�8yR��^=z��)lw�����=8J4 p":,硱Qb��Td�:z�F��+��krf��Z��D�DR�0Lb��2�b�W�"��J��ȄΝ:�b��ɓ��ȥ�I8��NOz���-��x����KW���W�8������ܢW��CZ^Y4�ȳ���a��������}�4{�8�O��Y��/����g~��݆��_z�� �n<w|.x���s���?��@p)¿xG/6����"S-"U#d\C��ј'��"̔�c�z>��O<�����G}�՟���۟���'?5�|Bp4lP�*E��ݯ-S����j����1�w��8!#ӑ�^� 9n�?|��3�Σ'`�֜�����g��@���bR �o�_LX�t�� .F���#J��N\�P�($�< ����`�#:KrD#�v�˚�J1br�Wi����m��|4�l!�ѩ�K��6.웸�a�S�[h=9��a7�>�G}d������2J�]ݻW��/�_3O'N��ܬ��ww����=�Y9��U��Φ��z>_י�Iv��'��v�	l�`��4���ú������>¤��HԨ:k���`.�P���0nz�W4zd���p��IH�=X�����AX�X�7r1�c�U�0��ް�?�JK���o���	�֘��V�� #ܣJUC������i�[A�@.���p%h��� �f��K�l��ҕ��FwC����bU���l��="Л�m_�ti~��wM�b?��}�$�6�h�W]�)������h�X�0��P�h{sM�k+��n+�fMx���tJ'`w�+�EZM�R���e�6w����O&����,8�N���JE�D[��khX�B���x���ǰ��#�>VSq#W�h�ˮR���j]���RŢ���O�M����jc/�6��x�_��i��0̻����U��V8��/�]T��e'8���B���xi��N ٭�݀�[iXB�0=㰅�"����╆Ch޼vUo^y݇/��>�PSK�ޟ^{�M�ym�&�χ�9g�5de(�}�:c�Х��i={���4X&���"A�7�5"#[6�����Ǖ��֣��t��}���vD�|�g�`�10��Y���0:\�,<��Y?��S'�Y���;��ޱ1
E�f�6��b�k,��l�ΌOxG���ӧ�{��w�4K0���q,��"8�� ��N��勯9:tceն�����1P��	�����=8����9�0c�j���MG��� ]�#��$�Iu[�tJg/����q� < �����y��7�������{��)��kG���7��Z�Y橨Mb(­p�;/j�+&b�a�?�I�Ts���0f��Yg
���������?{�ދg?���"|��Ew�/&�����Nn��{��:꜆���+�A�\�jrսG��rnA�%�0�29��'?�ٓ'��]� ��xD��:c�꽳�t�����t�̴�~_m�w����65?7�����(�,����m��$5td�nLRa�2��t���V����B":4�pf-�՚ai|��I��7��,=�{��޽~S?��}?��Ү���V����7�3$�4~�@x�}�(�a�M��h�C:�Zϡ'�'�cO��Z4���,Ԯ���0��&c�E�]3qqѐ���]9%��A�I����$g�5Fb�/�8��:�1�i�I�I*M��u�Rv�1#�>��f�b
e�0]�]34j{B2^���/HH��(u���Z��I��s;dM�5�U�z���CC��{FD�A(�˱��L���4����������s&
'�e����C!��{f��,.�L������Jő��݊vO�y�E�mo۾@�r�� �B>D3��H��X��D���P\#ٴٿ�J�Ȕ���̔�����z`�g2>H1�	�c݄�\��ΞV������1��m4����im--�'�D\�X�~N�x�(H(���qUk-픫Z�+yF�Ո�L�Z�߱�E�~r���ܰ���'9t|����Ąv�+/���V����T\5��T��\hf��m�nkm#�P.���R�Y���NÄ~r E��ɓ���z��5'O���Ň����'_;��gO*_,hku]�dq�]]\P}wO�O��XO�F�=�OjciIs�AXM&ig�C�w
�����517��ޖ{���ѣn�(�S�_X�N�
Î��h��u��[C�G]��d�f���D���O�SA~4��מ"܎��	$>��vX�Hʓc��i�f?z8��h�Pn6����iV&k�
(�@������'�D����Ea� x5GF��̡�ý���ԉ�Zr�S�!��10�A*@g,���}�C�eryg_){�75�J�[�����O~�S쩡�ܿ���u��j��<,��0N�<�LÒ���+�	7ˤfE�����cП��~,����Yt��ǭO޾������_� �$|����$��<����-��]D�=���'t|l�&��8���\.�����sb�Ly?��! W/���#C�c�H��~��"�(8��Չ Cg2Uy��k@�bQ�T}��LNiueŖ��6>P�����	�ᘬ�߼a�7n�q3])�/�5�0g{�$4�o �"�Ih%�th7>pK�t���!�	y��楫�˟��>�RyG��>�����4����m�]�����c�}���cZo2��f��_ڱ
2�fgB�:�+�����!K4��Qh����tT�W<���I�a�)�ceB�,n���x�;\�%��L�D9D\�H��C��'1� ��_w���V#�'S��ŕ�� ���*�D��x���GzttpD�LỨ6^�	1����p�H��!�Q�L
m'���`���F��m˯�U��g��}���ddavF[˫��ܴ�t��ם}%B����S���Zo�Ϗ���8�51� qh7��/)Skh$����ɘ�q
K{�[z9��{s�h��nC�A�c*�BZ����Ɩ�ї��{xX=����+ssZ���>�XD�����9�/Ř\�jG�H)�ɫ\kk}w_s�kj���$��ޮV�ƚ�kjC&1�HG}��\y(�UP����АR}E���c���Q,�Q,���ț�Z��-y� `[;���xͯ--����v�2�ׅ\&o���g��7o�ʅ׼�@W����Z�&�i����#C�p�5[������t���CC^?w^���䴿�n�0Sr46B����'M?��l+f    IDAT�:� �	�qi���}>�J34o[�L�l3�?�< �U+V%�|�. E���8rtL�N�u,�a�ta85&a��@��M�,\��jݙ��?��g�)�L����zxﾑ5,w+�&�i�����	s:��Y��ft��Ο=�� ,@ӿ���b.)�|����(I�|_�@�+�G����`�0���y?�{`��x��{&��u)�=�s�q��--�3�7����O�7:��PS��wKS{A�$��j+<:g8M���ݶ=�a&a�z�fK}���C��?�o��̟���E8_(����t��%%#=zxO��!E���mr�/�SO�G'Ə��7,����bR����d�v��o�ʵ�z��t���Jň�r��O�b�%S����6j&���s��VJ���鼝���\˯��*�2ᰊ�L�	2ɚ�^V*���#�����ßW!ݝ~��OjfmU�ق]���
����5m� F~)�Z= @Db�
�m��o�����G�s̓��������8����Q�����4�M�&Q�T�ʏ�LN���Rؙv���(A<���BM3!L��N(�c=�pg�Ŏ���	�μ��yL�%�F��!
<L,]�3��{HW.t��2		�7M� ���20��a��ZM�m\:�����C6�o�[j�L.�؝�������5������Ⱦt��f T,�gj
�4�8/򨠭b�j~uV/w�$�4��G��/�4����9�&iʀ����@ɠ H�؃��Mn��k� �*i �[�p�!^�}�PW*����=����Sw<�L<�f�jr�����]�˽���V;�(���Z����֞6Ke%����*���i�]]Q����\N�=E� mˤݨ2Ѳ�!�;�+�DT�Ξ��T�Q����,��& �<1n ���&�d�i4l9R#U��㾂
cG��S~xH�ޢR�E�!i���LИ`�u���^���>��zr��;{�ޠq<�pT֥�g�+�a�_�[=�|n2SW�n�wӶ���^��4�:�ݣ������'4�7��tF[K���㨗]�!e�����V#0��Ou[�ۖw���8&8�664��dLo��{x~�ݽ���5;�5ba�5���Ő:�9R�F����׫��9=x�PO�&Ռ��s��l��K��u�B��9͕�t��K�;ȞO?�� � �'�e`�?����E�Ƞ*�����uI�������4<�AZRZ�ˆ��3X�g�U�3Ӿ�![�d�i�'�7��o\�J�����ŵ�V7ֽWF?�D�dBGG�����9��p[���+��]��AC�D�E��0~�V_���� CP�x���J�Mx'o�՛�~1���O���E����������k�|A׮������N�鳇�}�/�ww�g����z7�"$�Z�@_Q=��hz��f!il�(��jys�E�ĩ�z�ݷu��9=}�Xw��ѷ���.t;'�����'�p-gJ���0���:H?A��n��X�ts��w�=���F�$����0#�٩�#7�m�t��C}���6C-0��?�f15�{kqE��˦���aBR"����^��;�o�'�`ȅ�:����TK+��f�}��06
�c.n��V@��<�6����=g"�HR@�A�8}�8Q2��S�5��4R	�Y�t`��r> lx�βS�76ִ���Z�b�"�j�zlsm��k���XT��>}$���:0�m>7����=uI�	�� ��@s��?$��&�����@G��u��Qvt&a&�ΐz(q��ަ]����� Ӊ*���R�%L�"@輾���)�n$<5lhn�V�W�����ֶZ��z�q]+U��t�7���LT�;K����3P(8�Z͚%C��R���j��׉��a��A[���6����1�A�
���=LۻZ����Ύ�p�I��u��UcoW�����z4�WTw.m;Y$%�u���"�{�9��W֋�ymV�~6�Z�����bj[�n�y/������OQ�����U��c��W��w�Q���!�i C�HV!�)j�}�n{j[ZXԃo�hciū V�Z1�ۺx��S���YkW�w�R�>������}z��w���K�\���e	U�6\p=�B�P�+�mY�� ��:�0˗���\H�[��Z�F�|8��jE5������޽{Z�[tW�����f������(W����An��������B:d���Meu��]���'a�Y�ܗ�����	N���9�-$����m[Qbt��iO��ӯ\�==�,�i�������B#d�z	����ߐ�G�,P7��>���3.-zEg�~�1�$��Р�g��>C���~�����{�S�'wV�A�p�IS�M�eP#�C�!������e"�m%���t������৯���_���ƷϞ�����kx_�|M�x�Iӯ^����mֱ��a8�wdxT'������v7�T��4zd@�B��%���/49;�H&�ͽ�ַw��;7�����B:���?|�����-�ƺ?BÝ�ޕL��'LMm
#�(
ց�Hd񾰯XЉ�����hbd��0h/��@rbǐ�e,��&����������sݞ��|��]8���@;����VU^߰-�<@��X�M Gyk�E�G|���N+��zzy9�\���ޙA���G*ż��^.��d:��ń��D��	K8���q�r@-i`��L��L��3Iy�.7bF/0�H�Ę1�m8N2��1�7�����<��9����NE2k��ίL����=]�!�P�׀�5�7�*�'��-�x8x�h(ju�=�60�ggw���c`b��N8�y:����,&�8�)��iH�"���:٣b�f��H$��������t
��Е�LM;_x�ù�^�+~-�����r����q�bW
�a�tǿ�C�Ol8��U�W^H$5V�ֱ�nP�����uF�ݴ�B_��2�D8��NC�S��fG�Yq��J���RJDv���Ry_=鄎�i��K�LRI�1�گ���(��R���v���K���/iO�@�J� �;��0�MpY_N�w�=TH+;<��谆ϞR~�O��~E�)K���~�#q�"+�M*�2@�}���z������Kj�*
�=a�Z���ɓ�~��n�������w���=���.��n���.�=}����0AX��5�!�4Ec�����F�Ϯ�D�s�6�����A���dj���1_
6��"$����w���²6V7�s��
$bf������O&u��)��x��e<HB����ZѠ s)VfX��m���t��(���W-A����W_�]����R)s'Pl�H16�N{��3=��Y^X�Nr䦰��j��y��4)W<鮮,��}�^X#OCR��f��Lkgg�(��ҒM����@w�iOL��	�2R�~�����qU�!���z����v=�	c�d�p��3,q��^G��دyw�QG*V� ��\��b�����{������z9;���k�����+&j,�����[���O���LiM���i]<s��J�`1X]�G� �|N/gf4���h6�խ-��y}�����;7�}��W���7�u箶I� �f�pe;g������)��a�z�i���4Uw.�������.��
*��}W� =�ܣ�E�oW�n���+=�}����z\�P9�4)�S0�PD�VH;K�Z����~U�(QL��@�SN��,�������S��1z��x�O*�3R,ң蠁sv�����.�-��I	�SO{�;�0��1_���f1i˻m�r��U� ����g�+���Ç�ꛯbP��Q"���@6�X9�����OCч,��	�Ə6���LR(��ց�ÇV��������B����r@9q��?�ǎ�sz��L+h2�A��혶�{�t�I�i=���E��3B>�X0�q!M,B7�z�g���2�[�����{e�J� ��Z�G`�v�a���)@�n�����k�=��ha�eu���M$4��h8������V��_+G�Âm0�L�}�'_�����7��� ���>�<���NT���%t�H��z��&��FD��i�DxP^\{u�h�Z���f��u�Q:P�	'��<e��Qs:(�Hp2�43	Ez
�S��:y��NY�IE4 ��'KA�� ��Y����T�Ӡ���\^����\ZQ�TV�gl���N���˺��u0�����a�Ǎ�-����K����M>n��u��憹��CZs|"����J�j��C" {N����c=�=������4F3ഐ�\�,	�Wl!eu���B1c+<8دg/����ֽ����ߙR�<�X3�\"Ƀ!�A���������L����O-);�qJU4�\"a����^?{�{E�v���%��3�~?��)�N�Ja�	���z��p�� [�?t�x?�e ��W/Mf���oha}��C�C��x��������?���M*�~}�͔�<	S���0�bב(y'����Ύ�hM,jAa���~w������7�����|49�/_�-^J�3���M�u�RѨf_M��_�ޝ[���*��"S�v���Ə�����ʲػ�k5�X��D+�P�Э��u'��
�����^�����oo�y������T��F�v.�C-۝!!�7�C+ܢ���%Jf�N׋;ԏ����L�0Ѡf��L!ì>�#�4�=Qjw&���Z8�h�U�Nݧ|�9�\��J� ��icnіw��Z�����w,7߸�����:ylB�v�Lfm;[53tn"y�X$�R��*��z��$�0�.LX=�ФS���J�����<_�`꫹����5�#zd���i��S����=y�<��V�{=XݵF��?��CO�	N�^��h�aV<�<l&އvUΩ���I'�D������9���q{m[���Ɓ�T.��epV*�L���y�J���igk�D
%�0��JC��֡s�E��T'S�{'���<�C�ƶj;;j�1	��2F���3�4�� yo�b����	r���B�F��j8�'`��a�A��;Jd�ޫa`���ܬ��KZ]Yv��ԋ���KD�)���r]nL0�h���*�j��K�}] 2����JU&ڰ�ܯ����Ե�W���6�U��>���+��M\�ԙ�QO��o��2J��wbL���48q�p,�	��p���9�L�}��z�Ȅ��<��bi���FZ����b:���A���.&L��˿s�'d��#��2R�4fav��I�֎�:6��WhԘ��?T	mȣ�IP��A�g��'1�z��>��aex�Hã�p�Cr"��"$&%[�[�}�y��
�
����|��~�{UPt��#��u�TBHzr]��~���yW��.��<y�-�W�T`�y��f,g�)_C�@K2ԯ]��;��*s���3zo�q�#�?'Vl^y.�����S4��uD�D�;�jfn��3��4�\_>~x$�]_���9��d�ӿ�K=6n����Ջ�m��������	�UNy��X����Tm�<Pt��8��|�wǻ���%���~���S��jv��"�����A�z�T����o�r>-�]4z��
Yt_�6"������?ob�}Nٞ>g�n���|��n\WoO��˯�Ч_|���y����:�9 �����}����UW�����57&n��g'N�ıq���P_w�{�V�����F��X�ӕ9ݛ��\e[��k�`q��fH�xFGr�$�"�uD޵;��f�C���Z�~5;��W�E����u�؄2� *�V�(ly� v��N�
ņƣi�x�bK���.4�@����8�!�i(�����ΊL����äG1���DMn-�2���e�,�;��ɓG.�x�����F�� ���&�����	w�a`$�gZ�
&+�H^���q8�k�=����7eP1�̎�(���@8y��N�>�޾>�:������t*�C6gW#�1���_���b�fm_��0���4�6C!�+���x��h�l�ݛk���E��w��
�(l5���a�w�Hu���#��^iw��L��V*A�^���i��u O�G�E��$�گ�����-��*�}�Twv|�>�����|/5�;H��=�9�����>�%%��t��[�}E���7ʪѰ���+�ʨ�k����~U���Z�<�^S��O������@��D���HF��Τ�/(=<��cc*�����'Oͼ�U�d���|P��EѡV3@Q�9�V��`�%���{��D9��o�q#(�K���/���Y����(t��Yɰ{)F_;	՚�T�bH��5Ӂ�t�<߭C:�������R�{��Y�xe�s�(�F���ȽJQ#Y�Fx�Z�Ԍt����׍��5<<hB�/~��>�����Ҁ��xD��d�Z��!����h�L��5��M���'T
}���������ٜ�3@�=�V��5	|���3C$�(�!�	�����Tr~:g M��㍆e�7I�����3�7����W�6#�������0;Z��L�������}Mn�h�YvX�����AgܘxhȺ6T��Tu��"�u¨#��;W�|d������?�ӳ�q�z4=��^�-^��v�7�޵��
59��E��O>��O M���5��9:Jk4�Nqŵ���ì_>���ʆ�K%�{=	�u�u�vw�����Ol�M$TTIPJq��$���7e?ā�_�������E�!nM��P�� ѹS'�4#3�q!�i����̔��N��ƒ�J[Z�Y�)��j��WG{�4�3�#]=�g�#˒1�jچ=[�q���e=y�B�}F��1���[.��d�0�̫���޴�9���~��	��1�@�%�AX1Ӓn���dɻR��t�}J�h�^�] F'+P�I+���֮��L��a�p��i�\W�\��¢&_��˹iw��C��@@�H,�1`�t���z�̞�u8�P�$�t���혀�;;ndV�����冫	iG�̨X((������������m�G����҈�$�1(�%�r`�A�N#r�Tfj�}f(��ZY�h�Zj��ԫZZ]��⢶W�=7wJ���~`�!RØ���k;f�Ih�ݒ�'A�j�IKw^&o6��O��$z�R�H����n�GX���0�ȧ�&���� V�z1���͠a������zyOU�����j�X��.{��L@*��%��gsj��ڨԴ�S��ڦf�6�^���;�T� ����a�0ۈ�Ů7�T����H��o�蠺)ty� �}'�f���a�Q�AA(¤��,�
�Y�O��Q���:�/�v0�h�Jӿ�l���˗=yQh~�ѯu��CM��;W� ͱ�R���M���Z��<��)�K�>�	b�y��!v����1�C*��I�"dw3�� |<Mw
�Ѭ��k344��o��k���*E���Z���wn(�Y?�懞��X`���)��E���[vic����#ݾ}[�K�P�'�ɚh��{��l������|n/tL7xݜg\Ok�C2�N�o2�WmA�qH2eE�?�g�h�l�f* 4+˫�[Zpd�e�ɔ_���ȧf^igO�d`�<~�'�/�?���U���GS��Ji�#�d���0�u�I؞"�h(�i S��Xo�?�n�d�ON��ww?��`��ϧ��.'�Y�u��^?wI��^�L��{�����x�ؖ�y���8ݪ}9>����IB)��_��Ɩ&g���������{z��Օ��S�>����\Q._��ɤ
���c��և-�����gz�౶�6��ID���hܾ�����������OjttȨ 4S�WOug��V���+��Z!=�3�'5�=�	�M*�+�����I�l�N�����ԫ}��_i�o@�_����ƕ�F����'�ի)��v��rȲ���&g��qӅ�34;�9v-(v!w�LT�ݬ��Tx�N���    IDATA� �LL�@9@��,o�&�����0vdD�x�2����E=�L���'�h.�h��ɪ�w�T��
�:<�3�.�/�ot�uFr�q�ZMX��z�pu(�
E�G�ĉj5���9�s�6;��|�S'O�l!��5PWi���������\���\r�?;.��'a���8�G��!0�I����L���ʂ� ��*�׽�B�e5��: y��09ˑ�m���2� p3���.kv���	|ł}\/���jjonk0�ёB^]��b^��r$jL��{>L�7����Қ���L�d�Z������e�j��Ǯ�;=܁�1� B�EY���������-͐�[%���"�d=�Y�`t=�R+��A!�F�}*�Q�ȰR�J!�;��	W��S�-�l�t�;gy�&]h­�G�����nᘆrE��J����Vf�nA�{M�!�S���� Q3��s�Œ�K�%Q�L�v��
j�x��b���x���l�Yi`�O�0X���L���4�k�
�¸��<�4�@�O4��+����u�Q�I:24��ǟ�^����+X5ID�\;Hj��}�.u��6/�z�τ�/_X��5�{����9�h�Z-�/ہ ME��f�05鰰� �r�}8Pat���`R��ݰw�� 	��3ל���߷'|��L���E&:��+�׏~�#;}����Gv�Zm�8�S�1�:��Z��9�
��:����8�i^���;Gs����ޏ_�ɋ����'��|jn�J<�N�MݸxU�dJS�^���;��G�R�3gu��5�)�ʁ+��%K�!�� �.����K���u��s�I���[�ľ�+����g&�����ku�ƛ6����J�@Q��
i�T�_~����w�:e���iػ�.�����u�����˺x�Lp=	����n���G�7�B�LT��M-�l�J���˺|���a,�}p�)��T\�$]�h���`ls��([.�����k={�ĻI��}O"�9��� �&5q���9��5��_���]��I ����C��[��Δ����/���A�N���'Փ*�M����>��w����ړ�[8I{�C�Ý�!,�`��v�@���6���I���M8�� ����c�IQ��z[���f[�qN�� �->�ǵ�*���O9�4_��5 ��Ҵ0�atv��)����"��R=ᡵ�������VVTZ�R8�\��p�}=�E��I� k�HX�t�$���VÂ��<�i�r��1��:9>�n<T�jkzF�f�:ᾮ�r��
=E߷���	��������l<Q����ˉF����7ٲ���ڒ��}����]t5���V4��VL��o�ii{O3�����j��}��X��\�Ƥ#!��:ܓ�	C����
c��UL=��ң���	�F >k9�M5ZĢ��������#*���4�)�Pcs[��n�.\��]���ₙ�t+[�k�À{���g}r�5l�1v�8���~�?& i�؁�>�|Ûl���ш;;=�W)�ܷ@��OA�=�&��$}ܣ�P��J�^���g�o��6�}�Q�Y��C�%$+�`|��xKo�D�>|�X��C�/��7�/���f�l�TV�\�󋉇�;��^����z1���?��N��ix�Qot��|ft|P�]H�6Nxa7�u���v��?��N�9�Z<�/_<ҋ���	GC�ƯP78/��qX�魀��{���hZ������|�?��?������W�~o��ϧ���J}��Ε���턿���9]�xQ�νf��V������(\!g�r��si�{.�o���+ᙅE��轷oz/A���+=z�@�ZC�Ν����!�F�;�h, $�{W�^���}��~��o��bc�X��-��T^'��ҋ'�������{Woݼ���.w�w+Z�Z׷/��〉���+�Z��S+���3�����K1e%e�H
�\o2�t�gisw_������}dx��ӗ/'�����^���{�dJ=�^����#�
�}�إ�gN��wnؗ�� :J<]�ǀ�����{���SW�S��#p{'�I �%:~�I����g������ǎY~`�)� ���|�>���;�0�� \���0�N^�aW�ק��>u8ɘ��Dv�L:5����h�iQ �q0�w��e��LF���5�m����\�t�.I�鹫ƒ�R�f��'<	S��b��?3>�.��i?���yJݐ$�7�k�_���
3z;�SkwiM��M�vJj��-޷AL�,�F�jӰY�̀pЎ�0��Al(�m��/��?�b������*Ѩix�W=}����@�	O94g�r��!���Z�tY���F���v��u��z���1ėL'���/tI}��O9RrqmK����]��������ӨPt$ p	�1�V��W���9���~%���W���P:eG,6�ޓBLt�� �7������^�+�B�栤1�,��i4S4$��k{qI;k��(��E������d*?�'������r��f.��)�p���EG[8��@|_@͎��yL�M|�	4��~������$G�~ќ��
�������{�H��Wb'���0�MUVeyo����tO���H-��(�A _J�A+,Az$ Wt���j��\ΐ��3=�1=m�My�U齋�p�ovK��~&Ѭ���̈��������%y0^��.������(�]�k:�^�6�٬pMG�o��^}��p�ӟ��{��H��s�;a�ؤ�>�W�k̓h�+�UB���d�5�=��W�y}�{�;����^H�eAՄ�y�m���m�Wh&'s:���6�|O��9ɟ=52"b�O������y<���N�l��!�~�׌�Au������G;a�'��G#�����7��G��"��o�����?_�ظl��n�XX���۟���Ϥ�d�(!i$��U-���ں|FE8���G<��E�����6V7�9�a||/��^�q��(��V�t��
GO���)Nvd&�v�zL;B��.��w�y���/���hf���:��?&���&k�V��ܙӸ|�<Ξ9yh��j6�`������6����p��F��BjpGG'098��?,�'ag"t���!�@�ü�>�p��m�����`d8��ح�M����`{wKf,D&�&u-�l�n ��EL'�;�΄�T|H��{zh�.#��2�0�Mt3S.�jie�#�C�'a���=~�����n�5���a�qA�$XdkU��l���<����l]A��R���D,8��7�[��bC-��剰��âc��M\�ދ[�qv�MT\�jKA��h�'Ο>� %Rp����߇א׏ё�>}R׏��m�C�6���h�O����{;�\�B�E�Z�N6c��(�fP�Ϫ�(U���al�pny��e1��ڼ$����t�ǘ�sJb�¥Ku ��,|v��p5j�Ej8��!S���DhP��Bvc�}���Q�UX�d4�)�� 	st(��Q�����~2�d*O�/5ʆ�C�dź������W��p7\���-�ִ��<pz�����D|t��4��i��X��A��j����t����O6��5Ԥ3��2�vKEX�[�K�I�5%%�]']'F�QLD�P��P��Eh����UK��:���pL���iڊMa���TJb�����Z�Y	Țr6�E��7��3Aݣ��Y�8��Y���\�ƹ&��g�o�~��'�X��<�X��/�j~����矢LRf�D:��1ם��r1�A�E����_�׿�5�?$^��ч��fS��&G�]�������43z�۹��q��Ӕ��0�g���m��Ȑ�"��	g\�h��v�@��;2��T�C�d�D��:����N�Ѐ���$[�ǎ��s���
��ob���3K��&}l�Ӥ5�U�9@���0@�z��ɪy��T 87���?{����ῼ���G���~�IG�_��W�>��˅�y|~����3r�p�4��v�*��!�5'a���Ćh?��+ais�T�-�9����
^�q�hD��O����nZ��Gt�p'Ș$�FMS����P�ȩ�;w��ϑ��Y�˫����`�fO�Ϙ9'0:<���05>n\�@�IM��Y�Jak��̿s�*��4��ܧ�#�ƥ�wrT����E1N���4`ҝQ�O�I:�����Aqo���2zhi=�NbtxLPha����5l�n�Afd4��7�3IF�
	��$I8�nFЊ�������k5�o�T:����olf�?y���d�#y��k�Hs8��Yl��hJ_Z�8�}�8�!�}���О�J��[2ٌ�=�4_/ah^C�s�j�ޒA ,N,���&Y��R$a����c��������A~dG�a���5��0	5���������&�p�!K��J,Y%�ƽ�P
�Qt�^dj�d��e���h��- �*:�����gqpQ:�l�Y��K�#��nC42���X�,�����bhp/���萚�g�������&N�L!EW�dL�t�&�ޔ��ag�n����6��8�]�5e�����y���pC_q�C_��7:��_:g�o�`~c�fe��n�N�jU�o�>�lN���GH�������$��0z?�7.մ�6p��v�u���.��IƢ���-y��L~vW�N�hǉp��ao��Ca� 1������x�Q�N.�I~o�T,&1�f�"~�I�j3HY��V;`�M��E��g[��w�3'��(���3�|T�٨Z������ه��-W7���պ >$n�Ax<7��>��ܻ-�n"Ud���aW�aaf������/⅛ωiMb�tY�y�y�m�s�\5pt��F��!�b�3�1�#�|��\�n�
m�f2�4��4$658z�mݗ���c�����F�/���G&�͆�:f�O�'rF�Ro�����5<�la���hCr98	�(m%k�:��w;��U��0�_�t��U��ht�w��W~��/����̣�������A7�<��/>������Χ�u�IL?F|!�N�"K�V(ckyE���&?°�p�Z��X�ޕ�o%�_x�h��A�K�̗�v\���ݒ������v-�*���m�mm`goO�?�0� �j4�F�&胃HD�J%1<��~�v��C���N%��F	K�]l׋�t�8�f�Gf�ݬGN*~x��PׁAo �Ǳ�1L��h��3	giiE{�p,��`Nw�jw�Qvy���<"�s��E�P��C���g����%S	�9s
��&N�4�32�F�F���<V\���3���8q�����X-��x�	��x�W�Ūi*�!i��d����[>�^�-J&�&V���2��-`S�{b��_![������)��iR���+E ��(� ��F��RI~��ϞW��?/�|A{�j�����#;~Tf�,�DH8��--acuM�����2�:�p1�+w�l<(O��#:�F�V�n!��BVp�n[�
:�2��"��:� �X�(�zC6�L�!�CxR>Җ>�]��� "
�zѴ!���1s�w�6�ٝ��uL��qlrc�	L	�⾙�����P,�tNOO!����Da#�X�%ܺ�����:Dc�TE�u��p��f����d��0f��F��Y'�ͦ���A;�J�H	Rd8�h:	G((�������)��b��Ă���N��ݢ��ՔL�S���-(�qqo	��J�����+��x�l����g���S�+\�ɻ�9Ò#�����	f�3o�˚0�+�����H�&���a!���ɜ���~�w��BAEV�'�&V��y�/�d뀠oz�����Ϫ�!�������~�[��H�T�T�W:Y�$UI��҉���щxL��*2�I�T`�t�E���N$��"*le7��C�Yύ��W2���7f5\':�K�"������Rn���b�8�J1nlN�$ ڃY�"��v�T�������lK�,�u�ib�u�I�#YT��j�SQ��|QEX)p>?<L�r a�g~2>����7���_z��;�~�����;7{n\���.\G<����y�9>����"�]��tj����~sac}US��'�'�K�e��܅��\����<%6۫/��P����EM���g�U��v1:/x���S�nnJ?\�4=v)�i�-r P�a�S1o	Ocɤ
!o�a�xL�/�>q�B�k�SG�[��Z�`�^�~���˃�q��,����gv!�q`���#�pjlG�#p�;�9�"]�U��Ѱ<���z����=���8�]م5K�]D�a�o��6%��z}D{�h4(x3��3�ޔn��Z-R�i9%� ��� �!6�lF��� ��Ϟ�ѓ9�{ʰ�I��Uo��c+�g��n�r:�*�b�q��fO	|չ[p���n4d�]I��%���o<4)�i��i�V�3nRMD�Q�;wF�H�`+�f��z1;}TL<���!>��ށ���CI=z'�ϊ)�B��,���ťÜf�H�·�$I�-��t�q�G��o�㰏��-�Ū��Q?(�����}%-3�ͮA:hɬC�-�T'ܑD�\xMN�]�i����q���C�9����L�����q8�����:v��1X�e<��;��`N�u�}ŘL$�_�����F�(h���krV��υJ؍�Ӂ|���Z�P!'D5�G��F��B��F�}�>è�<o�XX!!���z�>�ܱ��0�-d;��f�!*��e�^1�0��>��{����vZ�R����8�r��;qjt#q�29=+�vhK�c6O;{�Rn�p2��j��b��ň�;���`a���ܠLa��]�Q˱�P��p���/[н�bR*5-r*eAa�A)>(1��O��N��!_�Ŏ߃E��Q4*=���>�P�R�,�z3��~�+
Ԩ
�&�������B"���/�j,�6�Ja=J.;�&W�E��$1�)�����X�I�j� ��b5lp���
A�g"f�Z
�9���M92e�쵮�L��_W!fs�{��lp��:�70����JN.��u�1�E��涅o�����J9�Ea�Leh�p��]<���?z�o�����u���V_:E�e���x8w�~�	*�\=�qdd
��38�����9y���89{��#�R����/��r*���l���x��o���o"��`����Dr`>rd�k ��}d�������{��OLY������d^`�(^'��:��D��%D�Mq��qAx�D\>�$,[k�������-�j�9z���0N���IJ�u"�"����83y���8}���=~�ph �#i��S��������G���P�H�V1[B5[��E��i$cq�2��F��C"��'�� �9@�@��/����-�L,�FN�}N�Y�E�A3�3$�+/.����eɀ���ܠF&���,-�bnq^��'���%ԁ���$?Xkj��z`�S�&aY�Y��6Tg��r���t��[=ԫu�K5_63|������o���WW��{���`���!x�N���+����m�aae�hH�����Wp�'W���e�qtdS��$�Ɉ4Äϝ]��� 'ǐVG��������}:�Ѫ���A���J%4�A�FWa}��P꡸Jc��fQph�dҴ�+u��hA���d!�Щ�Q�gQ�g0>����(���cbd�HHicd���/�=��rdDV~�TNm![hw�Ћ��Bm/������|>�O�(�څn��6�-T�����I��������.��m&�ћ�#���8�o�^�:B&���k军�I�4QP�C��F�{W�ψ�����6�m6	2a��NѮqx0������&����"��s��)�,���'Y��bQ�Mڒ�Y^��t;Q�V�y���%��C���    IDAT8B���A���w��=0�|&hrA#"Y�����U���i8"�,΋���3Cs^�n�p��Bx��^O�c�T�/\�3���0�n�޳'p�E{t�dA��a�ّ H�Ib_��rC$2Ò(~N�v
�=���4�ύ��!
��7�˲õl{�$�%3 /@п>R�g�LY,"ۡ���/�U+	9"�Kr���ך�%"	��PZR�Z���&����nVe��p�P�Ѥ"�k�>�,�����V�Rf>�O`y*���?��o�K/�߽��S����������_�v�r�E�N,�-�������]��+�/b0�ă������R>���q�a�e
�<V.�[
�n2���ť�����/KC��a�OW��U��=z^M���sx�ͷp��Cao0���pt�M}Lmi�����ź˧"�.���>d��K/��^����ˉ�O?�A�*&�1�J'v	�I�jM�L	����;w�qqfg�u��_-���R	O>B0��kzt�f[�����\��wC1_D�PE�ƥ�1{�������瑩	��������DM��������m�Z(�xpy5#�&�ǁ������,�$�x]H�G�ռCޝ-Y���H��
�H�����JM?W�P�͇�?�:Av�F�k�eLRYQ�˽,a{³�bM� j`I�1L*��ٳ����jnܿ���9^�k$9�4J�Ν:+xm7���=�����������2Z�+����U��H[zdIf�6;[VD��`��Q$Ɔ��Pj5������M�5��	g�)͐��-1�ea��M8H&��g���M�4��l��e�-<l��8ba�E�F�\�+���D É�)̌�K^D�7�;�r�e����PC��E*b]:3�ZSA�"|���#�0Yh�JYK�R�n���V���L��wt��!�����`��e:ѢTm*62�Ix�5cO�C�Y����R�L���L�r��Ld�R��CE�W>��~US�Zy����<� G�
_��s�GqbzZ+�<pY�I����4��u%d1)I��Z.X|� Ԍ\���A��"����������3,b^����>G�o�}����R���TZ�!P�7�>�B�� 2��BzFI{�t^P1yL�3��ke�azdX��w?�����4=��L��L�|����#Q��t�0����)�*����,~
��a�[��j��]�i���oY|K�1o�Ԁ�ޚ�5��[v�*�4|�$N��IL���{���]�N�h
�*��FU��jE7DȢ�'=h�!�Z����D�z�	�p'\N�f�8�������������/��y��w�=����/��r~��#n�ח1��5J��X|!w �C�cx|������������X���
���k�Wl��|��M���;}!��K�XYZ�A�"<Es&��(���O~�;w`u}[wM�VC~���@�%Fe�t�?�9Ą�9{P��׿&��x,�"L��:���d�%t�������.�]ن<����(A��"��ҧ�fpbbR�Yute�p��=��>��'���sv����GOa}cU�q�P��(׵��$|db
�OnK�^fg�����ZV�R!��ka�ǭ^;�}(8�eHF�|� �'�E�#a����L�o�C��C:����&�s>�S�)�h�v��a�M�A��-��D��gXo4dr��8e*����DkL6$�.�he��tP��Uũ���Y��N��~y��
������O,��,����D�'�V�3���'gp��1\8uI!x|�|V�t��7�0'��HzV[p�$3��&���QO�#������a��p�) �1��J��dq��Ut�7l*��MF;�AYa�d�i�W��q�L��5j�	#��e�//�E�y���x'�M��Ԕ�XY��@(2�H >=���(^��p����E�{pz�3�nk���C�"����`=[�J��n~�#CLN�56�n<�.IN>�~N��QB����t�38�rb�AJ���h�(�r]�R�wʭr�r墊���t�4�s���q9�7�ˏ�Ӈt0
���~��$�x���;/�,�F<�O�>-2&�-~��;���^����o���؉��L&vǸ�qW�&���sx套��9��*WK
��C"� c�q��~���j�Nv���������L(���D��C�P���Rؘ)T��Ej(m�\:�5��9�`���m<�����a�rs��F�e�clM�&^+oyz|G��%W�~�	_,�"Y~ɏ^ς�vb!�u���lX�-�z6f�:\M)R�rϳ����V�K�4�K�F�4��CS2'pL�ynb���c������,���Wzm��n��4>"�Z��E�v�<�h�S�K�F�����nO��1�m4���������/�?�}���'�lm�f��"�����<��ZÓ�����wQ,�{$���vx�8��}	;�7�#{��Ns}uK%�����_j0�n>�kW���񻱼����y��c�*�nO�j�k�{�!��ck� NJX����3�t�Fc��E;I~�Q���aM�)��u��%��H�L�B�X������m�pY'@�-/��}��Ȧ��r۰���&�C��h<���}�ի�}��]��ff���wc7���8��AU<�:hT�9'��G$�C�]�ѣ�1�!�K6&�����c�,m�!Y�6��IÈnGהM�UN��g�+�WJ�R��g�ݐ�#.��Y�F�Ā�`x�W*r�bP8�Z,6��^�X	]�Q�MR�a|��Qɓ����I��n�`Bxh֚�+*:�CCx���x饗0}dϞ�?�)>��M�)�Q���ݰ_��$6N����S�C�c�;�51l���tE��i�3SQ�X$�H�O&Pj�5}�{�D7������TX�����wР޻XG�\E��z�6�,�l��h%&�sb��&0Js(�`R�c�aa�oM��.v����U�^�����0�L�a|tJ&X>16�$=���Gt����{_a$�QZ�H�j�~�n�d�E�nlby� �=�HX݁(|c��MO�5�B?U6p�,k_����|����#ᎇ:Q	2n�T�T�hMf�R�L��Ԍ9d&q�n�<���e'K�sJIb2�@6/�j���zC�9����Y\C~y]ֲ����x幛2S��̝''�@Ї��]������s�rz-�##z>ⱄ�ٚVJ���2�l�0=6�+.��}]�,��=z D���U����ڗr@`AeA���/M|F��5a�g2������2���ǥ�`��@Bzٽ�
��&�ѱ1�GF��?���U��6}N�q8H��U+�5�x�OJ�Xh�MDKPi�,ؗ�+�[�ėwX�/�6�砷��	����bO����&��ޞn�^�|�/�|]}s�Hma��$�������5�P�=�|n��xJkm��\��y��[ɕ$y$)�ׅ袲ȼv��Ǣ�����"����G�=����կ����ի��K/+�wso��ǻ��X��$��*�DN���m$��H�"<��)J���GjZ��N?�T���k�T�B>�-�����r&&'��r�1��6�߾�M�^RnP�nL�	k"q�l밤�
=L	��K"EȔ����rWC��iGf`�(�����c$u>����]3M��2�;}!w��B�%�jEjN����?@��!�=�׉��u<xp�KKJsi֛�a��(�J�6i����Ј��Jp��%�:u�C�ڟҬ#C��2s?�l(����DNTM��-9PjhP� bB�EvU�jU4Y�^l������)5s��
,N�wj�)Éx��&=nFF����wP�5e��?S!q��m�Re,}.E���պlk�~�up��,���Kbsr*|��>�{�=���4Ý�5��ȩ�zaI��A8��X*��㓈x|�ӊ�RQ-'y�K[H?_l"����W�*h4���)��ly��6��u�X4y NMO ���ˡƄ�|M�rNz�������6�|n�q+��F�b�r��i~�^?ߛ[.a,,��>ʅ'��F���022��x��3�9wѡ��x-a�|���%t�����M���h֙��~���LN��U�P�dޱ!��F�N�H2�ܣG���b��*�1��!��i)�t�FYL�e(Fk�HM��;uF�g���c�WM<�95���率'�0'�~���ȭn�wP¥�'��/^��-]+~�4� R�w��w��.���c?�����K������ur��p���e����<r�Ͼ���%9Z]^���b�i��-ޚ̬�_?�V6�,�������k/���'Oʰ���>��<F�Nn�R�#�%S�"=:&̃��X^_�>��5	�y� ��%T]=4<�"A��>�鍃�i`�Ŧ)��6�MV��SDd����灍��^eO��Y��u��l;䩘jl��Z����F��ߒ�h��Y`5H�{�������{>��m3r�`XD-}呓cdIU�Cȕ�7��Vn1�Y������+	�ٓ0�5k��$���"�����[O�������%hv��k�������G�k?�Á�#��i�8�6&%@��yc5mA�,����ev������;;s�hH��ӧs��SG�jq9;����g?���*e�ռhY^��P�bN6e��i����'3=^y����s��磏��񅂲{k����D�GQl��uPp�iy	K��ۃ�z2��B�/_���;	����pz*�G�O�K{�Y�O�bsc}�LV�4]�z�.�8ҩA�b	dPmV���� O(�Z*�Q�	F��6ִ/��$%������k�j���6x����,�^�>�"X\Y��DŢvx|"��U�"!u�$51=��/K��i��nZ�1CDPk��$�PJ�ǩ���iT�oK��!��w��#�I����񵗟W,e����'�}�[woI>DL��e�_�3��Cf)�ZE��BH��j㞶f�����H�!��fKR��nN���P��EX���{E��D\S�Z?�ޣ�n�B�R	B����\�6<b�tW$]ᤧ�	*nD$x s���+�|>�r�(ׯN�&�Db���G�G���K�p��)D�>d2�1��U�;=l/.���"�� �/�Z�䆦@�P�@�h�d��aG��K'�f���X�I����u�@���)h�Ag.�)6z��2�D��ڎ����\F0?O�:'f�98�y��&)҄��u�.�P��a��S��D�n<�
��꫸v�&���� q��^�ȅ�ݿV���ގ��3���ƍ�����'��k�j���^FE��j�B�������?���f��G�G���͎��2�,=}S���*���<��'ψ�E���d�(�9��9�%�%> �u|^����sR�Mv���2>'�cs�xݰO�At��_��AR$U2�Z_�;L�b̪�<��������Փ�َY�c�0�SQ�WV���>��w�L{4�pld��-8Z�zR���j��v��n���6�P�f_����6����$c�A�<5r|]]��(�ѦG�����B"$�z��#�����Oz�A|��|��=�����;��ɓ?�[Y��0�^�"bV"�>�������T�z�`��MR�K�� o�h�	�+����+S�ݭ�����
n\��ӌ�󸱱���%�E�85+	S�[�߽�x�{o�Rnʋ���6٣:S�B왽��vs�o��槉�`˄�K�)X�-�D��Ut�A�{���枆)!�9��X�EGk:��ɤH,��!ܾwc���E���~f~�s���(�$K�%��j-������Νq.w�d*.6&a��*���P�K=��m��n2|���h!gNd�W������H�����tP"��5��c`�����#'c^�s�[�o�"�����Qoij��A�'[�+(QQ�dPҨ>L� ڽ��N�bt+�����5�_�%ٛ��s�nݹ�[�o����:68(~ 'p��#k��~t�B�7��Vn���'�ImK�Lړ�7�!7Z<�/���m�Y��9�����!�~�G�k��D�kf��n�r�bܡ�ӕ���1Í�2N�#�ϖ�%	[�eb(���Q9����H9@�k�ׄ���Ňd:��N���s�=w
�XP�?�"��=��e��d�o���{O��ɣ����K��8�	�Cx�1��i��FR�f;١��r����k��[F"תյ/�N���-�ڨ�ܐF0{�+.��k��9�)�"LBV�֋^5U�0
�9�>^���&���bF��9�o��\9w^�==���O�8�@8 /����mq"�;�)�E�¥KJ�Qa�sM�X��ÙA$0��r�<��=��w�*��;~�,��*t[]��糉H��cqI\����Mѭ��ؽ��|P(�JU'2CC4fc|��������g�������Jș�S�4ӴC�N����=�ri�Ć�S;m#��*�e>³�M�U1�Ҧ�LSQ`�y 测���d�[�-[�dK�߹��Z?��2&��d!j�p������C�y�֤k������2��������)I,¹��٢V&2 �ҫdJ'.z�������D��?�����ߣ��G�+��ܹ3�x��=��|�;�kW���#� ��ǳg���PY����� M 1���=�-�'�/��w �+ �w ���7q��q�NL"�b{}]F�bNٰGgO�ۮ�'?z��wP�4�i����M`�u(���U}���k�S]^���I�3#�6a�$�)4Tzc[Q�{=�[e���UM�gǍq���M��k�p��YD�x����(h������ښ��z�o��������Q�ݞ��$Z�ԢLrJ�"[BI=�g�܅���}9�����Gg)���
�V�~�h�vKI���~(!6I�9w����
ʖ^2���4�����AF�U�lж��������Eo�zK^��r��L!Ȫ�u�m�O�����5��ۖ���e�b1L���[���^���c3�.����ǟ�|�&zO4�8mA�L�=����l���+��#rN�PC�^��N���'͵�v�6c� 1�%==���OބJp�B�"�6p���3���"zp�H�iv$Y"Y��ր�0�!h��a�;���o�dj�Ƅ��`@�d���E��p.#'�V��ωH,�T:��Gp��Q�M�*�����ԭ"�g�������]<|��B�z4��T���mӃp� ��L#�J!D�,	nb��2����Nm��|d�`�=�)e���kNt>��Z��&����+ݗ��9a�w�|� e�}r�J�CD���`��
�����c<>(��y��ϟG%���Ύ�3gO�`7�������V������`bjJ�F!��]$C�QڦRGr�r6zo��7�?��"�׃!�z��2>�a��R����=����^x�3�c3��۷���c�}���8���Z�v��#C"h� ��I���kk�v������������&�Y焸|Di
B,���w�-?�!l�PM��%[�e1�����ٿ��mdL�:B��������X��%��,�J��P�+=�����5��e�B��a1��wy/�M�דr�s8��������DN�M��?,钏!0���h$�����y�_��2�����.���j�\�x/����XDE,��ǽ����
�wvTN�Wm�Eng�U����d0���F���i';9<�!܁D�~�ll(Ԁ�N�x��G�]�$���M�-���|��.$9��~^EN"��a�M#�u:��&��Xt�e�T�����O�=M�2�~��F���̿Kj�ӭ)�ߋ�{�߉�.]��3�K���;?�7����sW�����������_��#���:J=�9Ш��nzY(f.^SB
"�R�k:l	�Ue`R��k	lv>o�AC>}&a�E��?L�+&���`@B:|UBٍ:�̎��	�q���8��A��BU&��#Y�-.}/    IDAT����O&�O{[�(zt��ĩ�@LR~F�G��0s����+86sã�ޥ��Ï?���O�C�.�#��F|hP������i����jE4�%8�M%1�(�!��݄G�����NLVy����BM8�� ��
�˹�����0ƇFD���{m�h���W�ڜ��#�.�Dq�W�tl`i�lx!G�V*4��X��P*��Dt��q a 9���a�ah4�x�C~���)��ۃ�O����R�er����4��iv���#�2������'=�t��3C����A��� [�ϼGx�s��Q	��l.''�B��@�F��	����A"<�D�DFY�}���B�P�t�ǽO�I�M�Ջ�𫯿��.���bw{[�Sl��q�x��p��}�2y�'i�K��PH�437�m�L{��`�����	��\�������c�Eoj>�$j��n���'@xS���G0�diui׮]Éc'��������w� D:�|�a䀔J$b?v�c*��P$���{?�YՌ��Љ��M�j�.��P,A��y��(r:s�[nO�:TLٚM��r��=9�8[��-�ѴL�PΟi�e&�@��4�o�y�M�q���/q����[d,����-�gl�����L`��0�v�RE{~������\��F/y�.�����/��������W��j��[#O?��ŝ�ߨ�{�|�"^�|�h}�~5k���@�Q5�F� �f�F-y���L�qH�7��@Ry���N\�.b�?��X_]�N���'f13{�v?���������^�\�	M� �{Ol_����� c,�,��;mOW~В����[>�PX�<�^�ߐ@�Bǝ����Y�-�4ӭ�9~/�W6���gq���������i�7��������%�ʡFQ]���mFm�S[{n�4��NS.��J#'����83���&i�O�'�\ل�����2���P��#�@�h<![��`���v���e��6�&��?~tF�u�^��斑��9�����Jt�^��mM��%����5�Ru�<�h����f���4^~�F�i$�t�
I�{��}|~��3��4J���Ht��
W!��X@�P�+����4Օ!HE$i-f��i�_�>�n-�[����q2��Z�l(s�D��3������9A���TP�9�^��ͫ`�!x�՚r�2D�D�h]H��ͥ��I8D��TR��GN��	��D�
_�}r����MM+�P��J�����W��JkM*��je���7�Df3@�id*L��'��0�dx��MԤׄ��D_�@��S݉�4������<�ˍ�V ���%���=���+L�=�j�7�*z��� &�&e�{�ӻ(�B�	�����W�(ݍ�0�������T���{o����jy����%0W���Icf�=�Aaj��R����_�=�S�"vq������ʺ��	�6��&�?��ikcS;��O�R&�����ÇD�l��?������* ����)���i�Ei����'�~��b�NC9荰�#c�pQ�F��"P�~��<����C�|</�B�I�&3���T)]ł��<�ڨ��lZI��kU�o~	��oň�g��"�����l�5-��>,�<�%���x��9��4#6iK{�>'�
�76ń6�i����lu{5ر��^rw:������{4>�o���WML�W��JE����������o3"����x��M�Hc���IbgE�=7�(�Fe������\ݮ���hOפ㸸�b �����rI�I�R�\���Y=>+x��?~��w�Q:���t���f
	�I&`�Fx�ӷ����p(�����~�,r�����{�u�ϸ�"���#����&�a�&�bOv!���C�҉s�p��%Meo���H�S82=�˗/"��`mc����xt��X���)�1&f"�sII*��йN��XU�������Ć�Ϯ�P(��#M�!1����\lǞ9�-�m:+�PdX]��6�NM<Hx���0�����L�y�$���0�HQ�Ζ��M��|��"�e3��Fk M;�IҐrEwbd�f�XA�9�ч��P�;;ړ�@G
�.xL1��!�u�hY�����ЪԐ�?"b�_ #��`�G'1�&w{O��Z��5!X.e<n�iY���t:e2B_mYR��o��.W�n0|�T�錶�-{��Ŧ�ð���HK`å�GB(�@$"=7�_l��0��>��[�X��fD�!$1��<pS�	�M��VK�ե�50�Q;?��>|b��uߐ�V��Ѭ3�DG�$)�'f��7R�`��\���x����f��6��2�XZ\��ֆ�qrTc���

Ӕ�`C�.u�� �����T��fs�l�|87{S�xr�	��w%��x�"~�[��sW�j��f2���;&�ڃ\o�߻�ŵ%�����l4��.���2M��ԑ�	L�09nG�&E���K��_���pʉ/�&��΁���O~!E�u����'ʦ`zbZ��hz�ӥ���g�� 2�r�

l<.Y���7|d'��b8�������ﭣ"81$�e�E�0��9��ueM�����Ğ&iς͉��_���f�k`���ʳ�.�bKsP����bn���}��gP��v�_&q�Lk��a�f�{����*΂�i>D¥<���զA�H�c�<����6d�kq}�lpz��'{�_�������������^5��_��+��=��z8��<[����N�y��%�v���x��`�<(�E(;��0��h\µL("�	3FX�/��K&(�a�4]X]Y���nN�SGg����g?Qns��"l�o�t�4X>�L��;h�;f/�縉P���n�FN��4+m�� �!�ɾ	�A2E>�V7'		���͟%�����{��5��z	�d���;2�?{��_���@��~��O0?�Tńא7�p�=lG 0�ǅ��&X�Z�h�$������.����x��q�%ذ�+���~�$��,eM�c�s*�p<�	8gSbv0$��u��Qv�NMk�����f$sb�U�G�5�W>�V�U�Y�eʬ�^��Y��'��i��U��iTj�3����p"�3�� ���m>Ԕ��sb-�˽��e\�N}�Z.��ujT�y�;=$#1��A�4m�@~��ϟ5����~��%�j��X�ݎ���#$�"�2��R*��T�]��[�I��p�\B�VL�c�p�-�-R� �0b'N�`i����{�k%�1�N����_N��z�~[Ey` &�V;�"h��=�5)|���4Dy���	�Q����ޛ�[�J���Ҟ��飘��Br|� ���l��\�.srJ����f3��$d��W��ww�4(Z�Kɡi��B�])�aؠ�Z�MLY{vzן8z��SXY�������׮����r����E��0,�\��v�6�->���:'Rj�y�)$;�A5�0FӘő�1�;yZ6���r'��g�����/�[���ӧ:�ǧ&q��M�LY���U�I�b�Y�rY�,��<��ZT���=9:%���(�͞���d�I�l����S�t�(��[ &ș�j��,l<ߘ.�)����~�&Pi%c�H~Q�M����V����0]���_�W�\HS�e�dG"��.���`+�\���ۺeZ�YgΗ_�a�������5�J�|1ڔ�6~�NZ�t3<���m�p�<���WO���?8~�dX~���T��^{�p�}���{�f�s��e|��s�ѕ��Ȗ��I2�?���v�E�J�N3�V[i�ܔͪ�N�
&��L1��<�6�WE��Eۑc3��9�=�{?����Ot ��E���,fv�����V��SJ���Ֆh��-S�j >���i�ϧ�$��;����K�|�h�da��eE���5q���E|x�n\���Sp}x��wv�q��5\8�X�>���R���؁��M��.5�A�<�F��su�KU�N��/�t�ѝ��'-����im_+�-"��LD��#!ԑd�dBM�7�An��h���,e
*_��<kdv�^�hb�v�KY��0eF2?/��M�-5�2��D=pO+uĭ�aDc"Ɖ�L.����ǀ7,N�!��;���a�M�� "�ZU��r6'�*�>ݧ�C�mٶ�hAd���Vޭ�Ma#g���0�Χ��n~�kT�5d��ni�m%�d���%��6�z]�sc������}+�M�OD�_O�Ә�9������؀pGL���Ť��d���Ɇ�׌ņ2�{�M��}��2�|��W*�t�Щsҗ%u��N����۔�dZUd�UTi��s/�a�M{�z����7T��Q6�&
>�
0ߟ�ljJ=��I�qRfW(���� ��)�����ਦ�����G�h׮_�o������﫡'7#2�������M=o6B�g��j�^���F"Q�o���plb�]���Db�g��B�s�V�@�{��<g�Ls���m���8v����D H�;�<�\�|���(�{kgG�8�RYlq~_��<@7���pdfF�p,�3#���d�,�l���^/ ��.�'�etfp��^�I��L�l8�]����BkPS�M�=,v$�ZE�.���ɢbg٩G�Hɛ�46Q�RkW���g��e�i��v��r�-ח׏�����ށ��H!U��r�������>f����p��Ɛ�S
G�������^�j������W*,,D?Y�����?��l��|�"^�v��U�hV�:0�'l0z���V4;H�exSБ���3RI@�>(�����	�� �҇` [k�_�G&�ő��8r|V���>��{���a�T��f����bTN�tx>��ԉ�%M��s�{�����!w�<h������jGI(�`n6,�2���VQ�7���@*�S�/��ː�~���ǫ/���gNj'�m7d0�/v�ܭkgm1�E��$���jE���Y���8S����o�~٤�&�#0M�d*�gvL�0p8���~��Șe�Mh��w;"�$<a������J����&�n�iŔ�~Ћ3b	Y�s
�V�7�8'r�Iʢ���u&�o9��0�h�2�����L%���e�IiJ"S!��C���|�	`1��)��Z�0�k���n82`)"�������^�=�,4N'�����s��"L� ~©Q�H��yOɺ�bs� �~�A tU����֨�[k��l�0栌������A�]2��sp��g�i-Of�G�2q5�bB{E,�
�ň�
#�������b��ҥ�	�=�/d��K4��`[�T,)v.�t�
���Yɣ@c!x�:���h�akmK���1`@��4��$L�ӸFԁ�����*"���w�jU8�I�����Q,Sg�G,���+��Ư|ׯ_Gv/+���,�l �����§����BlH�S/��~�&��I1��rd|/>C������{���5:�)������!ѓ1�l�I�"����
���͛*�$���x�tN*3�qP�KNU��������̴�|*2�ӳ'pi���b+���|�6��Z�`�UF������r8������"�q�нne�je�3�;�,H�#6g�Vߴ���H� ,v�ڷ�6�L�ӶI��R8�)[7�g��C�K�H�I�gz��:�t�J�����������π\!��s����!?�����c`���ŦQC���U���]G;����Gf��?�q���/��o~�"�����������³�j�X\8s/_���T
�jID��ՠiW��D�3�e�&A=o��)-��^6iv~��-ێ�O`bl;�ܾ��1{��;�����3|���%�glo ��ү��N!��)Ȧ=��|���W�� bѨ.(g��Vh6/�B���ü\v�hr��5됦�=�Z���~�����<a�);|(6�p��s��7~gf�!p�����P��Yz6��k�L�cb-9	�i��j�P(����,d�i�m�bl��[^�>����Q�N�/���[�����x3��9��=jux����)
ۇZ��l���J�n���九�0u�Y�$e&��$��V�^#��ϱ�".wO!c���<8=6��/��ˋ��m�����L,�~�ǅ�@L�/{ԩ7�8��C�S7p0�c��>N߄�d�iI4T��@42�BE�*T[A���Q������k�P�����r��f���&�Lx64W�u�ū`�=B����=(��l���=6�V*��0KN�;�N!�#�Nj�%���.' � Z����\��q�솇؎��L�twgK�;�k�H���1|Y��	�G�������uv��Li�eЮ7�jvԐ��sme�����$0Y�����~�����Q��!�dK�˨2��P��|�1z3�����eh�Fp��U��S��4���WX���1��W����\аt�V.!iꙩ��f�2��ׇ����c����nll�Ѭ	�'�f�}�̑dF�#>sZ�O�ّ�j<��[`<��~��m���"�W�F�rsh������X$�{��9l��#���3�^��RfO�D�T�]M�,.,�D����B[8԰9���8��xEd҄J��j"5)*�� �|�l�T�9�~�x�I�ڌ�f{�����8�pl��JR�Ό́��E�
��)?u�݋<��[R$�-jӹB��=��c~e���s9q<�a�o�ǜ���߼M�����Ix�tj��?���[۷��s����g�u�X���K�E�?8����>���W����4�cjt�x�5L�����f�k�=0/��I��k,�oa~~����>�d"�Ln��������BKOJ�4��1��=D��<Ŏ��,��s�,;�A���%X�9�<H� ��#�m�)Ά�y�	��c� �a�(��K�4!��l�h+ț�d3Z߱��l�I?�׾�M��~�N��@��g�RV)�]D��ecHhi��YŐR%�cdM�*��y��k�M�K[fKt8��!c�鉅���	�`����A�9��L�F�FG��	apNYސa���Y|6�=A�<L9�r�l��0w��7ޥ�֐(�2s���j����B�^I)�wa:��`p@S������xN��j��1bn ����$">c�μ�z����Ȇ1%�I ����`�N���{�8g�<*���"?��vG�~/�rۘP8:��{�C��>T��E�[��ښv~���
;`3����z���y�Ѹ��B�����zlH�����z�r�� !+��`�{��d1���E8cx0}(�c3$���N��SdT }�K%]WZ�*Ǚ�ݶ
�����D%?6]�N���a/��b㣚�y�6��2�'��p.�Q�m;�A��8Ő�J��f�r���n8�O�JGS�DD%�{;�C��F8�Ĺ+W���^åK���F�u"����_���ĳ�yd2��T8�Ӊ�hT����������b���(p��DK��׌���7��/�<�1��
B�D��N͎�ˇb	��9c�SAy���6�w�	�r�Q�A�@4�dl���� ��s�=��W�Hc�������m��n��m���(��)�	ߍ�6�ÖE%�+�	S#c8w�N=n�׽~i׉H��5�fiv�6"i�p9�	��*�.�m޷,�nQ�[k:$�����{{bd	��%)L��3���M�m����ʌߗN?�&�֢��b����]|�'?�����#|�H�{!b�v�&�(����m.4�tw������*�w����åg�M�P�;}�_��0���]�V������%9ɉ�4N�������4�n6�B�NSv�����g������=Y��=v~�{[x8��}�-l��"�#	6aY�TI�v��PY�����-�)y������u|�D�q"C��X]�����"�0�H:��Ԣ������w�q�g�]*�)�|D�Z    IDAT�����"�� ���*��ΝC<�C�R���<v2�����q�ZN U�[��	�RZ�GH�R-�˥�"��Q��)4,z��)A�S="�.0��F��+���$y͘�J#��W.�����\G�^��ؐ���G����3r]�0Y�4D��bf����A0�[[�(d��/@;�V $@ۿ�.��1@���'�}�ۿ���}AW"݅�H���r*c���VGS�������� )B�l���bKS��KWq��U$�)4�uxh�I�$���)e�?#&��'���!Vs�}h��Xg�ʒ�-��`aa+K�;��` f$"�DB1���k��=P��Y��Z���s���톟�����"g	��kS�8�
~��;2�V��C����	��9�#{��@#�?�sl����9�訊��ilHz� ��#G�T��$�Fu����7�����.�7�����}�=6'�ۂ%�q
�g��N&y;_��+6�^?Rl:�A9 I~�d^5S�rhQ����Kx��W��/��1�qbl��t�������`�'O�I���`����I��D>?�bA<e����iN�H��Zar��ȕY0(H����2�m�������P�Pc&��'+��!z�'��1:9s�������ԙ�O~�~��6�Pqt���a �C�1�E~�<?�`q"����k�0���|h���&1���I{���U4y�7o�}�##�3�Z��e�����X �XDB��Z�r��z��h��Ej�q�����ޖ߯�,p�K��n�Ír����-��;ocqk]*
N���?��Eפzy�j��<�Q���*�N�d�n��g'�O���I����ra���j���sx��ue�����G�������L(-����^���4���K��c�S`�i��2͘X�����Ul�HZp��e���t�)��w���k9u��@eWv���R��0�R��&>vXL��H�`'�cvj�jU�x�b�&�+;5veLᇢlW0)S<�i[:�h��!��8v��7'�@,"6��ֆ&an[n�x��+��y{���,;�����{S�uuWW�j7fgG�\��H?�E�W���%)	ZIDP i)��j֌�q�)����{���;��E�P�{(Twuefċ��{����k�	xqzr�O>���"�eu0����������7;W>�
v�մO{��>�ܮ�EB���-G*��$,�{1�Pk�=�b|tr$��lX�tw��}�v>���$��ch�������Ջ��.4\&	�S'W�q��e���z�!Y�D�r#�ZUH�-�lM&�K���p7���Q/V���C<���q5h4")��l���K�}�y݃
��z�ĠWzM0�"�B���&r��$�y��m��J�cYl��'c�җ�ń�
����t�=��i_L�S�h�3ٔ ���u���^�D��g�$!���v8�Z�Y}Vl^���y�b�?��<�;�:�70���lߧ���]�E���_�CNqbEӈ�bLa$��!M�eS���"%���E91�/S"�s��߅��A�z:��&I��pkGNj�vyO2J����O`��D����B*�J&g��LW��	CG�~�|�P#�&�fs��,�<ɛN&.\��o|��^���l&�]*u�L�����<�������#e�WVl�y�0.T�|��R!/��ӒA��]-a�PUs�r_���ѳ��t�g�yƝr�C��N��ռ,,�tub��f�,��m�Պ����^�u\�r�����O?|ۛ(:���hJJ��,])�9Y��܄�/*a������t�Db��}��.�
K+odJf�D��C�����"[�����"�Z\�(��L:�D�Wv����d��9�Z:�\ܲ�%�"(����&9�ю��A���1~��/�q��l��n�n��C�e�iC�iq�<#��Vq��F����&�華�I}�;��������V���d�����g��U���	���?T!��ux���!8��ˢ��"mp���bEW-�E�V�Y����XZ���i��c�:s�6?2�S�l��/~�c��o����&����\�a���@��aG�N����tx�x�ӕ�uS@l�*�4C�R�t��ִ�U�("4��en݀V��e��[�?�C��pif�{t��~�H)?�n�����w�곷�p�������Ճ�Ū�M��RU7;:c�	���pZJ��i7
o�{�sOD��x���-0�2��!� 9�p�(Ӡ�-�~uuY�?4�X���]6'd�f�y��/����������~�N��o�n�[�I��*�Q��w5������#�J�҂rK���W�\���)bEH+�t(�d����&�>���1��9P�T�?0�"|��5�
��<��W�b�l*:�����K��b�+X��u1�a�N��5A@V����Õ~���&`bf��I��]{���f���\!+��,�j��y�����:�eP¦�
b��L�P���C��	R�ԭV����T����a�=�G��j��KgT���x/�Y����3���Y50=5���HK7YSy�E�#6�G�+o򣃸���w��Ogdl�z�dJ���*�5�P/��������<nI�B��y���!��9��t�s��.L���7�����+z�D<��3�ךP����\�޼/��xس �Y����C�� �!Z6k��C��s�!�q�� ��zMӺ䃕�&7�L�Я��J���I�� "�v5�>؜-Q��)����>{���20�L1�O��o�.�wֵ"�3��E��M�����B�U�$�H���k�<}S���ǝ"q�J���f�҂i[nT�r��VmqAZ|�$!/I������NB�U�
���:�t�$8z�!���*�!�5 UJ%���w`��C#�x��[���X>�ŏ��{ۊ�%'�͔�<c�=.T9	�2���ӐS��v6:��q~l���嗒�x^a^ZP�q��:�"8:�c~�>��=�l�>��^��b
��DW�]��>�Si?#���UQ��p�H`��;G	���Mc���]Q�s	�~�.�wv�M�L�?�J>��nȶc'j%w��Vs�ɔC�Ƥqꪪ�(F�&ښѱ��=^��$@���	nuf&��J(�\�Ġ��B��r�b����~+�ϊ�E��3�K��&^�t�8��?�s�{pWō�51k4���0�[iT���|Aw"���@����i�e�RfJ�u���Ŏ�p�]����|�u���giZY]��ܜ)mmO]�<΢y|v�_,$���r�J�&�m����
x�_�5c����Ƈ��A�a���"4���A,��փY1EX�d��P��T��]c�]��~OW�����yQ�%�&g|���z��C�����ʹQ�h�8�����_Y�����xXj�.{P�L�E��h�GBٜ:�,L����Ԅ�`x�p����=+�}� �Y��m(�N&Ҵ=�
�pP�M$��c�ȃ�;�|:%])Mm!���>�P���T*�Y9�	�P#�T��*�&N�t`c澚��%�*@-~7�y�kl
t�*��`������ц�@/½�(ԫH�2��OO�H������UpX�����%ꃺ9Xy�Ke���Hʫ&I���ϭ=05�!�W��{{L�`�?6�������q��e�y�-<w�6���>��h2�ω����c��P�fDh�`�c�}xը
�.Ʀ���C�D�I�Ϝ����؂J*cM�f�#�ԨBZ֧j���s�fD�>ԝ5uDbx�=>�Ѩ�h�;���1B<��r����{����c~cU9��@@�,¼�[�M�br&�q{094�W���gdf���=�ݿ�)~iZ�� �1�yk��߱ȑ�7ꑰ/�{�(�7V�y��I�N���\��l�Vރ�Љk��C��?�+!���������&'���#��;?����Ւ,zyͨ aq'�� ��J�s�f�e B3��ь8=v�s�?��/}�E���M����������=��7�^��7�C7���c,,Ω3��e7��P� F��1�ݯ�7���H4�@�W�ff߹�����c%����p�����v��ţ�8:��Zh�<�ܔ?1s{Ɍ�B�fC'!����
�S��+[Mpb�Cl�Z�' �K50�7����"�Z��jł���&��o���m"�;d'	g����p/��"^�q� rg��ɏ�k�:�]�,+�]��y��O�qtr,� _��/��@{^_N�k+K�k�u�|��%ÊDP.s;F6���O;ѡ!��DºY9��on�@�����A�0��D"����nm�`��)��&���!V:��7�[3�]�������(#����c�#?�F]�eJ�(����ùZA�f�x[�E�R��T��ݽC$N���@�fG:[�g
���hu��IG9>6�3�|��	&��y���4]�)�ד-���m���d����I��'N����65�3���jt�^��q2%)kyiU��<\���3�Ta$Ȯ�nt186�+���M�-�<�RrWK�&#%��g7���aV��h��q��x�1ΰ�|Ap3�	���CMR����3!���&"��a��U�4��	��(��4�F*��@6?-�R��V6�8��!b�bYy�!NA���@���Ϗ�߇�ϧϗ��B���t��[��A(ځK�n��W����gdC�{�ި!�"����f3y?R
��Vj�>��L �>ֲ@lY��:���n96�\���)�$?�
�X�e�jɁS�t辒_qЯ�:�T��q��hgLI�
x(3$T�F�P4�]�GE����?���
����LƱ��~�f}E���?D.Ϝ��k�1=2�Z����M,>������0����Y�y���$o~�˨O�&���y��eoW��-�%��H^i�Ms`Ag������f?���*ZP���1B+-�d�T׭-Vn�)�C���s��ڰ�J��x+;��V�p����i��5�k���׭u���W�lښ!��Ϧ��������7:	/,,�?<���{O����t.|�������E�H&��d^E8�:����/փ��L�*^�]��;���1�WLߓ�8f�<��i����1::���S��q���0y���'89M0aC=�YZ���<���v)���p��\�r�j`k~��s0M�v���ֳ%�j�*�DAdI��"��v�MsS� ��$�LԄ��ݲ:�Gx��@Z�M�;�g�����zP�f���"~r�C�����7�.w���)��v�����%Ν7�`|dT,�{��ƃ{�4]�0s�u;첫䮜P�29	a��Bx8�H�@����+���K+kJt�u�<�;/9I6e~@����I����/��|�]<��!\ȗ����.��ٖjdB7���Aɯ�Ý}�X���y=|�!��Q�fP���7D�L>�|��@ ��W��C:_�I2�i��>�3�� ?��}���f��DZ,oN(DE舦ϝ��jKR�}v]��Z��RSדMR��'���i��)�U���K�����6�,.ca~^�H��&��ʲ`�}̩�	V�E�:����q?���0��z��?��ɩ��yB�D���n�}N
�<F�$�R+��Y�	R�n�ӂ���u�7�(,�z�%̆�ls���_�3\6��dy�I̟cw���*�,���$�%����i1��>����Y��:Y������d0A�TF"���֎v��X'.]���/��+׮�J?�2����ʎ����j��ҷv��$ʨ����ʮ%Q2��iݢhV�SX����*�o^;�S<E����h	3�U�e!K"iY�A_H;/_b~-��\"M�j�����Z���Y���Gx���t����c��V�JY� r�������iܸt	��hr��L�B�у{"c�%+߃&�f�X�6�y��[�;-�)��Vb��t�i���}֟�ĴB.x�����o�,?��݂�u?�lm�K���gA<5����R��{���I%ꥩ"�ˠ�X���̦e��W�ot4����7����)�4?p>���_ή/�W'�\�k�q��M�!R�4Vמ��?@��������^���b|x�<D�x}�rv��w"U�"�:�4�pq'T��Dq��%\�D$�"|������*]%����k�^\��/�|��������,�(ʠꕲ��i�L-���p�R#�X�!�������[q\b{� 0d��F�a!o2}k& �>�-%�>�A�D�j����� �فT��R�!W�ɩi���¥�ID�^�Sgx<��tR���$zb1�������VV�Tܹ{�M��K���B�����_���7q��+�t�b�6��-�s������[���cnvR8������GZ녥e��g?����Q��7���-o��)����ʘ�C4B[0�����熑���v���G��Q��^�+�e^E��yԭ���!�4�" 1��F�'�l�\�T%�^��w�l�I:���u�ʄXi`�)�.cA�l\�M�?l
Xp8	�,�PЁ�)E�V�`C�cRW�� r�j����`�	��'��סK%��x��A��K/alr1�^I������SF>�)�)X<�"��������مh[�D�Y.N,��JIbk�*P�$w:�[Zy��ץ���酻��)�b����YX�������	�uxt�
��7��	��G���ˆ|���L
gɴ&3}=�v�Zm�'l&`������X%�ׁ��k���,�^�0e��߸����ϔ�X��Q�G���k����ŗ_��J�>�J)��#E,�d,n�a�s���)	?O�j�m���_��eC����ҍ�VA�"�BҨ ��UD#��zU��4!V+"sr���-J��5�p�������ߍ6�4	b��*�?7������kH7*��,�Ӥ���W�͟G��t��Q<s��;0��)� 6<��g�׉��;�E�K����Z�g ��^|Q�X�B�������s���3@�|���'[S0է�+kuEf?af�ö�v�C��g �6��Fj�@�,�d*-S�#Z�d�4./j"N����p���� �8�N��H2W�^��m��,�D�(yl�{����������8�F'�?o6�~��/l���I:�y�^{�Y�'X������g��=����p�=Cw/�����=��pqW��\��t>-�탅�2���֎�W�K���B�����:>��Kn~o�=�Hl�r��U$���ؑf�����!!L��<d�6�h�ܹk<ȹ�6���(.+����C�����b���A��`e.���!ˁ*Ҁ���{��E�_`#�"|qfWƧ���O&���]�iڋ����R� �w���U$�LCj*olr�gT87�6D���}���\�|}�"N�Y���F��)���#���F	ހO_�?اf���Y���HS�E��@Hl�<�*u�?捝�礙|D�熇:��h6��t�k�
Q��2�I,�E����D��Wag�PF2�_+��]�8�C"�E��ό���pp�.������pQ�Ţ�f���1�pbldT�5�?��$�&=21����m�iH��V�������	IYgɄ�Ĥ��nW���#����/+��ׁ�.H��<��@P0�_חR�k��8�=�!�`H� �I&���s*̣TT�$��u�������ū(FNw�k��j�c&�i!7E�/�R�0������I�Wn'Jt$��%�8Bye�x##=;������%[�
|���BqK�BY^ D�ZE8�� ah�����A��#BY�&c���-5k.O 7�}w^{7o=�F�����F?m�ؑ�i X`�	`M�ʤ�� ®|ݚ�y_�Z��z")�FA�UD�شe�҆�Ns,�d��i�A��1� �RiАÐ:�^b�2��ȉ�ʮ�Ds��9E�lq\�./��
�V���G�t��d���(K����^b�U�����!ߋ#c�FO$�����_q    IDAT5-l���Ed&2��\˫����˦�$�Eg��s����l�lBY4�&�h12��牓���5"r���133#�!m`7ww���D�!��ޞ~=W,�DC��N�C:����������!V:�X,�G�r���0�3m���R�pm���&/|��|����Y�:�Qo6#N��3��|�N�-�������������8��~��ܸ�h  �!f�~�٧8��E1[Dg8�v�صŔ�JBL[[� �K]p��(5J
�fWtoa{�4�vS��^���.#$� ���5|~�k�Xu���N��54�e؋uT�cJ���������-�!�΍��<����.O܃(��N�EY1\|ht��l�4�R�J���H������0�Ȳ�!@��:w��6x;cp��a�y�6C�{��_�A��G!����{X]]�q|_�T���Ăm8�>��Ҋ�p/�E�"e��;95�T���M��
�`'��	���4�^�G�Ɋ��=YZTG<1=�����=�/.��>G"����e
H�®�2>�Fo_�&<B�
� ��i�6�hR��3�EZ�y�6v�,�������@���H=���:_M�Ţv��t���L
��9��/����
��^�`hj�9i�{��y��x?��Ʀ��<�������9r��j����_�MEX�2�O��D����)ߩ׵�$��ZN��lmnb}eUa�$D�o�x�y>�ڢr��rk�,[��}<p��5P��k�����x�8˦�*X]Ņ�	�7���w������4(�8:���U�Ǔi�gi0�R+}��{u�*%�
9�e���c"N�Dt:Pc
��h��`5����b�Ӝ���d�-�&>�&�h0�(�}�X���6rNBz��6�vp�8�J�ҥ���w~���*�e�QbD���V�A#H�jM�RVJNd&u����|o���n�R�
��R6f��W���iC;HT%a1Y�6e�:�h~�kkӤ�{QS8�Q='6ԩi���r��x���ټ�����el��qZ+�J6��n<�� �ܑ��M;�N�Μ[/czpQ�_���K�X��w��.cX��a�3�4��籷�+H��C�)uz�����iEI�ݻw���� �_l6� ��X�^�"w��5�������iT���5\Z]����ns,�,���]�U�"��,�1��U��=����ӕ<�=A��Q��3���o���~&�wx���=�P��s�g�$��D��?����w����|�E�����o����D�����x��MtG�����\�G}�����痦/�!���W�v.��mJ�*'��q�Lh��`�	���'܁.S$�I;�E������>�+X��c��������4�ӯ�.��������	�Y�l�(������eA7�F>W�������`i��=0���8I�|Y�ExdxP��V���s�d�ܨz\Ƞ�d��2�[2�k.���y�{B��2x��k��.��p�dB!	a�}���hﷇr������n>{.��Q�/~��t�CC�����O?�Cs��E�QeRY�V�/���W�cN�l$f.�`xtH�������2�g������u6s���{����ߍ��a�VIsH��rY$qp���`,u�<̂~��Cv�$9q
-��	��+��9����6�\�"�+����Y���͗��eK899E&���]�x(�!*���s�|���?�?���9P��I�H�J8�+Q���ZR
��v����"�֦����y ���p��L�L�[g����*��/��"�C�rh��r'�ɗA�&L�H$N�}�;;���Ws4�}qKR�&��[+��(~*��z0q�,M�kR4^�$D5��'g��֏��Ȉ��(0��Z��n��F{h4��|�VVf�%땺o"z��zp9�&D�J�j�+Z��H��b����n;�]HFoGlD���4Gh�5e)�\t���\G�(������=|�;ߓ���M���%Y���_�rS�Y�]#WA��6��$g4u)��~~-r�!�U�`-��9��>�����U}��+e3K�;�-$l"��г��U�\R��ۥ"̆�P-��׎���*��70�����	�+y�YfV�&D1�h���Y��D�׏������0:�AȖ�R:����alxD�z6h�bM%�����f��3����1��v�y>-����[ϩ	a�&4�F�����̿;35���5E2%b~��E죦��^sz�!T|X�����I��8��A���t��,�,ดE�V�^�j =.x&Ѳ�t�P�O7��n5-r.}�"N�_���?��F�/����~����?:L��Ь����2�����|��;H�&0�7������C�`�L!��g��p�ER"ugw_�=���ҕ:��(�]�!�xww����"��Ь�0�;���v�W1�ُ�U���ܣ���%����j�I?�����!I`�o�T�)W��y�׊0�bvĜ.Wɷ��;)���aBA?.]<������S�a�|���X��
v�i��(Y6���z�"����No�|
�~��U�}��/�^*c�{ �����d���ҫ���+�|������s|�ŗ8��;�ه�q~�.����g� �G����&��>�^��澁^5;{G��O~���]�h��Å��ۋ`$���
�wp �C������
���� |H73j�`�!���-���e���Y�f�JI;{|e?�D#�f�`�����HT�iJ���ȗ	�Q.U���Oѝ*#8�a�Li��i�֑�\	m�6\�xI��P'a���9���m�L�:&ֲ�3��Ǣ�=��ѐQIk�&Ӕ���ϸ 9��������Oh�X_���:�й�$l�����
 	��8�d��a�����X��]�����wj�y����4�or"W,�ׅ@0�����a��n���%WQ�w�t�V�OgQ�L�,'-=k�D�0(���s�2���Ҥ�.�j٘�	 ���s�uT���?,x���!�V�$��i��ۇ���{{�r����&lD�HB����Cln� ��`ll���o�o}�DR�U��_�2ￇ��x<7���M4�������^��H~���$-5y���B	��y�F�$M4=�yV��ӌ1H!����`o�z��AM�y96�~�'|�	�ͥkC(YNN�����U��1><�"���f�V�rz��Z%w%�/K\��ࢤ�RW���D\�	�ɛ�<c)����ds�s88:�/��BT�#�.�arB�|}������#����"$t�>|���M<��M5�{#o�07�#�I$����Q��z�h�͛75	�a]Y4^<�E�oB&Ldl3z��� ���'�ã#�$��'�y���WKs��
�$Ƕ���yi:�UO��:E�%�uY{Z��ɢN��C����O^���7^����?�����O�{Ȏ~���舴�qf}u	}�.��F�����F�TGaⲘ�GB����G�IF_=z���}�I����3����*��B��?���rv��Fz'�ӭC��`�>�Ņ9�����z18�#'��'Kr��Y}�YG�\C�1h4��䀻�O�����|��$ŰLd(.�}�Iѷ���K��Z_������=�{Qp;��Nb;}�,��/&G'q��%ܘ��NO�b����+�8����@���lAIA�l>o/^�D�Ī�p���;7-rw>����K����<��F�F�������Ç��Ĺi��廙��GGW���iRf�Kk��*����h׀���ޮ���
o:i�c [��w��Ed1k�#�ˋ��b&e+��	u�	֊�M'�L��eB!V�	�Xq�+9a�?�ry�O��f	g�d��`�-w_�"ҧi4�����������M�9a��}%Ř��
��4��%�N�,�ܥ��"I����ӛ�ʝ�JW1�l��%��*�,��e�@�-w�h� ������>/ҙ����.j��2�����������I�l���	��5l�X���Y$��G	�F�)�Y��?7P��`PM�`�����]��E�UF
sX-)�������bK�9:��S-�����niL�����5u+E�2��sI���N��OM���h��S>�,씼l� _,�677���C5�����˯��F�('1���PK|��G���O1��X*��z��A�#�|��\.��9�G��6}�U�iNC�K@c�x��uЏ�j;�@M�X8���.�6i��$�0��É��f^��T@eg$�5�������y=���x�*J����:�o,a1��x5�b��
a�r�h��Xӥ�PA3S �yj6\���T���+��,a{w�Rm�p��:�N���t#�I�p&+C��ǃ��NL�Mh@�B���ه����Ｄ�[�$�a/�m;��2b�ONNbu}MS/Wׯ_�u,���%<Y\Ԟ:�ˡ��:�5н�-?zF�r``;15���1��4�.�S�|��9��K�2��< �S�ߓ,6�;f���ZiN|&(�k�s�~9�3�������x�_�{�?�[[��d��ޛ�^A,F6�Ě&����;���8:�e!Ǯ�LJ���E�7�.(W(�4�ă�E<�9�A2xC��̳�u�:::ې)�`cw�C*�V�[�?�nw��K����1v7ֱ���;��W^R�e+F��S%J�:pt�B�~�N�:������P��]��K�΃��������ը�@��l,��}�;zp<�Q���Ӂ�ӎNv.;\� FFp��e\���Nwj�Qܿ������Z���.��
�

��m8��ӏ[Ͻ�חO'��q��9��>����5tww��g��a��x�l^����.�`y}��v�^*�2�Lp��%�b=����_�%�w���ڦM�CC�� �ݎho|�0|�6%߰VfW��F��X5�����]�Fb <p&`��U䪄���o�8>N�s�zWL���b����M��(��%�H�&QHM( ��!���O��gb��D�!��4��d�U�)�b�:��T���+8��f��'�S&���M�(O��]�Ѹ#�2��*�ZS,�_$ց��.J|ҩ�|�9qЖ�~�4�ozݚܡ������Ȁ'�@����Xm�*�6neu�ZXD)�C4�Gn��1�R�D,{�D5���P��P�=_��T3
&�I҄fW�g#��#B�MF��-�-�#~txc�����0�dkiY$�QO8����ĉ����k��>�F��zem��c��ҫx������;�s����T��P�O>��<@[�*�-�D+ч:\�AJX�{��ŸgC��;�iaLrb��Z�?z�D��N�y�d�i��������������Cp�vvt���4�U�X����Ң�(��t�E���&�m,a�t�F@]	d��Up�Nx�@�4���l�<�M'��ard�X���K��u�w"��4�F�PB�呔�Ŕ3�]=�ǅ�)��w��<�3�V��^�%Bv�٬��jjVB�t���ʲvݷn�¥+���"L����H�/���ɠD���5g����>�wwad|�c��"^O�����g��P���r�Ą�^7�~�U5;\���\����&v����t��?y��;�x���{���,���Y����7o�A{(�|!���E|��;�uFb��uk?L;4�8�	*�y9����K�^�ln
�>�Qw�$%x����B�V���2>��#�1@�Ql"P�!l�"w���aɣ#A|�508؇����m�wggc����n�(�,�<w�yd���Z��^+v���|��b͒yMȉo�v��,rү^����Q��'?�%�Ūχ����ύjȇ�ہb����\�p�&ϡ��5M�s����T"�f�"�/sr���>L����ū"*%�8=9D_O/z���W��\���6j�
&��1�?��'+�|��e����ܡ�d/�e�¹i\�x����i*��>x_y���pM���0�n\C�� �z�>�g�7MX��pI`k�٤�����AʝQ��E�;� ��d}r"�1
	&M�5V��U�	o���ë���qӲ5E�h�:��C"����\���-#w���~\Sg.�E��,f��}�9�k�=���a�YP4w�N�a&sJ��B;S;�ӱӊQE�V��
'Uv����{Mag��A�,�2�g���p��B��Z��B8C'���+��L����]��,|{���U)�Z��}5S���.���:�ى��>[Ѻ����BRLre,�4�������e�����\A�F�%t֘�����V���^PEZ��/�[փ�wN�-˧��\��&^˖������ө�T6L�	jwK)Z�"􀅎���7jM|���U�IEl��u��-O�F����p����ecN����,py]Y���dVz}���>P�I_bB��������\�I:�Y�>��{�`z! ����#��~����ڊX���>���� :zzQw8$�9N��Eb��=��F�D�Z=�Ã�'XI����5W |]���&j�J��p�ʘj�Í��_5~���ʢR�r�2ET�E4j��E���
ʉ��
������8�c2YYZ�Θ�K����6��KZ�M��ˆ���Pז�����kPz��Wp��E����K���c�	\ggjP3��x�J|�&I��C
3�����\�ب$�9|��.vsgH���q��r�v���Jj�tZ++a��'����TW����;��������~wnc����>��M���+��ɎNbok���'�:����kߦ�1�Kփҿ�i���e��y�X���p��!�+!_j��^��clr�j'������|�b���i�l�R���+�,ڣ!�t�?��~��)V�,b{w̚��s��K��x*���e��˚ x����^W1����ɳ3{hI7zڻ%�!!�7���z�q���PH�Ԍ��#[�!^+�YA�=�r�_��\?�g.#Bs�rk��x4��kˈ��|�1����3Wn�/֡��iK�w�b|p�|'�G*�{����T�N%_����I��h:Z7i�M��V�r:�ca��Me�X[_G�IB�C�E�����׃��Wq��-r�85��i�
5��rjp4�n��Y��V�������Q���Z�9�5�X�ym+�\H��^�;L���R��&V*��2Y�9��NS�>;L(��{�b6�)6�	���PF�m:l)�2��eȰ�Ӄ%g#y��? �D�B�D!�ю���ZrG�d'B��&�����*��DgZ+�Qe1���h��ށh{���������(���먖P�̖P���9��;���(�X��p��54���~��m�]�g�p��M"��7�ixS!��PZU�4�l��l�g���+��/��i����d6�{!�H�1V0���w�\k�࿲:4��Ԉu��Z����|@��ͦ�R���zm��;�9،�:;�̕M�{���+�bzzZ�&����n��ҫ�������gɉ�ߛ�AG{���|6+H��r�$Ս�����n�k:�>x������Δ��;�����ۜ�06����!W#��r�*FF���"���g��k��4�9��G�{�0}�d��:�	^/�Ο��W�[��x���'�{8�fQ�9Q ����s��}qmc˕��U�n��R�nL�`��O�����?~���2ur�t�L��	ȗ�����މ��1ܸxYߣ����Ɔ8+$]ݼ�ք�	9s��?8 �Q���w�,��n��)¯��._��旁-�|�
��S�c�X�pP�P�
:z���ۍ��q����w�ۏ�J
_,�a5q�c���\rz#�B��-Y��w�}�;P�L$���|ӎ����H{�������Ƌ�����������wx����[/+�d�����_�˖;���8j9qj`GM�"���`�&�<wt�Z���q2�T���u<�ҫ����>G�Q�$����w?yO��L��C��8M$�ߣA��I�=�0�x�6��vw���G��F�*�qx���Ɲ�    IDAT�qB�TGg'G��!3e�@Ns����oml>�Qa�:�.�`,� ��~���+��9���1ʮ��Ⱌ�f)�Zg�a �h�M_��.��B�Z���*�֖���TK�VL����ǹ�I�lN���!uql��#(��a{Gt~�xd�V/Tt�p2ag��Ր�5�[��yX0�.B��CJ}��v��hd9� 6@ɿq/�ۍK�����k*2�¼N#�b@�˩]�-AC�(���<��#��~�\����b�R�Ȍ�"��,4��And4�([��d�-�Ḋe!�����p~gy'*\�H�)�I�NW�	n�vv��}2<��G�4���HZ�bL���}�ji�	��P |Ń��0^IR�Sg�����5�-X]ߣP2��'�u�*��Qi�T��H	V'��׎];�u�RF�;s�S:]J[��z}�������-�����"��Z+��i���QJE���j�\Y��T���2�Xy�E�
��5kn�óS�J'-��4M��7�\+�$Y$>�>�uS�����&\���~��˥�-KUd@�#�.���RY~���"���gbb
}�ݒWr@"%�o Hƿ�8K�"����nT�c^,i:��&߀��,�,Ĝ��?�쳊�����_|�w~�s�N���yM8�	 l���/�e�o@��'~�8G��z�-�:���I[�����J�\�Bݦ���Y�^E�i������һN��������-a%���JU�h�<���̵�]��Sb6Q<?qF��H?�{���QhVt�R	�,��Hx��{�V���{��y\:w�&�dUk�׵�������sj|�2ط&a��ؠ����P@��%iA��o��n��}8�O?�D�$M�ϊ��dp�)�]E�r%br#��r������,֎qXʢ�u(���g#E�4�v�L's|p�k���S0ymv�磑����o�;k�x����ͭ-���Ó.�9	w2�Ex}o��/Q�f�m��������t!�E���a*�U7*�r��l���,��I��_�w��-LL��f�ci}?��?KȜ�L(����
��R�X��5�w��	ⷿ�-��>�<��G�J�́|����	��
z0B��C�,�1��J�����;ٖş�v)��eG����$�z:p����Ǐ�����_�E���2�Q���Vk�վ>y/^���P�j�+KX�^��;;vx�RAŀwL7a�ɉ��Y*&�˰���D�[���c$ɵT7!�d;�(��(��Iq�MP��b'k����C���*MITę
���Ego.^����u�pw�i��&��J�6��~Y��;�}����&���f��>߄TT�)��)�{>�-#�8�)衩I�]1m3�;��v��
��n,�k]Ab>w����>�BBW�L�h==�����dʩ�̼fʅ�d����D��I����ѼoZE�r	AH*�.���B�,ob�k$�J���$I���;���>��9Lb�6�����Y�rҥ�1#���!���E D���4�w4���92����"a�~�q˞�k�p���
*���駑+��l�bId-����
u�E-S
K��]�1��絑�(w�E��d:��al�Hnb�7�	'ϧP���&���6lTZ���x��� 
P�yS���B!̜?/r�řs�z*�4��s@4���KOp��#W�Osa��3��W�N�O�E*�j����ffp��U���}���"FRfÉ��ż�X8�m��ؐ��<c�Gi�¢x��-�Ǹ*��ޒg~"q&60�2����|6h�cpf
�ӓ��B����v���-�n�`�,.������p�00����&�ph
�Gp�gWF&1�b�x�P�l� �>I�\AÕ��i�[k��p�#Ԇ��nL���ʥ�z��ՠ<ian֤1g=��sA9�r�	�{͞�E��ͽ5	�\��|�U��}4��N=7Y�d��� �ˣbk��rh%��e�sSӘ���8�N/Nk3	�㠘F�mS�+"�<[�\�j���5H(��愻֤��󡎾��_����o������m,�w;��C7n���/�&8:�J`sm���'h��
Og�#\D�V%��Z?�T��d	��,8�88I�4����/��[o���f G	Kk���O�͝m��Ʊ�H�+��	9�lQ�F�nCoG���oct�O�>w�?���~�u������&�HH�D.f�R��J:�d"�wN����C�9���9tD�Tw�"f��,&]�h���	�G�l��wk/=�7�K�Ӹ}�2��b"�̮,`y��`N1o�4(�rU��`��r�|QBs���Nx��Ag�C)!n�8�&��'#�g���ܪZNI���3�HА�Q|�y:�}掄���̤�zN����f�>��O��ǩ��5� �A�7�>��ɒHj��a0J���M�<�rŜ:]�tz"�Xep�ɾeh�Ԭ��wƢ��do_����N��ds��P-�"JS
�t�b�e����r&$Y���<y(�SM�(6� ��YPfA%,�cljR��hg��V�����I?��L�78���ƏeV�i�߇E��B�lA�aʱ~]���M�s���p1M�4���;�pE�h���'b8�Z����'�GW��Uh)��i�'�|�jڿP#�^�ҍ,)�]��S����Ց�"����B��PE�-���*��t�$J����3�!0įFC��#�_NM6��j��"�Ѥ�w�L�7�^G����"��D{D�������a��L�tE+�u�YH�V96ɢ�;M�"���,Y�,������v��\�x�\��9GG�������nrlۛ[�jM����184��.�TԌ�""��ӕ�,���&"ݝ��r	�3S��'~x�#��|X;����*���4�(�k1q��
��&����;O��������+87<
�݅مGx8��rN;\��HRFR�����0D��hLŪ+ڎ�ϫ!&�`��,��H��>��Y�:�������%[�����k�z����[��ءm%]ٲē��=9B��ݶ�P N��T��012���Q̌O���!]+��Y,��T��^;*,�D�,�D�UlV
\����#�/��8�pi�����7���7^�����������ag/>B���[��#�:���2~��O�Q@_g&G&��J�e�R�"W|*�`'��EN2�<���0�����3���Zǋ/������c��$J�46�W��cvq;{�5��ZL����,�t���g��+����n>sM{گ�����u��y�ad�5lƏ��˜[	*,P�&JL0a7Dc�~��4mǵ�Wqvr���M�ڂp{]���B�P?�����������D6O{��n ��=7\�=C8?<��f.	�g�[]���&��g�%�Hr	o(B��y؊e��Uml"�{��iJ�B�yN�*wu�*�N�f"%�Ž�1v�Mr��QNb�@ZlNx� �<g��x������\MML��+��QWJS���[�'_x��CÛ\+>l��%ƀ��5�l)��2oYו��Cs�bQ$f���eu΄�85�x��X$�1:��>�(��(�F�T@�#��"ma��S/J��$C�-�N�S+I��;�S+]��X��xЪ�`���-Å��qt����@HB��!��}'��;�.�������U�{���y�g�ɔ�
<�l$���SM��sE�qjcB��g�H��x࡙�� ��F�
���&1�+��n�N:PJ�9�� �8�%!���Rמ����BANNz��[�x>;DZ(�i84��mK_dI�Z��;����ӠO��	ggBv�
�7�x`��E`�:?#�T\#�d����M�l��K���n|�\�O͆�Y
�|V�H��q8�[x�����|�wq�I�#�1}�i���g,&��ɉ	�~�7��͟�a��8=����J �͉�39>���ɀ��w�>G����Y�ؔ��YN�lθ�~��=���uc`r�Ã�B��PgL�8���-����q�⁊M�T5{ˠ��t��ز%��t��W���g/^�y{��=<~� �B$-ݥ�n��	錚V"[\�q�䢯��!����o��W$��l�����V��")�;D�TZZՠP|x���/>�T#�+ S* �0�8TpC^ =׉ �d;�ы��A�/�T���f�r���Be�I�����'%{i8����<��oBEO0_��,�gc������ML��򋏾������GcW�\��WE=��2X_[�O�CM�Թ��F{0"M/w�,�YU�y�2���T>`����N�&��+��[��f�M������>������������%B��
��+X���n;��z�V�S���*<$\>�e8H��8uf���I�ౠ����9v���rDb{WN�C<���1ɮlo���5F�\%��h�$`)ӎ�p�L�ǋ��(Bm���%<�\�v∫4= ��\~/*��/NA�� �G����S%�p''X�la3��7�=	h����rY��6�Lv�,��� �\S�Kbw&ͰfQ��r�t�{|~M �R~p��Ɵ����)�P�J=!j@�i���#MH2>�W���h���#[ȉt$G*�	�H�)���A�p	N��sZ/򰒑'Z���gy�'3rZ�5�����PnM´�k#

*�tE�0a6��XGZ�?�@���D����Dɑ�ý0{�\��B��Ⱥ��Q���J�r&!�md4>`�>:�N�GX�C�_���i�hs�I��w�$9�e8��.S؝f����or�CCp}ڹsb��)�a�C(��H�c	���IG�4!r�2IY4�!�	�9��M�-�2��Q���C���B����E�B�6�l:ihB?6Xd�Ҫ�f���9*���`��
�s�dFh��M�혮{�T�Ťx�g5	���ё�:T��v�_YYR����
����B�����h�N�X�$�`�xY@6���o�տ�A>55"�'�8�wv�����q�T����!�Ã=M���^{�u�=�wv�������ٛ��T��i'"@�6�rN�
r�Mg���m<XZP����(9(Н��2M>m:qա�o��`Á�h�z�e�r�9�'��>���Kd�C����^7.v��ZҐ�\b�����crNhq,kVr(c�o�C��!D�*勄^����阤?�K���RQ֨�o�P�E���I�i71����v�[/ML+4"]+��'sXN�㰐F��@ى�E�����]�B^�"̐_Ӯ"uz?�����"�����l���;{GcL�>s	�]]�W
�X_�/~��ꆆ�{156��?��%�?m�X��v��f2��}q���ul%?ˀ��Wo}�MLLr/����*~����h~�'�#2z�TBBN����vU��V���	�����M6Wӗ޵���e7��h����!�E�ҋ�7b�R�ѡ��	8�ҁſ˩^׺�ch'J�/�=n��Ş@v~M+� ����9ܚ����v�؈�b/q,h�Dݨt�)���v���I���N����P.@wjyA]�Ĩ�kTjbt�iy��C1{���ͼ�y��k��(T+���!'��/�������/sZ0�cS��a�\��(�����Ø:@Z�yi�����")�)U�-d%+��bϲ 2��]4���3s9�sY}��jn��E�GR�ۭC�v�,����(p�/�$"'���;i&����t��!~���c1�ӗ�:*U万*��F~��C��������>���2v�*�#����H�%C�S�af@=5�ĩ�0''Bvd�sZ׳D�D���6;JyDʷ���j[٬��Xh��ً�����i��1B�8~��`%)e��
S�h�X�c�p:�D5�MV4�j����Ô���ԗ�S�eB�[&"�RQ�*�.l�x=�w�Uh�*�������2��+�N�A�/��X_/�?�l���$�f�泷p��5D\>��o�����K^__�.uk�:I��$,iAr�=���;0�g�W��e���$9���տVc�b�I���@�_G6ql�)ա_2�N������{���W��-qr���y���s9u�D�R���\6N�W�/![N�w��Q���˛k���]��G��I�j�Ip�1ֵ"�j�9}�\��C1|�Λ���o `w����w?x�TB
�Ǆ���X�{�rC�F+c��I�ju�R�	�Ŭ@�8��0��Z��&�4����?7�P7ɠ>��PG��.8C~��h�l7�o~?rc���މ��1�h��2�,�M�R�<%�i��&�n�"x�򬠹I�8!F4�#'������ݿ�������X�����w�'��t���Q��w��1�������#*�8!�k�ȡ�ʎ�N8��$�q��Y�R���������Y��X�x����_bucgI
�=�����N�7w�,N̄�����EL��v�n���"w�ԅ�A����ÜP!�_���JG�����`H��R^��Jp��x;1�Y;}x����p*�(���OE�?szr
�F�e���iC�VA�Y64aZ��GpWG�P7�ݭ@u����M�PLg���	[�k����Q-���RL�!��\/I�K9�ث|�Ƞ��88��)��k��ØA0l>?�Y�H�\2	5�e����=&���Kh0�����N��1�|���(��L��B��B�t�x��͞���a&�*��� ?7_^{��i�Ű�!��$x��mM�,l����L�}�����"LD�60���(�f�M�&~�,J���ǌb6V��.�ptx(���^SRO[G�}��z� ��Ct��k8��W��9�a��ke]�2��/T(_?CM���՛z}<`Zd[��_��ܴ����=v�"���p�xd%��mB��P�ņ�Rd&kY��Dg�Ts9بæ4�E�%�
�U�n��_r4gSf��!�t�ǩ6d�_�|�)��H0ҦF��"�gL����ִ�Øv���ˁT�LɁ�ņ��7���~xۂ8cRR��@[D��[Ͽ�g._��\W��eC��o�W��y~�3��� HЀ�Y,�U�]]�mu�Z�R�W3���؇����y����y��5��V�j���Ѷ�-�N#u�7,=	�$@x���l���^w^F�PB�.��y�9�s3��}���y<�/4���H:�"���V �I	c�����q�؆{��������Y{3O��,����"�*���T�P �ty�/~�Kvj����RE�~��-}Of/��X�*�VB�.�&�!��׾f���%�G���{�΅d`_ /��Z��Ԝ����^9���zے��M���_����b�`���g?���'���f�rQ##�rug�KDw���nb�YW%k$&c���!R�S���:)�I87����;g��߯4j�?>.�> l}C�����������l�@g�̄&�GeD�r������=�l[��f�0�������������@�c��P+W�������o�����]z�������,�M�8q�^y�6�۫ L;��~�e@G�l��qK�ڌ�&`(��\\́�A�pmٮ�߳՝����,Wl�k_��ұ��	7l����������~^6|�;����IB�^��[��d���
���K7��||�,�O��7�xH���D��o�@��BQ�p�Z,Hf�/�j~�E1�E'u�����P��
��X�2��y��ٴ4�	C��ѸE��h-�N�U�?�sI�1Wp���ħ�Q���F1��D!6KAw>+Y��%N%
�A"s,���M�)x�n�������B�$b�/��f�õ�.�f�R1�w���atg�W��i�[&�w�#�Y岲n� 6��5$,[�6I�Pr�J٬�����gN���8:���: �P�� !�i]�)GC����k��YϘ�!yE��8AJ�D-��	�T̃9�_x�E��I���	�@�&]�x�1���S�������4�go�tR��{
����r���gIB PD��&�w	�əˮ�} ��CZ;�cT    IDAT=:iǟ~ʆ�S�=i4��oTX�xf�u���`�`�i��mQ%�VEnb@v��=�03`�DI����	�$x��V-�x��9>-�~�YEp��C%V��yNz�ՒHiV���鴒j�!����A�i����\�]B���Ϝ�N�)�����h�������]{�������4?�*���m�JEs���!̈́��_y���
�������)����v/jmR��^eёAȂ�1���O����e8P�T�ڍv��%����`�N&53�Ym�mko[�er�}������⑘ݺ��x����g���f	k�BVA_ɱ㿋Ϗ�;��Zv|�}��_����Y�@�y{o[hd�}?@���p��<����|�e��=�� �� �DϳF�*P���v��������[	����a�FF�4�����U����~�PR�0�n���S/����\z`˹]k�#Rs���Di�s�w�k�Z� 0��$�C�O������o��ԁYz��׮�����V�	¯=���X���l%bT�F��ء�R$��=��H��ا�5�\su�n���Z&gۙ�e�u{��/�׿�u;<9a�P�V�tpb~����ޮ>��j�u�;�-���R�a�SE��Yg,�����0\B ��] �����LX�]\1d�|���L���Z�����?$��F�W* 'ڙ�0q�v���u����q<���,&!�i�km�rQc4��p�p��6���Cu�Y���84� ԙ����ʖ�����T�jǻT+��kO�]p�n��o[[�7}P�j[m8��jqB	�6qH3?u�5#cXg��8t���d^[}�6�K`���NR�O�H��qhUr���9'�pM�|�UU��&0#�P}�ݷ썿��ݾ=�k�K����q����۲�S�3�Դj�h	|T�8 Q}sRWk�e�I�[��g�U�|������=[�p-i�qLh����8��O%8�wo�V�}���
4��[VAh!�(�5��W��˭3��Mݨ;7�!�I��>m�Ϝ�xO���H����1n �(����� ��6�9�܄�V([%W�8\o� �@|BSc(�/�N�y�x�&�L�E�d�f�1���)��������+U[͚T�|�B|�-i:8� ��ez��*nT��I�>������G�J&	���׷��V�n*�>���ҽ�N>ٝ�0T�h�ҷ��=������,����9�[���4c#�
��6����^@�x��	�!�P�����ٰtO��և���Z����_y�^������ݵ�>|�~��O-Ӭ��c
6X��<�"�$J�,$��d��}�˯ۗ_~Œ��fs\Vjeʹ�վU�aΝ���q����Q���^�!��Ru�����t<І/9�D��Ѩ��
Ѱ���C�f�C��u�+X�wzy�r���6�yn��v��]��8oŬ5QO� ?K7%&Zg�J��x�0A�=�J"Z��v���у��{_��[�z�/��ꥻ7wnqy����}�3���I�Z���w��~���X�#ԡ�5��ߩ�#�����pP������9[�ٷ�s�������v��!������l��ڥ��X>W��'O���D��aPk��rJ4x:\�|<�1*b� ���[��4��!3V0�?�Z��R&�"�@�"�!�K�^�+��5ᤪ��@��;���d���.�d)x����jMHZ99�1���<��D;�%�mP���%�1m�p#`��,�>�Z�������g�`'��@���ґ>���Ă�:Mu�,�N
!�-!�B�yF �=ҡ��%��)��� ��}�_���u��Z�O�#�������Z&g�lN�B�q���N^~����o~�NM�x��|�g��o�쭛���K@��i1� ��>&���*U�� �J����4�5!�^<{����x��=�/Q�IG�s��8(`b�����nY��f�ם�9sCGh�SU�9�[�<ZR���P_�>#����hWSeT��Jm�!��A;��3v�̌�	(&�/���*~��%�Y��;�Tp�a�r՚t2yiSS�8F �f��OӒl�fi��.�tmY��B���=>% ���y�={W`7Y�0�!�@��|�It?�t� ��<vLr����P0���I%��W_�ހ���t���o���as��R7C&��K�t��yu�w�L��ތcz���~I	������o
�nY(���YAPv�`A	�FH�����\b���w�֜"�nF�K2����a��TwZA���Y͜�}����+�}I'��{�����w�PnE"�@�E�&/��!uU��;-h���/~EA�`��bpA�ټ;���z���Y�磂G���+~$C��~�����fvNv��x�}t���a��GE}�3�W��!�CN]����(h4���>?�`̈́ז,�k[,$n1E�$O)f���,�5,G%\oi=$bkWꖶ�����{_���O=���}�򝛿{���	*��~�&�[�U���N������>zL�`�8�BG����0͢�}.�lj&���g[ْ�jf�����W�ԉ)��Z����~�W�J��ɗ����9sV�wUU�}�ȃl�e'�G���D�1` ���k��d�	����8�
P�Z�����72�Fk���T^�!�bӡ[T/���*B�ZT���l�0߯���Ʋ-gw,����� K�O��kB��y.*5�hc0_����r� ��@��ׄ���C(7���VsY�>�;����yU��2f�1_��?t�t�#�Ñ��{���v��.C�v��)�#�e*o*\�����Ύ��@~��Z�����cD`9c�p�����B̃���lsc�^{���׾.IA2m�7������[v��=6Z��}��5
��� $N�u�?S�,�B�	Zyl�@Kh^��#l!��c`M�ø��R�tg��1)��n�*'��9���a�`� ߑ�A�o6���������<dk�붛��^.+A	�X֟�Z_�J۱3�������a\���m�ú�  Q���ܴͭ����]�m*QNX9|��+�"W�J�PQ	�:�+��4ZjK��4sGT���I��j���J7~jzZ^�T�w��)��c U.�`K@�J�9�f bO��\��`|Be4<0h/��j�����oh`��	��G}h�_�Ю\���θ�
�D_�3u���.��D����L���C>�V>_����{֍��I�gJ�QCf4�}��E{��9�	�PI�zzm���~�e��$�x�k��_�����ܜ}p���Ϳ��zY� �<r`����E��*4A�.�|��/�f_x�e�t1y*ʚ��S�Ӌ���]�~�Em���4�?��ǿ;�w�ꄠ���y���	��n���*�GE���$��
��-v��Se�W|ڥ V��dZw8oזl��{̭'kd�g�@_��7a%���jK�w�����~�;N�����/�������z����{�h�$T��>���cᶭ,/�_~�/$[9>8dgO����N�� Q%ж�2Ug�ɡ
E��ڢ]��oK�{�_�Z�ܲ�_���gO��h�iK�쯿�=�3{�bє}����le|d�,h��`Zr��������H	Z��VH,}l ���^p��Dq��Ǩi�j�H0������\��5) �dӏ��VK�b,� ph.�n�G�l~oݶ+N�G!ւ�B���!q#��3
�-	��8R�v�-��m��m+m攽%��m�z-���'�!x�UA�K:�]&�22p����c�ܰN1z���+�
C:��w�jMGܦ X�(p��!�����E����e�`�,�p^�♇�����Oqk��9 k�\-�5�K|�s/���{�Wu}�̞��?�;�n�r o�͉�_ɘ�WT��Q��uC�\q�1]�x�O �3��̮�}O_�*Ԁ����Z�T̡04����3뢣���Ea<� #�L�Z�{�>�.-�yp��9w��^|�����[Z�;swlcc�Q���,���1IL<nc�����q;~괍O��.�Ҽ�ԇ�y�n�n)��_�/ܱ@�S�1����-�+��t )˺��DL뙟ת.Y 
��K���)�����Sglj���&l��]	��"��x ������- k�D;V��0C�޹�hf�k`j���^��gft�"�jt<"<�w�{��x�-�t���7�-�g,��BHF��U'�vx�:��D�&?qCx�
�g��r�7oж�4�wT5�#YY�q#�� N�C�~t/��0)�����TŌ��7��u��k�i=?x�h�]�h�w?��j�Z���p�NO�ׅ������\ޞ;^̿��U��V�ͥݟR�Ut�)�:1��Z�P��w���.H.$�����tgB!��0�0$e�s���J���H�G�����m�T�Ę`ׁ+�p�e;��;[e� �:_Yߜ����.�k2ޗKm~&���"����?x��?�����?w�.�����k����ʌ�Y/|^B�X��w6�G?����)?u�>0)�d�C�h��fMU��}ͺ�_\���nٕ{wlu/o�r��2e;s���9*�x�i�ˋ�W����;o�`¾�_�D������j��=A��� `����)�T���*����F�Æ�[#2!W[��c���H,���!͡�D@�G�p�.�AQ�(�� �e<���/�����1�*�2IF�W콻��a~G�y*Ḩ9h��֩(Ua�GGY�=�	Ph�j_*6*{�[\����ś!��Z$��1j��3+ּ�-d7ǎ����i	�Y3-�F�v����= $B���RD#�f��2$��f7��ZiG�ʥC�����h��y�MKPl70��,�4�->�9��LA�<m� �RMN68�0��«��9��l�O�S[]^�̉�"\Z�t ����z�"$��A��MpH�v&���q�����$��2X�z��G2�H�(��t\F�|���٨����� $TqT��x�]0sdf�AXn.���^�<������L/޸l�~𾭬�*��dCk��E1�{mt���:3c��A����b������@6��zM�LX 82�L��Zy?g�\���u\�!&p��o�(��.K},��d_	�r86����kǎ����Ӗ�첥�U�;7o�����G�-�j��3)YS�ϻYI1�T�u)�7K�HZg,eӇ������˥#����˲�%�j��w>x��z�m	�E`�i�p^ϴ��ԭK��U%Mt�|�o$c�Qr@�3na?�O�k�L���1�3�1�=�o����hع�9^?��u��A��bQ�;��׾� �z]Z^E���7
:����p(�x�ɉiH5d0�(Ul���Ɔ�l��ϒ��L"�(Vu-0å3��\���t$? ?/��$��LQ�{��R��Q�c�
ߝ��ءS���!a�q�P�U�;��_ݫz~��Wr�k=q��|�JH�Vs�_�(w�*ш�^�YN��Z�[Π(6��� �g��9���?���t����Z�o��wV)$<q��1K�:��3xg.����rs����;vg��kVn�l?W�S'g���<oSG'-�������S�w��a���_�gv��sʊ�H&�ֵ��()�B�v���5�
C�G�<QC�W-f����c�;ަC���/F�W�l��Ӈ�Y��P���wՎ����%e��
L�R��
�}o��2���~�,틯�֍K���m9����������d� ��z�(����jy[@���e�.�[}+gi�X:W�꜅���T�\> �J�-hF�\�_�:��R��kCG<�A�*��pH�Fy���D�/W�1^��4 `c�M��I� �����g�В�A�@M�۬6ĝ�uhR�\@`uS
G�9d�F�b�^�ݭm��Q)b5�sN/���S��-���<F�������JK���҂�o�8��,��	�T�PQ�� �!���N�/��K�5ь��f��h4p� �,(��Y:-��g����]��ao����,ïm\��L?��4����\��M*��T��`NM2K�o&�>&xz�^��Zqg�j���5̓Q�b���	\|O��܋�
�� U?�F���ѩi���Pe������x'��jr�Z�1� �%f�$�$5	ǜ�C�'�h3(vo��Dr'Z[^�5�b�<�|�}��E�t���c� �k2�U j;�	�u*2�t�p�b7��W���Rg�p�;^<���`$ V�O"f��"Rѫ�CACE�9X�c�v]X�>��N������BJ4.\�b�7m�弅RI'��@�/�'�)]�m��

XP���"�b$`-3\�sb�����FV����&*�{�o%��㽶�F���H��J�a�vC"3�Ξ��@e$3����_�%�$���`j�x��]�VC2�/��uG;dO�A�]��I)E�n\4$'��P�����o����}�S������O_�u�����cE%L��CV*f��ޱJ1/�сa�T�/fpN���) +E[\[��+K6��l����!E���3��s�m�Фu�h�l���?��nZ$����߶��3q�s���O��G�U�B��A�ꊮE@��D=�.-���n��Sq�}%��{�#�B$���	�~L�p�M��v�m��C���V����ԏx��#�:@Eb[)����h�';l`h����-��W?����Q��ʢF��T�U�Z(\���τ��P�̦�;�y�f���������l�����o�*C�&s ,��wJ�9���Ϯ;�x���t�ZD|V��_�c{-*e��E����4�v43`cn�+�w���Ц��"��4�X4w��6t�\S%���Ցhy9�Ӿ��d5#���m2*��WXy �ki�+�֔�(Px�y{L!�8��a�豽lƖ�V����Fl��a�3� `5e{c[*#��i����Zo��	wt�8�Oba?8�y�����ܼ*�N�A�I�h>d�F��|��C��g�ˠ��<���p@Q!>rԆ�����!��Z~�*m�:48ZN|�Y�[	0����Ѵ�^���᭪�y��BI0 $�HX	��.�A�����G���P�:$Ź
�c"�J�bI(oTԎc
�Vҕ	V�HMZo��b�� �1���ĺڮ�Һ�5�����#���-d4��V����U6�̍ <��H�moMSI 6^������j������N�i�؂�VP�u�N5 V�BbQ�x"�0+7����[G(f�GI#h�]Lr:24l=йBf��v��U�����rRI+�E�2�=I}�hm�� �A�%Hk, �k$3ҝ�>N�>~͟����'����j���<*��:��� ���qw��i�<=m��ٯ^�����"�F5IS�?9��h�����OtC��G7�N!�U�EG\End�~���I�;,�hx�����#���~���|�A���w�ڝ;<;w�*�/�����Y4�͝u{睷���W�����>�M���
�i�#Ps�2���m��
P�L�v�5�GϴR��g��W^��M�hFG������z������_�S�NYG"fW/_���yî~����T2!C2Mf�����"R�:~���?#��`<H��d�JE--GMqU"т����xԆ&'D��4�g��jcC*]T&(�����yQB-J�6Y0�����İB��Y��f/ۭ�e�o�ew�����dV!6�`��iƨ}�DDX�l ZI����V6m�����-RA�%f!��2�pmѶ�ɑ�.Aח�Tu�3���>��A��8��h<ꂸxپ�X�u���v)%I7�fp����C6�/1`~A��8*V ��e+�
BD�y��ɬ	�f��>
S,d��BX칄PmF�̓֕L�`U��SBG���?{ �.1!�����{J,wr#�GL��3�%�P�5����OM�� C+��h ;     IDATmk��T�:I���̜;`v��Iݿ��E�tᢵKUw���X"��B׋/�d�+��Ï.�����I�J�� %�aZ��*dJ%?�(q�CAqj��h	�x�y�7mh0 hJ��źC�����'s:�I`iG{*F�{ѧ�l��[��2s[�4a���D���a[U�u�2`"��(zNe��>sW��8�p�D��q0�@5>>j�������>N�������� @⿄��W���ޡ�S��e4_(���C � ̙"�=����f�������?2)1��6�6�|�z���
(1▐�	q�c�{��9�mm8t�o{ż���I� o�K�/l>ɀ��Ǩ�P�����c
�����J<%�ޘL�':nrz�2��E�f��yRlY8� �T܎��L��/;ߪ�#f�o	�0'e��ģOQ��&���
���u۪قU�Y��B�xh<B��3e]C�nVlm��֠�;�!�@8��z������߾�ῼ����w���;�󟛚>i�>��t�9H7v������L�U�(��%y���#��1��z��M�q3���
�i�i��v~�}��svxd\�,�?��mv��2�_��/�铧��3e���ù����f#Ãd c�f��0��޼�>hG=uzFAx`tX׳�����U�W����<^7�G�RQ��z�v�ښ� u��������!��!�Ws�"6#@��ݬ�����ĸ�N�X�*6��HA���e�u+��֒{���ʠQ�!��ޣ%�܄���{Ô�������7E�O[�"�x(DHZ^{��\U��&���9|���������tGqld�:���-@ә N5��u�A�����Y�'˩���;��������70�9RЩ
N������3\�b�u��vt��I����uZVf�uA�Q�kM�Li�zj��Cxr��s@2Ao�X���+�����lykUm],��=vhj�U�M.��?&U!Ѹ(Q�@�9z��AP��*	Mf�'PU�ݓ*���js@��������r���ns{K���ͻ�C�$5H����+�יp���q��5Pu3m_O��J�^iu�Ƽ�G���!kK7�b<!u%�d��H�ũ�^�#ǎ)�#@��@.�4\�P₨#�$I�t�{�����_�=#
�؀!�w�tO�{�9�'c�Vc�.�	 �%]#��¬+鳇]�@G+SUU�!�9�f�%�Z;��gNw܆�o���-�<��d��� ���G�^�YJ�2�!3W���%��`_�"�t�E$�.[�D�3p��n�s��< ��%�1!TдyI
@�W���tư��ѝ��y�>Tmd��� ț��Ȭ��Z���3e�Μ��6��=���^�k@+�B�g��oC|%;�	���"kdrf���f������#T�fn_m�����`$wP��G$�)�p-h���������G	�߻���kw����{s/� 80&���֪]�v����[����5��^�F�����J�D�bj��M�$b�,ڹ�g�;6qHY,�6o���-,>��/!p~�D�WPq�X�n��#��V�L��*ts}Ӯ~|U(Q����3�k�Jb!����ҌP���,bi$�M�C�bf��&$�R�Ж��Y�U�U3���R���2���� ����C)J6y�;}�:��,��ۃ�e{��%[���>�TЎh� �IP�H`,�Ӛ�z3���V�����`���ֲ�]�#A��O��6���1!>���Ƨs�lߵcE��ޠ:�mEg  ��;�:�?�>P��T��Ħ��ku� ��y� �n�P@�J��<㖂1|`�,`��B(�D�j�y/όM)�hȺ��֝�ZT~Y3.0d��#o�Tň��S/h�Zӵ�&��Kn��3�Bs֣A�u��{p�BH�R-'�@����Զ <���%u�c��	p�=�M9b�[�%��}G~�,�ӝI;:y��y�h�G�RIk�� L�T�� �BA.��>�deM�h�?�b8���$�R �`$h�h� L[Se�K�\A����M@��%PN����5��-'�a����{T���Z�#�%mP�ۄC�"�9GZ�x�RY�)f��έ�4#��L�ì�ψ��������s�I�X+�uI*�,��=!|9����,���_�"��djy�-�)�^�_Z�`SP{��Ʊ:�oW���<;�O{4��K�%�^k��dqu��ڃ�GJT�P}Pl��`)8���լkh~b3���"����tJ��%�cl������)ºT���3�7<ʦ�}}xY�R֓���vh�"�G�lT�	�f>cۥ�m��C�#&	�?fsx���u(ԩ��-�[c�*��lמ;��li�|�m[��0�G,��+���)y�����e8\�����������.�����w�x��q��˯J7s���U�q몭����ڪE1V��j�7J5���J�	4����'�twZ(��j����I{��Sv��őj��U&GE�����ã�Nu����ڲp�i�&ɥ��*#׋��{O�F���(n��:E	h{sS�E�-��1{�z���F))����uxH,��l�n�U��m������D<mC�c���-�hKp���S�NX�U��̪�w㒭e�-[Et� �:���2T�6Ί0zSo�w� �\FJ�GήnZym�b��%����e��h�U^귎$��D@@	�E�,@��_��v;�d߂L~�I�Р�fc�Sy���W;� Y���k����Ek�Ϛ��}�~cx�rm��ة�/9�w�PP ��ǧ����74~j?��9 ����!��ݹ5kk���R4�D̞9t�me� ����O����P!�,ִ�����<�v"��Y��G@(�t�zA���{��'�B~��`���c�Ц��ǎY%_���e��A~`{�����@�>+Z�J,������FBU����=P�/��|1z��%H"%K��q���a���ZM��P��OP�!b��Z�a�x��������K۟�Nz;�S&�w >*J*@��'�@���Ǻ�[{�h{�0�(�:	y!��Y$�I8�T�^���>3c���%�=�����Ċ�\����]�r��PԞX�?�P�Ev�B͖�@ͮEU�Z��
^�J�o�|����O�c}��3������+\��y��z:�&?ia�)D�Q���������tB�=�g(�.�"W��=Zc2]g�$K�ϛ�@x�=ɍ�yѸ�N{mo񿱍�+�j:f<O�D�"��e��e�̫����=�Z���l���Z"lt@NK��1G���\�#h�Y:�V�(�{_"%w- ��]�P#%��@"�������G�,�G,�hYo0v������s�q�����MQ�����7o�э;w�v��q��&������a��^�G�����.�d��T�C�q�ҨDA��'�
/�#a�XX3��c�v���L��h8d;�;v��%���T���3�ڡ���D���۶��vv��ꖊ��\�qf�i�܈�h����' �CiUP&�.$iȡT�2���<��c�Ѱb�j�Hܒ���4����B�(N�^~_t%�n�����E�#�i�x�b���T`�:|�N�<n��+Fk����ms�
���[��`n��7� Ԃe��x�J���59� �g�K5��ܱ�Gk�[Y�P�n�@Dҁ���P�^P���~ˉ���9$9��������
��� ���j	ˑ�Yr�\{��}��d)
����{����9����Dϙ��A�����%A�j�Ҵ�@�#���O���3�Q-P����Lg�#��C�^Xxd�}�U+��&��k�K���z�v����>���0�=�kx��%z:-�ե�6��F����94 t�u��EĂVÙ�޲��a;y��=}zFZ���v��[ZY�Ÿ�DR]!��If0����M��P��/ ''��l^��T�ܮN�P�|�2�eHO����3T�o��8M8���ѧ�ц�+���n��X'�����ĚB)��+sdڵ$�$�B���փRX_�S�j:)G�aUV�g�Qoi�0��h�c��*F�R�x؇Lx3Z�9�
���e�
Њ 瑌���%��$�����5[:�d����%]x]'Uyʒ1���;9������ɀ��%¬�_����i}^�E�c �A{7\#�Ͱ	R���Ҿ]��M��Ob\��p�Lymj���Б��P����^��0	���hDi�Z�_���}���m��;�Z�A0���Ϸ�*�Bf�./���ΚeCM+�LjZ�0��B�{���@��9�{�I�f�.;<qPIt��rA�s��g�\/�,�!�����u�7���������_�2p���߿y�M���=��M4���}p�]{pN�Ն�Qɗ-���6�,0�ghl�z�,�j�V�j9�+;1u��?mgO�(e{o����[�\��s�<m��5���y�ݻg,0	K��\������q	2���.���km�J���������e�N%�q`!���UmK��K%ThE�Jym6���}pᢕ+lR7Q��&&�r��Q�>y�����,���#���E��ߑ.n@sD���2	��tP�2�.-��c�t�2���J�(��(��-��²�<\�v�l�&iSӒ�`��$`�'��S�W/�%�{
I�y4:n��eNˬ�1�	�W"�3�y�Х�N�9�֢��}�g��V˚��y�HHk*��p�EH^�N�	�3s>�N���|h�PF��1
�5s�d-,9�`/�G܁�����bթ��[���͚�f5S��r
¹f�"])��v���9diWv��d8�5IT���//>���U��{�b��}vv�=7��sE{����W�7u���kޕH %�fɐ��c�H�iA�sBM��T��Z��N��9��=��N� ���}>����'ڦ�:�J���!ϝK�&�G�D�}�� g�٤�`�|ˀh�5���t�:E�?��`8�Y%���ѝQG5c,�Mص�ᜣ.�H�������_�3��$�S�Sk�_O52nQ-W�=9��W��*`9M���i�{��0�6p���q�.�	c��gN �[H�	���6@��]�\_E�G]����n������(����_BGN�A�]��'nf2ˁU������j�g�����~��v��X
���S2��4���х��_
��Y����vec�2���"�I��u�ydfa5D%��gj4�3�yH������f�d��4�θ��_��2ˇ]@RTo�ƞ������~�b��裾k7���{�<u|�>s���i��]�p�{�`�ʹ������R5jT�e!����<n��C�����6~��m򶰿m�F��M=nϞ��3�'��w����wmimI��8ć��v����׵�V��X� O�#���a���������u޿�XĆ��V,���,��S�W���N"4'c�`�WQ K0j�Ŭ�T�p�AKj�Z�?��67w,��[GG�8(�ܟ�>sƎ����C�-����#�[���̮\b���l[��b��8v�mٖ�K�Y�����f����/��I<�ְ���YX�V�dI�d����H{Ź� �Q���F�а-�" Qu��#��p�A_|���e�������C�)e�q���ţ��0��V�'a�6� ��ô�\($���X����T�� 'W�A��0ɕf���f�R����_��B���d�yED���s���9@Z�s�7�C&�L9gk�]!7U	3#OD�CPR"a��8dG���~Z{;���m�χ����Mi���֟�S����3OYi/k����͛7-Sv�c����CR^��Mno�x:���̛ۻ���b��#�gP׃���=�p��s�}:��
�6J�9	��h���<��Z2�z\I�2s�{ȸ�T�ݫ-��]�u����[Y�l]��<w���T�	�
鵋�U�Mt��]�|Q%���m��p�	���9o�#��Е���灳T�;c 7��j��IZ���p��4��7?�'g��x%N�O��r~.
���0�BZ�U*E�����+��{���F[����*>�&u}jg��ϓ�F"�$ʛ�!W�H÷��(���w�m�z�up�v�	��37������K���e��S9!y��$��O��*Dr��=,�ڻs7��E���V��E�˧$�|:Mā���s@{h���VJ�:(� Z��9�.�&�0 S�|��b͖�FwN�����w.>y�!����z���[w���콹_<>}�^y��6:<����ݷ˗?��G���V%���%� �*��L���i������){��e�7�hZ�V�Ƀ��矵��O������G��åG���g_x�&��F<�u��޶{W�Yng�
{-L��y�̈�%��F�Ri�UF
��#�� `�	o�Q�~�1njV�K�R�d2-�t�1M�";�`Go��$�q�=ܹs��®o����`$��]>82`��M��E&p�����5p3<�8!�F3`�
�����S��1K�X�#jŨY1زF�U�p7��7EU
�B�A�!���0sk8^0_�9yU����: WP��v��y8\��fV����_�w=@U4� D�?W�xT(o.	Z�S�~eP�T��2��#s��3��N�������_�n[WGJ��iO�S�F>�U@B�Q:\/_�Ci���b�N0��⋙�ڝ^&�&��+a	�[t�0�K�,=�o�g���"��={Ξ>}��;�V*l~i������F6�$����?���!L����A���sV��m��=�y�me���<qlJ����݌���JD@asPvB� L�M:ܾ3�4��
ר ��?��T)�mf�3U�g�$���LdU��\�}�n�O��C0CA7����� γV���G���u�l�n�{�f��R9C�����s�����~��F�N�7Tx8�nd����N�����o�k�k-�5�J�Z�D���<���ˠ�$8w6G⋫���P��s�؅�+�KWѱ)�D�u$8�ԡ��!�g����}*��C�����mb��L�s�4�h��q�s bO��#���r����9�Ɯu�}�XU��iE+(#!�}ٵ��@M�~�n�g����5��(�1>:�I��E ζ�I�YJ��k��Aq�ޙ�iW��-3+�Ú	�$*���u%Oy������*�����*�liћY/�wh�G#����[�8�0��~n��?��?18�[���w>���'_�s��^yg���7�h�޽_8q���K�0��ٶ��X���;��p�J٢5�u�9�i+r3iÍ��� ������l�J�K��>xȞ=s�NNW����mo}�����^�����؄u��6?{�n\��ޚ�r&�P��d���:�s����(+%ب<Ģ648�kwc�J�a�z,|�!�;҅���ba��NZ�Zr-NT��szx,���.�Lu���m"��ٷɉ1��C���,/�鼉�q��m7���kv��Az5�*�
�^�[]���=[�fm?д����z���NY|���}��"p��������f�V��,��!��H̊uO�O��U�>7��Is(�Tu�a跒@��=�b,��0��G=P���kR)gE�D$��p�:�D_�h6@���jC�`�[+9 �'y��C�$���2��^����ż�!�� D��: ��+����*a�d��c�l-}-Z&�Y;0��,	���m�N.eՎ��8+J2�*��瞶gff�U��=����~������d���i�b�1�=h�'��s��Ze?��~���$8��:{%/H�:��- � W�d���^>+
Z�3���hFº6Q��u}�/g�k�$U����:D#�ٙ��4)q^=�Qw��\�T^�i��Pϊ@)%:O�=�{��g��;R60<�%f��� �ǣ�WRdC_��Q>5�d    IDAT�̏�����(PS�� *Q��j���:k����d��JU�'�d\�V�ɵ�֭�������Ob�p����K<D�7�g�PҸ�'v_YM�C��3��Y��
.T�b)|r��fኣJaL����ą����{z]����z��Δ�d(�[��R�]ZZǝ �s���X��(Ja��Jֿ~���P~rO"���
�(��I��T5���P��GG���P	�w콇��ޣ9��$�	Z�V�LٍIܽ��5�J�ٻ.�f���č�~�K�|A����p�H䲻{��'��O�d��������Ư���a*�k�n�������<�Ͼl�M�����.��B[�R���Q@�EӇ��V�Z���'����H����I�,S.�
���8vTg���lys]=��^xQA�y��{w��ŏ�Ү�� & t(=�|ffΨMԨ�,��5�����ʚU�9U��1�F9����<�!��\P%Ò�+ʢBe��:�ɠ$F����f��M4jv�������^�=Y�T�
����$���C�	Q��x"e�H��͠�f����kk��jT�Z=�P_��>f}�-�B�n�+:��#	K#V��-�����a���*5d��/W��7�r�!�*<5�:�&p Ti�Zu��|�Z<#�g�a��P2������@z��T��W���_�C�[Z���8I��H�V�Rɤ<�G������ݼX�Me��N�r]O?���������W�&4+WE�E�Ń=f�e�> *�<�s�i�JѶr۫-��m=Ã���u'x履zƞ=}ƒ���sr�fneo[Hw��4pkj�{�w�N<���sq�=���LfO�o��rU�*j�Z��TR�~"GKs_�1��@� �¾`�c�]7 |�0A1!	��Swt5�D�!U��f� �bфC���z-C��ހd�;�_w'�v)�,(�R^S���{����x�AO�գ)1w�-2�란�5�����ۢDěk�cy7�t���O:�l�gwձ����ꗵ��4bB��{�Z�/�0��y�z������%��{O�# �嵫2{Ba��5$K�U�<su9h��c
�C#Ú�S	�� �9�����H>��ڊ��������}x��RE��W�KM�N�� O���xq����p�Ft����K)Tw�.��X/|�@����PؒhHh�3g�(q�B��?��r��W�K�}��t�>\��r*�p�oCx�`���;�O2�%Ѭ;� �[��Aj{��]
��HBϚ}�yR/;8�tL�ӭ�����?��o��S���ƻ=7����nޝ���S���ӟW��hgg�>|�}�׃4}��̧�s��Ӫ653P�~��	�Zz���c��LJ2���	{j�Zm���M{��mekC�g�~֎��ގ�-ܟ��.�ͫ�,�횤%i�V��9�6v8вAh)����hW��3�\�����B+�I_:O\f� (]��BQ���\A�N h�b ���4ԙ�bfǚ��%#;21j�i8}Q��ٗbk._��R^D&�m���࣡c݁Bª*�m�em�X��p�]�F2� |��6~jں��ā�l�����+u%+�xl���/����#Un���t��f[�`i�x��j��9�
��Tb��94�c�ɱ��YT��3� $���k�}���t��x�d$W����mon�"&X�)|$��pKzGV.�ܹ����a+�e�s�قj��R��8xi�1��e2Z����'pnt8�/�C�~�N�ª�@�ڢ5lf�-ۨX�;e�c#C�� Gy��9;7}�ҁ�|iWv��?���-�[�^u�M���m�o؎�N���g������ma�r��C��V3����ͮ��cQ+�JBa��p�8y`:ޏEAأ˸`��GO��=�8	*S�9�9���LIL�n_WT���ۑ{�ڝNŭ��3��:+�3�Q<�4�]Ã�=�o]��j���'Bׄ�F f��{��)���!�����sb��ͯ�� u�3��$~�g~�@h�셖*��UR�bL �G�����ԸG��R�=V��t��DA�iG�q��rk��)��B�]��D\I�ǟ���I����ú�{���������#r��􄟿��bo���}�!Q�_7�w֋�8�&[�>����"�&��eN�wE�
�gý�iPn$���T�ǎQv]��@�O=��t�ֶ��]\�k>�k٘Y&�g�Ź��I��om����\{���5��{B������:8 ��4e�w��E��1l�m�l�����O~��ڴ?���ݎ���,��_����w�G��^8��M�.������'���#}�Z�Z�unX ̆����6���uvX�����{$Op����x�1z�م�licM?���Y;sdJ&	�؍������Z�T���� ���#�Y
�]�.��щ���r�{BFSi!0�6���.Q&�x�;Z6�E�]�J�ʥ�T��X7t��.;4<h�f�zQ�IŬ'�f�,@s�]x�+U�5���HC���*�u�,L��s�*�h6�6)k�0J���6q������ʚ-=\��֮g}�L�6�֕���&�̥ ꣓=^���K������%ҡ��� a����[R#�(s�|�k	�z���AnX>5�
K�HܢB�Z���a�kC�\t8ӎ�gjl`Z���;���t�C�o:Su�Q��^����4�M�P ��ߡ���U�K����=�o8d���6��8iI͡�3{B�ӎ��X2�J���C�mfz�R�t�يW	?�^�Ij�*��=�vx�0��������m)�q�e1����I�xsH0G��{!�Nɱ
�	F��P�M��B��0����s�3QF�����,��:��� L5GNE��#���
�Q�xO B~���z�`��P� ���I^���=�tʆ�G-��%��R�bZ��Ui�6�:���?�~Dbh?�2yI�6�%}��x���$hZk���|�?�I����j�����U(,7�p�8$q�"�� mf:����r�7�}��%���	�*v�n��y��:%��h���j�{B��3T�Я��������	;=3�{���Y���{pA�$��5����<77�mxɦ�n�{���S���&|"� �}�t�]���XS�y3���P0(Eħ��R=�ֈ�l���+��ң��O�a�T1+�����FD�BJ��t3��p	.�Hi��	��Z��ך���mM*a�!���������7�{�& ������p�Rǥ���+�f��ġ��+���?6%�����������c�Ri���C���WMm_��!7�A4��H_�|S���<l/�y��;�m�o\�PA���K��'�n[ZX���Y�3wWm�l./�(d� 0>��a\�[G8bcvxhL^���J͵�%_�K���&D��s,	�1yA{L�[l����K%b�ۙ����v'�'�a�=i��LYG$h�bIp��E�X+�jV�4-_��YQ8��L�Y��V��9 �O��-�R�-ttlx������C�����Ҋ�R�7�%推;HY��R�"�]�Il�X�,ڡ@]�/@�ِ)`hN�y}1��؄NѰN�⚂�KJ�9�L�#��vh`H�yÛ-SY3�e.�f����>�:��x}��d�i�&��pT*Kz]�m��H0ƛ��q���i�Z�z�����A7�θ�X�*	�'?Hі�3��5$�Ќ8,$"R*���f��Y,��do�Ei�vt���6<u�%�f�r�V�7���}ۖv7=��Zfr����6u��}���ݜ��.Z&��(.��8�h��s���V��=e:]긂~�9O�X�Vo�}dT@B�Q@޵⅐������U�֦�cG�*�v��?|��戮v	K��D��<ɍ@@H}zjM��q���x��D��kQ*�2Wٹ�C����;��ŬԬZY.Q��dqc᨞c9_�(�/��`6ͶuF�+�ֵW�� �(J2\t���
́��C��ଙ-�$f��6�yU(�VA�V� ?Qg�V�l�;���RU&:�ks;�J�Ni^&���d������'hd/8?N���jMv�X�N�ͽ=�626*~�ݻw���?�;���VmhC����^N�ʡ�y�$����RW��*hVM�F%�#���K8uN���Z|�6�L<�>'@=T�>s�&��[�;�����y���`����tۍ���a���V#AV��^c$�p�.N�x~\�P�tAK�����m�"W[t�x�,���9�/�����/>�J�ͅ7��]Y�חo���c�=���:1� ���!�T�r��AGX/*����kOϓ���q���Qsnߒ<qtʎ����=8��o}��-m��=uf�N9��+�����>���ei��KV�4`Ɇc�sk�,�,�hJA�7��v�q�w����sb�bq�&GȠ��&s��%�i�ұ�%�aK&�֙NX_w�F�l��Sx��Ӻ!$��v6�����py�ֶ�V(֭ܠ��u(e�������v�b�`S��H�a��TLݣ#6|��9dA�0����Qk
"�\^�+�c>�D	��NX�O����PO�^��ղյ"I%�^�K����.����� �͖u��m|tԆ�-�L�#��[�j��.w"!ʛ�ohE�ګ�eV�����Ʉ~��:��Db����(8T�f���|�jǽ���:��_���u%lFG���l��L��TJZ���}��E~�a�����X��:�]&��d4��pdhКͲ�x+�jG3����몦 AH�ډCG�_|]�A�.������-z�d��M1�;�E������4 &�I��D�>�vf��v5��G��ha��C�&��> C7$��.���꺒(��ylӶ�x�Ҭ���t�e��*�>�kw~2�u�Z�B�.����c�1(�fq�Hcʨa?�6/]_x��t��D=�I�S�s�K������'��#N4�_Ry��k�kv��1�%	CG�	� Rì�.
~�$o�坑̰�R���R�z�,�k��:R^�g%��7�&s]~{ׯ��� �U�q>׍��+�߷(�u`cR)=�G�����:�����grhe��pؓ�z"eO)K���<K�s?P�8�y�?Lq*��S�{�3s���Q�V�XG$���`o��B-�֭@���C�U�~��-5����F��._7sV��)ΤT�U��ZӲ[;
´��<��Z�n�W���W��O��S���;;}0�_^�q��8�:w|��͜QX����¢� ��dz�phU�umJ
(t"���R<n\��p��1yR6�?`c]}��Z�^�l�ho�-��*� /7up�z��mmmU�� �!i8x�ea6B$��ζ���V�۳f�dHvD���n�X!W�H�	�|#�T$�P���a�P�:�XXEl�Ö�ۓ������lh���{R֝JX7��R�ʙ��wˏ�mv��-�gm;S�J� �e��b���i�ctQi�sY�Z��ښT�\�$��>y�&Μ��c�m�Z�m�-�lZ"ݭ6?`}}C%0�r-,|�u��`�,ݑ�b��c���^F�Mk��x�'��"�!P\J~@����%jU=]���'$t-���є*mQ��n\�� ,:�?��7U��RE��^��eɴ5��J��T(��H�O�ǀ~"n�FK���W�;�ܾu�fo�t�]S.D�� L#���A�$5���^1KvvY�����ɩ���P�kR�)�**p�x������ۏ~�whU��י Ը��m�]�2���o|K
t7�ܰ��xC����N�C�fT� It����؈S����nmo��'8�� LU�SF�<'q�确�qmS?����ёUр���r�l݉P(ك��
g���͡���φ�J-� �Qm�ݩJ�F�]m��`#��}��Ʉ�0t��8=zP�{����{�,�A�,G������}���	�~����y�����N�'U�R"s .��ĵ0�m��sH����\�>�u�% ��2�����*��,t{ֵo%r�N{��m�l���n�L�T�r�adz�� Dk���Gb�x�*4��t̐���S��P ���T�Q�Q'D�w�y�k��<:�<q�=�XȔ�.<��PHcA�bkU�_�΁Q�	�@��C=�����\, _v�:S2�P&���}�̚�ٰ>�q>J�� �3�hsT/T-�nE@A��]>u`�_���+��ԃ�o��0��?\�5�o�&v��:iO����&��e�t I�AKn��y���$��=���d�S�p��]IKXF���0+7*������ʒ��3g�ԑcB7c�v��{��f���vk��p����d-��M�l�Ƞ�/�m�p�o�l�[v7�f�T� G͹�T���N$,�xg�����H������h�����;M&V�%��b�j;[�_���meiݖV�l'S�|C��E��H�'��� �Ył�%+�K�8�">-$6 B���'�sl�zN�v�b��Y�ް��?`�ccV(�ʕ+v��E�9 *-e�ڈ�yŵ
�F�� L������,�U���hA?ªhZj�0��L�A4��o�]����H�2�	������]Vjv��1����gm��=�Xd���Қ��
�IH�%J�0��E%��h��~֙�ˣ5�����agW�~��~CH�����29��!��&] >�z�Ƭg%�!w��9S�HF����	;�̳6}��x�� �@4 .e�a�@�6�{������?HoW��=�b����i����+:��n���y�e�y%v�z߾����������lR�LQ�%Y�D{$�@&H`�LL#^�1xl$��1�d�$�x$Y�$RII&)���}����W�����{�9�{�;F�X@�Iv�����}�w���������ޔ��^l�p3㓈G*��RńW$bA�:quc����>Tѕ� e�T�n�!�H�`�w��$��ڈ'Ff��<�闹�����b/Ґ��xp��L���3o\���v��94U���f�
2��FW�,���v�T�E�VךAn}��ds��F6�~>5�]?�X�d�ڰ���=�S�y��<`�K����q�5F2�3�/�O�aD�A�p�Fݰ�{.���L��le���3��j&MK;E��_���rO�g�xI�2�VZe�q�ޟ��m8.���@�Ū	B1-B�f�R,��\g_'L�31�V:�晭C>��{����c��AD���0s����k'�TƟ��Slh��R7�'�Eޣa��gˤ����	�H� �(j�v�%"�.#O�>\v�f����M�"2ed'�����tNb�i��T�Ґ�Q'w[KO��'�◿���ѿ��=���?����&���Ǐ���#O mE�8(FS�M�'=����ٔ�c�pM.��.t�{���(�غ�A��mcuk������
��'���# ٨\�9ܸw�܃������"�Ш�M-��hUj(헙+_ۥ.g ��'<�i���j�������]I�b~��i��cht ����.3��-UQ�-"������`}m�{%*M��|�~�=d.F���Po����sY�?�@�Q,E$N�j!I|h7��{Q�C��G��� ������H�s�!kg{K���n��e���Y�4<P�M~`��)�Lc>�EB�dTk
0�>��@�~�L���������^w0��m$E�,����L��߸�+��C��`?n߼�ٻw��Y�6��S��F�R,�C�2e�
j��e�Å� Z�z@�%9��ĳH�ݍXqk�˫Қ�{���k�y��b6>$��6ӱ��uv��@H�a$Á�q��������Y���	�����K�&W��ƛ?5�n����/#/�'��ٓ���(��[7n��w���ܼ�Č�G��>�tNR���e~�,���+�kذ�.i����M0x(�XE�7��D��͉�$y�q~-Z	E��j$?1|����urA�By��AG?�O    IDAT "ߑ�i�u�2�S��:+���Af)D�8�0��^T?Lh"��Bj�	� �����U8� bh h>_��<��+�疚({%�Ɓ�?kM�������?WS+#�����;D���-�='iH�?�e�]��G�1��iLL���m~��N�[�lP����mxvSe������h�c�0i����j�!O�8�����`{�hV:|_�\�P��Á���BG
(�� .@ѿ�R����@�4l�)����L�Ō���sa�SG+�+�;��#;������繣���L�4J+k�O�良@�kT<�jK��DMy^��F�ʤ?�|lp���~����'a~����o.ݽ�Ͻ�@v��!1���C ;e���bl�=�v�9��Љ1���q��G�؊��:�>�ܬj^YYӎ�ږ�G����L�jo��[���2���=��]'�����ֵT�GH�BÆR�0����i�Mvr�
����c�_���B��F2D<�8w~�-LF��e��k�U.�������ͭacm������ڠD���W4��*5�<��71;Bn�XX6n�hXd(����4��Z~�R�.w ��-!B��� R�H���=��y�..b}su�������+)oHAn��v���9QУ�,�4F�l+OYI:��y����L��f܁�2pw�d��a�^�1֑d��:\"�G�04Ї�7oj�}+�L#�H�eQ�41�`^^˞�e'G��B��P��qjKR8y�0�D���U���fҢ��ċ�~Y�.�3�#���΃G�>jX��+A�%7� �����Cةo<q��hH�R�g�<	 d��h���_ZY�G_s��	Y����r7>40�3'Oዿ�E%�ܹ~��3�//Ir���˒�{g�:��s7V�F�ncB2�.]A����%X�6r[�ɭ`��4����ȃJ���97��ܽ�^��_+wj�u���I��$���'������EXM�}����@E�òF�x6ݶy�M�CCLcNOmN�*���d��`�ec��y��u�ٽ��5�u�(�b��� J�rރġ��.��t��^E�����]�_��X�Z�Z'b�/]?�V�ۓ+?S4�gfZ��"��	Pn8/�V��`&P;��.̂�9�W��~�J�7?A�W��� Q �8�T�Lm�D�fZ]�������r�[��v��q9�����C�Y8)jl���RqYdǆAg�\��F���0Fp��wO�
��1���9!#���dخg,O��K$�G���2��Ǌ���ql+׎����ғ��Gg�ړ�sG����wfG����|���έ?nt��^й�5!)��89P|/��er$�d |���|�l;�A�;��	P�ώ���z��v�zYlgR�}^�x�ƹ�#xbhJ�`�mrvlc��b�<L�j�=Xt$щA ��m�A�
%�z=�E
Zw��jT��6Ѭ�V�G�V`+"A/�ɨ�f2��i���}h�	�屳�"��{��`ua�k�D��x�M�o@E�I�{|��-ྒྷ���"4�ُ�a$+����Z������=p��F���Ȍ�`h|SSSr�!C���p��a�d!��"�o���XQ�B��e+-&�_u��Õ��$ev�$ݐ���b�o�'U�i5��ԟjU�G}�'q�����Inp�ׯ^�N�1��>���I��w?�H��� u��C	�9�b�:�!����=��M����=2eە��0'�N���ۋ�l��m$k,T��I��w�8x�z9�a"����14:"��X<i�ݲ04�0��^qO����EM�|]�ܦ�-,�p��=��d���翤�J��������
0M�GL�� ��HT��^~_��N�Q��5;L>�|o��`�-lmoŢ�^�d{2t�NDj��P#������0�yp+��2іN.���A7��	�ϱ&f{:�t�!.C6�"���2E�mg8;�����Si�	�����Ƅlug�lX���g1T�`�s���A϶?TCeQM�6��iz�
J�����!iu�B�Y���r�p*�F�>��)��f�ip��o���&��I��u�i2���^�)y=�ܱ,{���%���u�/���
�������sϛf��߫u�L�`,ou�ѫ�ps�T���~6,���v�����P6W���!FJ�}�3}�"M���XV��0z��1�xͰ��߃��D���`�����$N)י�ym�]�	Ż�*���pvu�"��;:�nȎ���o�Ӌ;����{�?x�?�������n�<��x��IE�Ad�J�Ё�����K��V~�O�	,��>Ī�EIE<~BЕnC��:;o.��:�0�9�xr�0.LƱ���͎I�	(.��m2�"������R�Lm�!�&�zA:l����Z.�v7*hsZ/�U+i�|H���H!����J�7onF�m氽����l-���W��n	�j]o m��D�2ݝ��M���H��l�k�CpG}K�Z�����\�cae;�j.�����va��D���ءx��I�>}Z�Uժ��=����J%aA��R��G�44�X����@0uxB>:F������{7N>���!$3���ʸ%|J͟􀭮}�`ѩ�ב(xp@)A4}�C;15�Gcdr\��?{������O��/d���q�K�7�� ۚ�d$�P���(��=&!��Pk(uj���&��B:����݄g�?%����1���D��f�Fq��N�,���O*"=��B�	i�i�et�����|�RU���/�����E�~�ɐ8	��?g� �b%�L2+$�e�~�PM�H��ǵ#H6#a�MMn/o=(ómP��u�l�D6wcC�R<�-�(���v�|>��g�E�Dۑ�l0f*3��,"b��)n٤,B�2�`���	5�����eT��N�&�+Ru�0�?cB���Cܙz�lr��(�@��>�f����⫟eLj4h��qM��n�q��&g½��~w�(�Iڄ0�����%p�g�e	Y�y-��M��3�ƶٕ���]�0��9��oas�X����N7-s��}��6k 51^�~gL::�y�s��%��+����U�x���̛�iұ(�r��j��(�EX׮V7)|U#��D�rK���ky��a�%Ѣ���b��Vد�\�g���aTn���&�ȭ��4���p�0�U֕@�����9���ә���^�P�9���߫��+��o\�;����Q�]���
�&�% =��O㞕I>�l�qB�c�Ǘ���s��=a���zY�H�oM~-�R1��ϩ��i���cxj�0�����O�;���������v_�Td;���n(Z��U���)�U)���mBp�z�\�
<=j\�H�CH�"�&Bpq���Y��J>���
6�����Ge�����]/��z�j7{ܽR��F�U�n�7+!f
�pX% =�KM�*$#T� 2
	[�ܨV��&鈾�L�aQ`�9ܠ�wdf�y�y|�S��aI!6ED+6�r���5,l�`s'/�������0��7���RT���r�^cw�f�B���vK�ŉ@g�Ӫ�?�Ӗ$"��Oڐ�i�R(�����	�����
#2��DvpH9�\��]���rY�N��t��>�LΈ�D��"�d,��4	?<4���l��ɝ�T+汿��'r@�6�
C4�i���������z�,v�I<�'��S�̪���E��(�!�$9���$��w�@��|��X]]Uc��/U��{_y�,-��s`f�>+^��Id�IA��tM��4ҙ�^7��~\/��;�����٬P���u��T��<i �=�x$L2��_;uN�+�*�DIX�8�U�T$�w�2�0d,����N���[f'(�#��f6EA�Ǧ=��v
��GQ�,��	fߨ0Dֳ��3�;E�;v5L��y�fp����D�U3՚�)z���}y�;Z�]��)���#�|L;�{��2?~��ִj���$�YSH���M���u��S�V,�%SP�}���5,f#)r�z��ku�xa�՜N��S���S�h�j�	��/���>� Hff��BjĆ&��"�J��_�$��M8\ȁm=�5��AEr�P�jY�] A"�����QHD�d(��m4�wwP{�
Yh|���Ӹ��*�R���p�J$뒋V�n��TLs�3bS�{V���˿?�����ك���/^d�����*¿��_|����?Y�^���j��H-w�v��3x��B��F��B���Z(JF�Vfno�2�$�p/����p��Ut�^춪��@��#����8�?���a��P�?,�q��.����_ԞR�|W�߃�E˷� S�]�H��Ь�Q/ᦜ��o��0ZyzHF��&0З����m!���.�,c��]l�_E!��n����At=,�*�6���y�z��k�z�}*�������q&��,�NW�:j58���g�9�^O ^;�U���2&�{�PgΟ����x�駑N�ǰaQ�|��m\�w��n��w~�J�.XD~��v��!��Kr��,��ӕY�z�&Bn/I���S�@*%����Y�y@����.�~?¡4Ig�2~Q��׋��	L�L!�׏z��wn����5������A4=s ��8��G�K��"��v�,^"�hgg`G�lL�Aܣ�L����ۚ��Ǝ�C^/����I�iX�<�+=���;T���$\F3��: H�kʭ!�h��;�����)���_}�UE�����/E�'���G�0�C�H���n� t�[{=�n��P��~�ŝ�c����6M�2��vw���'�������v5�ΟGr$5�ԣ����h@��X���6a���
�~YTe�(,�M����*���%�F�;|�(����;_B���n_,&�\�(������g�R͟+p"F(hc3��F����*�Ho���F��~p"��VD(�8'&�ި>���ܘ����y��fڛ����l��h�jyD>U�ӝ�9��*I��V����ò&���"\���ȵSv�iN>���b>Sl�����&�Fd�A�6N؉]vv��v^�u5�'�ƩOM�mZ�3OS�}��=���05��XL<���aË�|�h�}� ˍ�R�ʖ-�ʜ�u5��2K{�v"�i2#���?�)����X���.b�}������ϼ���+��w��^}���ҿ���pb�QCl0+�f��F��Ԯ��Ѷ)O��"���{�W+_]�����5F/H�B� �C8���Fa+<�lU�Q+�L8&�(%�6�6��LË�TV�":(ED����#4�Q���p�X[Z���"v�WѮ��*���6qa�4�"A.���VB��T��bn�|�*i�����$v�U���ѥu~��B�}A�<$y#��
�m� ����B	�e]�v����֒�41s���o0�[.Zt�#@��� ���x�3���C��P�A�F�^jT�oVq{��ݺ���%lR�ͦ��@�������@�6Ƅ��2��Tq?�N��D�
arhON�`0�A6�.т�u�.��tV���⢊-�R��ӟSNE8�E�����a�iS��1����b-�*� 'N��ɓ'q��1[�e��|X�6%�b`�v%;��<"�Uj���M�*Jn�޸��Ak��x�I*c{\���Ȥ�}�y��bdܐ�2�s��;pJ>��3h��y{���"�`_�&h��^{MF4<����2�_ZYV^�{ ��&��Zm1}yh� 3)H�����h!	,r���)e��^a_"?�KX����i�a��d�<%C���1���:�..i��vhrz���pg''�3g�	�ʿ�05�/�u�jNf)=�R����_vLb8M��<̋�z��[0���8�-�#f��j�T����l3�t�ӎ�W6;�6��zlm�%�4��-	�ѕ����P�c�bB���㖠��y�;�W5z�<*r�������122�喜M�;s�KLa�+F����Up��(�z�@�|�Z�Ab���(��pRN���LCÁj`�f�0>>�T"���aC��5b��4�Uz��YO��p"D�y�(���mxE�#/��'��D�Ȧ112�ϊ�yw,�}p%��R��}��Y	0^�H̨�
��g��)�3Z���ohE ��kt�L�Y�)�>鄽��d߿?5z��~��7>�"�g7�yjn{�_][����&�})�Ը�4�T��(&�R�#��!��8� �rY�u��:5w$���R�@u��N�L�tW;�
w�Pb�K�������m"�H��Ŕ�J[ʾx�4"^���a�����V���~+�g�b�o���_��Mm!��$��k�H��jqOW�ۏ��v�s���T��Mƕ��C"[,B8�)8�ˇͭ��_���*ַ��_��+cڸä�,�pOŹNRW�!�4�7�u=�%���G�/���sHg3��(a@��{ɮ����yܺ���WK(2��Z���T�왉��X�����g�}�C��ZM��829�c��L�@���Uln�iO�&$�I+���ܼ�cN }}A���k����a`�K- Q|�ooaqs�;ۚ�I$�!��S�e:?=9�״KwB�]�K9��)4A��hl��?y��<hTj�����&m����.�b��<h�;Ib��l2O�;PK�9'�h2�h<!��P�w���J��v��R������b{��-�o���+R�"�蕕%��X���R���܊(��(?�vr
 C��j�.r����ƹ�%�b�񇃸sKkk��+��4#0U�I�������#)O����եe�'g���z�w&�ܪ�ܢ|��h���kg���2�[=�v4!�m��%n�!�f��͘k`UN��g$��&a�jQE׎V���"�a`�c#C�{�Zk����m=�%��l�o�P(�~��jBFX�Et���UP�n�{fju��Pe?��U|�"�����2��XSS�7�a���=�ys�ʵ��ʺ���r��[ϿM�li��3+�e��
��)�p�ц��|r+�!���V���Џ<�ɩq$bчtA�JS�i\XX�@�N����i�����l�m$E����3�"l�c�$�L���>erA/��.�V9O�����O�#�'�;5�6b���xv
��lH6%�ȥ"��p��p�yk�����������V>�"�Vn����g7W���[B�
8Hp�� �ª�����*T�+��!�_ y���<4��t<"i���#�T��zQ���{�:��y�06�p����XF���@,�G����E��P����c��ټ��#e�J>���7p�㏱�������L�C�^A�YQ�s�V���k�A�=���:�C��좢��.-�zmD�)D�I�NObxlDQv�X ��j�Q]ݯb~a_����K�*�2�:1	J!����_�:w'm4���ͤ�~-�J!�?������p��L>q�l��t1�:�&
�26���za�C�.�����;$�7�}��u}o>��G��h?L��:?;v���l�0OcrhǦ�152��ۃ�7o�NA�sفxAܹKHհع�d�'2�
Ţ
G8�T\�+H]tG��v����M]g�h��8~
�ΜC&�U*���wѪ�PN�#ݚ���Y4E�ٟL������XCN�*�<�zQ� �~���IS���i���Ј��I�V
��y��]ޅy�(&�G%���P�{w�?���C�t�|������ה1��_����V�V���~K���Tkf��x����4RѤ��غ��U��ln��E��v��TV$�щq��B�(��`e	ۻy��`����Y�ү?�E&�Ԯ��L(bCc�\�[�f:��:Cf���#��>z*
��&gD�-c �Lg:�).�bro��}8��c�K,Ԇ����nBT��c6>��x�FBf�94Я	����ϲ��D�8i�*�m�ml���l�)2"\I�������"�L���~��w�^���DW    IDAT��:��ɦ����JA�Z������op0����2`a��]�ݻ��%�cG:;ua�i6���h׫��fKE�^5Iaj�ms��Ƌ@~^�#d@����(��(։��p��AĢD��|fSb�eF*2tn�K�e�axw�d���8f���@����H�Z������8N��y�6���jU��n��"^�c~t�,���ڦQ&�����u��A��jή����4�0S�H��N��C��o���|z��?��S������c�����s�������-aQ��(dp6<���J�����!��N0I�:�MQT��:R 2W{^��m<+�A9�TȜnvt ��P��e>��6�"Q�e�pr� �R��a�	O@�	��q�Z,�����.ܺ���e��X.��nJ�&*���VU�f��B���eWI��X(�DY��6|����76���1���H��S�g0�JE4�Pl尼����:f�ֱ�SB$}�F�X��#	�ŗi�nNB,c��TZ҉*���ظ�fϞ���Au�4��Β�/�Fy�n�ɍ��1O(�ˋ�57�{�KX�\�Va_1'{v��;�'7:?�LU��J�_���DS�#xbb
���-�6%�D�Z� �ߏx_��>Pq��A�MR�,hO^�|���9��#m5��}e��"��6&c���8�)Iz��6"�;�L51�tQnT,�$mq�<83���!i�	�2��4�6ޗ�`Qpl���&.6\��,*9�S1p��}ܺ{�K�2A�����I�N��#c����k�}�B%`������n���W��ʧ]������=ܽ}S��ןLځ�>�c	�����f�9��W��#�/_ӽ�v���H&q��gl�D�g�ɝ.�"l1��~0�X���B> �y�E��;�ƢF�eCξ��G46�
�<�Il�,��H�dM2��D�t��w{���i���H�j�;����1��P���"����btlP	mcc#�ǲa�}#�%�u������=}�����&�H���S�eT-ڷ��.MUn��p
y�V}����DrP��A�E��3�h��h���~�|TD�χ��}���oi�%�M��?'tF��#w(~��B�iT�V����tR�$oc����c2�)K劇�=cbl�N���I>��N�.y�s��lj|��}��8	5�� I����NVN��s��f8E�� �`@�hO9,U �Y��y�5�ȹ(��(G}hD|h}f���/����l3��ღ;)�gm":C� ��:���*R���7G���<7s�w~����?�"���}�Ե��wcu��j� R�ʈ?�Pσ(�H����D��B�o����{٩�+�-�i�p�+Lq��!|�P�w��d8�lZ�%,�P�U�s����1������ax���B�
#F��kU�lnb}cUZԥ�y�VDS�[Z�t@%	Pnt�54�x[-��,��1v��ei�����H6�h&���rz�k�,[)��k�E�Wװ���͕�\ۻ5��ĉ�pYA�a�8
:��'*v�<P���	�k���H�pT��#cc���ఁn�Y=R�-�����5�fF���KM"9�w�2n/.`a��xj�Edcb|:�ёJ�nO&M�	L�`��Q��3�7�e�;*���>�}}�f2�ԣ+�1uʄ��;��h*!/�ͽ<�67�W�(Qk�{8�%(o��ϝ����_PQ�w�&3��pg��JB��b��v�͓��y��1}�����	���I�a�Bx�a(�c�J<�k���h<�X:)B֭{w�Ə��.}�?�T_�&g���TV�G�cc����r���$�b��~ 8���k��5}��܆&��s���^�}��A��|݄��îHI^cp<.A��s�$n�!Ǧ���<0�@4�+7�cuc���:��5I��ćD�ZSnBR$ԛ��s��S΄��@�i�uL:�l_ZE�DDG���C�[�lB��1yr��$�qU;��q��m�'ኑ'9EF�О�59j���E�!_�̦��p��)���(ؠa�U)�da�*���Y��>�'�)�>��cv�I��bu��d���e!��{��!�i���%9	�a	�/T���Ko�s���ȡ����E�0EQ�R����ʕkX][S�3[daۘ�F�u��o��?�X�<�A��z]E�v��9(nRf8^��v�p�a���¹���ɣG&	}�M;X����q�nݹ�B��������$Hj��(iI�-�^[&,D�d�i�1����C019�H*���r�
�v��v��0��^t�����*�v<���xb=+~���%͝p�,+^fy3���l�����<=s����g�>�"��n�������ۻ�K��"B�(�0R�w���Ç�˯�4s�u�S&�;����ŚH$u�e�������3��-_�/�Mzt�lk�;X�m�)��l"b�����0K �P^�B�
c$�9m�q�p����Ϊ����D�X�����/Y�2���Lk�wt��.�#�����cuâ�U�d�'F085��@
��ш��"��_����߼��[w�zoŽ*X����Zh8�� Z��@"���";YG,HB\��a����db�h\���	�T�uM���v˱d�O����{N�SBO� 4�Bܟ���������9��1M(�%-���]��p���!ң�m�Cau�9���蓴�s��[]�NnSל�jfxX;iDLOO
��}�6���S�013-쥭uܜ{��JQ�|�n_�鲷!���ᩳ�����Μ�q7/_<��DЗM� kq��v��̴v��pDS'�Pܹ�ɉ_N�:s�w^��IV��"�oBKX�H�#�K2���2�~�]���{�1'�i誴w�Иd}}�F��*v���$Kq�������:��"�SngKE�����3t��aM�������~Qfl��s�ϝw�L|"/_.��nG�N<���)��oa���n��,�����2 �lr���+��b�!��f������A��î����<�,��.Jt������u�K>�,�^�J�2���H�loz;���q~|��sCr����ԉα�g���CS�T�����cƤ�e�h�B��w��>��MǺ�o˨H��ШDǎW���5E��<~߿}O�ɳ����fX�"���B;>��g�Yg�q�d���ʰΫ���.]�s��5����eַM.�w�"e�(����F�ar,߭-�����Z�RJ~��Nd��#8w�N{R+G�6=3�a�\�|W�_�$,�O;:Uar"s���0ƝFX�o��Id�z�P��������C��7*��Q���F��rЍFȏV����M�3ϰ����0�٬/�(F�(���A��Q���%J4xb�p�mu&���yz����'��~�E��������z~{}��Y���PN#��R�^��Q��)�O���f�#�!�f۸�D�������)E�t |�9��M�;@�TJ���ҶwwP����K��l8�C�I\*T�Qf�B��Ji�ۛX[3f;;�������P!���;f"{�� ��,��.H@�,D,7�3����2���$ID�	R�h�m���ͅU��/cu~QN]�T�hR������v�C�R/� �|+�����4*2 =u8F���(�?�d�W*�պ�_@�w��'���L��$|��Y�8�$�GG�����s?�t�&�s���7�����U��!�$h�-BSANC4@!���0�FK��@2����F2���cgc9�yK���"�����6����|���c�d��081���-5{��&{l�Z2{���'�h��}��}�ݾ�����HS�H�5���A�R�ufjR)@�x\���"k�˲��{�LY���*���Qs���#�<bDd�G0;7�b�އ!_(�Mؖ��ܵ��"2� V�J�#<y����lZE��k��j��~�T
���v���Π�/�*rrlpX�4#>ז��N]#?>��PP,���U,o����l���uM�/��簙߶rc��L���2�-�y`�U��),��dg��
��S���60 K���q�<tpj(��܎��[�o�̺����^�D���"�9��C�q K�ސ���ȶ]�l��WH&����҇F��q��!�<~L�`(`��eXB�/�L�;E�σHEԟ*��;'�L��D!`���H����&w�W�>6`&c�pe�51>��~�p��A�Qt�5�Ih��b��*~���2t�����X_:)B|�*>nc��0������J� ��&V93A�(k���H�p��i<u�4�=fǝ������v�,�|t	�/_�fn�V)0���儌M���-�AR����SG�50:���)����������z%�Y^�-�=T�e�I�y��/'EN0�m`"F�\�\��^�a/<�xU}�ׯ��x�g����t��[�x��7���W��t��3��/H��ƑD����B��A�X�(�`�kX�s�i��I-M02�����5�}�׃D:�=��2�P]fx��"�0䞇�����Э7050��?��B6<�YfZ�fn�ul�sb52�m�<;���F�+i})��ni���3�v��H�1�MbrjSG ;֏P:�6�ը!��wP������5�H��vd#H��	��#��B��qОNͣ�u��j�EX_^���i��Éx#��M�4���%���ɘ5ᛱ�)�;�f&5� ���.o�����i�Zx���\ƍ�Yl��s�P'�C"wBπ����;���s�O�c80<���!����SgЫհ����{wM^m8~�H0z(:aj����S��dE��ەK��hY	+��CX�S��q��I�}A,ߟǝ�ױ��(�eH�p�d\�rm���'K�B�B�M~kK���w��!���Z�y�������p PA��������{�kz����%�p+��.�������� �>uJ6H?z�u\���`����We����V�{��&�p ,�MʔM�(S�����w�:vjrh �"L����.��y��PC�H���O�}�<ʢ�-.bk;�	Z�׫�H֤l��M��SH�z�v�7��̡G��߯�Z�Y���u�8p Ǐ����^���*��dM���el����]��Mi�Qkv�a��.Nv6���)���nOt,�j��O&K�e�����IT
3LOL����x��)��@�4��ŉ�\��1�^�&�s�]S4�mӜ)+���m;ʶ�d���M�3��I`���e?K���>��<�.A�G�8��^z	��B��ƴ9�G|l
H�{��wp��Ui�%ݲ#�8%+F�LЯ�1�1���)U�k��*�}���������я����_ʆ�}'N���:�_ӻ��f������K�%A\\^7ӮMܢ��?���x�^�t�O��%��>F�1r`
�3�(3K���V����>�~��������Gy�ԩk�k��G_�&`S읾]�i��0������^I���@�����y��'^�����ח����NٞdFD�����B���n�Q,kyM��}�\L�`�}d�Z���a���]l�,�d"f�8�,�TZ{7�zyC/�����*\�&�fZS��.�{���]lnn`ys;�]9{�+�1;.u�z��K�:1�a��C�V�6�7h"N�#��ġ�����)��Qj\(nJ�����]�a��V�/csi�bCŗ+g/��ii�	�P�t�#7@�g�����uX!�#q�KG�fCE���>�H���:Vs9�5�H�rk�����V�-��x�����?�C��TL�����(����.ݾ����������n�1�=�k�Mຓ���%c~rz/<����Vq��\�q]�9O�<!V4��E�.dO��Z�_��L�r�}�F���=��Y{��;�����*�BQ�[�c�H�;qi�\^{�3�O�(� ��t��^��CڰUm �~pTf�х-N����@`zK+kx����;響
�c��\��aww.��d
�dF?��'�\�>�Μ9���ڏ_S&Q��گ�Y����;��kܹsK�u�|n�VO�=��I�7�M���i�D�ذ јE��^�����٧D*#����]��M�Xmr�--Fjv��dK:��{���:��7U�IxS�m m���i��̅g00<���erlżu��صp�V�E b�<u�tu�3���C��^��a- �v��?�����K>�ԣ��*$��o w�=�,8q��y�<N�<.� ?e����[X��λrt�^T�5ga$�ɍ���p�|*XAE�2&��Iޙ�U�m�
��5	�����?{�4^|�E���a�7�N��4�]Y�����p��e����s{,��N�V��4��e���0ҍ���|:��,�b�s╆ڋp����������3i�7��T�8�%����%�K&l����6�� ~)����v��4���M����A��(�S�(�z�w�j��Q/��w��C[Kˏ.mOiڡU���x8۞�N����$�F�����2�g
!�Y_��������~��O���O���ks��t-�3�����X��8�� b!�W�y~'gL8���k���o�H}_7�ݞq�O�I�Z�
�,��Y&��ER��!�+EMΜ\P�"��a$����T�6���I�Y�ma}'��ZQ}�V)����ͬ4!��T��)����w�b�4����5=6�c����K �E���.��,��xp��kۨ�VQ�4�������Ӽ�Xk��i�	���h�������A����Y!Xޠ�V��$��ew�����=H\`�s�~�������v�jMZe"$\�b	�{��}��$�eK�2FN�����x��U��wVӮ٤�x�d���R�Dv'�"�<_ޤ���#	�=v'������x睷��G*��?ӥ�%,//c����q�앋�|��&5�|�[���Y6\'t�x��i<��y��z��<�q{�-5b^"1��F�I��d� �p��y��e �sc�{�uݗa�������L	�2���H:b�S�''T�>���~�]�������	��^��5�Nr��!��Y��Pp�y�ǯ��+(W���_�5�������/���+�����f�#*�$f�ll�ޝ;�3&�"&� �F�y��ӡ$�T*�'O�oxP��;s�p~�{��H����
>��`� �jFU��)����m���U6=Q�������O=��{�9;��v�����za{�o������Q7�l�}l�Qm�Ԑ9E�Ϯ&;6�6d�v<lНՁ�wͿ�x3{��b��}q��<��gq���#q����m"ރ�9���{x��7���L�r]ڻ�K]�_�S���f:�7)ir\�%;Hs^g�@�q���!C}0I�/|ҵ�T ��z� Þ�f�.]�ի���sV`��R�z@֠fv������yV+����y`17�H�G(�������_�2fL#��)���&��4"^�y ���G��_T���D4�o����DR�ڸl�9Q+ͶBV�De��Gl$����|��"�hú�6�=������8Y;�f���4U�\�d�J���eݞ�Mt�k�_��*/��Н�c�����?�ċ���/�vi��n
��V�X#�,Cq�[��.�l-�EM*�hX{|��th
�k�q�X�L�Ӎ�	��;K}>�����I#5��ha_������Y�����P��v~��]�K�+WɈ):�#�gx������d�Y��.�;m$�>�%��dЗ�`x �h��&*͚L@�
�6rhr<��N�����C�7@��A��D�זg3	���X6,����Ѽ�\�� ��F�XE�RC�Q�{`����=^�
%
n���Xk�F�$#3�=D#x�#ڣ�U����j"��#=2��Ǎ���3��:^�D1��IBW�XBf�¸C'a�:<�	]�$?��V2�œ�p��qd�1��ӟ�o��,�� ��H:E;;NǱhO;"F/�ue�    IDAT��ł�Q6-�m���(HJ~^8��	<{�F���q�2�������'y��C<�Ȃ%�ǝc:���e������?����ð�q����W�u���i�R��UM$��\l$}A�mn��vB�!��&�ɖڜ9sJ��/��Y!z��_~�e��������kW>RAv�}dӞ;sV�.'ҹ�����S���3 �u�R�~�"d������"�]�uU�\[��m��W)?�TH��Ra���L� +@ԿXTnc�v�Zt7j(j�2��Y�1���g�K��EC�	��G��ljrm4��ߝō+W����BW,T�f#���;#K4!毶{����b�WӦ͐v4���2�Ф�����>�O�ۨ�Rc�OgoJ�������
�7��n�\IL4�K'5�p�~�/�pɖ�a�kՆ�_�s|�l����E�����'��ً���ŋH�b&/���N�ٻ�i(�K*ro���]�a�05�.5��bg$Uz��xhmI��f�!����mw�����5�Ĥ)�� 	�Q���ֽ�Sѽz�*���ܻ{u��L��=s��#�����C0��4_~>����<f��&ыPrw�ݪc�[G��B�<�^�~���$�@�I"��"SE�q�"�ms]:�
R����*�Vr���f���'���g_�ċ����_�:{�_��+��2}��U�3� �t#i��ϡv����܇�|E��,�BQ�:�8aq�R����[�來��:��r*��dJD+2�<�;� c�AX�3u����/a����¤$Z2��!�DL�@�W��_��hR�0��W���~/R� R����7���q�[E��J%`w���pB�^�|���N��d;5�5J�1�D�.�3�h�eI<!���^۹=llnc7_��4���fM0t�2���������a�PF�Vq���h�l-7�OB%��������Y�ehj���C������be{[��*	ETO�z�#�l�љ8�ahtx�dBv�^ʅ��M�H�<rs����^�G�/c��Jjj����Çu/l�T���.��ܻ�]���Ϝ×^z3cc�~�c��?RQ '���9�����Ζy��r�>� �����;ylon	�q܁Bf�1�hJֿL���`F����2�߼%"
<B���2���
�ff�v�RO�>��������?ԡ�?��W�*f1�o}���}�:6��up����RnE�isc�[����l��O;v�b���+��ˈ�G�:�C�2=�?���2�p,!�<��cnU K�h�R�;��\]��:�k��W��H�D�C����_�/��sl.�>pZ���UFm^���_��z�bY(�i�K��	�m�${�2;a���5�����2F)���\(A��Sm<Ĺ�x��������������gے���\�v�������.���&���cճHڡ"u[z=2��G�H�i�M|mNlnY"�Q��g/�>��!G)c�i$Z#��S�/_����ks����VD?���ai70�4�����R�)|~}�m�av�r*T4���R:533��~�+������vȊ�T)��_�w61��>���=����eO�j*�Yo�r���P����gB�hT�f8��+B��3��^Ef���*�ݠO;�1���+��G5���9&l0�_�o���� ]��Wc��B2��g(���������������/�����^����ܘ�h,���B�;�j�F[��eպz�Ʉ�u#�B2���׻Vn�O&j�>6ZG{��F�3�G����_:��j�t[x\�d,\�"Hl{+���M��՛h�(�w�M�C���4�p��|�(W��,�
�3���7��<o�v�r4�E�:-1���rB����� �ޒl���Yl�Q��!\�����M}٬�GjG3��8��R&hn#���e,-�aeu��:]�ܦ���$<D�$�`Ba�BA��qk��b�Z$4M�-�VDN���NX�_�K�4�I�?#�<�w.�"��s�D)�!��!�=�!�{�������Т���~.�����	���������4����d���:x��������"c�� 1��S���=~�l�>}�"~�K_������;��_W��d�Ӑ�E�ؓO����I@��80=-�!"�c���$��L�NΔ��n:���"L�I�|n�#�$iq'LM�۷m�˃���&
6�V)�$�ϟ�W~�<󌒯Hv�$�XG~>_��������7�3nߺ���EA�z^!5q,�;��(����Z�OS7�ϲ�#���A$���C"M�fL#C=�#^�m*�X�Q#2��Y7�p7{BB�Ѹ��|�hO�j�T�-o�dJ�N|�3�x��TL�x6f�v�0�����q������X_�B��t��	Lb��+$E�y1�l�t��k�a���b�y���@~5g���U��vf5ߋS�ںq�����4���M�,}z��^a��39;�f�3�%6l4�q�ht�0��=��t���<��y\�pAnTlM�50��q]���dO.},āω�t�$����`�]��v��4+r����ux���5��D�����"�˿��*�1�]XT{Ҙ˜�6����ˆ|����Ѓ��"���G����v�A5�d���)U�e���υB��=4E�jҦ2T!fnr��u��c��&�s���r����"�g�7r_:��lwټSQ��*#�D�>+2?�?��'.��W_s�������)J��빫��w�������^���4bfl��8�]/b]7z<���"�C��B�Y��aR���M�_�}q_�g���/q�ף-dL�^)c{u^�K�2���S]�	C5h�A?�k�=��T�j��Pj�P#�C8�ٹ�@ah�n����o��BAB$��T��(+�G�X���uX�I������aAdCDk�2RN��c��v��B�(�&���K�/��^��@��ɟMG���=X��{����`�fQx�K.�-��S:k14��A��M�W�6.Th�FV��'�^`l{�D�u��T��,�D�n^�:}h�,~&�,Q�1L�R6�1�x�3�/�������l�܈[��<D6xX2ʐ��(�?f$��h4������$���<�iP඄����l�.^�/}��'�7o����lo������&�g�"���q�����BN�t��ye��줟�H�;�fk���o�UT}g��VX����ʪ�r9�qb��I�S	k�o�L�LZ$+�9!��.`|b?|�5a^���: ���o�Ƶ+XZZ���EM��a��D�.s����i1H~4"X:����HO�̈%M�3�09���� ��E��	h�� �A�o�D���ʚ��<]��𚦀�<<8�?q����p���&�������bH�kkaׯ\Ǜ?y+����/����Ҥ�(����C[���:Eٰؑ��c��a����AF"t��܋��3�\D��4��P��xX��� �������?�ll�t�Z��y3oX�]���4"��t�<$N���� �ɏ�����xY�Y��
��V�f�=-'O�}�I8E�7ƻE`���	�X(��������B8,��|�),l|��Xғ�u�m��mG��GM��=�����cV��D�s�b\��OĬ/|�8tx��>��춈���������᭷���ڦ�e��+��s�1�К�C4�nd���7�/te�����"oi��k�����d�x�H ݐ_C� ,�����N3щDU������{�+R�zv�t�����jMx*M������#�}23�=j>�����U�+���׷���B��HĒ802��pB�t��P#��"��Y���#�Mj{��=A�H�+��&��)�@�{r#H��f�2�0� �~s�h��ww��<��"c�Z]�s8W�]��(�*��F�u��\�[d��i,��5����I�C{8ހ�
:�:z���8=��)�A�pY��Ё��E��{���"}e�����#=8��0%1��A��Qk3% {;�o�h/���"*�с��'B0�D(�p��
`���/S�s
$�O�%�(�����mQ�	I����a���ᾄ<�irk�v+�w��N�}9�:>u��^��d��s�ZWv3� 	+ݮn��XX�����nX�c}̮M7��}�5p
�*��;@����v��>�/��ұ(���x�W�|%����|~[/5�J�QJMD:WM����J�$�J䌤�'�UT[g��kX�5Ή��C~�{�s�6���4a�u�2�^����0¡�+����Դ��s��Q�ko�.&)��|�+������˿�6�]���C�}���u��C &)��(Ж����~�%��H���5�M�9�1�G��y��~-./�Gf)?c;��#��w��Q�sG�������1�JFmr��g�ן�S�N������'��$�TÿU�s��z�*~�ڏ�������cA�co�zES8�c7h�^���񽳸�>Ra;X����"O���=0=3��|�Ӹx�i5
z�9�׃����0;aa;W�E���#����#�t�i6h��=���'�p�f�Yِ��,��l�����?��tF�afP������WG_�|E+��~$�C$,��/�L^�x�H�c��GGu�:�=�p(�4D.f�����|}�x���q��A9��M��7]�<z}~p	?}�4X4rH�7�g�#i��W����PQ&JC�7&��W���;a��p��*��xH��,�<#6��=[zx�������b��<%~�����P����吐��5Pp�$���V���ֳ�3��&�����;a~��~�������t�RL2]b�o���Rio��[:4�T�V��h�RQ�O���~ƅ�7�7h�j��ڕ12�N���̯t�Q��5s$y�ۂ�t��Z���~^�(c�^U1�6��%�U�����̂d,u�^K���!�}C� و7x�MC���\���;����=���G�>��/�ofX���l�!dƆ�@���}qx|�t�'�Fy�����/�c��"�Vs���W$Y��|!�I)DRicI�����u����C�c�'�3��M���4�~&d��������JÐ��~7\A}C��#�^���͌�&ev*����Y�vp7�}g7lL h9G�)�P7�Zj'�}�U��W�L�9a�]�CȐ��Tr�w�)�vqWo��.�XA���������֏�W���(z\5ЩHNDѨ���)M��ZM�I>���"��H� �i<����e^�q����@[M^�߯u�T	[J�TLb��������{��r�����h������/����w��||�#��wp��#�y�� �!�_<8Ȭ�{�;)j�i��k����a�M��L�+��_�*�j�$[�%[�˵�C� !��'@!f:�&���6�IH�TL���Nf�$�L � �i @(������V�7ɖdm�������9���J����y�>O��Ⱥ�������=�yρ��0�@�ӻw3�x�	y��cr��%���u�Ra�	Y�}�ml3+a����x*	+J��l�a���[n�W�������
NY�a/Q��2m��E�/��U��_? +:G$D%b�>H���^q��������ܠ�hV����zt�I�w@:$��T��ǈ���9rZ"�G%��O|B����ת�R#;xB]7$�������oT�H� ׋�����%^[-3hAi�햛r]@�#s�.�^?���=��I��׾&�?q��S��f����Y�G��Alxp����p=XH
�~2z�x�+�D�V�����ˡ����cc�Tu�k����ۑf�.{T�q��d~a��H� ��A��o튅j�Z6Ќ��u��E&�8�X�;u�'/�@�8C}�#���]e�uOz�a�*�N}�-E��4m���S����l#1%�2b�����������zރ���w��p�?W����l���BI����7��0�A�o��*|d52oKaA �@%�����,�0�,<h9b�U���QV�&��&K�K�R2B��k������A]�&ҁ�Z]��Q��-)�j&�q	�@gYY*���8������\3�aH/�Pp;��$җ�J��Ȁ��^���f$�bFzK����,�R��MCb�'N:��mJe�"�s+2?� W/]�k��Ҭ�x���+N�W2�^q{�-�{��Q$ϣ<%`��1;�E�fr�|��!�� �(�2�pn��l6x8c�	�d-)����V�;WVe�Yc����j+�*�
$.���'�w-7����c)�|1��4��q!��Js���1���0�J�����+��l3�-VKB��j�?��W�%p�+��?�9q�鴄^��P�0�GI"�ӻ��S�Ƶ��O� �Z�G�J'��d�) �f�v��ՙ@ҽAx
� ��B���D�*�\����)H.\�@a�[o����Xр�V��^�:�mq`~������=Ġ;�c�<�u$��@H�~C������`%��5YV�U%m%+T����<� ����� M��`�羑���yp�L�DS@ ,W8�nv� �]��B��z����w}����d�Q�"�+bV����������/�>�k'�#n�@>@�i�-T�ZB� qW�[��G�AK��y`a�vO�oaa٨4��f���S^��C�}r�E�`���� b��sK\G���5*Ciέ�o9V{�Ng��9G��u����5�K��W,i�#8$kUV޵j����]�\��u`䀴
�Z��kw��ӧ��ѣ���Ӽ�b��Y��j�_1 mT�`u�@H����s��XW�S�U1�^�Ѫ�8>��Yב�u��	Ȗq�5ʆ`�:��D������#I���k�sި�UX@�\��Q8��mޓ�z��H��~GfV��ނd��.��6�hX��� �Rtf�(��I�R��p-H��`1���{1^h��K����nyס���|ރ���G�Փ�����Z�T��Q�(0��lQ���HוF�������q�2އ�z��e�΅!�i�;�*O96��D�'�t]�%���hT$naD������dq�m�����~$62��^���ȸ����ŗ���#�c ��R�P���A8HI&�[�"�cKy�I_1#�c2��lٹU������@pDTH++�t.^����ȕ+�R�0 S��E)a`0(�R�8�^	@���-�
w)K	�οa��lp��Joi@J��	"hCD��nK�ӖryUY��?H$�_�������ڊ\[[�J�)&�)�fr���&fI�`A���V�5pA#�	T5)R� �B@�K8��諩Q5��n=�_�?L�`�Z <vV����+�~���W� �Q�����!�Zo���dc�@��ò��6n��Y/^e`��\�PT��
�L�V�'�C�A��		{�L��%���Q��X��Ͼz�*��/}1gi�VFE� �p�0�t@�����ʃ>@q �o$�Lt��AP�X
K�w��S'T)xfx@� ��v�Y���ߒG�8!Ϝ?��D��!�!zrt����%��
��Z�E��tZ>�=�� Ÿ�y���N�~�!ʇ�*��7<�:���z�Iy�cr�cO��p�C%��Jr]w ��Q�\1�dbj���QaS"�ܐV�z�N���+5Y����I����n����%�_�0h�kՔr�Bb��������E�<T���7�4��V4m A��D+\#GB "܇x�9���5�x���'�F�(C&�Ң�Yc#���Ũ$a�'?�NWN�=�9��'� �	p4�0�@����f/#yo���3k3�CСXԹ��t.>u����{��w�)7߲_&'��D�㓉��*@}miQ~�ay��#�\���9�\��7�>㚍	W#b�@#��6��;J    IDAT���m[�ot�:觯\��ZY�R�G���)d���c�c����p�ԕV�)H^�J�B�;�CWLx�BN�e·���zWoٲ�?���7OL(�g�zNp�o���9s��*�j}�Y�?5-�vF�n�@Ŭ��!�-��a�_���V3	��s�d������t�@�E;�xP��t�ff*�X��
GQ�g����~S����D^G�x:m����yenAj`G�:��-����ӫFK�Xڀ�;�۬�������a1ef��D��q�c$�?kJ�Rl�g�c�둩�mr����"=�"C�j�&@�,/-1�._���k�2��$���4;���-`��K��+�B����t"��V�}�ѕ66�a����pm1�/�f�LNy�"�F/����ģV�J&�G����͒�Z4��U���a��l�.L���-�1�&�ꂖ~���;D��Z�?f��*}n�G^���]�9nD�1_exO6&]Δ���9s�6�)�0�T�W���_�jټiD�����׿�e��
 �% �u�ّ�C�,z�b�F��⽩Ċ}
-����A$:���~qʜ�c��6��yM�z��P�YtF�z'��!�~�w��~资����X02�*A㗿�ey�駨[��Z�����~�Ǎ�������#���}j�3ۏ�8.��x��8~6	9hÀp�D6���b/e+�s[F�@��B_�y�,����k�嵯y��-��@b��!����O3?t�C��R�L�(��l�����U��)��*���G��ZF��a(�1�[�$2��h��d�z��}$@톓��S��xݗ���s���:����*{�	`Z:e�R
��W뎤+"oJN�����2Y�+�o�.�#��p�q:$١��^�'�b0Q:��o}KN�>���|���K6�^��t�J��z��Nd����)5C$��,�2RȫF�!�F<��n;x��yQ��h�m�~��	��IH�¤�4�HcE.T$: i7��]��Мf�לB�[�t7:,�k�ryyAf�KC����z�M��?F� ��@��]#nJ)Q�"Iʂ�=���4I�~N���R�Lt���~�����jpY��z=� ��{?��S/�A�^�E_n��n:�aBפqd��Ut���xCgf��e��N3j��) Nv�	�Q���.�e�� s�$�>4��`���$����:�4R�����5�30����$�ۧ�_�&A�����識]�LU,uln_�+���%f��`H��X��Hш$'E)0�b����عU6m��/*��E'���ۻt���]�"��5�WZRE��s�W�B���Z±a��Vo�
�%���C=��]�^��o 5X\L�w�7i���v$�p���Cq�oErT�\���[5i������!	.4b�,f�<x��6N: ������%ͬh���"ц��u"TڇUU0�� 5g+�L�ʘ�R$��m�P��Ҙ�y�+erb�<����_�O��Y����r�RJ<�Ԫ�!��Q�橤��W���Pc�����7�����+�hQ�� V�$������NB��z��{� �讻H`�ܺM��巾%����~5���H�ʕYN�����D�(�,
�x���'��.T;�|��U#a}2�i�j_8�!+����*��ǽAr�ML[���9Ͼm�f�q G�'\ʳ��*����z�+�5��A��X6;��	q�B�����c��o��MY]�J��_z9�d"8�����W��:4U�c%ՓO��p��d`
�>�J �
����z@F�	����(�1�TD�O���JAx��Qt<3+(pqNX��ྥU.Зjm�p,*;$´r�ȴ��Q%�9�2�ρ�0{�X�a$�%2�wNNqL	Hu�i��T�H|z�MP��  �
j���հ4��iO��d�Zf��F�]Z*�u��"F=�DV&4�0�P�yٿou�'�mU��P�3� �!�g'��Z�L��`�ox$Z�gfe�� ���%�*w��#�7<�3kf��\X�� ���=҈|�]E��9�XP�VS�!�9��O�|�^�3$ꠝ��k�y �0Ȧ�Ȕa���7:�ǷN���7���<�����l�[�o|��������+7�=88���#��A�Ili�-QKs�X��ʖ�1.*��\����U%����۫Rx���l���Y>,:B� MaF�ݒ�+�Ҭ��,�de ��h�~W�pE��*�Wgeu~�Tr!�C�GF����
�֨KymM� ��[쩂,�4T��7��Ċ�#�&}h1�ԗ�K��0�
�U�<F�2�4T�ɉ�2�}�l�<*�����#�	���̌\xZ���i��tR�$=#����ߴ��,�U��� �knv8�>1��l�!���Eu�]�Vu�{9�z	��σ3��@,J��+�%��Q�Z�-!�Kͨ%Z���F�58x�!8R^U�q�E=�V��URdW�WXat�bW�
�#�!�恦*a����p G"Y�|A^v�]r��C�zZ.�{Z�����'�<!��$� ֚f���Ce�7������x���S��.� Z�^���9f�g0��Lb�_W�A�E?+e���*3d��'�@�:x�~�'G�|�	B�Wfg���[�����e1 'j{>�lUҀ{��@G�V�U�Ið�l����*M9��+- �o=p?�p:������g�
-�B�+d�4 ;��ț@%�D��^~?Hx`�c��Uw?Y���3�#$A]���*����Y~�ޯ�Z�.�b�K��@��&���h��X%b0i������,S���cֆ;+��*hsFݐ��ۨ}�o�.VTx�\)�ȩc�Y���g��*�S޺NV%����| �Mq��Wdye��� �MV���n�d%�^ɻ.�)��s;����,S���X��R.������f�t�l`ps���"<���8jr�.�R��t&ڎ�qc��$hs���uHP�=�l��;dzǤl�:�m�g�������������E��Ş�꥓<-�0�j�&��4>A���\����
�xH�'W�Krf������c5��MI�b��J-K�l�ܧ8�P<h�o�d�Q�'i���CA8F.�{F��r�ض_��&v�?۰�W�I�������3�/��r�^��XvN��M���\��b֦|����t��	><d@W�H�yG����U��|8F�0`̮�U������9��S��M�ٵA�puaAVg.Jcu�F����
}dh��DV��>�"T�]��Q��p����=��p�����ood��3@��D���H��H1��@_����@I2Yh��҅D�ߖz��B��J���qhI6�'��+��
E	����H*-��)7�� d�"\Qr�Lq�C�#G�� #F����#t�Ƹ�jY�^���+}�}$n�`�w3Ʃ��CC{��@+'Y"+�	z��,��
�X>�`��B�$1\��p}�7����Z�k��B��H&0*�W*��J�0�����!(`9�[o��_rHn?xu�1G{����47�BZ��N�~ ��<�s����q)A�L^-��n�(T,Ӵ�ş���H�#�Ԃ��POB%��t0��Bf.���)����³�g�!4��dH�u,s
C i�zux6�/G�p/(r�U%3��|$z��7��������9G� �+5<+-����oߺ�����N0C�9y3��y���8��}/y����Ioo��/�g���ZBU��w��%9����}]ʕ�Z��#�;n�R$Jr�v���29+&?<�q��ύ�� Ǒ Cy��b;&?�a�zT�\��� cX�u|��/Pޔ*o);zC%��>�}��EY*UeyɖI�Z��&��E^#� }}��,B�3�yշ޾u��J�����H{�QB��'OS���Y��u^d�U�W3��5��x&at/�~TR��z|�^O5ң�
�@ ���˖�����m[&������!�l�����/\�!�{g?ʔsVʉ4���y��� ���D�?�g@v`82�iX�^[fW婙���Hio��8��LX�VMF�:�փ.n�`
�%�������$�ML�A7��́-;~�m�S��o��#��K�~g��(��PF7���歲�X�f�%$RLZ١7�c�vj�"KE�Cc8?��$*�&���H�&�""{uaaN.\|F��:�80b!�ѭ�e�3đlBVY�M��< ���UY�vM�����pEǲ(h���>�ApR���M�}���E0wu� !M���<67�([���*���ltۄ 1��H$�g@�l������o͏�
��V[�����M%��͊ED�M@�j~U- h���W} *cs�}U� ���Ijs�C�*&'�a��E���A��Kg��Y ?+���`��(��T�}^�'�����bI�Gt�cG���s'���"� �WJU|OV��{ހ]!�D޿��ɫ��n��ҩ7����2;s�kOU�*��X�v�y
A��7�c~S�Nu�M�%*1 �UY��hEHM����z��i�>���� Z�
&��S������y�}��S�<M�2ƙ���P4����K6?�/�#��1*6��5d����K�Z�;"�R\�:M� Y�v����?������$�z$�$�V1��j�E&�6��90E�x�K�C6QJc`�V��*�����|�|�[��j�Α;��W�\�뜕��� 2���ϐ< ���8%֡(U�><�p�����b5���3==��A�"-�:�ˀ �����5��c����G�D�T�Fr�� ~hp6Wϑ��@B�� �vT_8CcV�@�rY�[�,��6q$(O��4�R�#؟9���}�i�2;'v.#\��sY��Q��ӦQ
�v��#�:SZ�k+��pO�҄=���2�
���ϋyٳsZv��� ��ʢ��\�W�r��S��y�?�{���_T���'D�4i��W2��+���&�(�BeU./���ks�E[���>?���r`{Մ��
n^��D�y�ga|���>� ��-����.$���vzl�z��=��� Ŭ���/]~�b��kD�̝��mhT�՚8^$v�g�x|`H��e��������ua�7*SL��Y
g�Y;}hV* .�K�Z��k�+c�7���(I�%�JY�^�>Ӑm�r�A0W!H��H�RU�	�+L�|��3�rռbu��@�"6= f�8@�{M �����2\�H>c����z]�p�MV��%��H ��!�Q�LOI;+u?��zKV������Rmu��=H"^�׋5:ל�8�X�O�s�
�U)��Sz�
�I\�A�MB�g�������Re�9n�,�|tN٢i%��Q9^�n�}#�V�.�cիTN(�NqyPZ�e��;C��u�=���c6,����eS�_u���W�R��%�P5�P'!;�ٲ�G��h\��|fz�D-5��z�i5�$1���ͬ*a���5S�
1*)� ��)H4�d����������]"�f��׎~���[�n�t�8\�[d�Hv GS�LLP����ʗ�C͜f �i<��B�ZW�xv���1��ejw1��Tp� mt� ��qn��x죣r
`�ޕf��*3���=r���r��e��1�ύf��5iV�v��<��r���Z�EV���J2��,�<܃�.j�Z���h5�0	���	+b���H��9"�	fn�	tƱej�$+�];�$��-������p�v��~����ߥ7�JL5c]��q��<aX�c�z!�s?c�~˚������nE�_w�`^� �^!�1#u�]��������+�j �'[��X�XHP�Nk&A��,`B�!X�7�K�0�	ԅ�� $���$���~���d�OMNR ���XJ��i�y���䙳�R�����Q6$�tqR^� �*�K��P1;J����[���̵y���(�ՊDYE��ș�=z1SZSBL亁+^�5�{$�)MR�1��k,�E�-�S������7���yL>i����/��4�k�z���vd��&��3�H�N(/ <=���P���0������Q�q�i���Ք�å�	| d���j�n4+k+���$�{�O�%Ԋ�5)D�L��ȶR����d�D�����t��т5~h�����/����a�&|``�r.� �4H"q�{
x��,<@�k��� � ���Q*I�W ��`P沜��D��h�M�,��!�Z	"�qM2[�jӢ`$����tS�>��i��"5_p��V�:��^U	�=;"3Tګi�H�UX�Q 	{gZ��b8:�g��wR�)�lNt�D���� t�5L�Ϡ���	FT����h�`�#CW��J���>TZ��a��3�W���ԏ>�k��LG	�lp�I�͔�(��]kaS��ٔN[ap���*�T���;�{<r��Iq�;�g8t�~aj萣ʁ!:������0�H�� ���W��Sg؛��+G�T�UUZu�TJsʃ}X(�1	�NaD.to��o�c�Ki_h,"��f�����E"�����$�vL��9bP0����*uv1���������Ėq�DI��1���;{iV}��<��q�a�=[$/u�e�������+�	�Z@��H�
P�z��c%
�@?ۆ^���~�`��t`���=-=`�C���J��?�A�ر�i,���d�,F�"؊�*�Cc����A�\��O��E5R��7�<���^�c��аLm�*w�~�l۬��|&��I��� ��~��I9s�izCc����:#�sj)�B��Ң(e)cM��y�jU<F�0I��P�jئN�K�Sn9x��ܱ�#}��l���钠��#����S2�{W.��F������PgT"K*�hE�2>���6hQ`���nJ&48c���q�ƸF���H�ғ�)�	Xx.L��S�-�#��K�x�Н��!EӁPUes��Ϧz����������|��O]����z��5��0�+�v �0��b?��3��)�,p�i�B%�DBe��A��#���XB#��K����e��c� ��O��I&e���d_���CPoJ{�*^�M�mT8��`��NJ��K���AHh�*�A0�q�!ӄ
��$$p� �̊�p*e��,X�h����� /9��V`[҅~j�-kݎTڰ��
ܨ�H  �Ǩ��5��(9�@���P��"ԕ$gr53�8�2z�Ȁ!��*e�^Pݚ"m;�L6k�&D�%X�8|�W��D\�����-���p��*T��rA�F�����fP��I����{`��D\?L0(�	�h����,��Ƿ�In޳O�MM�-���UT���8�������A��!�s�'|E�Qp�� �{�,aq-F�lZ_�o
�C;b/�q�
��
��h^mY�K�|�DhB�N@J��6Ǟ����9j�O�sc掃�k?`�sz�|��lC�.��A��`��<�WJ�1����<�d$5��쬌o�}�v+�ɪ�d�ZY�V�Nq�RO��z�ٿk���m����X!�z��K���G�z�C�Q;��b��u��Ġ��Mb��^�PGá��t�b
C�j�������{�0�z�A9x`��z{h��A� �bq����1���Y��W���k�2��Y(H6���,./&��8����d�����s�/���w� �ͩ��;�b�>:iM0$b�Ԕ��%�VSN>yV=���=��4�'�H��h(�>�_�����|�p�N�� �kù��q G3������9j3����q��r� QQ��la� �D�s�'��0F����۔0�3K�����K*�A�c�@�V7���ז�6iJB��T���>��6�"f���Q�SO{����3	ׁ��1@D:jH��;=f��L�]?�����m �y��|3����/x�tb���,uZ�V�m�y��������&��$��: 6�Y�    IDAT�x�YY[2�<+�RQ��#�=f��w�X=�}gݾYjey���2��H���+�c,�<�KS���d���bחb7�Ֆ�ِ~�AH"R,j8ZYk�ey�%�NH��+`=�������/23-��IOĨА�����%F7����+�C����Ƒ,�k��Z�5D0ZFDMS*�p;��4ɀ8�������d\E*B_�R�jS�`�nH4VaZGc@h�+�4�ܕ���@�-<�R"f�� �Tg�i��yKX�E��7�)�٦� ~@��B-A����2�P�hM���sڑ�3��"�(���W��X������&(�4�TAϊ٩Ƭ 7#ت�[�|����t`M�R�փ.�HT��е~p�B�8�*)����j���o�?c_,w�?,��a�H�	��R0!�p2���N���g�!�ĥY�+ L&���V|*��/����� r���=�)�L�;��/�X�J�%;�z򐮄���@?Ek ����/�j�)Gff��c�?!{T�eJ��z���p�`�#i �ι�n�ɋ�gfٿ�duЩ^&��ɨ���)�p��.���[��n��c1XXKvb�Ѵ)���O�W��5��M%��;U�:�l�d����H��ΕV]�ol���'�5�R�@U:��}%�z�LMMI��H4NoE̲�Y�'?��3��1(C����+[$����Y�,�S���z�^��w�����S� m\���^^ i���̴4G�I�	�HB�|v~A���0qa�Y�.IT���\�����5���F]9��-O�q$�`]cv-Z���վHQ-a��H�ya���������4��c״'��nl��b�r��nA���=�� �|}�A=�����]��E��Y��m6+#�z�!/�ER�c)�"�ZK
�3π�Č�'����X�=P�*Wm�]A�8�8cR%�ڲ�mȕ��,����: ����ϰdߦq�Y�Bۗb�+n�+YT���ݎ4;M�)T�k�TY�%`���P=0�].Lm�%ʨ��ze��F�(�=��6!#E� �V$dH�fH���Z-)C>�ِ�v��m8� Nr�W��n��+�� "�n]CE�*��F2�kx�kЂ��Db{��k�E@W���<HVOQ��P1X��[��
��nDQ±��¬�e�K� ��Y��J�沯�f�UN��*��A8(���s�>2vm��|�H�4�X^7���66T��խ�f��S(�C��}� �^��
׼~p�kf�)�]9H�#R�<(��m&Q���~�B 8A4�e���P49����i���"h�$4T>��� �d��P��(���4p#p�׍�VA,f/>g�2�Wb�q�p���3��pɰХ��[o����"���IL�/5����ȥ˳�У��7xH�VY�!1����ډ(esӃ�3�Z\CW,�5#Y�+u��Z���X��ic���r���:8�'p���{b��ܜ�:}���h��_ H�B�04���m.${ZZ���p�p_��3�Ԭ�le��Q�A� s�/���ܾUJ�>1�6��;�:�8��e9��Sr�Ҍb�#xQ�D��������� �G�ք�I`�@P��p�P�R&���N�d��I�D�z�h��L �_�Td�PK�я�gT�'��ty�(�z�d3L� �@����8��I�
X�V9��RM�8L��s|�0�b[]�0=1L�4ͮi�m˲�b�P�P�X���-�l��+q�����җ>k���s�Y��m���_���ً���r�+��(�n�a���ё)�0�R�H����? ��N��h�	[��A�؇h4��XBd3=y��h(p�Q�K��+	9��=�-��#�n�.S��b�k�Ԛ��z�L�jK�U��ZY�W���>s�F%-�7%�Q&χ���6�U��G�s:��C7�E��1p��G/k` �J���4dcQ�2��&GV�
ʷb	S)\i�,N�E\5j�7� ����_�NK��X�M��I?)�[M{LX�j3�t_n�|�A'y*5����d�����Bt��u��^_(i�4�QL���ՙ'�:��_ϼكՕ5�A'��ԇ'��8:9"&.��ŧ���V�^>��4� ��@�V�J�T)H!�H����)�͘�U-�`i��<��{���*���L/�}),�3vݍ	/�NM���[W����lثׁ��e���<���}�����������~�t��8��Ĩ���
y��ѾADH`c�lR��G���-�һ^$�6�S�TB<'�Q�0d22{eN�=v\x�QYXU�%���5A�����p*'4����p(B0��w �1���A8m��s��{Ӿ���>)��Rꅢ�����-� ]�|EI��,St#5�7�Ɂ@�S�;E7�r`R�EE(�B+Uh���+�<)Z�u��r�YxXk�~�Ͳ}\��額u$//�	��\����/1S���H&��K!b�mi囎�qAK���RZ=r�(gl��ЪS-:L���:���;��z�Kh;\ge/U+����V`�W���g�&[)��q.y�q�8w�(�3+��)Ɩ� ᇑ�E�4lӎaĞiY]C�iX׵�f,]1��'k�i�MC���D,߲�Xvm��$��ˊ�@`�v���(���r6�y�+T�x���{��W>�oO\��׺�BՈ�>��<GE0��g��c����P�/q�K�gdǩ�N��j�P �f��
��1&�s�a�Rn7d�Q�7/z1A�+n7��lQn�>)�=}bU��6Z��)�&�W���܌�\���ZEÒR��/ȫQ),b0��z�lw��~�+u��A��<t�A������ ���r���@60'2u�a��q8b�(��=	]��ޯ�\�1�&&���?���\�V��m���d;e�*e&�� �E�͝Zu���=�9:�di�x}�A�Vl�TY��5����蓫5�wZ)�}��n���!�8\? �j([}��������t��)EI���Bz<�@Nkj^ξ��G)4Mt��v�+���y����H�E���dH���[_9���$+8�lx����?µ������­©�nj^O]k]����P^:��,#a �I�וt�`h����PB���J��ID�)$�轻�� ������$��.��Ӕ7�:>�9\��0�)�X,����S�屓��X�၍�`mw�6��7��D�4�����ڱ�� ��	!	��ϲ��>1���#��y��Q	�A�_�x�V��O�תf�J� Q &!�ӧl��t�12��z���T�1���i`KH@��o�s��d`��I8+Q�32�/^�"/^��/#�B�6)���$)���iR��ϴ
f�V����-""��2)e�}�f*fad	�LڒQք1���ʪ,,��}��Wl�rs��f�q���ܕEQ�q'�����ZEu��۶a��ql���g'��EQ+q��i���FbZk�Dkb��m7L��l���ذ�ؑ$r�$��,�;#��[�l�E�o��9�_����Փ���b��[�}�0�˲�d������Ȁ�J10$$���`¡��`L #�������*�
H�!M�+�c�o�[������n�Z�m�Ɔ��3�Y�J��R�b��])���eY����ʒ�kel���<\>��H3H��8�@$T�0o����6lF?־^�� ~��A��(*���!h�\B72Q��V�?�8 �B��iy4n��C���=y`Ce�1)Vz
�S0�
�)�"5(@��Щ��s�dA��K�!+e�����C/���W�ER@OE�H�3�4�z@�I��F�L�u+=eU�)���҃)�M�i]�]��1{=+F�Q��H��t?��^i��U�f������!l��CK�aT<����@��\'f��d��	piO����(:�hZ����AO__g*�������������[��� �&�!n��AW���8��]�R�E')�*��F�AXM��C%E�`����#qѐ0�֫$�7'�7����v�<2J(:�� <?8�Z,�Z�&O]�$�N���!��� ��B�q�/�����U	�gC�M��H�H��a��eA�{�n�(�1�i���}}
�`F�n8��o�%X�6��5����G��{W�P��I�C^c
���{�pו�6��g��8��<�`�Ax��V���g�2`r�<�.]�� �2{u���c��#qg�2��0��i��i��a����0�8���$1����U�#K(
8o��bA�2��|!�X(fAh#�j�+��}py �tuy�J�CA�gF���b��6�B0���$Y��h6��k��sF!��|N(���׶o'ۏ�Q�$ΗJ�J�������\�ޘ��Y��_����r�ʅ?^���5	���:8M����ۋ$%R��t.1$�I-��2�t)�eW�� �z���}#a/�h4�fG\ϔldI^�><${G�eK�G���U�|iV.>#�W�H�w�����߯���+C��u�VVde�"�F�f�p\"�be؋-�Uo��6G�u�tpDi�R�"����6�>�]���I�O���y0�����INM���@+��S�H5J��gu�T��l�ཱ�LE�XGUw)��h(��*��ϑ=a�B!� ��=Ĵ���;z��`��4��s�K\����v��%%1�>�V)K�֫2�5A(�P���ji�z[	c`���@���}��6�%`�þU���f�J��:Q�J:`T���J�9�E�M!8��WC�@nF*(s��Y@&Ԥ0K�{�d�c]�P�H&��u/�_�(�d;g��������F��X�*'3K?3]��t�RY��{��d�!~���J��� 	��l�^ed��O&�F�!����fl&��#�,!�L��tIx�Qa$°��h�^o�mF%�N�ـ��ϊ�_ʍ��	�h��l��@x�w��KC�u�'��a>6�v�I������ |��.�U�f��9M(6G�`b��Q�xa5�(�DQDn۱I��5�j9�a��i�͐�Ү�!��XI����z�PL�6��As��$�IL��@p=aF.�?�_/����$��İ�b#�l{�rl7�� �-�q۶�cYa�~ 
SA�4-�F,Y�!Q�$θ���q\�0�n�S�8����-�o���~ ��BA"m�u��V��$a��&K++�R��g�'{��>�Y�w���5'k�f7��}��ް��Fލ��*�{��9y��W}o�m&�8��-jX�{�93�I�+�X��Q�X$b�a�AfA��� G2"�=��x ^�uo�'����A�Qd��$$}�q"c}%�=6.���2 ÂZU.?yZ:�I:-)�s���_�z�����do�Κ�\mб#¡n9$����4D����A�W��^�ГZ�)�����U��i��6��ɾp���W�U�@ "�z~�}��0��a걉
ZWE hQ�P)��T�
��J׉6�ᜒqt$D浖gCU�yE�<tc�R�* �]�k��q���x����������u���LBT*c��1�������z`O+bt��윣6�����U�5��@������6>O�����8l�����*g-?Ib�%RAW1/��0�"h�Z��*tB�� g��c�\���]�8���?�|���6֯W��~�^�1��{O�nM�K+�t�x��i^�4�%;A�P5�˪[�z*b���L�lz��q��F�����,���d���>B�[�a��H\X�I��qBy�!�Οg%\i�9��`.�H TC�!+5qH��F�>�� L(_W��b�z;�Q�3��g3�0*a|�V��G�r�7X����Sg�[��}���A�t��3s(��>4C3��0�G�_��p���Nd۱�Nl�Nb��$2�v�,��7,k�4���#�&��؎�M�8c$Q.�Ɍ���o����^$8���$�0Ƶ�=u�}����=�V.t:�hxx�Yq�0�ضm�[(7�QǶ�|���F!������g[�e��iők�nd�A`Ʈk؆���Y�k�<3�ǵ&6�~d��]�nj�6�dikc�͆R�Z�փ�J���K�~�K��Ե������)��K��'g�d-�lC܂��F�`��$� ����Xp)�#K��i�`���I�d�+YXj>VhV x�����d�����۾�>�JI�ٮ�{d2t���ui/-I�ۮ##���
��QH7���2�C�W�Rm�ă|!�T�nNJ��J��K�h4�E�}_@�Уi7<}��.�$���HhanM�:` l��!��1 �Z��9��7V\�`��W����(�� �g�)���د� �����&
!���� 6��CXgL"
 �f�	�W��@��ΐ���:L|=��}t ��}�+eUE�0o
w�
j���_'g�s�N��i���d�(��J5�#k�I�(�-����:�7�<A�W'i%�����(�^��N+̍�iʦƟ�
Z����n�@%�"�� C��	��f���*ɹل��b�>�����j��N7F r�؟	�a��a�I!�3����@T�f�P�4"��8��(�#�l��@n qB	^2�ˊ*�@�cC���N��iu[k��_�-�)I�Cɹno)_�7\�����m�9�B��p��"��~�iy��R㌫)�a���1�u306Ϋ���+����9���I�J��!Fմ�eY�r�v��RO���-c�ݻw��P�:��ksb�pty��:w�O����B߅��?p\����ÇI�8r�@{���o��w�0�;���q3�<ǈ�m���m|�w����;��B[:��}"�j�g�^=u�����<���9R{��������ã�}?}`���2�m{	�|�T.�ݐ��ީ֚�����WZ��~�#)����{�?� �����g?�������r�d��=��R��(�&C�$%�(L&:Ծ嬟r���jV/
���#�Jb���bu���{,[
`Cz��x�5�<�'�2 �G�"�5[^]�P��>Q�W�lN
��
-��{Q���Zi��(R�b�~56:-�:I�"檮H3W8=�1P� ��ԕJ
��?�aZ��h8�a92}m��5�b�	�+`�t�Uy:���Y!��3��(0�!=ͲNGuTE{��<=����l��(��t>sc KG�p�i��tvr�^��F�����u�x;�d�T�KdԪ��\��p�DqlYVdF�A�q�Fkr�?���l4�E^��>�|����o�fbFlFb�f�D��8�L3f�db�u#�2#ׅ����@5,P�݌�0�?�</�汉�o[60�$�f�.b�q�	L�B��yA7J?���:�vXO���d,ò�l�qr��i;�'DV�@(�mB+2���nl�~DÈ�$��8�-�N�c*��#�.*K#ä��FM��z�O,+,t�q��/��@M���;��~a���?�oz7�,��
�U��2�ku9yF�=vB�����ja5��*^Ek2�}> �b��W��R]KZ�i\�S'gC?��Ī��c�0
��7��a���oڽ{����#��C�� ���ry�k���O>�;����?r��ܫ_����C?q�]w�{��d	�J襧I�M1�Zp�[>�ē�;y�����/�u#��k_��ޭSC��gz������� @�	׃ ��	�yҺ~�Z�|pq~�7��г�����F��s
����l��T�?���<xd��Rjc)�O 6L(�vzVQ�")d3�u���1l���!_͢��Vߣ
���y5���`�%f�#��%��K2��+#�W���P���[�g� ���+�|���g������v�ZoH���  �79��##���@��JqE��`�"<���ɍ02�۴Z[g��9Q�}U�6m��k
s�S�B@ F�r���.]`g�$�کt3�B���@�I)�D��p�}ɺ�@�@�Ң!<��E�*0��[    IDAT�G%���b�fP�R	z�6�ㄭ'T�`�n|Eq�a���0�"?Toj�)b�h&��Ab$�e��i��m�!�`��{!P��D�a�Q�N��n5ڡv�(�"?l�nP*�z�8v� ������Z�U_nךK��[��^a�ŠrF�*iA N�Ȋ#H�Ȋ+�]�1���&�c��0I";�c��e&��QB����^'LZF�v�0��4�r�'�s��-�&#+#�B��1559rd����>N���;t�P�����5���N�t�=���h��B!/�vG._����|@.���r����7�(B��� 	���#�	�����hEQ�D������y��x��G�2��#���|�7Ƕl��]��i��}���џ� TR� �1�����Ǟx����W��#G���E�߇����s�y���7�v����ΝS����Y僘E��Nb!�an~n���ӿ��Z�ώ~��j�>ϯ׿��=�v�|�];����pH'$Eq��VE�:;��W��?�8��>��/=ϗ�]��S��O�s��"�_�v��(��T@<�i������Ԕ ֻ{I�95g�#$�*@���Y�xp�d��y3f@ajb]��1�����I�����Q;AW,TǍ�4kU�9���*�K���ĖC(�Ro	�`�C٥5/$ hܹ�t�:+��c@��R�EP�D�<}�Z�h������eUդ��C��!�_j���< ��.�a�v̶���H�0L E�����d�|>oerY�qh� :��$�M�NȁL�������f�^��~��~P1��9�����u3�i0!���U=�	P�8��0P�u:�4L��P�-�5���՜�gE�����j�ڝ���h�	
�.C�8F,}��Ac	p�3~�N̸�b��a��[��fԣ�LT��8t�؉3q��b7
�����n�f�I�ٌg��dde�l���ˋ?��Dg�	垿3U�]�ɿ�.��ٟ��ݻs���NO�R6���6����љ�yy�أ���Krm��X溕���>LV���S���V3ʭ*���$��y�:��='z��ѣ���t��wۛ6�izώ_ݿ�-����7��&��8�`\��n~nq��S'���j�72�y�[���7�r��عsr��1�'�h��--ז�Ν{�=�f�Ф��{���?ݳ}���w���3c�Fa��@� b+���w)/+յ�̮,�ڧ?�����ھ��s
��@�O�f�ȋ^�TF��X�bf�$�DAd����ߧ�=��Z$�A7Є-l�m�RG@��P�9E�A����-Lь���k�q��mw �w'��d|�_��[�]��o�9��E�2V�V��~I����JjYP�Egws���B#�c(�qǉ���0�01�@��|? ��e��u,+�ضoZv`���A��i��i����� ��@��P~�q�*��iZ��8�l�0\˵m׵|ov���r���y'���;�2-È��"\��q�~�����N�_	�Cq?0����f�~^&�8��fb�mbҾ�I;��Ј��ءaU�����������v�b>oD���^���wu�2++�\.�l�t���ğ�*0�G�>�����om�������;�`��}����Hb d�( A��h���Uy���ev~�Z�ڬ�a'I2�1��hy��w��2���=yB F������֑�����G�~[q����?�c�ԯؿ�GFȎnCq/T�&�0*�k�K�Μ�͑���s�=Ǽ�ׇ��?����}2�}r'*a�0!����n�,./-�=w�߬��4e?�&"���n�����?�yt~aU	+8��n�V��?_^l��8��d���O��7v�=�L'�9b怑�Q��q���V;q��Q^<f�B�!��"�C}�c0����%v8��J���6 t�~�L�^��t;�V��w��$�H{�|q����knݷg�h	J^����$ݶ��$�.��`@S�#Q��5�	6[��6�Ql��3������l۩5��z��Vkt;+�c4��Œ�)v-1�GI=
��$�r���q�%��Vێٶ�@R'vP�Y ҤmY��yqӶ��HP�6r�8�hĮ�&�2�1�[N����M>�@D�==�`�?~<�Ç��WV���9�;<l�{� 0а+v"���Sv��H-�����?bi��O_�����-o��=;����NnU�"L�`�ĩX���:/�=~�:wm��f�uΰ��(���p�e���Y��%A�� �<j3��v��ۭO�ڝO���/}���Ѽ�o�mjr�?���[Fǆh9	�cX"����k�dy��|�ܙ{��G��F�7��-/޻��&&6�U�{;��Q	�_[X9}��{����|��u���,�G4?>��v����[7�;��Ƹ������ ��x~�������>��>�������s%��?�=_��]�z5�K�l�� p� �jݮ��zq�����4�q"C�:ɣ+]�+���u"�ۅ�Zd8�cDQdt"�:�ԍ��;����`S�"��:ݮ�8�U(�m~��7�����@_l�f�:�	6�ﱑ	64��AU�)Wk��v����r#��ӞE�,�-'�3�X�J��n��u��h4�NOO��y����Z�����{�|�;��Ç`�����[���l��c(a�sV��R�+�Kr��مٹ�O���o&��o&���$z�H2���8��>��/�_�:7����ڝ��z��9��~�s�?G·{��G�4�s��o�t��w�oanwથ�-�9C�\Y�����|#����÷��3���ͣ{��+v���UU&��gΜ�_��/��7�g��׾632:���;'���։,f�Q��d���;^P�T>��^��#:�1�_�q���x��n�s��|�`!'�Q�%&��N[Z�Mie���jˍv�b��<��}+:�DV��v�Q��{�B:��/�v��^�7�>|�Ўɭ|��7�l��F����臲��*�N��p�����{-��-y�%�����7��4l,m[\U��9n�0����V�h����/}���Aw�7��c['����}�96>l@���GP�
C���m�W��S�N��������{�U��7���7��֩��eb|/�h�ѤNT��!��_[X;{��=Q���"fa�j��ݿ�cz��S۶0�f9��:��l�9o4[�ry����g��?���X;�,o��]{o�7[��߾i�o��Y�c\�լ�߳5��4����p��v��y'�(��逸*��|�?ˇ{�M_�ߣw�o=|h���?9�w����!�-��GC�WM��Պ<���sK��R�~��8fd��-�zu�u�2Ms�v�dQ���n��Vo�m�[�
���k>�l%�l�w޳w��it���)p�3� g�r��j����3�����9r�y������w����m�&�MLLh8Z)�9�\�#TK��s��}��s���g?��0����~���~���aǎ��Ln��e�4{��4�sɳV�E�����:��G����x��՟�OG�ހ�{�ύ~lxp��\�����u����2���z~qu�t��|�.2��bL~�~���;�z�����lzz�O޴��Ѐ䳮֧V؅�I��Ғ<��#�\�t�=���Q���ձ�C�i�K�d�m�%�2]S,t�a.x��������=��>����������ʦM�x��G�����ë\�t�<u��3�μ�ß�̷%z�S?�Ç����mٹsj�h�U&�:�ߴ��C$0�������Qs� ���[��Ν��~g���~h�ÀBM�(��C��j����gf~��G?z��>}/���A��o{�������=I�H.�*�ˍf����4^��KK��k�^�o���ڵ�Oطl�_r��(�+3)����~��c=u��wO��g�~�H|��a�S�n�'ŀ�e%Ih؆&Q\�h!̚W����s�O�T�������������`��?���Z)W�O�<��3O_��ȑ#@�n��mo{ۋ�m��Ў��{FF�HF���f�C?��R��/^������w}�c[�!'"oy�[������75�m ���ѥ�s*�j(��Z5^\\�����#/��|^x���w��; ?�S�����5�'�<�otS�d]a�+� ��f"R�T�~��ٳ������/߈[H�ҥ�~��}��i�p_��W�	�J.µZ�s�̙?�4;�������&?<�mb��Ѐ������X�-�^��h���|��ճ���|���B��O����?�}	tU�����������.����(� ��Q�Y\gZeAQ������eDQdHI'�wUw���n>�o�
���[��$�Jݷ�[�S���h�dJ�fM���h�ز�����4
�#zUu��=��~�����ۺ�F����*��.�@}D H��sZ�;�ݹ�
�=H�`¼} 	C�/ D���ۿ�z��ǖ�|c=)���~C۵m7��A����؞�":n}��f,W������~����޽{_԰Q�כ5i�
H؞�n{�`W��c��z������OҾ�}��۴i��͚6·9�x����lx�c@µ�ڷ�.M�Ѥ�l�E�"@@�}�ݗ�ݺ���k��\�9�r�����7�c�m�_~�s�#�_}�R�����޶mΙҰa����\[���u��4d\Ւ?��������+'>�~��-

�4mڴ]AA&�'�q�A�0�(���UTT�_���l�}�hڴ�ԦM 	� [�K���A�5�@�X�C�������I�m]\�z�uqW�M��b������g��{����� �ˉ�Fc��L�+�.���~���;w�[�Ҋ�� �{�w���Y6h $lK �*oЃ�c�j��w�=?���/���ٳg����U�7��A�,���=��L�5�д�G��~�Сq$_���ׯ��xF�F�=^WF4�2	�I���fF��*+�Ö,�����$\o���8E��A�O�>͚�j>��λ��(��@� .�ׁΒ�_~���]ߎ��h�R���sG�sZ��BQq��99���	)*6	��	��}����.~e�R���ѣIAA����E.((���pbp�<N8`�zEE����c/^LL ����WXX8�Q��B�ǉI�r�0�'�)��'>>ZQ=rɒ�ߒ¯.�CI�.�
��"�_����^Բy�gο�>� '�tK�2WV>�C�0ڽ��������ٳ�B
���{�Ժe˹E�����eO$a�7�ط�?�8t��y�'e[�>}�y��7��
�����ghce:�C0�
�����tE��U�~h�Ćax�=���S6(*�A'X��<�
kI�g�I&S[����_xa3)���:����P�(���~���7�|�EjX� ��L�=�ʴL������B���~��-_<Kj<䐁ojР��7l$��L#�۴=�X<��Vݺw��a�g����v<����z� ?��u�A�Ԗo�Gb��c�V��w`I9r�}�sR^^^>�k��Z Z��l�Jx�4wUW���5k�ۤ��P���Bm��#0h� �ϓ;���֠� �0L��"��P���O�c{�7#�Oy��牌�1t�u���4,l$���3��`�7�	UU�>|�r���7�ڮ1cƜ�p8V���ր����X^��j�( 	G�q=�����4i1O��G�:��pL�x]��B`�Դ�i�Ў	g$k�#�k-���X׹>�����{���<��ߕ�g=}�Y͆�qY�>����U�<�U�:;x���`d¬Y�@���w���z5� ��]q�S��*��!MM�����Ǫ��|�I"=�p�O<����$�v��EB�W�1�2���I8�В�Pxu\�F?��c�r�O>9��,I3�Ng��%�.8��S)he��&��4-�X���mq�zxP���No�"�{"���e�&����
Y�0�e����C��$*��?O~��_��N�=�����-��������'Q�D��ސaY��D55�﫪k�=����:O=�T;�g�t(Jk a<�Ĳ庱�!c�z��F*�����1�>�(1��	&�&�����!��9�9>NHԨ ,�	I�,~�ǣ�<x�`ȩ�%�z����)�����������=��e��吅IH&f��-��WhG�Ϋ��ybƌqVO���:]��9��?@u4x冩#+*OS�T��_QQ���?���]�ƤI����FQ�s��!�� P��Y��_UUWEc��dIxz�����KJ�b��-L�IM�hc"��a�'��j��̤��dס$|�H��(�ӆ��)���<�$���f-{v4�L�{�.��UVW'�ˏ.JT{t��iDԀ&O��tJ��99�K=�M�@f1����L�B��Б�Oܾ}��7�xč��1mڴV@���VQd��RHׁ�lO��v.�3TU}3�&G�5�XNxҤg��,�Pq)��'�	�C^��� �����c$Ѹ�Y��	���$\O7��6E��D`���JE�����܎�$H���ͨUUU�W�/9V~����*Q�S��ɓ����jn��J��k�p:��K��탖�`(r��f�۷�YREc�&�j�9Л�|!����4�:6�}�$g�[sP��N(��C��<y��k8�Iq:��$��v�H���</�i��4}l2�z§����)��o@`֬ٝx�� 7���R��0�'�v۞�����#K����Hx	�\�����*'?�8	�킗�8a(��"�X�CG��ݫM�5k4���g�}������N�%�,�X$|<��pR&a��E��G��!�F������t�ԙ� �yMR���%����|k�X�q��0�#�i=�iu�)�LO�P(��瞛{1ˡ��\Oh��x�	@��	 b8j�k�C��,)��ԩ�߸�I��T����P^��|rs}�HpkMFf�aָ��9�(�?9v�X"��S�6�Ei��(���b�����h�eRL��x��Ph��ѣw�ԍ���&N�xÊoȲ�Wo�|��E�ݮd�φ~L7��9�\<b�"�g��O�%h8��CJ/H��s�,:״ҫ�s=�Bu�,��`ǴL��|b��Ƭ(/5�=��#��ŝ���%�������<p���xL�@D"r��za<~�?v,����3g6��uI�Dc�M�m]�d�IX�4�5z������O?=��c_Wd�B(��3�f� 䫧�d��ìJ�ƤX̵����.��%���v��K�/@`޼e�S[�s�.�A�I�'*�)Lr�C�R(FG++_�	E��3&@��'N��Pd��^��kN��x��c��$��j�XU`�cՏ���	�fM��0ť��ۑl�$�i{�'�0��@cs"�
E�<����H�k�'On����,^�G�fH^�cO8�F�aT�>!�,�$Lj��:� E !�dɒ�dJ_��^��ٞ���0��7��XUVV�E�<���D�N���"�e_���n�p4xtY��,	�a"���<x5�{�ᇉ�ʧM�V���%�t�[���|��h�M��1 aUU�F"�q�G� 6�k��\)Iq� &�G�"dvXi�z2�����"Gӏ� E�"@��K�$��b�anv:;g�Na�<a �D\E�TT�7n\%	ǌS�u9���ͽ���0��4��h�O�4��X�����0R�����Ҟ�x���6	�H�mOX����a���I��&o�*�|{�<`{t�te�#ܲ{��z��0�G���tb�'��A�P2,XP�PxϠТE<pX���$��E��h�;G��HxԨQ�>�{B^n�}yy9<Tg�<�� �d2i�<�:8<d�?�P��������s� Q�Z	�
������Ǎ�৤��S���L�N$��T/ a��"-�pJ7ƻ��*:1���u(� B	ƚ    IDAThٲerJ7�#ɂZ��S2!�)`yC  ����5��`RC'ƍ�v+��rss�5hP �W$�s�!�>UU5�Uլ
��C}��;�?37bŞ�X�(�b6ך���2-J@v��m��ՇG���#��'>ۀA����ތ��p��ǒ�^q�3�kZ�XYޣ$Lj��:� E����lqq��,kM�9��q%Ӳ�V����A������p\�o���$�5j�R\�?�������Q�����±�q\| Z�R�p���ꚱS�L!R�=�?�1c#Y�'I��:��A�����/��5M�.O<����!��1iҤ�`��y�� �pV���RD;8��1�����S%R;DסP(/~�&�Jm{uXT]ۯ4#5t�0����%�tȀHIw�1t�tw�Ѓ ݥ��04�p��{���������[����|�LKp�C���e10�+a��Pi��KB��)C�%8T�23X�՗�ˠ<z|,bP�Ϭs��C�M��ni�?w����_�^Ex�S9�c�H���ʌ��}�&����[/��h����6s�涘��1}۸�AiC�CX AA˄�|V"o*ʰ�3�J�?�6��)}m�l���8�$�������W��Ep�݄��L�cn�E�F��ږ��S����Z�Jց��u|�ȸb_�@�	�,�����]��븩{�+��b҆�E�|�.����Ƃ��>�����2��������I�,�q3AļsE�eM�3���yő���C�c�4��I׭��t��w'�pƚ�y�fz�6�"���oJ�Ԩ眝�G��.mq�P�l<&'��ɸ��y����K��#����k|�A����M��:��|��M��{7�{x�ߣ}-��kc)�J���2���&�L�=�x�29�
%��Ւ�ѓO^K%�I8�w�;D�_a�W^X���4�a�߰��N������;S�u�&m��iP�����h�U�>H�-&^>��f$"��o���z�K ��5/�U{����[����.�s�پ&�d�!C���B�#��^'��K�d��bi�Q2�����Zd�ú-�
���X�)��v��l�uP���B|?��m!�U�x�?�y����K=� ����?S���<^��(�$g3�p����X����
�f��NL�P>�c��ri/�B��y$ԺJ&�� �Z)�H����!��2&�ӆ�Ѝ"7������"F����(�pYAYl�:ĳ|�~��5���/����,{>J�]�R�ԡu��,4W��llߛ�9r$�@�2M�a��;⾴�~��+��F�ڷ��^�T�aY"�x���'�;ϸ�������2�Xtgn�I�*o��K:|o�f��`���	��>��uA+�^p�:N��flk˩��D/�9w�'_9E�o!7�j	̭��bS�8B��ZR`R�O9�I�ޥ�i�|�Cm�g�/��2��cI�BT��E]2� �
�.����u�����	���P�
�#�3 A�����hO�TqX��ƹ`��ۭ��(�<�!+c�04M�����E�>�8:M2��TH5���p⊖9�L��={��h\<���/��o�U�Ԡ��lK�w����-����(/!�n������f���s��w��Y
3�O�hL9��z�e.��l:�bh\60N	�}����	Ș*5�RNJ8qI櫓�v��dQ��4���ɂ�EE}�jR�͊]Ɔ�ĩ�����$��������/���V"��iW�}}��ǁ@�vO� �Lo��7}��U8�=��ޟ�C�Ⱥ�Y�.�h�ŧ{Oǥ��/:v=����>/�.�2����B�k�O51��å΀����\\;�P�M~���A�-Țn�	�q��,��v�B*A��;�JCF�r/=��.�Yś� 4Э	>��f'��˂<�t���l%2����G�;³Ѳ]�8�tn������Ǳ���}zJ��θӖK��I��b�f���&���1�N#E4��C�ۺ��IBQC:k�)���b
О����e���Hq�'��Fo���%���A)�"0�X� a?Nr���,�	;wtz%�U�����_�Xr�>��|6�hKhm�6|����)�� �/h��~�+2�q�Zs�]��O�H%Ԭ�Ȕ`��!���Rd[��T����������5���d0�4�i��fK�������aK�S[�VB�������1Swd��`���[">�T�������s����
�ɒ�W��g�L�e"�^� Z��'�Q�O�uSe}%͚��p��Ȁ�N��k��&��ߞ=�.�RT��t��/��մ,�ˡ火�(Vi�UK�=Q�ɐ�ETI�gL��Ao@½Ǆ��%)))E����&W:�q�o(QZ���R�H�:�$�㶮���d+�3(pч�<T�Ǘ^�E %�`�I��P���%��4���Ms5P:ʊ���E�+�LQ'C���jW�0���a�8a�-Y�7�H�n��.�m��و=_�'/{�	S`�+���`�1���VuD�ˢu�?a %�o~�0�-�T@ԡ��+G�Q6�Q�i��5���ž쪦�X��������Aܘ��f���b^��9h��n���U��_�ig�y�����.دi�`c��}d�u�{Zj)�u�#�xoME�p��g/�]�j��X3�Z]� K؉�'_�<y��{?�J����9!����_7���s��7��V�q�����hOnj�3a2��M�G�)Vה/ȶ/ZP/,���.b�_��w�׳�h�$����&�	|1�M�L�v�W=��BJ+�J�����dG�nA���ŧס�* �4,�"�W*E��N��gGky�L���jKt ������|~���F�ܘ��O��s4��{0?�Z�(l@� 	�&��M�Z*d��w�y�R��tF�}�W�������6�����e�[������.��\u>����X�֯�yI]�aV3�z�I?F�$}�"��R5�a܆��.�ԊA��e�'�l��;e�fu*j���x*df�n�K�Y�r�I����=�)�NB9""l��(�?gS"�A��Վ��#r���d�ǂ	��4�>���T�.���T\����}�y���&�
���[r`H���]�������w��J�!2���PS��Ȭ
�m�i���NK��ǎ�클e�ڒ\���z�}�K����(xu������CpF��7�gIr�͡bPm;�N9�0�/X�)�q{x��x?�cNĿ���ݹ�Ta�����VN����}��{�/*�~��?��7�0�c.�w��|,&�� ������MzX�S>���T�<��:;� 7����rX��%�A�U������p��:;�4dA��m˔���+5�s.�����Y^�>%�aW�I`S�'Z�����3q������ӏS0�=QJ�
!2a��;�y�-�~��L��o�����9��F�l�#�'h�k�J�A�G�W�5�׺l��^QdPl�U}�聥MN�g���"ǋ_S˷?R��x5?t�\0^'���;[�<o���������朥�W�J�����Ҩ�Ϙ�x�V��5N��k ��AƳ��J��l(�)��j�8�|D>� |s,Z�)bgzs�]�&ȣ�2�}�� os��Q���ݦ�����e$R��#�r�ߡ���^��{����+��	�$`g%盝 ����8M杫���_]��6T��3�E�W,��G}��j����LGƀ�J-NE	YN�3�>oϗǳx>QT+�qn#v�V�`�/�Yc]�v�
�0���MM@'��eČ4��^*hy�M�n�М�C����|j#�?��Ë"C�G���BL�L��"w��y��ñf�<�y�%�ɶb!:		-�p�]8�u���	0/�M�V�����G���b�1�o3���܏��	z^Ї'�+�D�f�������l��i tQl[<>�_� 1x�F��~��6�<�y�9�5M馋'�%�0��a����P��¬�V�� ;�5�}���]�W�Vv�q!������9;�F��ҽu�����
�x쫿	�����<Ol.��|kT2� ª�R���m�ܣ-��]���� 
�###�!���]bY��k!�1n��H�)m��'�kʉζ�x�Et�`F��w��� 
ٵ���-�Bgk�ޚ�v_����#}�`O��~�j*_X���U{��6�2w�ޚr����M,��|��'����:��toW��!���w#S�93+d�����R7?�_���������?�o��  j`u���<<n��ex���@���u+�j��w}�C�l7�{ȝ"tp���N�y��|��qh��Xz��3~J����S�_���ӣ��gO.5�a��moæ���긑d����,9ɾ���5����FY!:�t�bGܓ���n_�05Rd��GN�Э�Q�li8�WP��G$�]1 ?��#M(���l�_[؟��=VT��zE�g���9C<z	��������w�]���.xH�:ۇ(0��H��|N"|����nS����*��El&q	X�7��?�2��\.��$.�f���]@X��{c�/xh�!�2p5�ht^��iE�5`؁%��';�B\ T�1�^�3a{
ܒT���[_��P�������~x���V�1D� �w'X�h�� jM<.�֖Zj�t���-?kX��$O�ŸtK�L���E;��v���U'J+����3"�o�}��<��h��4�bR��h��SW�<\�����Jdޘ�\aFV��չ#"��i=�oR����/�����ya����sc=��}F�?���4_1�����d
w@#���xP�k�ep{���R{��V>���g9�;�.xPw�s��E�a�)w��r�kfcK�/��d�?z���<�� ��B)!"���O�M�P@1� ���j�I���TT�y�	Ɯ����_��3�b>��~�;K�WN
USS{��3�=��H�%����4zzL�&�,�S)f���R##�WQ�J�C��B��*4%�Ƈ 3�l��X�f�o�	^>'�w�����1�Q0G���ת��eQ/�m9���sT�P�*�2��:0�嘓9$�V��;Ttv��h&���K���*�\��m���M� �*Q�ؚ��f��ϥ(�S�1�b����G�ht���3_@�]贮Φ�V�"E�P�C_�5�+��h����uS����T^^{�¨�sێ�5N�����I�ns��rĽ�N��׍��0��+c$e���S���'(���|��� m�zh?���XZ���=X�@2��B�A5?���j%�T!oN���4ʊ��yt8�ȝ���-����m��.����U������8�C�6�3�#�p��
���X�s��^P��.�ꝺ�j���&'�j�tg��K:�PH3�B��*$�,S��MQ��	O�:~�s���;��Z5���-��T�ms\��*�X�Y���7�\*���Z�o�Н���U��<�kPR��UI(]C���L�o�YM�+X%SG;�ĹUz��h��x�����^��W�$K����
qJ�Ž����YY��W�r�����ۚ�X7ښX��e$�HՄ��T`!}���L��͞���j�E}�rYF_UƄ3��x�|8ӑ>;�=C����sC�I����5�
�����W����9�ҫ��;���Xd��i�d	�b�%Sϐ���W|�+'5��enw�7\ST���F�	[��b��DW������|�`��*��u�2)L�^���Ŷ�!r�	5��XZ4ɌGW)XU�w{�Eߌ��i�hs�%�)B�D�&J��J@$�_�}Qnv̑[QW���~��͢���Ή ���ѺpmNů�6�>�oU �P��?�����|=�45=�x5`�����-{��oN�i�}�c���\�`o�h���^\�0���~��Ųۀ[dE�k0�
>�+\Ʒ`}�',C�<[�v�ؾ�[�F�K� 0n�ο �y2�T��4�"q�l=]Sq\�9dƀF���w&�!��%}9v �Ʊپ�`SZOg�1�ȡFo�x�}fzZ�QE�-#���'#��g����Y��d���~U{Av�[IU����� ���V���y���d��i�N|\���Nu������u���ȑ����s�^������a.P8!�&˗8�� T��0�ҶrL<\�w�'�:F��dtb2�q�<+�c��P���3ӱT��Zt�b��K3n\ y��vX�͑�`L��kL{c%!i��T<Fq�kwd�3��{i��[5���W�#EP,�蚞����9��`�G��U�\ d��I�ıj0��q%�[6WX����N�Bȇ�4������׼ѓ��+U��1�g������j?6��+ߘ�O��N��f�2�`��e����T�,��;,_�x4�Q7
;�		��"k~��
^xwr7��D��v��;S����.f*TXC�@�&�r��^C|,�:q��y�����S�����flL4T�L�B4���0��Hn=�.x:㊣�f1,��N^��Цh2�c:\T9�P
�qLs��IRZ�)�~:ZG�~��G������^O+�4��u2{���"�vyƺ�ݼ�H�ObK��ku�-���L��򯽥U4G������})�%�E	�G��ǆ�����Χ򪛩K��tr޻��GMįq���3;X y1#*�"��dbCxP���b* �S�
�Y�ut������F)`Zu3}#h��Nti5y�R'��u����Y���{�H��[pPf�9:��2Iއo����.U}�3�����8p�����{B��u��5H�N�bAU��js܄w뎫�ł�����+�b�Ĝ�ƞ��|(����ք�]��O���t�dEǎ;����y��Fв��6�6B�=K�Z4f�L��Ɉ�_n�x�_�y�:�[�-t\�_(��VVV:����j�3 ���))����~�ν	�F{M�e��N�KѦ�|�O��э>L�	�~G�_��ҏ�2D�Jhw��e�Ww݌���I�ظ�g��o�k���<���0'�j����i�]Y��CI?F#s��u��P����S�'�B
��ӌ8}$����C���l�8_u�Dۧ���`�kG����4���X:a�[HV5���@Y��o�&��������5`R�I(��S��`��YT����Jx�D��&�N&��o���df<`����P+Y��
�I����^y����R���		FL�.fx6����Gf���[�bo�}RS�ћ����-�<�r�(%KBz���N���h:���C�C\��I�������/�&i�!�r�_"���g~5�j�����6X�`y5�b�i~b�sm��Ӳ�Y�Q�{��M=I��2i� q�Mg����Hr־�[�&,�����Gu��Ў�X�kl���k��IN��)�岎-��!)ԍ?���AW�e��^;��zc�ײ\3.d�:* �g��&�nB�p��@>K�`�Q|���"���'F��G��XЂD������>[=��p��X5W�,5wg����R��2��i�Q/q��M<|̐��XH��=um�3�cƎ�z4�[\5�@{��ZK�;�&��$!�z"�n�,���4tu�;zj����#]F���S�rR�GX��V�e�&c΁QJ��/�_#�xu���>,g[�e�qX�V����{�n�j&��jSh N�� �f�i_�Բg@��>P1̌�I��:��,�n�L����%)MC(I�A����j��W�����٠�ok!�^W��,��b�<���n=V����-k��-�����;�c$��O
RBY����L��T���a��G��/5zb��<� i�`m�QA�~���7��]b=�k�X#�v|���������ٗOc�	Nq��~���O�J`�qL�:;���js��3��?�ď@i|��8���!��R�5��(�B���ddg+�dE[W7�Z��4�o3������'>�D���ɔ�����?���>#g���p��pӼ�͵���U���B|e�oznm!��������������&t�Ii����+\�:��[�<=���䶹x�؛7�?n�*��xOɊ���/��Xpp�	qj���p05�쾱�Ba��I�^����s�1�j�d�8�V��y�����˅ɦPtz�RHƣ�����W�g���)�BL� ����������:��Іk����I�x$��v�U;����(/���(�aN�����ղa=�Hwi�݋-���sj�Wl���Lσ���2���R ?�\���.^�*�U���v7�'��R��k"��em�Xeu�[���@��o7��,F�����>GC��������.�<��
_f�CɄ�O���8���d�J��]:�sa����0��Ȧ�	�!��
�js�e���{J�>%��6�r�al�-��O��j|���	"��+�L��Ų: j�w�2���k��4��K�yzq�kߡ*'���΋b�
P�w���~�@߯���>��(�"ԕ��K�*�vY�������[d�@M�l�q 6�6��b��C#�Hɛ�r^�~���G�?P~#H�brtL��f'����/[f<:�r����s3G)�� 
�Ú�+��=5'�`" x�RD?O�
K~�<�U4�2�wrN�r�����5�m�U���s!=||�r>x"���:|�w����x+�TZxqØ�IH�;��iqY�ײ[n(WU�hK�)ff�!jC\�sZqNWVi�g�*����~;X$�j�F�L�@��2�[&�g��{�p8��wE=;��qefݦ_����+�:�J�Y����!*���:YYM���5JG�K]ٝ~�U�I�lQ#o���rp
;�\ܪ��K���!Y��U��*-U����r�i^a�]l��ny��D��m���ʻb��+��x3哥?����n��dʇ��V~D8#���)�"�w?��c��7g�W��wR0��w�x?͢',���-X��e�hAA�Q�D���5+���N��~��k��� ���5/1P<n�I%-p�l��W�-����[hR��9VJJJ�Y\�Ï���zK��f��[f&�6ڿ5��z����������;���F0,+��f��P�f��S��	�:_`�� -�65���Hsf`s���<�eP�]�T����R1P*����J7e̖h��A�+Z��۲�F.�
N��ó�oU�}�Fv�+m��Q�~G�:ߗs��Uq��~���<���n���,̠u�� ��%�mJ�r�rK�WwU��z�5�A��e�֣J�{��c�!"y�m�,��N7T�����Zwt���9��t�Ѵ=��k �`�^RR���|/W��v?�'k}-��J�t����F;
��R�7�7ٖ�?�ḿyN��G<�%�@�耄=��������'�c|���e��YA�vwU�4�q�*)KW��M�t0�����ϣ���29ӊ��ѳ�������^���8�b�=C1�D��P��Jg�����ސ�"T�~&�ǈ�|E��X8�����2O��s�
�d] 󶱸�)p
�6��i�m/N���_I�N�>�@"�>6������	�l�p�_7CU�����X�=L����m���N�G9��D�q�Lص��,j��-�r.���o�G7�*�G����U����:����++�훏f	���O`���L9��Ѻs��s��ݕ�Z�2r��	���z���9 s�����]䁏^�a#���n�����W�+��Jؤ�������P%g� PK   �<�X\ܜD�	  v=     jsons/user_defined.json�[�r����T�p��8�xʉ�RI%��k�WeЀ�=��=��HJ�B>Xظ������6��^����z�_CLy�t6��U^��pF��j횥�������.�{�g�xa�Ǔ����:^��WX:��N��~�M� 7X��!A\Ѐ�3iϹ4�Q�\c�\^�E,��7d�qtk�u]��k�q������������EC2H$�7�!�t@�q-l�:�]p_����&e��TH$��cg���!�	�\{��޴��]	��
�]�����˼x[�r��۴X/����~=(��S�	���U�o��_���Ψ��\Y���u����U��u�8R��\������3BV3*�!ltc%_��������-���'?��x6�>ۍ@�xB����C��䟝��� �κ!X�!h�}�c���Y�}�g_�"�i_���t�> 6���� ��88������D1=(fH7�H����ߧ顇}(���	���ߧf2Ծ��V�o�t�o�Y��`I'@[�j��n����x��	��F�tT�V�/�"m�X�y���wG?MN~|�Ԗ���b+mZ�O?�n�Ҷ����9�&,���`�MXڧ��E̼���OӃ�9uz��n�>]wדAīӃw��6���U��%��p����2Vu��(>4��o*����.&G+�/�.�!��Hس�1J;ĉ5ȥ��Q�8�]�iwgA��Y8�t
	�t4!g1A��$�Z�vg��ʉ�H�ЎX�՚"�f�')L|vg!3	/�����bR�����ԌgL#����X-��.zb|�>�h[�d��K�s�؄
�yB�:!�{i,JQ�z-��YI�%{��K��F��8�#�d�	+n#�I�Zdc)RΩD˦��o3��xF,�<=�l,�J)��l:cP/�'t�Xf��L�4���~��e�]DۚW]�w�ǧ���O�����I\嫁�LB!�Id�&�8���44fA�iE_�a�[���`� �K���H'l�@Z�)D.#��#.�3�8
TY-"ф��f8�ׂ��C�gZ�g�(l����S�@�Ԓ�v�t�4�T������v��d�	���*�n0����r�s�І��Zt�H)8]&�G$8��LQ
�dTq:�^1ZDhr$� &0͉��QH���E/��$B��1 �u�-�F�L)���m �Q�I�]�eD�!����������`�g�y��X��5��Y�ô���z9���M��w�vQ�'�x�K�d��v�6(�Wnv����X��7�~(�o�����S8�+i,/�f�m�i�dS�'������rT@H��n�q���f{����7bܜZ�9]p�X'��u�;��`S�����"��{����#��v�8^�>�u]�ŃPqzi�Oi]�Fm\t�;�HY.P`�5bU4q�H�C�WLy%�IB=�A�F���"�)���/2ŉ�%|�5I�>�6�*��23HmZ���dL|k_l �I�A��}[����(��޴ݽ3�3ιĝ{���y�}|r�H���C���Y/#��t��)�"�18丠N.C���n;�}4�G�}4�G��'���3��'o&?�a�j'v6�FDʭs()N'$!��ELR#�#əݍ�3�r)Im�"+�QCK�as<!	�5m��t���F�f�g���"+���0&%~v#K��Zw�J�TZ��@�bg�9�&S�_������O]�g}����� t��]�"<c�s+�����h����,"���9$�p�:��G�n3ST
�k��V �al��{�Jr,�`<҄%Ĺ�Ȱ���p�"�D�l���@:����A���x���1�LB�ꑁ�S�=�1����ɶ'���l�|���;GT�E�X@)�Z�H3E��Qq���+�B3��� w���*�QZ,���vv�so�!>AI��E�aH�4+�pĸ�oH#��D��M�'FuF�"dF��`�S�O4���c�4�5�<o�#�__���~�v_Lg�-V˼�Ӹ�:��2�3@,m��
�EB&�<냨�w�n���M��AB���@{�8E����n��u��AA����<	ȥ�ӆ���n���*�ޒ�]z4�Z?��g�t����F���~-6��9�G͏��Q˼k�9�n�\������.���+f����$Y偤8MFS�}`(F��j�h"R���K*����xÊ��_�*�����vC�1����W�>�s(�`�E�?M�rC^��^<�w7�� ݹr��x���[�M�"�<�F	�����㛍��tǅ[hg����\4Xލ�z�y�L�m��;��4��v�+�}�4�T*��4�#�q?��G�5��j�>~�s�ވ�:)��d�o}�� ��j�>��ˍx�z��y�罞�z��y�罞�z��y������PK
   �<�X��6�g  ��                   cirkitFile.jsonPK
   l�X,qJ؏� �� /             �  images/278ed6c5-ad12-4b42-b098-da68003ec988.pngPK
   �<�X����7  �  /             p	 images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   ��X�}�R��  ��  /             � images/3fe24426-b06c-40dd-b590-a579c31a1c4f.pngPK
   Ŧ�X���j_  `_  /             � images/43e0edf9-5f24-49a3-b78d-83485af402b6.pngPK
   �<�X'(�5W �@ /             �  images/4737cce6-ef6b-4e79-82eb-dab57378d86e.pngPK
   ���X��Y9-  �-  /             > images/4fde46ef-4620-45fe-a6b4-d27a85e18129.pngPK
   �<�X����+  J  /             �J images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ���X�j*�o5  �5  /             <[ images/5ca6391a-909f-49c6-8bb0-8f0a302a1c0d.pngPK
   Ŧ�X��~��K  yK  /             �� images/7ac84256-6e9c-40ba-9a9b-c812e48c1c94.pngPK
   %�X5�3$ �$ /             �� images/8251b1b7-c97c-4929-9682-a545aa133660.pngPK
   l�X��� � /             . images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.pngPK
   ��Xq�q�  i�  /             [� images/963eb574-430e-4d09-a29d-074ae2ef552b.pngPK
   �<�X�&�}[  y`  /             / images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   �<�Xp&�[  �  /             � images/9d6941e9-aeed-488e-a8c8-e310224fd4af.pngPK
   ���X�V�4sE  iE  /             �� images/b14b5b74-4377-48a9-90a5-00abeaecdcc5.pngPK
   ĺ�Xm.���  ?�  /             K� images/b2b92e47-5c05-492f-ba01-c47f59068786.pngPK
   ĺ�Xq#Q��  Ț  /             �� images/bb187b5d-1fc4-4a4e-a882-8dc83b4f659e.pngPK
   �<�XF��-$  ($  /             �6 images/d88a5b0e-66b3-4edb-b452-47f46dd40326.pngPK
   �<�X~��a� ٮ /             �Z images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   �<�X�J��$ ?& /             � images/eea7d5df-ba1e-450a-9b5e-b26e568e86c8.pngPK
   ���Xg�	�;  �;  /             �4 images/fb3f2d9c-813f-448c-93d4-6d887e4d49e7.pngPK
   %�X��%� V� /             �p images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngPK
   �<�X\ܜD�	  v=                jsons/user_defined.jsonPK      �  $   