PK   I�X\.ŋ  H&    cirkitFile.json�]K��6��+�kQA ău��ll��qGx�s���ӭ�*�V�r���_@��HB����]��f�@"���Hd&��f���j�X�������u�Z��}�������n��X>nV�?���ϳ��ܿ�ͯ/UT��_V�j�y�)˪�QUgq�T���83Q�d�yZ^��xv��U9��S�4�V�s^'Q�*%�V�������-3J��Ӳ)kf��Qn2%��le����qZԲ����9����s�gSe%,1Q��:JKGڔ*��e�����*/�$*S^F��E�%�E��ʜ�E�d��g�e_���I}f��9�eNiYPZ���2���0.=���d�,�H��NS�ʵQ�fҤ�Y�3/@�X�*�qT�ʲ͍���0�`JSՆ'����03	���#��$J�2#U�g�2��*�/� �}���f�\Cj�S*��،�4,+�겮�,��m�b�HVFE]UVE)$���r�ʲ���PYh&��W�Q�V{�\WEb'��c�S`���H�͵���E�e�6\ۺ��yQ�*��̋�ҰR%u��.l�Mjm%�2��2K�"�Յ$Ma���i�4�@-{)L	t���-C���{�D����Jˤ��3���wi���Wf���UW�A���i9cu!�JFYePR��V�ˈ'R��3/��e]'���dm'p,S�m-2����g*Σ�$qR&�*4�����µG�����bڼ`�X���
#�F�+̧X k�X��,��CC�!J�;�FW��gpܠ��,N���8M9q�r�4�X_{냫�����i'h������nHFp��^�n�9�@�hwˠ_�в�Ϡ_�вo�e	-�\��_�в_���Q�^�*8�nYZ�Yh�N�вoz7-�L��х����>݆#܂P���AM�mRЙ>�h�{'��|��(`�aq��.��!N�<�t�I��(�ƊFg0I�~L)VO�51-d�纎��k�ı�
��q�4��24��Q�De�K�LV������"��o����T�L��=B#�x�}��q� Tz{��+/��/c�^�Gh\/�\zg �@E#���4�� ]baf�aȄ�/`�la�%�x�~��%�Y��y��=!:�<�
�aP�à��A1�b�\�!ӫ���eؠ��T�����q�˼�1� TzyAc	��h\�]���/�h��>�\z�5�@�׺B]�����u	v?o�u�z�/�	�_6CPGo��������E��a/Ku���k�{�g]�������=B�G^ޝz��lSQ�z��m�Ξ�N��T`��J//�S�N%/<�J���;��Tz�v�]�;��Tz{;��T���+]ةG��;`���
BE�b�PIà.xà���/�_�,�Y�0fa@� ��A1��à��A1�b�<�y/�a��J/j`��J//�S�N��^D�zt*ax�ذS�N�wZ�N=:��I;��Tz&ة u��ۋ^ةG���ޙ;�.R��zt*�r��z�W$ԩG���#ةG�r���w���.O�qQ�2��n�e��^_���*��պ�ֳ�JV ŵ��n��cR˞o�����>�� ��Ii�w�
f6O�gZ˔>�2�����-@����e0@Ci��I�i�rd��������:{<MSM#���Pޢi�k���}N�ᴖ��*%�K�'��Lѡ��GG�����uc:��!J���2))z��_�S��$D��2�$��{�O��i�kMɨaZ�'��V𩆔�)(�^J�	�;<�@�47e�i��2�^-6�@'��%)�3�j��,FX4h3�Dc��� "��C�	���N��4FIFp���2q�X`@h��A��T��[�JC7�e0
9�@�Q�Z��10*N���4��Iـ#x"�#������!\���W?W�c�,�B�����ǟ\�ӵ~��e`2	�{	� �v'��}����a�Q~:�`��7���Yp���̂[d=L��1g�1��T:Č��@#��#.2p�4	����� ��_��&������j��a���Mr9F��� �25���A��ó���!f�\d��	�1�I�=Cp�$�(�sx���$@
N�AAV
*��}�8�<��&"1@̕�3@L�m��St�	T�1 G�.rp�t��{A�EZ�h� ��M�I^t��^t�)_ӂ �rDL �}���`t�Ya�-�prq5���g���6j`R��f!�!�t-�=#f*R=E�$�P�V1e��iwӌ�5��PB����<�h�jF+T�-��<�>�"�w��F�1 ς�!L����<�\ .�˷�G�����xD��a�d��&�>Â�d�_��&��%=����8m�%�g��m�<�(p����w��uo��z�@|����·4�y$_?� �q���4�ylH�B�9�5�L� ����W4�Q�1-r�z�#)��bǷ-F�-h���B/0��|�A���R����Xg�K�<s���)��&�ї���i �|@�/��U[(����i���}
�����oO�%�TT�2*����$}��0#�bj۰%�Q�V�4z��N5���SAͩ��^~@"���0��|��^�
r�]Xg�K�<	��A�z�i����ޗ� ����'4�Q.��w=�U
�Y_��`��*���k�Q��m��g��-���7���?�mǼ�^��`Σ��k<҂/`����Р�A>|%&{�n���%j����,|m�Y�����]��NfQ:�������[sv�0s]t'��O�Yğ�^�n攜ӛn�ܱj3�GtN�VB\7gl"v��ͻ��?n�v˭3��vyڪ��R���V�l�s噫�#o���0w5���]�jpW��cdf��xַ�RU&�*JS')D��yU�N�`��Ã���i�;��,��ْF4i����h��eq�sd��T���m7W���M����t����*�Z�yt)�e/@
N���<¿�Go�(����-+%A2S)�R�7N��`�w��A�퀕�M׈HJGh�tP���$�����)R�B�#�ӑ��c�v�t3s�s�ێ 3ԣ��>3�nq�{ۉD���趃�����ǉ0L����43�C��.��'�;B�ВD[b�-��9̵��"l��i{����5�)˫'�okh>���{���k���_��+��ۯ���h���W��*ٿJگ���j���W����_���t�*m�b�.����bmQ��<X[ � ֖;t�����bmq��L�����1_WV񮲵;ɶ^=>-^7����U��6�i������K��,*璳�_V���b��d��1��rǉ�c��s��a��:�g);�~[�,IYde,�����9��Q�r���:��^H]����X�_�M���b��ɖŎ�����K%۱;+W_���b]<U�>>H��m�{H?��Ӷ��6o�bu�d��b.��{�1m�c�^��$a�%���0-�3�H^�Y�xTUn�P5�3�ۉn�*� 3UV�\ hS.OU�i�%b���f⎱�I���2K�\�$��zdrg�xnE(���Tpy\�s�d�\�(���q�*-YV�������Oߥ|'7��ߨ㛘{ޘ�*Z^h�y!;k��ƈ�&��8ٍcN�T鎹^�&.T�Eu%�&��ίk��(��fIl7[�[�����T:)i7�S�B%sc��b/��N[�)΍��ꏛ�K�[�0kJ��<O��Xx�4<9$( ��m5�I,�V�?''϶��شܿHE���"9y���I|�,N���s��,y|x��OZ��vu����Y�<���;�����3{v=�?�;�������?�$����D��*���Q-H�6e�X�- u\����Z�֢eY�s�hk[gE^��Y��,(|M���w:�B}�`�i6��ş وtgg��9����xE��C&�L���`W�Ḓ1"9��r���̚�\�(Mc+8��F�deČ�?V��t��~�Aq���֋�>{�Ug�5������m�=�.�ү��b��ms�=�J��~Ξ��/��s�S&�y�?�-���>���~[�+������J�)[/6��?�t$�˞�3�ߩ�~^}�~i�x�����k�l�nV?-^�9��â��b��ñ�m%ˍ� ��i�z[�߬�V��ޙi�y��w��r�߫���=�j�P���H�mZ����=���]�^-7?,�]uR=�<岗���	k�����ղ��[[祊)k$pf�]^R5?3-i�Je�̚�V�9�te��g֐Պ�54W�p|s���4'j m�皟�̚�r.N��T �)Uε��5ൈt"�H�̪k~��@�2:�����.�U�v'������Z�7!vV|��ޘ�wKZ�se��{�3�o�Dm�n��%�Z�,J��J�_�Iw���-eS ���7���v��|�ĭm���iTQ���c�R7^$�V��G0?%�=�y
�Y�.�漻\�#��:��Q0��*�9Sl��?�y*�X��3̥��I��Q�����Y��e	k��:gu�b���l ��<AJ�o0vϒ56����`��w��5�Y�Tbr���$�zm7�gr���(�4�3i��Ȭ��9����m�pk�r9BYG�U�.;��e�t�W�n����`Ϲ���0�{bۊ��a�ct��V������bv̞��[���u����i�w^��� \�C���mod��=$�֑s�s��o���2K�5��ʮ���٤vF�qn�����>��J>��Il�⻝8��T���@dv/�ǉ�&CM���Y�~[l���|sulOBC&��JH�J�\�OE���]����Z�2�x.�8��Z^Yi-��`V-�J'�[�4!�B�Bʛ�ޢ���v���)�#:q�-|6�7a���Yl�`�ε��]q,H�s�͗E���(0ϭD����j�����t.t��]�Ҭ��y�"������͇u�������Ow��-���
�n�>��?�������G�lm7��o��i�Īey��W�%�ξ��5K�?�q��Z�-u������Ǐg.V�}����a;i_ݯ���p?��qk���^ߵ�4̮c�3���,�F�O���n�D ���b� ��b k (p7��x�pN�YL	�5�V˞��JM'~�ኔiA: İ|lbPzv`��a�����@�8�H!��NP��H�b-5 >ا �4��3��P�_�l�j�'ީTDc�BJ}��(c*�1���40��L<�X�6K �I�$�` k���9�BT�`6K�s7�B/��k�[�I@6��IA�d�R��@��҇3����2��U��s�3刍�n����+ز�}��^����L.�W��5�֗͐�B�Mv P�_��[G�bo������l����׍R���<���؇�[�LC�>��1�Bl wC!v�L��F��s�����e��<j�4`1�/Y����.8b�L���G�����8�
�q�xr8�Ig��:�ʗ�	�l��vC؛l+���k�n�<'/6�ZĎٙD-`mR�x�	�sp5KuG`���R��+���5	��6)��S9�!��R�<Xc�� ��������X���l�n7R�4�jS-����8_"�R_9����ٺ2pD�XĹ�E	E@�U�A�,��?h0�� �:��3���v�T{ȿ����g�j0pw�����Vj�\<�t�p�<42Ҡ��:d���KM�20``'�N��M���+5����ر���o9p7ԡy+� �Y�����;'x����MSw��W����(��4��p�C�#m k�v��:OE���9�ʁ�@�LV���������������A��f18���А��I�X5�W%I7��g��:�p��a����É;�q���;���4;������s k���\3���߇�c�5J��x����rc,�X�o8t������U�H t$}�r���nî0t!@`t(��e������wo�]Q��æ[!����)��p��h�h��=_44Ku'�ʳT!����q��g6GG�A�Y���v��,ц�g�R��6Z��k� ����g��)c����A�K�Ǯ�	=�p�� ������Q�;�IA��5J���f[<=}_�m��"{z��;��n���wU~�-߲������Tϯ�C��^֫����ߪ�b�xٟ*7�� PK   l�X,qJ؏� �� /   images/278ed6c5-ad12-4b42-b098-da68003ec988.png�zeSL�5��ww�ŝE���Ⲹ��ݝ����ު��3S3�a��z����1j*��HDHPPP��rRPP�|����N.�=��@�k�J@�ΐ�AAQ@�K�ky�\�<':����>�������w�«P0~�o���b���F��a9�5E�5�P���H�B�V�Z 
"D2�[��B��^:M�r]��/6߶:�Ӧ��a���X�9�lz޸0���W��L5HƴSʹ߯��l��4d���}[%�7u�[����;;KW[��1̈́��0�7��0 �LN�c����UP�ǒH'�13���1���#��Y{�Y�"[Bźq�kL��ʾ<�p��������#G��	��Ṧ�aj\��L��T�6���)e�矌v��������P�a\�4��Ԭ����ŐyA�^�pMZ.GZ�)V�:�S�J��		�t�¿E��!�Ӗ��}��}s7~!�t��(t<H�У�H&�K������e���qҭ�%&�8�R�c~ꉑQO��DE3'��t���k�{`��>�'.�
�1_,B6��<-�� ���m��1*���s*�{�YuK��^�w�B@z�R��&ed`?{�J��q��L��e��P�U��v8p����a'Af�N-��O>`��t`zi#������ap1�Ę'�pB$�,Qܜݥ ��ՠ�����K����H��������l��t2}�*����>ZM����u��=�~>�Վ��ih���!�y�tt2������дd���>�kL�E�W�X`_O��N	�w��3�V��ݧ�}/�-aDX;ڢ�{�Y.f�/�����>�
2����!���(1��H0/��D����(����yA�w��Op�׶b����(QQ��O��Ó��������
��|�5��a�a�<jUMBLp��R�1��	$~�������:\@qj_X��М�7��ɟ��PL��58��_��A/]j��R�RcG\�e{�ljS�?�H�+�[�$lz��X���i�:0����}����C�y��33�]`:sd�] )Ã૞6CTE����6I���֪�I���vr��;��P#�]�P�[���,2m[N�Ay�JL��4�!$&�b�2�HE�DŊ8�TVI�Ǽ�K�W�s%��5�gz�(��j��晎����O�A�8�/,4�ح���H�p*z%�Xa��p���]$�M7��8l�[�c���ӗjt���Q�������V��G�F����[�7�4���InM��A�;&��0�[&�ޘ&���(y�DT>�x���iN&�hTw�$M[hb��:�{�[<�F���_zf�FB*���Q���=�0���Y���.��\%7�h����#P��n��PmUҬ|��n�O>�{�5���4/J=J`��� ��f,���<H���n��*�������U�*
ć�#!y#�1�6!ӧ��R9��y�3)fH7��2�����Z|�c�����}7���t�u�`&Ԋ���p`mG�l+���O�|�,W��R<���o������lV?�ʈ.�� �犣��6=<���_��153�3=l�ѵ!�:/�[:n����@k�����zhygm9�҈Vd��O/�m��R�+�7���U��m�v*V�8�e�v��G��p�5Zr- Be�|N��,M�	re��ҝ,��s��7���C���8�(�jY��>y�Py�%;���"�u)�hq'}p��'��N!U����֐��$�Paˈ��&���?��(:�{i���2��e\( 6�>��%'�g��� ��C//��\��U+��Med�C�g1�.I�v0�n��5��'�â�F*�f�J�CqIcyKJf��C��%|�ڵ�r�w7&c�o���|y%%N��Rႆc`��f�P�g�X��~�[3�;�����"��2�>E��2���Hu Gcab0�k�UG�ӑ��2SHAQ���!:�}�Ӣ�c�}��<A�O��Naz�T�kB�:��Z�HV�j�I��9i�2;d�=*��48�:Ρ��g��ҭ~���#�^W ~'�T�������p��Я2����U�Ĳh|�q�`קJ�b|�D`b��g���'��fZt`��%���c��bȬ���n�B�!|���Ma���H���"Rc[������N�7�I���C�M�q�gY�bh.g��88�2G�w�(s�:��X���9��$�eM�.�\��)�9���03܌�2�m��9B�ƫ{X�%�vhe����u�z�3i��!f"E�L�-G��XL��RFE�����\^Z�kUy�B�w�-V�V��%[�������:~���/9����X���ұ�ef;d�w�����O����ݧ�e�s�1u�g ��
��.�
a
7���D��[E$%̬,��R��p�I�bȏ;����aP�lJ-*����h9�-E�Z�H�!*է�/����~�e��[@�"v����9.����:4d��w����5L���K�˴
���a5���Y��M~��9����f����*�Z��X�n�u8Vd��C����I�.��e��|����q{`Y
�eRJ]mW���K)����������c3�Qu�����w֟l����T��B�;���^,�m�[��`������~��"�$f���euÄ�";�Ƴ���`J��7]WU>b��Љ��>�(���qf	����\]ܪ��ԣ8x�fk�h^=�rN���B�WK�8��ɰ��.`Y	�#����������b�_����-/R��cdiS#Rd�n�Ǆtq�i�nQL���S�!0��n���^5�s�󕫙�6�{�q������S9�g���Jl�wu�|�]<IݎL�{j���[ 1��p˪ҏ��  ��3`�3�ײ���1�݊>w��Ȩ4��D{�.�|9*�
"��8$�-�j�$f�"zH�����!�,�^,Q��x����K�]%g��Ǒi�j��d���j����莁�f}�t尿�-�����_�@>���5G�x+�P�_�,u�:�Ao��
 f�!S��k
�x��$�c�Kt>1�Is�ؾ�*I3�Dhpf�8��0� t �Ķ��)LH(y42�9sbZ��<��*�u�%W��R�Km.�����f��7���\��Уc
����1��S��e �:�3�'t�VqT!�7�us�a�^^a%�3v��d<����S��Ub�G�x��{gg-,���6��!�r����������Q��a�"��6�Y���R�����J�5b�kP��k[����4�:[�&�2d&�]�h���58f�w��$�]�g�h�R�!OU)�����D����x/<��{�je߱~��3�%�gmZ��'K<�@��*��N,s_�u����F��S�K�`q�U1���?1릂��MC1u�bDj���F�	!7���߅=0{P�H5;[����r��e!�}EM�jqT�1�$WS_�,N�ǁ�B#0q���wfh<GK]_=�;s��I��m}Y%�jG@E_Zo(�R �3�2Cl�]��IN�u�;���"1�M� �C��"�Ը�W���h_�+%2�Ѿ�*��43�4�1�-�(�}D�W�-ڸ�E�rS��3����U�Q�'6.��H���; m�"=.�m_���^0z�F�������@魈5U��� �u���a�g ��[�Q4돿�DXg!*��~�� ���kL[��>0�`j"�ߙ��b�X���j�9�� j�#s��M��r#��`����n
��oUt,�b��/o|}�)*6p�c����0�G%�����?�{��>�wRK�I��)���E�K�ze2�@?��+ͅ�@��/�,�"8k-�U�SU��t��Gd��Zr��)�ޛ�臆w�(��t-��m8��[F�]��?��gGnH'1� R܇0)5�j�F�X#��bCl?��H�Z��T�nh��]��#mO�=8�����[�$>,��5)���Yb��H�z��]���*�����u8ߪ6��LV���[�r�)-�b=����Mǖ�*+�����5��,��$_�u����"��Ăa_��Dj/փ��{(�yE�ܓe���G�����ť�i.�j;P$�%��;Rx0e��Ss��d��u ���)�XF�t��K\�?���;6�2�I^}����P
J�b�J �F|�M�&��K�M0>)�����P��6����|�J�\����YC��)��]V���ÏLS�[���h�Ȭ9�Q��#M�Cӳ��~�3/�ஔ E>~�_�]0{Q�ϔ|�����ǋ �	���O�/��h���k��?���g���|ɕҜ2�w�i
N+�o7d�G�z.�2)G<�eޓ��-�L�ʳ�g
��fq
K�#&��34��O�� �$�H�2�>d��p�W�r�_�on��YlU�a��,j���)����<e�CWٰ(C]'��5�M���;;���Y���f��G0�.4	�63�	��:�bT	<Ys���BЌ�c��H��>��Pz�-j�
?�10�T����e~ȳO�>����r��]�É�-����'�oX����1W]�=~[����aZ����f}A�d�n��V�S��h1ʢ��+��lq.����>'�ʴ,(�Q���V�:{PynolNa$�f���;�352���2�	��.PPB��UζGUǪ7��$a���=ll��Q:NZ��v�zַ<&�1�'�(�v���`o[��2�b�:��v5��:��𚧰D���Ï�á��@�M����5i��d�<Q*8ci�K���p.L^��u�z�VWv>v顜��K�>=�/��!�`|jV:�E��!;� ��pAx�U�.
��9��񣄞m,��P
Y�1��xґ�x�Mz{_mOM��Q;m&[8�Nq��W��H�-m~[�y@H�i�'��!��p��O�&�P, ���A�T$'�T<ݝ~�`��&��yY�F���S�?�Q(��C�+�);��d1n�8��^.L��Y#��W;�]�V�T�V��..�Ջ��}6�VF�C�t���,������m�׉��*�q� 6D�@��7�{�ő�@���V��J�t��ƅ��� utI ���ڂZrw���)�\'N��s�#��.y:���'�3T�-�����&5�><$f)R��s�M�p[}���F��F��X붣�$���%��XtCCF�m#���5O�^�+���e�~���t��c�umYȘ�}=����sk�R�c�<�����3\�� Q79�3�~��XP%�rb�RǦ<ɐ�#"�q�PKw�x����h(1����!8�S]�˱s�ӵW�m����K�$Db�>���oy�rA<�Q�(��#�>�5B���u^���m��&f��E�4#�E�7�6��+šR�0$pLPAX"
��8&�h:�D=��-��&-!�����]�l�܌�!n��Y�ڀA����j�,m��FrQ�X�92,V�TF�x(�l�v��X���G�%a������\'J�+�>�"F}�y��
�k@�7#aJ������:@�їK��>|�%�: �\ª�	����`2`��޵T9q������vʿ���Nyq���o�����dhS�ȕ��}D�]e��@	 =2(�?k�n�eA�8�5�:��L��;!>��p�SO�[�}Y�_7��4�`��/�� 4�,�/��lMd�'>O�`������xk�����g��a���
�x�sd��5�㟕��6��[���k,k'N�16�{�X�БF�K���?2&�	����N�[�	�҆ �}��)k{r3#� eg�l�-���RH�{?2W�w�Q��ڡ-|�h����]���@grS��k���Ԇ�^7���8Lp	c$kZ���F�y�6����"���hBry�j	C0��4��+�DoG<�]7�#DBe, pcߕ,9�`k�e�\:��ΝN�� �Uv$áD�I����p�9�,���M.��s�S!��p|��R^�M�t����8��u������^��j`ð~*?��� �4F�XY��M�ǿ�b#���ic�?�P
���VlL,"�pw��6l ���U�(�L���cZC8`#�N/�,�y&b�Ջ�`��S�p8�1�qRϠ(��aAF����=}�UR�.k��i8�����W	o�E��g�|�6�$�}3|NY�ӞIST�=�����Ѭ�w�[�`�r�:I�Օ������^&ͺ�'�[�(�06Fa����������6��j@.�����v��A?��e�/{�s�}�i1�[?�W�g�v���R�EEG���QM��ң�ux�Mb,َ+�8S~6 mFy	GUS�`#=�?�8�>�9�'�)����T'����!�(L ��DHp�{�m|�����2��<
}�����i#7%� ���+J�Wv`k$3
� `�� d���S�m�ϡ~�؆"�*:��4��F@p����ɦ�	&���x��yD��O�IH(���vo]�}���5i�Z�{�v�{v�|J�[bQ��`#�Qd��r��fȶg��B�A��U.h��A-I�jki��	>���|e��rm(#�V���:!.<�����	���o�	����:��p.� ����vX
�[RE����� C��?��T���(g��߮[#9�8f�&qz�����uc����Y���	y�[7�瞟�sFqxՆi2�{J�f���0e�!">��nF�*y��E�[&)R��F�sR��D:گS������l�m�ibh1��ā��xo1L�`�PG��;ZhSh���ֈ5Ƒ�כ΁r�A�[�3Գ�s=^������������p	�3�/eX��������{���#k��,����Lo�P�),����|�AAe�J'�,��R�E���u_�ͤ��	/FjN}x`�/���]�_��%_QN�;����*�f�������N?�L������ ���W��'��|�F�f��Ws�;A<-���H���$�9��]	x�լ�=�/z.D�XRK�(\�N�ᓖ!%gP�q��b��鮣C���N�&,����"2�vCCIxh�)#����~�zU�#�}NY�X��t������R4Fd��"�	@�e�ǢD5Tm	JC�5c�p�Y���g�?BX���)���^���9�J �O�w��˛D߱n�P�3?j[����3��tϞ�B�(�N�����- ����>@7йe�lߛL���TO҅X�C4��&g&�k(��Nm�2�}�-��Vg��ʂ�<�1�RA�L�s,=C* �q��`�p���-L��k��~�WO��C���HI`�]�����$�Y�����Ƭ���W�+b���&I^��`���aKT���Ǘ�<$��YW_���8�fAҟu�w��$bo62��������Y��x����{͉6'�����'�\���s��a��J���ݔ(��_vI^Yх���4���I�hP^�&h`[��u��,QZL�r�����a�T	A(-Ee���	�W��gà�����ݞ�^��A��D�����>!z�[���e����z�Z����'�k�-����HS�/Ew��)c�= ��+[��!Q�[��H�����bmI��U�{~�ϡ��:���^�, Z�M	)���.�~`��s
$ܧ/8,��O�3�P�>%w��m�W#P�)z|.ܵ:�g��+'������Ǖ�fÑ��@M됺�����ŀ�uE��.�Mza�E�X����ҏ��Wc~3{��!&�V����՛�&��r��N�VM_�Gi.���8ޗ�J@s!S�4P[:]��O�n��R1.eܨjX��P��
y*�,$���;kn(�Á��ո�@Ʀ"�z��|�e�}���~_�JKH����
�e��-9�G�4'��U�煮z%��|W7P��""�NG��u6w�l͙O�3T���ޛq{���������*�k��wxIP���	]ՂaGR�	{���}�#���9��9:ʟv5"�'�S��%5�x�&\e'5FI4ƾ~�_/ ��G���g`�43A�C�ߪ:�|r�x������/�746��-�s%��JwbyN��H܌or����v4�ّ`�#�g6t�ҏE�W^L��]f�g�r��sh�v'�p2�;�}�w��T��c�wA*KbٵޤX�<��6�mm�WS��4e��R�i�&MD��x��R�+��	�҈���0d�6�/A�fS��f���� ��Ń�g��ܐi	X�Ÿ�m���`Ċ�ǑM�75�O֤9�A.����}��~p@f�/�����:O�E�MG��9hGB��p�����i(�]Z��b��	7����-Ɩ�6��U��8��?���|/$��bSlձ�:Q�a���E��Ö�	��G=�+�
z��#
P��H;�����]���y��e���ρ4݉��S�9᲌�i,��QJ$�y����~\N�P����$؈ ��G|��qs�������N�ȣ���o����Q�(�xYj%��\ACb�=ew=E��G�Ţ���'_[}OC�O6�kG��y�?x�KɆK�=�ܥ玎I<�B��ަ�e�lԜ�5@��D��O������������r�S�=�� �� ��KYbD����RKhMq������e4Ҙ�憮(���rMJ�<դ{tR�&�P�~gx�>̫�lS$p�Kp��	\Wa����]�U�*~\����I0**!�B��}�-��|z�����f�T��+iד����A��l�r�
{k�"��b��Z�ZP�4b��������'��#��S�v	6���A�d��_1.bz�uGp��݇���d��g�g4��I���%佰3��ɉ,8�@�.&���ed�S	�d��*�/�$�Ҧ�mJHf��0��Gq7���#u��=�9�d-J8P���K�븻4�[}��6�FԘ��gbU- {MG�V)�<�:<�����3�5&՚���"�IE����*��ߵ��B�؂J��M�fH���2��b6d�R̃]��e�!��s�B�`@��mR-�,�|ʳV+]�_�F�1�|����.݂z*'�չ�~�i�W���-#PN&dS��n����hW ~"�EŠ$w������:��"bn���ߗ��*��j666UN��Þ�:϶V�N���HXv0:�?9�����p;��d�|5�e�M4CN�)D��&�����=�A�r�U^9���#-���3�u@[p��`����ҟK�6ϧ|�q���.`+,&XV*���v�Q�|*cU�-]���C`��L�;e�ўvt�Hs�3� ��ըe-�m�� �J�ƵȒ�`}"��ĵ�U�^dzL�y]l���4�I�E����=}�p��z�+���b��r�T�rD�y؅V��ٵ4���]�G��|TY�h�V�����n�ƭу>y%!���UXl�AioP3p&9�ݪ�~�2�G�ԵV�9�ӏ�Q��N�Bs%�m&���(w�h���2&�=��j��zK͘;f&D�ߐ�>N	KR&gO
�ʋ�B�y�@y�Dۮ�����Siw��Xj��ƾy�vJ�DQ�Cu������B��u�����2qjR֥�9��?�?D�!eT]�%�L����y������9P�=*��S��s�X.����55�*�q#b#[O��~|�l�Ӣ_+���J�D�ea�e��lvn��n��R�.tR�Հ6�`�4I�f𛳧��p]Ҥ�(\Ԣ�ϣ�խ~�Ⱥ�^��nu��r�� �Ξ�h�
EӮ�k�\��ҟ��d�F�����q�Xٍ��L� O�<��������7u����cOl�_���-�8��4e��zZ�����.ggI#����
��'�bRܓ${���E��OY�ѹϐ& ��pC�076d����,���^|��A~��5l+�j�?5���h���˳���؎�b�R�蘆�8(��/�g��H��f�Dퟕ֚�Tжs~�,]���}�w�
���y>ݞ���:����������;8pDGZ��]<��
��pʬ�޸Ҽn�x���謚.l\�#n�q&�q��7{�w���n��	4y/�6��zbB�B6�;�3���DJ�3�g,�M4(<� ��S'[=iϊw�c���ѴPY,��n��&�m Hb{@���䕴JN'��H��Z��=k7�50�!�s��@<n/�3�~�D�s%��!���Mپ�#��S�+N˿�Ke��ւEM�  �5/�?��
���R%��FP���8c,����	v�!!Q]p�iRP{�|GS&�FA[#���޹r;�`���N�]h=�& �8�1�nP�2#}�)c���OYnkʚo(J���h��^����g$K���m�br�ո���e���M��M^��k�J���S=E��%@�^�oVѢ#��)�[�6����s���M��}y@p��'������-0�<�2�L)_�ԻB@�ګ��%�΢f���`tV�b��4����xj= *�k:���	Nyܓ�+~�Qo����*��H(�I�b�©�PG��tH��=�Q'dʆK>�!o����Ysʃm<!D�S[@���eֻ�����	�y����y[b�y�e�D�d����SE�6/Urt�g�SѠ�Вu��E��T��ZL���H`ɀux�[葮��Ǒ�T���$��z�4T��K"�V�<")|UppԞ�\���MI�����^�{fn'n�-���zHұ˯���%`L�Q�p�W_(����~�AlW�ԝh��{]
���J�xe�1\����Ñ#v��'��<�$��j�����?��3��ߪ/[԰�.O�"J�z E>f�)���F{6�%���y�u*��;��)�I���ImĐ"15r�1��-)!�Y���`o:��Ǥ��Ь�F��)����/��ì9^y$�)Q�'�ƨm�t��V�����.�3�>J*����K�R?�i��9Lca���vdz��3FB���-���tU�ib��6�kP̉'_E�:G�I=���$r`mZ�mR��OC>M�����<"�͢�m�	�ߛ���F���,�g�5E�$�����ߦ%�D ��Ύz����A����"�0B�������_}�z�;�"��m4BSR���J:8�2�?�d2��8�|[��yҢm�Qo�zd�W7<mP�mc-��n	�T�����E��#I�[�^!�X�Z��<#}�>��&
h���0�TYjsſ�x���\�;o3}K}Y�O���}x��
�	�:���۠�_�Z�֑]}�G�^sjm0q*!\Q_ą��/��g�c@��˻0������/j�n0XKz�������_.����t�
��_/�(�&��v�yG�<��䤦��aW.�"��.�!�8�j�D��K�R��4��RG�������Դ�t�}0�
�K�j�����hm-�[�z��#�t�Wo��փ���D5}`�@��κ2L���XA)\r���J�#� �+9a��z��N�bL�e�Fp#�!�:�QO3��l=�I����=��[Ðf�閄~�\{R��
*�J���P�\+ts�O�j==��iqh6y�����F�)�`R(�Ǎ�1��b��t��Ϯ�H��fQ����}��pp�P�f���c�2�[�{CM�5��J2�����&���(�O�-ۙ<e��g��)RO�wA'nԡy/�����ޞ�co��k��N)�Y�܅�\��s�zcjtTn��#�UL��KR�UV�ne�@�a)���C�Y�sg��`�������T��4�7Md�v���1��df��L
�L����忐�3��	��=^��j��x}�cP2*����A��͜h"�m�y$�8�q
�q�����`�w��	�T��=ȆL0胛�w���)V������i�J�9�f�r�)t�rB=X̧�m���Z$_E����2�U��,̷�����)n��h���o9ʀ�")�06�|�y���qi��?^)gG�N�^�#l|��h�����7��Q3YH���:M�<��駒�e�b�%g�#V�\(L��Ǫq�n��?jw��$�̭w��n�.�~�͝{���JX�����+PXY�������}58CYzare�z��eI|�H���
��a�8��-n�V�C$\"������-<�X�Mf�{�L�(�R�}D����/+z&���Tl��4�[����nw6d@%�;��\Ke����ie��a
�qr�t*�OVՎFp$�i�G��{r��l0��"�~��}ؒyۘ尢�G[T�WH����b��<D�y�6Y��Y�x��B�O�Y	�����qԈ�|��m-N�U�g��S��Ë��;Q7����IKi�|�!	2�qK��~�������YG1��v5�ONT����9��$�ö����l�����G���Զ�H��zvP@`ȸ-�u��h��"���Q���:L6���Ov�A�	e��P%	�6M[M��df>�|+�Y��n�������)�w?:{��6�˅��ף���?ώͧ����Aɤ��p�%��*!������kve�aվ��Öx��I,0d��)҉p�#/&��B
��]`|�L�.����i��W۩x|���~�z��Ԇaw��x�Ȣ����>��v�?����g��}��nQ(}�fl^�3�b��"�Ġ��Gwr�7�j�c����yH�E$���Y[驭"F�َ��@���_�eb,#?�Z*�Yi����Fboh)�r�W<��k�h�Ƒ�؈��$X6��<c�ה�h|�c�Ƀ��o���:�!D=Q�#�b��X�"0�@S����%�uT{�̽��BQ`�\&Q���U����]%�N�z���jQ�M��<��b�*�M�g�](/�ڹ��Hg .)itԴM��Q����(�<ơk��Ü��\ٴ��Cw��T���:g>9��?��g��/%���^��u�<�y���J��E[��-�ķ]:_���IuF.��]mIi�,�}�F�ݯ/�b3<R�{�/^�"���'��U�Г����KB�%��*#�Hh�)���V�#�+:d֗c�g�hg�#�����巸H�����|\@�5%�����o?x�pߖ@��[Hwn�h�Y����:�SA	P�{�X����E��j,ݻ�mh�we���n*����d㥊_�	�;�L9�%���u��������0B�&�n�
!��K�Y�3�T�{��>̔z9C�m�=�1�J�9��������������)��hm���05�-����p`'+~���������v�:��&բ�g�tũ�Tz0�%���,p<?�ڢ"-yڲR�c,K[�p������=4���yo�^1�c{�ƛ[�ᴴqʝ��)> �a����;a��=��p��ZB��B��<�C�u&G&05���� ��N�͞U�zȝ��@Ra�%�` Q���&т+�=��t�Q�!	��FE>�H)Q���mg媜!���q.̏��%��UWs=���+{;R��w�ԫ���v�&o>�&J�uF�s`�GF��,j2=Ƙ���ՆF��4W�	�
�V�1�D���)�Zd$��G	珃����+����y�ZN�q87���LvO����˩��l�$�=]+b��-l[ �K�K:(���MD�l�'�}��}Ps0	��1*���Սz����|����8 :ls��f�³��S�t	⁨�Ih) N�3RYS�!C�o��C�.����;×�����y�m�P��Ϝ��C�d�s�Z�LـV�a�N�!:�1�����/�'��Y�c�9eA�DπJ(����YU޶�#��7Ag�3/4��.��7�����aw�|��Y7�� J�+3�$��ܣŶ��1Ms�b��G}�tm~\��Ƽ�^3[�G"rL�dO�w�zc�����[xcO��4���ZM�ea��z���������T\�
~�#ϒ�S����}�c�U������w�������؅�����V�ʆ�����!y������xg�"����Ӿ�{x��V����i&*pN$DƓ���5fp�=�V���2%5��ؤ���w[�N޼�`�M������풚.�6��T|���t&`�O����R��eK۬+/�Y��5z$�JJI��][Ӽm�A���Ɓ���(!���P0&q"���!�1Y�����`�p3�"ʛ��KY�t����_!�,�k���G�~}�?���������Y����$?f�A��aa=���:,-"�"�|�����.I
��>��hmcc��^��_���~��O����!�h�����^�9��mw �]�+O�?��;>�X���dŶ`��>ȫc���6��Y1��b�����3(O�47�@6�U���o�),$�� ��Ŀ����e�|2d)��Jј[J����X���J�/M�����-�����G�D�����<��Z����C�b���hCK��%E(c�d)7�$�ٓ�l�NR�\��dHl�-��/d=�K+<�+�7�;Ɵ+."�e7g�O]ooB��q����AW,�Z�	�Y����H�p@�[�k�_�>3�r"�r���%~"v��c��a}%�MQ����ZM�mK����� �X#Ų2��6X�)7�����c�h��y*�u��7�_���{3q�謻�$�B�Z�]9O�oL�?_ĺ��}_v�:��[	 6�-�H���� �L�+8��d�˯��mm�1�v#t�c�vN1�h,��h"i�JVW
1%
}�;�g�Cc-�Df�\3Gߤa9�t=���qB0�� �&a�ɳ�ce�♼D��U˙m�rf�?چ>������\�S��-7�s���~�x4o��)=6�Pv�	[���N�0G-l*�<�D&����/��(ntb5�dB����,le˄�^Ka��]?�^��=��T;��q,���X7����������9���`�`V��bpD�5�`J�:Su%�s��vpO-�S�ؖ7�������$�K�L,�eP(��hjB�6�c�ĝ��v��f��T���`��w9���ܷ��=�,6:���EN{���Y�XE�=v���`���>z���~�G��������2��~�`��J�&����x�7Mꑷ�1�B��|�i���W3x���Z(A�6��.7[�a��(�*w�g��mz�mm!�.��w[���]!\�`��[Gk�t���v��\(�\��²:w���#e`��
#ʥ�}p��������5�A��S�8y}�~x=�Շ=g�:8�O&³��e1Z:�9f/R�6&�W��}��'�D0g�����N�{�6f���jc�C��&��It�=����_�r9�k�!�-�[�C[��V�e{�F��l&��AK�|�:�e�1�a.8�D̑��M!�WKo��T��_���G"��
���j�����0�D��e-��H[�{�h��A�{mkcV�~��ؠ���7��7�K_�k��&qNE��x�� ����x�L�m#�r@F*��F߼ no�өA3}-�������زej�$��
���'st����z2�t<cz
}s��9��Ҕ���js"��r��EĢ�t���T��;�y��ة�,n��*N��D��;[z��e�4�f93�D>=�'��`�*I�L��K�ʌ
���v�5H͕�+J��������O�aQq_q�7�	��1n^�J҅1����}��W�7���נ���V��Օ�<�v!�u�uiuU������^$r�H�d���ŝ�/ǋ���z��`��;��M�Ŷ�Ah��>�
��hmx�$��h�Ãnњ=]%ah�`g�_pDRI��[j�Z'��`��-��+���þ�+�5p'�KJVB�3Y+�m]���]���ʢ���HB��QZ����>�P����V��+�#��{���|w^㵳��1��F����U��S��p`����=�
�����;�a{"O`
����"�:��/��/RS�vQ�~�*���u#���0�yW����֥�pR���=�4R��� �齔�N�.��[
�:��^�$��&y�M�wy���p�*��f]v�A�n��w??L�w��T��7��rף$l�~)��$�S�3�e����=��}��m���M1��9�lL?X�w�@ eP����� �'��o+��Xs�TV���RY_l���)p03�ҳI^]�<C���I.�������3O�Gb��+w��C��~S;��F@�|I:Y�����"�ӵf۬������}��Dz���� 1@ο�;=�1`����c���T�i�˄��r`�y��Oe�ܕ��]yH��:����Y�2-+��p}���dݙ��kJ��nwZ]IV�;�
w��3ߑӚ�h���L��\4�5�:�jq��y�������cL�q��IS��O���;��10鏥e�k��X۸�R,���SI�	�cW��6�[����&�,����#�����i�!s���'�h�䐦�������P3;I+�X��R�{&��J��=R�-��-P�R�̽G����x�y�h��s\��#t|ԛ-8��Mְ#�k[��vĨޞ]!� �E����}�L���Tp��p�b�T�4`}x.�@��J��oon}�o>�S_�����õ���9���u��/F�8p�lm��s(_#hT4Cd�q���>i�L���vsʎ�˲���M´|6��ux����Qw_ߺ/��茦v����p:�Q���ˡ)81�8Y-����Ǜ�b�����^����q�\�<U)*���w�Z�«���C�L���{�5�����������}Vl���s�ŽWi�ￎ�J[v��ѵ��LlPo���:w7w���)�V�]_\b<��jʟ0��|z���3\\_����ɿ��`��E�ՕҞ��%��}I�sAt�]���g�$;Z<(B�v����u2$�����4q#� ��*b!��aW�5�J�*e��?>x���P̙�1qb2�.]Wy~u6>���L�,ӞU���,��N�|("���q�eXJp3@���il˶ly�T-� l�z��T�҈a�	ERp�)�Y�zP�1�-�b�p|�z�%̍�� �1v���^�`�ݒ	�޴�h�����d����	k������h1���)N���f����l�[�U�à.a<��W/0M�X����ÚWǃ�=���2K�]���D�t?1��PVJ�����l�KX�L�p�3��H��������&�G��]��R�5T�X�D�i4�ۃ��M�sDi�rc��PG$����0��pq�Τ����MRAg�M ����_�����z�_��M����A�rt������h�x9���p�qL��j��:p��&'�)�hbx��ܑl;|�.�̊�ƀ̀�'V�����������a�ޕ��/�p1b�/�9\&�)%�T��1��H���=��w{����x8�˃}|z�/  GȉfS���MT���/�1B?��Fc�j���yI��/�p��g�n6����ob��$����O^��WR�J@統�[����AMy]]KW��Z���kaTϏ��1���v��Z�7�=�rZ������-�7�k��{��3���c	c�fx�H;����߽�Z���/�^�r0��Ύ4R�V��67k:ЉR�V^�""5�J�z��'8��2AT�1;��ϥ���kzy�F�RYa�ͫ�	�l��{|F�[����Ķ��c�h�L�ڞ��b#O��x���s�h�ݰ*QA�	��n���S_3 ͳ
WI4Ro6%�?q�N��l�-Ƹ��5~�J����6�[4��<=�x0�>��Z^�.�F��$L���֠sN��k1osc������&�-���z���|"YҌeMܘ�|��0>�4A U	�)AcG_�_�$c���p����Q)4��1��K�_�7��H���U&�V)�0[�$�qisʁ0!�y����]1�S$��}`B
i���J�
�＾��k���@��?|��s=���U�[�Ѹ�jr���Ø�o�wK��&�6�[y���Ow4�T1j(O@,%�fI���T�Fû0-PI�������lW��,��#a]l�2Չ�/X�u}�I��	,��'9�v�xsW ��x)pqy���H:,������D�w�����XX��ݵM�t7��X�8����?>|.m�x��.���oJ�i.��� ��G�/ğD��kACt��;w�t̯Lf��ȫW塿��S|J=lp-�D�erf��&��k�wP�*�__b8H��n�%M?S�����������:�T%Tz�{�����OO�N�B�.M���S\�_���L���������T�'WG����^�₭�L��dΘ!c+w۲�Z��x�s�^�4F,����!��w���b�Up�Nג�-$\��5��d2�P�]����dcUa�`����D�	��U����Q.�	�&@<7�͂��f�NN��p<���'#aml�?*9��T�fҊ���Zn ��8�?D�^ܭ?Py"ِ��N*�%��}���5����f�c� ��:��"��o��qӋ��W�)C�A���C��l^J�լ@1#��N�W�HB��ͻ�5̮G�'3�L��.�FM����I��<�YE�y��$�x��D����5y=-H��G��U��V��[�0����Vm���_�������s��'�4ϣ�o�����.���h$]Ab%�=�s���
7Z,t*]�3��Y�i���a�L�&���� R#�2���*����6�����z���V�q�	�;}!��S�Bmw�k�{�6��Z]�@�:�d&�d����Q/� ��:��h ;�﹒�����쵷Џ&x9���t�����0m0-'�^��O?z��bd���x�է¢Th2W�qy/l_�ؕ�P��>��j��NS
����T:�0��f���0��{xc�.*:������P;��z��[��g����ở��Q�/F�x{�~j�ZA��d���K����ְ��`~�Gc/�quy)!qX���֑��o4�j˳h,����pM0��Enϣ`(X���]J�2�g7������Oi���Y{�(��2��C��$������[��ye	�8��sL��Hv�`������P�\.F��ߨ!hTE�=�>�񠏓�DZuIa8=��t�H���X����i���K8r(��cs�l��D�o3m>G�f6�~����Igvz��E$�iN��YY��<7c�Ô�zF���Ȕ��3.7a��p!�$K��2ֈ�����P���N�0:�����]ӛ-���D�	=�7�&�(�q�	�9"�!���f<���A������I�BZ�qO0p��8���Z�ƃj�{o��~����������ӿ�pˣ����/Ώcා��:
�--\�r0��B�V]2�L&�NA�����s��lG�m,�V&�b�2i(�l"#�R� 4��^[��z�s�I;��1N^��Sn��7/��:!z^U��vg����Rq�3���Z]����O�H2a(�������m�6q���/�߿���ev���|��t�:h˽L��ы����sb����1y�>�l졃��k9��o��@T����3<�:���J�X)�w�]���|l���E��5�om"��G��>� ���]����:�n���}����s�fS�}9���@vJ�l1�K]���Sn>C��ss�FH���!~����j6Ģbz󱽻l[&EgCH�tT
����N��nle�?�����˹e5��	���U �tE�tK��*yFn����sY9∿���an�4\Ut}ScJ�$��N��LF8�8�97wCI@�<�z�38�0yX8u79LYk�+����34�r
�#�,P�d��4ղ�9��}�{��\$�ȩT���I2;N2���27nӲ���(�۶Gc/I��<J���<�?�3�Ј43]�<۪u�̑�� ���@P�ʜ,
�nJ�:�o�T/�@Hd��}�><�Ǆ��f��WE����$qƤkg��To�ۿ��'�s{���vpv�+�@���dc|����B!R�ML�����v�NK:10����RGl�����#�1F�p�t��N.a)e�y*��{Ua7d^���*\��q����L��~xy��Mۛ>I��w}O�{eVem]��t�,wB���	k�`��+G8º�[������1B��_����$+l�Ax����vO����^�U���9'+����^�2뗿�9�y��OMv���L�⣮��VE��Vn�)��)~��@H�+�S�����D��vqqa��u��vQ^�W�����kO?��o���(������w�^\����ݳ�����x�l2/$k���=�i�+%��"@?9ۗ�	=5�+���׮ʜ��-۫W����+�B�w�X��jG������������ V	�oo\��Rզ�����dz]��E �OE��:F��4??�P�B��b:��G�/>������3�n��C���u>w���r$��5M}Vz6�-c�x�	��QjI[o81� ��?�4�5�뒨\��XkKN`�Kv�a���·޷ʠ%[�Z&+��A�X�8����5���M¨��H���N�AcG|�`i%��Ap@�ՠ�̶#�,����mP��2+<�A��]�𺰰k�E�4��!/��c4�*6�H�T�y(�M�͓v%[��+u�QY�� ��J�T_QO� A�(:q��`�SY��V�V�>}j��<�l����t�wϔ�|A-+&���ۍ��>�������g��O=s����������d���~s�y��^�έ;w�y�[o�,�l!c�U�[M|j�nt�
J��dxp�q���,HNL�=����
l�z�����;�h�Q��ΦC;���"nx3���3�����^��H�Z�� �1a�B�r-`� ��o���О0�8mX��B}W7�m�\Ӵ�i�̾�졝t[
nd�uTPJ5���>oEN��Hgt�軹AKZ|[�{;7�V��������$����S����ީ$dFc��_ߵ��	�e{���<)|��6��t>��?������m�<�[:��I���+7e�c��u��1e]�VmhCWn�����MJ%V���������o��Ak��Y9aX̭Æ�Oh0���iPџl��d��PI�g�OM����s6��X@�&��h�qoT�z�"��&>����eϣ��t�r�50O��1�����oF@�֏|.ZR�AO?�k�QA�e�6��j�a�8D�m�����q��A.w.(j�~��)���w��P��paZ*���2]O*C~�L��6�-3�-c�3O�V�l��������	WJV�V<H%��P�ɢ2y+�+V\�h_7N��G���g6Ȧm�����frj��s��K���An�V￻u�K?}�O��zp�gO��{���ͤ��~�y�5�[g��07"�rp��^�UEX�/�I⡹1�#����E~���,�zR������jlr�w�m���Sۿ8����ڙ�d�Q�e�6�d��B4���l�*��&������^�r��k���i�JY8���MdO���M�zi������d�u5٪��j�~���Y5U4���L����}���eN=��Q(~g��X��?�e�ESYJa�j�R��zf=��.-@  �~v�����c+��={�����P�v��u�n�[����g��}|O�[]BA%��[������,��<7l��ܘ�0�w�qq���;L��i��V^����e��ũ���nO{���ՃŌ�'�S�q
��u�e�W��(��}�����k�od��bQ\`�)+d�xӦ(Ie���Unl�ː_"�QZKG/@QD�p&�,AO\�\��(�����b�F�9�H���̡lf�M�ƿ�B��C{���y�;�$�-{�FO�נ0�Z>d��T�
;}���y y�$&z�*cCEC���U�O��&3K�'�c���X(&V������N~�nml�SU��Rъż&��*�N\\6�/H�%0>1���S���c���Sq�KW����	¾�7U��ٜ��i�,�޻S���O���۽{��O�����J�7�݋ݧ���`���[6ҍ˅��R�����.L�bp�E��4��|�Eo�((K�	MJ˳��O	lL<1�`6;m�֓��mHi�^��|b���f賱֧L�
l7�v�&��vW��F�a�~_�
)��o�����Ll��'/����v|rfk���]�ز���(g���}�����q���@�ҫ���;�Y-[�Q0�x��=y�J�}ʴZ�lw���[ۻ������R������Ǉ���?=֔�MF�d�٭���E{�쑽x�L85L{�67%�������s`�
L�����[��C����ྮ��m�V��������za�^_�\*+��׼�K���i������٣��53��2*����W2$zNP��b��4ذ�u�V�xz����R�0H[�T������,��+�R&EO�^Q>#%W�����oJ��yp�8JWB��rm4�0f��V� ai��I-�x�S��w�d�l�R��^�zMݮ~Ǭm��l	n��y1�&�%���+��D��x���!1p�%��iT>��彾�_|#܇`8MR�?9�BH�3��Ԭ:q����۩���E��	u�\��C�D3�ǃ�`2���3���S{L�m8�Y!#�n���rI'���2����M&�y|�\��nm�K_}����O?s�������W����׻��%��ſ�x�1��APɠ�&S��M�de�@pSO@^wE"�qr�`" qL9y{s��"�e���xO�W�4�dl�6���Fт���~�n�7m=Y�).��;9>8�����5[��5�F�����>}bGG'��n�\U��^��h6�����)��������Vϖ� � j���H'��Ų��sU�Z��|6�fk
�B}�Rٜ����Sp��� �+HO��۪�Y:���/۳gϴЮ_�f�[[6��=�{�^�L&+H�J�h[Ud���yt�v�B��T��jkO�����v��#a�nE�@3E{��]�{����gO������n['�����i% ��L�Z��J$>�>_�̺��:}e��|��u}���q�Z�l��ғ1U�X2��D!�jp�3.�E#9D�n�����x��Z!��4��u���V�L� �����Lf(�Cp��*��+���\A)������#��Ȭ4h	 �f%���Ւ��Tt�O����WN���1�I�t���?�}�<�kZ<n�lr޴d���2IZ%�l�ꅲ��ܱjP��������:�/ټ��};l��G/���TA��%�9�U��!1Bb��bN��Ap0l+���V�Fe�����/���w?������T����L����ō筦��ܰ���0����b�}��nH��|=�QJ$�+��o���YR��Cn$YN5U�	(�G�/���A�&����k������,�tO*m��M��@DO�
K����4}%�^2��/m���:���nn����j�DN���2���틆Đ�ښ��{�n�6�bN�o�)�r�"`ϛ++V.�,��Xo2�������)���Y>�e"ŏ��P�L�X4��kkV�0��������+Q���^�,�un�g'jēa0��	p�HRYk�έqv&���ښe�EM�����/�X[�)J%M�߿q�޻yW|�.��sj��ߴǭS�ȑ�QZ��+��+��6lw��G��hHB�Lm��ٸ7P BuT>
�Y�5��P�W8-�\
K����[i�b�M(P9�sPjP�e/Y�ܭ�
{���	�����<0��~�28d�N��;�E��RY(e�P���:���b��(���C	�ó� ��lC0|=�-0�� �~7��|T-�I��n��$�LiE��n�L��,5���i��Ya4��$a��D�P%A�i�ه�`�*JIe;����ϥ� -�y1o�H�!��Z���abn��2|�����5�Q�}t�����៽��V����%���o�x�n��~�H��Ʉr�Ӌ�V��� iKӀE�i��.�n<dw�* )-i$��go728hX�7���_��fv>�ڣƞ=9޷꧅�����C�%�Sy�-⟺&���̊\�糱�_@\��-&F}I�<}�\e�c׮�fm�J��Ok����m������?�ݏ�    IDAT��sl�J��ԯ�-h9�Z�t�"�Bl��ן�ub���E�ey�U�^]��8hm�"e������p>g�L\�n��P�7��ڵ�i�M��Хs�?�MK����tfG�"ts0mno
��9�o<{$h,2#d�y������Z>Q���oOG�}��|2�pS�1=���tz��Ï�sq.!�ב˦��_�T������Lq4������C�P�W��]��jYN�(�LȄ2>���v������ԱoHt�}��s��ÓЮ#(RƓ�!N�)^�yώ�}|]�t��J<�%KE�D��dT4��De-��A����Ofn��]�{��NY��>j1�ʜ;`�U=��)j�d���C��T��׭� "��T\o����W�x��4�T��0DR�A�)�6ۓ�u����!x=~f!o�\�0iF��B%��'?����n�
�땕��������Sn��<�����c�L�_�.n��l�}a�	^��/UA
ٌ�֪��Y����An2+�d�7�w���ɪ��������}k�nW���@ے��Ɂt���oQڅ��I8 �����.��k�_��$J�q�X�f«�5/���L�X�Z�nׯ]��lA=	&���Oͬ9٣��;x.&��tz-SP�x��%����"�U>��vl�qb/����Œ�^�ت��	�x�;Q�΅2B��{~�g���
n7�w����0I�@j=ܤ����z�H/^>a͹+׮Z���W�3���'��t3.Pɖ$���7߳��!�ԜtD���G��`�u�|$��Eo�`�h���葍�=�����T�o�խʐ�P�����lw��j�a��g~A9��)n�Zm{��Lw�~�ǰ5$�*���%,]n����)<w)X?W�|��=k������ީo��E^����gM����#�L2�%G{�w�A��Pp���7����1y�l�WXܖ��(O5H&<��
HX���.�LPP�-"�y2�`���K�!�%�0��O���O�����I% ���AS*4�TJ��3Tq��1�1��@6��DJ�T��G�*�_�Ͼ��o&���o�H39���^��^�#O�J�����V��hj'�>
4��k�d�*�5 \w��E�^A	Z	�D&���d�:�<���t(�Dq��hel���/��&�.2L@��¬#��J�
��[��&z����Sm(��L�0�EE[�'�*ɤ��=;���e�e��;t��f����)��nyU<�Z��^*g��g~�{a/ώm�����<s��U��^Y���8�lzרp4�62f�"���A��:L�,a��]�o�ݝ�V�3ov̗6�F%f��ؚÞ=|�XN�4�77������.4����Q������œ��ݱ��{j�����u2�� �K
)�h�ƅuON��՞%F#e�������BS:���-�iB�S�X�B�6g͖Tn���MA6��ٹs�j�����n���VP�V����{�ܔV"�226���0(�@�n�Q�COL_�G��9�/ q��;8�����h���@;tR{ 6�+ý-�0�~n��T3��ϋA5NKcp������ z�ʋ���	{Gz{�Sw�S��h1�E��Nl��I �i�7�~�).8�f�Q��}�eQ(j�,!Ӕ�$��)2ⅼt���[=7�U�&��zꗯ�3V�aT�~�������7Q�����o|���$��{��p�z��� j���~!��hܳ� �ɎgpLK@C���ݟ ��H�i�G�"糺Qh\1ES�����w+�R2�DF�*�Z�s�k��d�V���d,��y6kyyZ&5�d�X!���r�j����K��p��˗�PNE`�k��Bߧ���w�۔we��%�̔{h��ȕm�P%R�N�����u�a�D9����K+ꉬ�V�m˄�Y�.t�Fۿ8���c�L�j�۸��,��߲'�׽��I_��b��7k��Ǝ���=;;�
�^iqA 'S��y2����u�N�w~n�t�6V���ή� .Wl6������yOFS������<?��GGҽ;��P�P��c�[[V�ٲ����x�(�eJ�``�,)8�)HE3ᐹѻ�ِd�B��|��2��@$��`���ܔu���Hg(Cxb-BB����xZ�
As����yp#�� H�L+LV�{��Kp��P�W����i�Q^^[�v��s��Kug�G��#R��rF3A���0��{e)�B��L�:��2�e<��]!yz���~�A�T%��u�KYe��+���v�˿����(pC~�޷��Nj���������u��r�W+�� nk+��q�����2�މ^�2�FzZ�|	��TdH�x��oJQP�G-�&�0`c�'��T#nzy<���3����66���@L��~r��5<�,d��JZ>�����{�C�a8��2�$�
,Ӊ#�	n(w�n(�rȣ5��  ��@��8 ��L�k�^D��Jq����h�R�g3N�W_$���k/Ϗ�=�^�R֡�x��=�C
W��ȏ�RE��R� jپn�Q �d��d�������3k��x��a7vw�R�u}���uϛ6도�ÿ��X��ֆ%�Ee�4�_�ۣ�Wv�n[�����6��t�R��U�.��^2؊�3��d�72M2y`M\=3c={y��Xֆ�&m��8s�5��k�ܖKWk���I��-�����Ջ JR��pp��\V������G���U��n����<���Y�� �i�hm�Z�
��0����� ���o�#����w��dқ�h�(��͞ڠ�'jGUk�čj���\���_x��?}(�7?����~�e�y�aK��[n���s�,
�fD�+.4q�H��X�R�B��)� �Ç�3��^� S��&��FV7�4F+q
��2=�I��_��-���E��wx_N�Мv��Ь���4��-k@�%<|6�Rz�B���gs�;�=�$q��']�&��	)��:��)1�ZY~\_6�.V#�	ƈrj0=6�g�ڔۀ�O9_�s�2;g�%�&�Z`�Z�)�`�l澱i��E!�3wK�.�������l&S]�ܺGG��+؝k���R��Ǣ������u.Z6���͇C����2+�n�k2��'��ϟڋ�#9���5۸q�ҫU7���ܝ�����x��~$�
G����0\����^!�$�*�G�wKJ���bƶ�u�;ۢZ����2�͗�c���<^�p�XJ
<#�%��⥠� χ�����%r�t糀!T�($#*i��cȒ�x�#����k����q����=R���F@=I̠ӱa���G��dҮW�>����_��|3�ۯ���/v��_��]����B�Gdn7�C0�-fnL�(����J��dL�K��ƓџNtJ��)�D	��Z9��]�	��[Ӊ,�Z�!��I��L|�s�@�`��Ef&g��Z��6����sH  ���V5�q�m�Wx�HQ�l�z�f�f��.�fZ�L��o$YXj�R�4Α���u����5�p��YRT3Q��($�+2�.�c�ϝ��]�$��Dod�Sl�&�5�;��p/��aZ	r_���c|?�#�����=4�l�Z��ߺmwn�Tߓ���ɹｲ	�2n5����v���=�1�~m��v�,��"���<�{/�˻��vc׊����C�g�M)W�5n���j. ������æ���e�8�:�| ��O�F����9�ָ^����/��9k��q���!��Ep#��L�$*�D.i���n��Czi�����we�P2(���Qr������8T�SoK�"�����4��W�!#%�-2lwl�i�`��YM��Z���W�����O�}�Z)��{��w^t[�*�!�Eb}n�<P�� ��` �x	ntAbp��wHi;'�Y������.C�s9e�}T:��S_dA?�HTQ�i��W��O��C/#��c@^%��F't������ד]�A�Q���U�?\�g�	���� ���"��h���G$�+�I�~y����d��?�e��+����Fb3@Y�u��@�Jd�D%yVp��F�fP�:�>|a��~�k��N�}ї������ū��ڼݲ��U�»o�{o�U�ot��b'��3d*c����3�Cύ�v��;��{E��?��=x �YP�U�^q�s�bz;��=�������p8����r%��:MNAHA��Cv�9_�VA0��ŀ(���I����q�iMj����������	*�B� %�IL�إ_���:��X�k�-`	Z� �yJ�4cŢ�F���a=����ٯ�=#��C��"X=&&aD��̍�k%dn�g��9�Q]���捯�������_�˙���+�ɇ_���<�+����^��
n@/<t0_��Fp�8_�VZ����$*b�R"�SvG��G�o4�U`�M\�%��ZɾI�pSq�̐����দ/Z�����m��ZY��!��g'=3~&:Zj�� �R>�Ұ�>���1�]Dk���`B�h]'}pH���zM����QFb���UpKӌG���1��鋦�I�.�!��ӐԀ�ޤ֦�_E(�b�/��S��������(��͊������O���9�Q��]���;�{�>s�m��v�����O�uz��-س���4�����{�_\���Ͽo7߽+�>����c�F��%��l���k6+ᰞ�YƁ����:���+٥?L}�\�E�_��$<p�W�3A�c��Ob�X���=�p�}�z��kn���Y����t�	Ϫ"4�@�,�Ḟb�KҸ~����D=f^�1������E��bJ��g>'TD��M=D�<Z4��q7Ț�������� @J��;b�$Q����e�vce�[�n_���}ǟ��B������{���^b������}8��t���̓��J�H�U�ג�� ���Ybp�&�nP��\.�7dqN1��`/$��θj�^%�[�)J�59���P`�3e)S��ēe�+�����\jƬ��C�CH�lU�y)�����]�pJ�ᩅCp�e0!��P���R���F��oi����%����7| r*�ۚ�G"��r��@��B�w�l̠������"���e��n�l��{B�^�Au�`3 �V�����疄r�HM���[��}|f탖��ֿhJ߂�`L�g
n�Q"[>ew���v�;޳f�o�|���{��>>8��0�p�nZ�Z�I&�iZ,K_�ܔ	�m�33��,(
4 mRpx�@�*��R�y^�F��$��	�6�qd��� ����$s
%�4J���*�r`:�gnq»Ȭ�����%ʕ�WC����дN���!H�
K٧$�F�T�x��v�&Ke��h�-��AIK����&��	l�V�R7��<s�ƻ�׾�s_��O߷��k|�[�ѯ�L����x�m��L��<d�p�_��m�Z�M��-�iʨ��S,N�����!�r����!4d/�� ��wA"�=��d���,0n:7�gt��4�r.�u�	�`Z�Ҩ}���E��҄*�I@��CEj�9_.\JB�GS& B�M��W�en�#����1�dqp2ҬE���{�R)����c W�����%�@��Y�&��ܖ�Zn�Ә<���3��b�0n\��6<:�D�k;+5�������Z�ٵ����:j�Fß��i�!5�'�:J�6ϧ���������Q��۷�?������֚]}�m��G�D�@1\h\�&�y��X�A�<$��kǽ'���t>�L%��k�S7!v�m�U��*�82]Jϩ̓���#~ͳ/O�o�<�t[C@���|=sM2���J�޸gD�Z�u�����]�{���� =�X[�[�5Fd�.������!�ܘAƌR�W����8�dճ�S�X��LY|��l��Z���ۛ[_�����O�����[��}����Ѵ�|K���2����� }<�X.����U+=zI]�r ��8�Ԋ�B��>=��s.8�+>��&�JЃ#������#HH�؅����b��喔fy��3#"��x����M��Ұ��׬�b�.'��bZ��`�MP"0�>���K�.e�Bb^�e
� �G���H;\�C���Ү�e�%;Yn�<�&�9��X�Bh�G(L,a�����=ٜ?`�0M���wtj�W{6i6�F�n��}Ǿ��w�]?;����5�N�(l}7hq#�c�O�jEKW
���[v��M;h6��)���;�V�n���6�&m�v5�jy����o*�tA��I���I��Jls0��7������u�� �5� ��*'�����F�~j(���m�����O�/��ƀ�վ�ղ c
<"ԇ����1X^քQ!��!�\�f��&��7z�E|Ո��d*C��+�b�Z�A�x�$�!3��j-���B���T�
���z]�6/�yrf��Ȫ��frv�����/������܆��h��.��^�i]���c!�fc��V)[?�lF����m,����JY[8U"R:��:pCV��6������ƿ��}E9�M?b����22�%h(��5fz��U^��Q:�9c�L�\��3N�������Q�,F��!��{t���S�#��N�O�`�e�^3?���"�����`1�)&�l�2�� 	�u�^N�dY�Cb��)�H���3;y���ggv�Z��o߲Ͻ��U�%kv�l��Nl�ș��6)�MFC�������m^ߵ�kW,S-۫�c��o߷��{`���77l��V��!�xA��@��b�L~U��J��~�2���A�L`�`4�X�`4�π���0���9�B4�t<�y�sܴ�CSeY�S]�1�����(�,0�����U!�����4�X�4�����Fp#�f�E�a�}	ؼ�>$>�Jh���Gց��� �X�|�2x���Y��N�VRܣ}��J�$�?�ҽN���;?<�$�-��5n_kc�K�{~��bL����c��~���<������'��=s�M�Q����6�v|�\�Z�l�\F���c)�pbVG�Q�o��4(�ˆ)���nUl �������e�8�W��IF�b
�I�.!{�Âۢ���~C�;�|D@�� P��AZY��`26��K�4)�1�d}���O�FD�{҃���
��g�u<4�cpW�ʧ�-���侄���_|*K	`�ȜC�\_f8�a��Ξ�s;��b���\�woݲ��mˌ��:���k���l8����ӱ�77�Ɲ�v��Y�\��;<������gr��_�j�wo�����d�Mh������~D��&��HO�� �}�@bK"f~����ʠw�����L���<���±�&{�)��*��Z��B_VW�G��<_>�MH����߅��⿝����f���2�K�9�����2Xv>m��Ot�f��>��=��c���.g������&>1�9z����8�����p�W�{����;�������}3=��ѷ��|6�GG��_v��-���7Ce���JE�~��Cp������N'A�8��P�."�aI�A,��5}2��p_ �f� ����6�����GMl���&����"f.ң���� F�C��c�B���+B�zk���%6�>`n8=J��5Ђ�LB�t��K�j�ZBp�%8��{!�r-*��n�\��Q��3��%f�.�,�2S������Ȧ�d>mw��Ş��,?��nm���ݵw�߲�|UM}TB����8�a�e=)��Vm{{ۮݺi�ׯʆ���P���������Œmߺn[�oX?�SdD?)�����a&�9���#鵮��'�g�{�ed�� {aヰ�����M
��F�GhDI�0�Jk��t�z�/+o�h@�:	�i$�+P�Q��奷`B��:�?�1\�(Gcv.�Q�;�|��L����^c&���{�o%�0�    IDAT�����NK�{9���h������Cѹ�gg�r��{�������o�n��������{(p���Ϟـ���	n��u��I.WH�sٔm��(���(K!ד�)[�	��A�a��a�-���&%�/)�.�C-��K�-D '@ؿ!_ȱ���S� ��)�`.��ʽ�3#��ǣ>��7�`x�8���<FJG��E\�M�gL`�Ld��fR���?�l%��)f�
�K�����׵�	-���i��M���/�P0/�9.��Ѩ3hv2�~ߺ۸ѰJ6k�k����v��!-~�A�ٔ9����t�v��X}}�Vjk6��%��t�Ց�?}n'Ñ6�m��v3	����y�h p�`E���@�0��x#��ǀY�1.�4
&h�+k_�*p�5qV�^��K஫����{�漃�cOX�����cЦ
tSX)����k �F��dv���,��'�'y"L��^����ơ������A������TZ3_2��ts����)�����р�ZK���45�~���؍���wW�_�����o�~�k�}�b<���Q�Ͼ�6l���_\s$�|S�ꕊ�d�M (�5�Iצ�*24a
��%���rOA�gR������)C����?i|\\��
���@]���E�QX�(��M@�c�"��8�
��¦���E���A�}ye�d�Jz�V�-�A�����M����cQ��]Y����(=�ˁ��#JZ/eǱ$�����6�g�p�����	���+���*1g����u�ʒ��D޾~�n�^�+�V@�+�p��WKTB�=���Ɖ=y�Ҟ�|a��^�)x�\֪�;�~u�*�����1cc�C*� b����db/�R�B
o�>��a��u "���C�i�(���p�	�(V�}f�����KߌCl�8Pp�wy@ꀉ�~i4ٙL�Ճ-�R�Bo�C1��lKx���ˈk�ZY�f�,�c���"k�~ z9���	h��%^&�6
b�>:�+R\"Y}N��CA�2Y�����L��@n�^[�����?���������[�?|�1������;g�n0�D7��V[)_���
�i�0(����?�=7q�B�_g,CC� �:=�������U��ei��2��9u*������,��!����v,P Y�g�B�1@N"�1�;h���Yc��_���L��Q4�q�� �Tt��8���-�/���%a�*�z����m\_���w	ЌX<�v³
�zra
F�IT��u��:x� �*n*���e���H���kW��΍[��Yw叄����|��O�2T����e�DS�\����v���* os<vK���������+�'����c���$�"BVM��Nc���B�`Ʉ�ҍ2k��.�l��=F�o*%��{�\B��D<�*h �a)�r���_)[�a��Q�(`��P��e���
�:^z3�->�����Q�Őt�Oh������~	�!�f1N�I
�풵��!������oPia>�
�M��Z�xxgm������O_ύE�;��9w~e����dn����g��T�e���)[-�4-U㑑5zN�U�%�E+bc�o�(f��i�J���ͣ�E?�Er�CRf�Be1޴es������2�t�f�hQ9�xh�E��)�xH��<<(ʘ$���(A�D���IY
�)p27Jt�^�Q ұ.], B���o�,�`�E�/ �������^���q�
�}�����̘Ž��-�"�/��>�\��+���<8�&�Ε-�zu��[u�y��|�8�B����� $O���
n��"PY�ش��W-�|�4H��/O���A��z�[>��p��t$�F�����@.�������@b�r�e�@BPQiK=�el���d��9������D�_@�s��S�Lʮ+���P�v�-���C
�D�)E���?������C\!��+"�ju��ʩ�3�P�K�zAǋ�"���}�kI�+��̞ܒ��K���A����2әU�YqKo���nm}�o}�_�_�H������t�?�4�E�̎�7�S.xhBͧ��V�Vv(���s}��-l�� P�<��c��ʦ:C/B=2nZ֋�<�U��K�?��MҠ����4��o� ��G�
F�yd�L�u.�� �%�SS���=�X������&%HJ�M"�$�,�4��zw(���*$�45������Ri�����&z>����������eE�/���@#�$��0��f�a��D�)�W�Ҥ�#k�:��}\�mkc��;�
n�ٳ��m�t��B��	���	����{2�)Wk���mk�ۈzO7eγ*�����F�G�CF�+}�{dݐ��y��L�1F���Ñ�;=yAH�k�'FP����L/���V,S*Xf�$@1$��̤�t(-�]��׀&LK�n6���Z��p іp�\ē��Q��^Zڃ��X�Z�	�'��Ik���8���
�A|�6�7V´��oCG�Cܜ�+ /\�%U����vvp�~-&�8�ߨ�������������F��o?|x�h���G�������-�*p�/�a�$E �����Ven������
S;�T!��iq��)W����jn���.M>PXj�Ƒ:�(o�_^�sC�� ��Ù��*K������~hDx�rI
�\n>����F�q�$T W��=E�m�'P�h�r?������o�qPKe!�z`���J�B�/e�
1j���@A�1�8ڏ�M���;Rsh�Ee4�%�8��xb�k�ڳ�鹭����ΆK���1��yhzc��Ȗ��e�Ik���CM�ʵU[�޲����Ҧ))�6�٫����.p���ۚ����2����[��o�??�n�-E�v�S�YHbǁ��v���:_]�L�h�k;
�����R �\����?�.l�D�/�}Ե����b���5��o����Q�\88�r�>��W�QkE ��¡�8ߏK��װ��W��F��Rp������M��w�C �g �Of6���Xx��t�Ꙝݨ�?����տ��~�y#���ݻ�O~���ꠇo�X8#` d����WVl�Zu�����P	�-"��8ʝ����F��Z�,����zhQ�%6a_n1P�����ˆ��X� ����Ұش耬�H���}�:pbȀ��p�7�-�0����3M<#��ņ
��"Ǿ���=Ì �8Q^d`l�n����M`��?���D�����g�1���U|G��,0�ܦXz����liY����a�d.E޳����׬vu�V��,���X�i�&>,Io�Xd~�_�:я_�۰;���U77�0͂��*�q�(�QZ.ʦ��E&g�E&�x"N��G6j��}xj��@" �R��Ŋ�rY���F�<Me�ݮ7έC�/�KbN`+��Q:C��3�	YSQ������ x������Q��eq��!�8���� ��$��}R;�"��z�6&���3��5&Z�A�P�6еbO�nB�Z'\���I��?�,�m��׳���g&[�zV������_��?���LY�����i$���p��K��~�Zӑ���8�K"e��x�R��ZUcp��h�3�rnd�u�s����}7��!���[���B�%BA�C��=f���s(Y���r��l��*���k��ظ��)�B��
%�f�����Z0Xp�鿂CP��2;�0��>c��Bv'��^hRD5Y@T�K�-�L�,s<�x�%W<r�Or[�=�@M�����W�.��@�D���Ԕφ��pz<��ށ��ط�鹭��ٴ��
�6v$-2?�9���RM�X�4e�/����+���kV�r�V6�%�I9:I���\��5�C�>`D�sh�3�
�9I�2;�6[�?���E�*�]��Y�#6�J�ads6�~^%�Ս�䘎��i���Cy�V�r�Z٬�N�=�M�6Ce;����5�eb<��S�����A�
Ce��{lj�Kn�:Y��L6-�2�x��h���M�.�z�ڇ<�@	n�PՒ�[ƃ(,���{&�A��&M�#�8B�&&�1�����-i����9�����z����?y������K�������IDs5�������p�y=��܉�R��O�tc�2��SϘ�)Sa���?(���zm����Η�S� ��uOJ���QElZ�6�~e�z"�`�d�X(�;�t����R�$ʀ���XP�6�`��l
T�s���)���*>i9�LEb��P�ohH��B�F�r1��\:�JT~٥z9NK�i]
�Ll\]�8:�+��:?��:��ۿx�o�W689���u+�lXi�&��<�� ��l���,� w���"��Zmc�6�]�1�����i��Z& �#OWc;z>��32�.��	 �V׆gM�^�,��J2m�\�n�����3o�ֺ�} \�C:m��TϹ?�E�k����<:�g���G�3K�3�R�&]msݲ���������鵅��Ӷ��NS�̸�
���v	�mM�CpS��χz�J2����r���r	�F�A�.ZHA��&�|�c� �s���N�@�t�2OhX?�|Ђ��oY)���b�j���V>ڭ���/��~3=��x�����ˇ��?��рi�gn���R�EP[�,����	���N��1�ի�ORGb�Z>"�'��h�bAh��S(��R�`�� B �T����A�~ɴV�HȌ�Y.#g"1���-�Tl"p���K.�3u��c�8���>b(9�A��AC�u�Ӝ?E
���)�i����ؗQ9A��~��	�JV� �� �d�:����52 �P��4i �,*Sڵ�������d�\��e%�S6e#�N3�	�Y7qh<�0KI����+;z��f��hY��+�ו�����9=����F��
Su�D4�կ;/�ٸѴi�mU��J5{o����ڶ;W��Z����#��Ƴ�@���T8��hl����N��H������;���V

n��U��Lz�Ҕu�lH��x���I �j��
 @Č���s ؾ����d�RY�a�Y8��쇣��9T�s}3��K$9Tj����e�� t��1�p�D��PYiR�e�T �N��TZ*̳nOmx�7d�7�����������)K�ɇ�lLz�`o����s;v�5C7ߧ����s�9<7����@-Z��ďL�d�@�2D�X�.��1Ê�S�(<Xŉ���Xp��/�'����,�.U_��
��4�tr�ƭ �.�G0Ҵ��	���|J��r<�%ϕ�e�(A�`Z�97�1%���2UpY��ʢ��	JQ�
3����d�;��C'M�Y!���7�?k�/��w��.prl!(3\
n���in2��љ�2�<8����ֺzf��Fi7�v�L�Ge)rn�T���徂��ƺ[%��dI�vc��)�L��B�h|2:a���ڴѲ�i�2���Y߲/ܾk_��m�**M�Aw���1�\�q���NXG��L���v����\��t��V���+�ʖ)��3�\�,�a�x;��]���שHS�@u
�X�&��M�B�_�a6���-�G�3jé�;�"bq8�Cm��co8������Ak��3���Xդ%������2۴ӵA��Vsy��NӒ��/��̗~�ߏ~���,�ߺ��ab�K����?G�wam��S��T����JE�W\�[=9�S��A�#B���=�%hT���b����z���e<c�iX�����H�^V��Ȳ"4%Ja�}B���??����)fNy�|rm* �����$I����"#y�e`�$|�[�f?|�@�T)�˩O���BiA�jv���:�^�/���Opk�����H��<�Q���b.�kl��Ȇ�9.�b�dqjf���	�g�Ⱥd��{ʝx<��e��a��{��?�B�j����qmG� �	Ls�!3Ar6��,���utj���*��eW+���!��>��A��L�ik��hOe.�M�
�������Ƕ>I�F*g�s�=���>oo�\�N�a�'�"�c�S-����6K�,�8
�ٜ%s9ktZ�vf��_��q��:���
��5���-_)�Ӕ��S5�=�:�.(�(�
Su��z��!N��^������UAɇG(�q�k�Ԙ`�׀y��uE�b��>���UV8�n%g���Hi9y>t'��`J ��2��*8:Ɠk\H��Wf�<	轒��F>o�d�6s���j[_����!���x������G��_~�:M�.��*ͽ����W�@A���F�*��D|�Ȳ\~%�2�i]q/	$�`O��+�[�j����7?]P*N�TN�t:���?@%� '��q�������G����
�|κ��BbH�=����^*���.��b�J�L����^6'�9����ﹼ7�{7��:�����r,�EIr(%�5=v �C��(e�_j�E���BH���R�'1�u�O�}�PZ]��+��DPp�i��+�4��+&�)�}h�Mgv�w`G�r5���Z�VR�n�NY75�)P�� P���(���>��t&Չ�Y˦'��~�gW�Y���i����ݾ���}v|b���ey2i���]ͦs��RE�Чٌ{��X<����+;k^��yÚݦ�Ĭ��H;]��?��#�w�f��R�2{�#!���uf���P������epsO�~K9̄��[R �h�) �������e������89ȓ�%�%�����P���H�����I�o�ߠ�i@�KF�"=P�z�yBÄ�L֮���lm}�?���pK	n�I��mn�skL�b,7��
UP���b�!�6)���H�W�'�1c�1��x�pɿ�ZZ��%B|��8-�O�F�F�߇<�N�y��(���P!�#H�?�pX�|&�y	�T$l"��`�K��OT���>�.��y�g�k��ط�e��L��B/��X΋?�p!�8e����-�=zn���[d1뙰p�Y�K�v\8$��-�Q�Nj���3���9�Ȟ���-9[���N_�[���V�׭~m���Rh&��q���+������+k� Y��-�ZR�6�g�#��gY�:����U������5W��8���6<8��q��*��w^}˾��_�d(�c��Tr<ku���U�%�� ���7�������zސ�j�Ӳ�V�F@D�vS`"�T�l;�SPbMh��l2R�«����	�XC��$��f�^��0�CBa#��΄��(xQ�J��ɡ%aWS��6����:�AȪ2��9Ӹ�J�
�@�8H���5�ւ�:������j�w^�θ��}t"�[<K7��^Y{����/}���|x���x���'��st܂�rd�s�ep��k�m��O{Mb\)+����=�8���2`�t
���O-��?z�"q\�`�;�%�W�b�*M6���6��1��2D�J�(�%ˠR�dAfH}7�SL'ɘ�
n9>I;S�^��<
	��V��[�u�qC�q�<c��:Qf7��l0)� �� ���x�r���` � ggS�>*�i�Nl2�R\d� �$!àI���@��Rޫ$��R�A�)L�
�Ol�^��[�mmg���senP���2 �Iijbv�����S�y}}�*����n�(�i~��9���<q٪����/Isx�`l�Fӆ{��k��ݱ/�y�n�n���vzt(sh̎��u��Vk5����� �ƕ�S���	i^���hbpb��s�6Ì{D�S.m�lJ"	4�a�`|L�C����5�]*�� VI0+b�]�I9���*�a�Y*�-����?�ˈ�J;��M��1��d�>Y��<�l����S���tgؚ�̥mF�W%��Fc���$ ccVD?ήS�!ӛ���[!ܷ��xF9��&����,3�[�U(�
��������Ko�����ݻ�N�����1sk�'2~��Q�s�Y[]�y�-��1�ɍ�q �^�~�i�ȶ��E��d���    IDAT%xǲzO�� ��zX����ô���\��c�M<�CL��,�2B
���(�޴e�'CM��Wd��I+��V�:O�L2$k��7���m0���)䊖�h �@RtO�D�ol�^�� &�W:m�NV,b�H�ޥC�(H&�7�1љ���h� ���NF֙e�,S�ࡊ�=R?�}�;28�%�pe�A�]��Pr��,㩥(�)�jk  έ��e�+���4��Ҭ#{�xi��uq������Փg�B�W�l}g[�3�M@�rz���ax�b27�	��KYy4��ѩu_Y�ٳ��;�{���` �/^���
E��*2/��Z�^�r��y�����Z�߷��3�h�����:���_<?����G����+d�V)t�&���3�W����1�D%�Br�(�*��e� �^)�J��k*�
zO����rYK峡A��A%a�t�JlKkvX;kw�9Zk4�TK ;���ƛ��)��V?.���E�MK����Oң��d5!�9�١D�C�	�OC��Pb��T�6�y������ͭ/�ܛ����\k���h���g�$���t��dgSvk����rU�8� ��pWS4�2T�@�K��EI��[/27o]F�c�fC�z��^B:�z�8X����(2< L�q�,�����H�f��mVj�^�Z1���ƹ�5,X��������U�y+���X6�'�	��U�z`����0�$X���W�E��8��TFY�;H�3)L�7,\�F�N�6�m6�>�w�5H���ײX�"oN���o:�b����^�&v:D|�&��@��o��L-75����N41,l��ʕϸ�t �$�x�"�Ϭbi+'2v�乽|�D���zݶ��X�ʦ�)� %A
J}'-G"����L���y�f�A�p��Ƈ�V�������}~��T����.έ�R�r��u])�ʹ�����JyŚ����G�������ҧ��6�ӒL�8��e23+p8%R6L�6�J\Z�U�>0��T�I��g*m�l�j47�**V+���Rԟ�H�3����>���;�Ǹ�&�@�&Rf��#�h��E��Z�ױ�f�·I��(6���l�d�BQC�d�ȇ�VM>�����Hj�)�L�>�We�ʰ�=k@���
ȋl�n�k��޺��?�?-��ڿ.������ÇW�����p��+O�'��fc��Ƨ���e*�mu5dn��Ud+D��PS���� UM�X܁�A�Z.G՛����g�IQ��
u<�x�OqA�5$�p$�lz��1�!��܂?!x�:I��ɰpߞά`�8i��n��������t58`�II�� 뢔�4NuE*��RK �	��M�f!�������dp��"�^(��ZD:��\N�R# �� ���U>4�=���"���:ӑ�㛣�����K�u�r�E���>��ٱ��^�����\���əӯN�mkk��;u��3��R����#��k<��<��~�8��m�붵�c��d*K���:��IFJ]�#��;����a�f�vr��Ʈ]-�X���c�i�T��b!��<��gtk'�����8<<�o~�=/��A+K�Dq#��M'*,M�!�a�+clCx�T �=)PAd,K��y+���5uK!�V�K�J1g����V�V)��R��Z�'��"��[�=�K��!zod����Zdn����{v����E�Z����c�M�Z((�3��\xm�B����K9�W*6�g܍\$��p������x��`s�������QI����;�W���ߏ����7���ۯ?x�s��݃A�=i�������d���y�):BA(���D���U
�B)�K\3*�/�@���ר��k�ޫ�}9y�����8/w��.�
$��r���q�Jl�ғ�{�f�.*H�3��%s�C�TɲVN�l5Y���v��i9zOé{]��V�笐-H6�EE��:�FQ斤w�ʦRҠ������[��ݨ�SsU
�tk2E0�8���.U���tt�P�AV�i��:}.��%ď���=ꫴ �#���q
����M�Y�1�zt>P���s���Ȅi'F������i{w�j�V�׬G��7��9�!��:[afVIe���{�̭����k
���\����\_Ӿ�=&���6h�1�[�շ�q����Yݲ+�T(�J�C'������+��ʦt��
`�����h4v�޽�lA�
%2�R�P?�Ih�Q�F㞳HT҈�f�8GW�����w�r\-8ZD����I%Xo��Y����r�V�˥�V.�m�\�|!+s9t�J$�� 6����l�T��L�?��2�s̳[=�����`]�J��%2�w^�-W.�k�P)Y>���}1c��$?�i�ܚ6�f>#C�$�t�`zhhTL�ܮ��>{o��O����;Ϟ]9�������?m���_�X/��Q�T���b榆�z5#97qCT݇M�8�����Ş�ņ�ӯ�\x/���JQ�6� қr�4'�z"t�u�?���(y:;��f����P�w��A��6�aݞ��
��md*rU�(T����x8=���ɸ��	��Kf@#f�����E�o�S����*��	�v�c�aϱB2�ť�UW�`^6w�\QpC��+&xm�,F�ܒv
υ	+Y���Tk:��^�.�;"�9�1zR���Lσ�I�c��
a~<��{��5U�n޸*U��q�� �{n���wcZ:���v���5�Ҁ�˧um�9�x��:%�M��sj����gM+��v��j���3�.U$���u��m�� ����D��jY�?�~x�fggg�p�`U�#ę���LlZ8��Mq�
�|��)9������AL�)w:z��E�O4�LNY�?�Y9�}��N{O�TT+D�R�9�N����1���|no� �m8i_��3�&����	fꕩ�
A�
@��Y	\��
���W�V�	��r�晜��A>m�b��oy�yd0�8<9V�Cp[Ie�����w6�����27�������Y�,��uf�\J��(%�Z[�Z���$��G?aJRN���WI/%R��r/����R�P��!��`d~%-$�����@�9�>���d��h|�r�)�ԕ)��POe�Lp��,��m�PUp[�V��
�4��P��B��B:��Nw6*��� �ٍ�OK9�CZ\h�y��E#�0�0�M�~O��6Q�(�v�-�� ɩ����\AGc����c#��U&�	)n�w�-�Q�A��sa��s��۔����`�MPSF��")���������Z���a�wm�����LuY'i/-ūM�\(r8մ�a���g�o��-]�@��B�Z�0�lR)��	|M��T����<�v�捖�[�NV���&��Pxr���g ��G@��Y�^�oϞ���Ź&� �ONN���H?�P sJ�{}�ӱnD�=5�(p�="ecJ^����5���pZ��%���(q�)5RR^AV*�z�E�4aʹ���B 0�eq�6��G�Ɓd	�ѝͬ��e*7��G(� �r��5�	V�j/ŁP&���z��ڊUkkVZ�Z��f�"�(yW
�^�[;�� �I����*a���!�|%������ln����s���HY�;��_9���Ѹ��=�4�7܆4f��i:�(�M8ͧ|��IJ�IK\�e��,8v �#�	u��]["�������\��$��Z�Vx�8�2 ��)e �G0%ԟa�`&ʈ��
ɤSi+�3*S����T�6
%����V�E+1k��jڠ��b���ɺ�x�M/D�;���S��dVx7M@�Ы	�5-L��Y��O��& /(\ɤ�2a�8[�����$=<7l�8�.����R����%5��N��6$S/��un�A׎�m`%�i��2D>��k@��3ff��#M;;Ƕ��i;��Պ���kM�
n��s��GSKC����=}n�fG�m��U��^�Y)��8J��1?S(zzX�樯�ĝ����Z=��]�V�mm���D����&���� �wi!PV��C��N��N�N���T����3!��Y�wB��A84��L:'�Jyɿ�%x	b	��1<�&�Pt�R�ϓ��lb��X�nR6�-QR����2���O�h*��dB�}�h%3xg{ON4�OV;jED�<�IK��N��0��?�ڪ�VQE�X�T��j�:�������u��n|ur�-�TƊɤ]�֟��y�������	n��v<��$��ʎdf���
�`�ŀPe��j�:w�#�WC��4�4n���X�JF����B�Ʀ	�:�Z�'%W��0S�9i�Y9����\4]��jジ>Gb��BY���z@��np~�PZ-���m=[�j:oID�#AB8uz:��EeN2���H.W��i���F�֌r6��
��z!���@!(��^�0���GV@��W�^�i���ܸo�L(��NOtP�*�E��|еT�h���m޼���������Y޽�y�s�]�]�}�����&G��(��Hd	%�%(����A�3E�8XQ� E"���>>=5�y^�<D�����E�#�J�]�5���Z����s?���l���0������S.R0�)$bJp:����l
oNCq\\i{oO�z����݋������7A���z^�x�܅���:y�R��Į"���v�*�̓��
�����`}�V�H~����*��\�uF~�r�^�B���(��=�&�O�4�M��<�^_^s�[��P��7��PI>C�>�&)V��`Z:�8��d� �`s�����<�p��7�R�r��v�f�̦.�\����+[��ёZ���p�:Y��{�7tmKMaF�	�/�d
�عqbF��;��0=1*CU���A����*�*��U�J��m׵h��F͓Y�hp��a7XE��v��z�l�|����������ڊ[7����ɿ�|p�{޻��2(�mx�6��j�N�|��Y���]��z�����M��"i4�j��p�$ܴ�.9�eY#s�p��_���V2U�Ug�<^B�l�����ڬ{5}�����ZW���>�����tl\ J��+h�^�v��������C��b�?�I̅�Q��ظA*�ڧ�ډ���Id:������֖�{8����gKG�2;��Eȅ-R-$`�aC�!����t��	#�ƹ�T�����/]�V����T�ZE�J�7���+s���1f S��>(e£�/Ի���ޞS�_��+f ��S-T $��@��G�>���4M�
���j���m�c��q�ύ�ր<b�hWo^#N!��
k6����F˫�r����E�Sym��&��~��E�G�F�l�.�8���Wn��'�l��0nbĽYKՊv���l�+���$�K~��w�M.r�-8�u:�D'G�;�h=+5��D�����ۡI`�Yi>[j�h<Y�uq[�5烿�I+vN�o�A�����*`n���.eyy	����FGq��)U�ʗ�~��V�ZE����2��&��^�z:�������(2���v���_����^[q륗�j��e�p1U����0��e������Vf�pAc��ѧ�`���J|���IcĴ�zt{��W�A���En:68Q�:���v���U�蠒�2�r>�Z��� ����N{]�&#��b����%��FL�- %�wXRg�-����5rZy��PI��+Z��-�`#�H�8���8l�ӯ�$"� �=_B#�> � Q�5�E��[0�LrF��j�>@uԍF}0ٔ�].FnF�ӫ'cwc�N˧7d�|��q���aj�>�ijm��@����/��g���w���:���˃R=�͚�:(��ʭ�>�?}����p��Ζ���U��xc�g�.��U�ͻ!�d�����%�':���n ˫[=�������խf��F��8@������+`h�����y��&���á�D��w6���JV�%U!��h��3p���]��[2<����<䵔Z��Ȓ�b�k��ťJ4b���ឤpZ�J�Ɣ5���Қ���.t<1y�bF�-7.����@��:D1X"�hOVِ�ˢ�[᜛�r��<&%6��RU"�'WT�VѢZQ�U�׼���/&���OM����REq{g����O������������/]-ǿ���&�7��G
��V��v�鋂Ԧ�r�غ4�(p�Y�=����Qqta�0;ڸ$x۝� �~�A01��\^;����5��E�kt��T`�Z�� ��[��GR<��n��3b���*W�,��кQ@5�i�)�\�)"A7Ͳ!gAζ��r��~�:�~6�o{�h�c��>�К��Y<��d>t:�R�H�D����8�-y��DF�]���7B�"a�1GFQ��c3��sC���M�6�az���)�kTUh54-�u3��z1V�Q>R3��=��]�������7���k������G�a:��r�m2:����3M�5�;��s��>0��^Ӳ4�Ʊ��sc�DT�&���B�ۑ&'z\mbi��٥�X�.������L�9�6�n'>W/s80���!z챽�/���;+WJ��:2N���*��>&PQ�x^���!�N�HG/����`L8�z��z	��-}H碸��c�kF��,5c<��Mo���=d��`2�-����xj#�2˥��5��i��,�iV�J�R�r��^,�SQ��P��ЪTR���fM�jN�ӡ^n������\*���[{�?�K�k,��~��Y�������٣Q�{��۟��Z��{��߁��'#�z�&v��
c�#��Ŀ��]\�J���YT/�	s����c�LN��*�ݯ4�](i+_1�ݝ�O��bͳY- })pZ�r8�y�F���E	�M�RQ=_��75��H�r����֬2�2 n9#"xl��.DAYh<�߂��tgA�:.F�N|:`:4�4ِy���b��*!�Y�<��{�h�����I�T��
�i��E�S��l9�6��Y20n%Pr'�{nl}�]���U�}�r�nS]�z���b]��:�D��������Q��5vw��l�A�ơ��J I"�7�N)�J�����?�[�ၚ��%h�Vt�ɖ=)�v�g�ǸeHJ��lb��?����딚��zG'�2JӜ�G!�L-YJ0��&v��H?_�ͺ;�`Mŵ�8F��QrV��$ �֖_S��9U+Gbfh���	�3F�ȕ�����ɩZ`A��s�Bv�N�Q�8}�QU�VU�k\1�l��	��L:{:���lK�T��ӹƣ��l����nG�w�'S4�ge��p�Ԙ	�,�5ꏔ�t�)�0*��ރ|��r��FkK��m�;��mwpjT4�t4��]��L>mX�A�u����?��~�����ҹ�_Ϟ�],F�l��/{W92�٥G Z u�Ro���o����)"�î�ݜ�lt�.�}fcd�ZG�[�K�CmtԵ�<NQ�n�*�]���	=t`�P�꛴�rE=,V�����ZÂ�'I�[�������`���9ԟL����M��`n� �v��ra�{�j�|1�1_	��kLg5��5����bv�c`W�DN�E�|��Ä��p��V6@a�׆�M�����8�1�-["]�5�;:�@0E� ���.2.��*-��M����K>��nW71S�f�\�> |��U1����7C:1�/�ya����y��;�L��g\������# 8*���Ͽ��O�i9�������=s��)��V�E3��\踾�S2=�������L�5��ղ7�Ÿ��fk��c�{}�Y��2���<װ�2]'檺�`KUx��
����h������?�	<�K���F�������a^ʶ�XP��P���|�W)�R�XT�V�v���V]�FU��}A�$��~p�裯8|����58��-M�g�������uM��bn������ڑ��l    IDATF�"J|逧����?�tV�JE�ZSͭmU)p�;ʴ[�4*�I�t��ߜ��g+���A�����?���_�B�+n�K����`0���d��rz��#}��;z�sߣ���J���Y�R���c)]���7KqC��
��@�����3&Z��d���+A -@ҿ�+�l0��9�z�.�q��7[=����3��y����JZ�rʔ�.Bto4p��؆���-�%��M|�&!�^ �}7��=���0bXL��~���;�&H:�``ƚ�1=������I�����1�9P��xQ����r!��^GRM��_��ō��OA��KW���GV�t��hc&r�,#W���6KI��T���]�h:s�JaoK��{.h��"�����y��lC���?fm�f4u����c�<�7!�m�ӳ��c��i<�|���=a��]oiq}�Yw���3s���~�".(�������7���h�1hD<�¡���c`n	$k��֒�3c8�l:�c���q@��8�nX�Q ���e|L(����N�ZȩY.��@~Usq+�r��&t'�$�$4�����B�w�ZR\Wv�@z�Ot~���`�.�\n�!ov<���;�2�U�PpJ��1���bŤ�r��ڃ�Ju�4j�Z��r6ԗ�+����&:�j:�����o����?���������<�p�?_����{W9��n��0�ֹH����7����t���<���ӗzys��:\��>��ƺ�\�w�M1s� 9+踈��r���l�s�Jg�\����Kzow_O�����g����u=c$I�r����{*�R*0A�J�	��[MK["�|o�6E|�l����ڄ9�bЏ�Ǥ�xs�!��j�yW� �˅#��+?�ո(_�e�l,ls2����()PIԠ��c;7��d�0���K<��P�
L&�cC�焦�c�A��v��Py���I½�X�RI�3�f���k�Ƨjݬ�~ת��rD�����[�� 8{
��J�������}�˘ ����g��
���֎���e4���鋗�^�h=�X�����Z�nW�����$7���VK�rm/��z>h<��Α�gջ�j6�c�@�� V
5�����pp'Uc����c ����F���+��Vn 9&M<�1Ai�
�ze=�b�DA�{t
}��������S���kCbd0��f8��hh�m4v�c�H\��(���̏�ժ�/�1)[zOV1p����մn5���5+u���x5ыލo/�g�Z�f��>{gg������3�' &tnÿ@q{ٽ�!�eC�xӢ;����Է�xG��ﹸ_��ӓC��44��W+���nE%����\���~Ҫ�5�BB���Y-U#iF��Z��X��T�s}���wp_�Zm˟� ]�\��������hn����VgW�J%H�,�N���w�7>ӨVT�x�Mr�kE|���B �JRX�� v��J
Z2f�q%`j�r#��IW�/r��E�%9�걐M�#� tfI������<G2�&l}^Gr��_���ⷵS�F�Z��	��4vt�`q<�_@��kA:�	|����ty���;;ʳ���tzu�'G���H%���Z�r�NRK�,��l��^@ОK�TV��sg(�/����5=x�P�vǣ)#1 P�U0qOGR7W�Z0��mo���\]���X�^�]ܬ7�0i���4����ļI����ӥ4�)�G���ҹ��d�Í�<�]��|�@���c�ό�yl��l�Mc�� *,�q����J��bZ��m�h��l�����j6�v�0�bI�R�m��Dn��|�$�dþ*5Вe*����R��ܘ�xc<��q���a�����X�UJ��˪�.U)U�u.V���r$�U*��j���f���B7����}=�:�l=W��|^�Z[�?������w�����:��l�ߝ�{?KqC��O-�s���]T7Y}����;��ή/��ٱNz�v��T�I�)��	7Ϡ�I",�hml���R�����s�W�&3en��]u�����w���������N|�F]�2����֞Z�m�<4{z�e�+,���}�U6j�^,`-��bθX����@����P��Ů�R����4t|�ڇ�#vmM"}#)R���(����tݠ=Ei�S$/�~�CGyVI��8��������L�����}k2ICφ��߅�i23&�g7��m�4��(�אׄi"��*͖N.�����=���(��Ъ�����Zj �L4�i��S8��ip~���S�&#����uv�T�j��,g֨�!ڹ"ʮl"�
��V��F��W:z8j&�Nf\�j>�����D~͔%c�����ȃL
���ʊ�
EJ6��x	}���U.��NGc����{i�
�M�n*��B�d��riOh��ڊ ��1�d�3�p�I٤�A5��� �/C��>&���Ɓ�������R4��MQ�~�.�I0���s�\�wqkTk~��"��-�ku��U�ke�y�汈�.7K���P/n�5[�U�e�*�fk�˷ۻ?�'~�5Y�ڳ����/_��?�t���ōu�f23���{o�?Փ�{������ͥI���(<fF�$E�i<�,�,���t���W&dR�36SԠ�..�*N�J]w��KUGs��h��ֶ�:���f�I���?PFӝ�=x����0��`4x�U46��ɘ��(�CM�x�$87��X��z}�dDD�tHN-�~���b"��T�X߸�=���9O"k��%J�d4E�̩o���yͯ����������!�x�y�&�󛍱3
�����Ύ�!3���Bm�fП�tj����J�m���������~�}o�N��,��ɬ���5˦5�nt��z����1w�lr�R%��zcO�I��W(��lwt��C8��7�IG�cU�l��BH����5��5#p����|� �E�%�D��TL��ύbu��./(T�Kc{�l5[�J����ت'���hhY�5���e��v���-��#��%�Ю&,�ت��Ce��B�5�T���*[�<�==�6��>�1o�����
to�[��w�+��o	Gk �JDu]\>�.<�K�[�Q�ĢzE�fE�zI�RQ���b���AWG�+�5�v)nO�[/�lm��?�S?�������ۻg��_����{�;u5X�ܞ�=� ��3zo�~��z��К7nH��*lĒ�����#���ѹ��6��,6�$�--��׃[]z�F�S
��S�ϯ4q������E=h4l?��l�La���0[.k�࡚�]�M��hn�Cwn�z�ap�4?����<��nGc�s�(�l�f�E��[.��ᱬ3�R����=,-��,���'�Q/��K��k-��K�/����)�ɲ�K�W2(�-�/�c�r�m�郅_|O�	�^���sP]0Q�2�#�Ya��tg�5�N�wp��i�qoV:[N4���^���A���R�rA�4��Aci��������Z�>���0�	v��w��B��T�� ��C����^:��*���;�9 �|ecz�pӺ7Rf8Ѫ7r"=KH�[��c��[p���z��X09�w�`S(Df����8
��j5z�N;o-,�S򙅭o��� �5CNi����\N\A(l��J��`G@$�is�-�|�/e�L�B ������^�!�R=A/��*��m�뀶2o��_D_����r��u��i��u�)5�I-u��{��B��	��X���:z�����������T���WT�������=�-���l���{����F��/�Ҥ����@?��;z��c�q-�e��Pɉ�/��s��e��4^�|rY�Mڔ�u�#]���ɱ.��*u�JsZA�=9���Z������u�6�z��ox�|����*S���h�Xj<�9��+���;8[����1V8S4��#_$�����H
P�o��q#|����8.��Hw(jh)l��S�3H�d��$�.~�}���2�*�@x��MC4��8%��0Ʒ0tG����t�`s���Ł�āģm�T������p���z�@b�x�0ª(�����r���@]���e��p�l���7���R%l�zC��c]�!��J�j���*;m+$�����U(+�0y,��[�� �@�	dcwX�N(v���e�%vG��,���-��w��י�8-�
�����3�'$<���ó���l�M��茭Q$P��9%rQ��=�-����b��&���vqmA=�^r� �V�Yc}	�F13�ď.oΩ�2H�fPB��0�A �.n���A��?ds���E.�A�sN.��;7����F�m��ۺXҬ^Ԧ�T��P7���z�/{W����zt�X,�U��?�;�����|'�����������?߹Z���t��F�Fq��EØ�-��/����y�T_��D��o���a^.� �gDp)0��	a|r1����R���PSߜ���K��\��WSj�P�;��g_h~t���0��t���O���k���㲂o6�~�ӵ:v�GO�&��*�u�2��-�� >��"vW��k�"T(6�67[��?�Se���G� �
�ы�+6�����B�+>�ŝN��pS�����{IA��%��p�Z%_��X��4���W� ؊Nq��Ԧ���Es��;�1d�G���/d��P=�Qe��ϼVŬ�thٴ� ���n�={�j4�g�)M�����/��h��ənN�4���q)ת�vZ�<<�y妔�.��l�c��q��ª
67��%利fd�x"�l��d��n�ZGZb�>���G\�S2j��0U�{�剢6�Y��^S�2NL��9�
�
K�H�t�k�4��&��mf�E-�$cuT�a����1��<��'zf��b��j2��'`
��@Dk�f�MG�h����Q�!Q.���&m#όm�J����m�q���j�a�:���6,��zE�v]g�>���G�ϴ̬�f��eQ]<����[����?���!\������>�l�������;�^��&���u I7�xX������<�� @i1�_�tc��� �So\�����8|��ֈ7��*��"��k��}�w�S��z������ҷC�+��].������R��<�X�YA�]p��r���(7lFwL4�Kiwxr0����6�[Ŭl2�V
@�al���΍��{4&���������w	7�3п�)���[�h��td��DRВ�3[_-l��	�W��е���\���x�����	��L�W�S� v�z�8����|V3���;���H���Y��C5B�y�tǛ���,ŀt������۞���CYf��P�����a��J�M��o;���`w��) ы`I��r������,��S�qAM4�,�bhIW���avN+�`X
��Z�v���bWb��k��RC��t��;�9���+4)��Ì�b�U	|-�W��W��S�\��x���򵢱�D[
�G�Yg��s����"�ko��x��|��􏉺�,����C�����(L�w���^����{��r��j�������FM�zY�뙾�]����6Q��R��tPk\>�t��{�_=��o}���8=�K���xy{YDh�-�Q$Q����A	A��F�{m��Ajn[jˮ 6cn)w��>k#�7��\��1Fq���V�Qr�������ˮ*��Z`e��;���_���}O�zCk����n,L0���a,�y�_�S�qf��Y���^W��(tM����F�i�:
��{l��Q��5L�>��oouqqf﯄�pВ�l�n\锂CE � ��p���d�`�H��ݛ�?jU������H���5�iB@�k�:#:���d!�Z���sH�8�1&�ᠡ�Q�y'*uW�:�5(���uC~Cj�ʇ�R�x����*d�<���-��g�}��/���`d�o�L����c:�c �/~́��ҹ���(�rQ���᪍f.v�Ñ�˩?_;Ҙ*���7,��roh20B�lp[�h"ާ��l�������j�iJ��=��3�&�|64e�1f��p���U��U/�\�y-[J�J^�r�!1Iqs�ÂhJ�H�՜��+��#쾗�&&���X�Џ"�1��&����v�!���]�S��أ3�"���To������ֶ��\��U��I����D��W����f��� ��h]����g^[q��}Թ�.�|6��7eS;�S� �%й�����O��Goy]Nh�秇vq��e�f�4xe�(���i�CL|��HK�2a��^�%-:��լ�{~�Ï>��gϔ�,���l�v�����?�o����?O��\�:(fr��^^��Mۛ��-�����o��ڧ�j��j�;>��╅���$:3(wY���=��Ҩ��$�h��%2.�W��牄�d�LT�٫]X��%�c�����k_��l�L��_R�X��"�U�Rqq�d�rw�PI����	�hS!�*_��������T�B�4:�g�k�,'�hU�?61��l��>P���щ~�{�����ڽwO��U�M�ջp m�9`��ۮ�h�+`G����ޗ4?{YD1������2�K�!D��1q t��[t��B����8�T�9`�tp`p��]e��#�|�1,��85'��m�����3ˮ*�%*� �jֵլ�ި(_�/p�L1g:� ϳqiK.�J�cvC�^1{�/�Ď��h��e���K����N�����<��%
��8���،�tr��
�����w����SikK�vM�RA/��?<~��z�%����ɛ{��{[����2��o/��/R���d��=���b5�%ǘA��9O�����׏������-U�}q�\��L�~��]�&[2&�;�m2=-j��`,0&��-��h�L��x�������O-vN���lC�E'�{o����}_O�~[y�+���~�-h4#L()M^��泰����m7#�H���8V�E��2tT�W+�H`i5p5�0r���J���J�		fFwh�-$�h�H����#� y��Dݤ�s�-�(��	��;�o4�L�IGI}��O�����5V��1��C�e:f��A�;M�.{p�TJ7}�W/5;�V��zI�\��|>��l��אd��_n�O�˰����=}��'�<;�뢓�wZ���S�QW�^����,>y�B���4 w�t��F��FM�̘�G^0��U���X�P����6K�$�
I�E#�28�еQ��7-����1���{�	���Nӯa~*�K�)U�� ��UԮ�`(�L�U�U6�-�3E!��#5c�
#j�)'hgIU�� ��r ���MOW�������y[��p�I�M��d-�Q�#��N���ƥ۪w��8�S��ֺ^Q�����Оn���2���I:�4x�����z�����Z���{��y9��٤���^V�I�F2ov�G�J��=pq{���UЧG_跟}��IO�RZ�R�Ft\��⚢�q���5��ؕ��m`��0��+��L���g��Ï4���f�g���o4��O����ꝷ���+�e ��}�q���N
�
''p&�k%2䖲H������ُB�`J�tN�������P����^Rm�zr:�񥢰:�D#J�Kp7~?�����$I#Od`����4)`�vo�ޫ�Ɗ��������dc��P�.�D�.2����6@��b��.3���KEq@n\2JŊ��nOǗ��ϗ*tZ�=�����~��P狉����X�[,�E�;Ś��[V��}}�ɧ���t�;?=�V�����6�luڦ������G�ܵǑ�s���r�h�iB�TQ]�2�(1Ju��zc�@��#�n{Zv�>�+dI�g�Z(A(�ټf( ï�WN69X.�m�pnf����2�2��bN5�9/� �Z��1���	Da�\�v��"�RȻ$b���7��x�;�E�� �c�4��    IDAT���ʤ���Q�8�-��7�Y{����*��J5���
�ͤt��t6���s�s�F��v��>y��������^Kq�_?���[�{6�����u�bе�^T��v��o�����޹�X�lA_>���>�ɴ�~I�`�1��-�R:0&H[�����A+�� �J[��Z��N?�\�~�Cm����NVf�?���O����Otppp7�����k�w�؍AFğ��#t�nW�� �-Q��8�moo����9�3�\j��[{�������<,\La���vwQ���Q��C"q���L�����e�n�dW�.�:D'&E7K�d,�
�'e1�ş�������p���N�+�c�c�h��@�i��b����e��=�ז�l��u��l��4�ZJ�l�s��9p�B����YK�V#]Ri�sdos�V�	�7痾��q��tT�5c���I&8�B6�e�+��\m6�l���q��LNE����.~��_�V��6�ㅖ�}��W��q����L��+�G	q I�J�`��m�A�dܣ��қ��U �B�&(.�*!mib*H���R�=�a�`��Wo>�UY�@�K[���v8v��{u��f1�k���=����%�8ԓJ��%y�lKk��-ձ��a[�j�̮\P?�	ҫ�D�ӑ^�^(U��j&�{������_�����[o�O���������?��F�d�����u�i6������>j�����zzp����#}v�R˱zi�[k�	�+d�<�(�-7�v8aA�.�?��U
%��ʺ��.?}�����!]�
�������ӧ���w���Ύ�Y����\�S��|��0��	"twM$_��hŖ(��|F���vvw]�z���Ł!�n -����ΎOt����s|�e5Aj�?�1o���K˘Ƅ0O���M�L��#'�P��X���y̤�s]�]��%�*��9������<�&K�N���.���1
���)\����c$�H�ܕZ`�sB��@����d�/-�F�=����hXH�6�Q/�Ҡ ��Y�
���Kn�V�{N�1$ܥ.^���\���!��
T��;8�����gG�{6�P ���t��v!�Ȧ�&���Ik�#�9qK/7gifC�6<�Pz4U~�R��t�!.d@P��b0�D��c|�/���ɇ�5A)��İ���F7��J\���l�j��q��0�<@��ۗBO�dk��,�L�
�s2�j֨6���R0� ��zc����#�o`fe��4�Mכ�Z�_�J��f$��2����#��by�.`�sqۯ��5�~�O��|�&����*n�������NF���tp۸�Ldy�t�ff����Vs�θt3K�.�:�hQ"jYH�$P�eNH\<l)PX���Ʉ�8�|�l�q�ⰻ��ku�U�婞���6�T�^p|󇾥�}��ڿw�r�$���e2a�*U*�:H�n]0�\G�zw�$��J����5Z-尿����6���/R�٠W�>ݬt���w���}�e�7k~Mv� >R)��� �r�o�rqF#Ov
�/H��0�X�Hh IK��$y<^a��(~e��~����rH����P(��^7V:5n�5���WW, 许б��:"��񁣾���s-W����V������ 2��!k!X-q��a)�c��ճ#�|`[�ɂ�6�ፆ��T)�`��G�0�,qg�d�W����w 6[w�-�,W�LC�&���ŭ�N+7[h~�Uj4Qi�Q��r���|�4{�>���V�p�r��s�����M�d�e���'Yta��gB�K!�R^K���RU����Z��>�N$�B��8v^�{��+j�Ӗv7�	
�� �=8�.c�����iTH{�y'��Xi:H�q��-���3ثow���4)���gu<����OϏLq<`!��j��qs�����o���{�#�\��������Ϝ�z��I��A�F�!����k���dzTn��WoX��Rޱp_�����K�x�h9���^a�����^(��/{�/g���-&���^Y�k)����f�.z:�͏4>�v�ս{��#?��z��wT�C0�j��+���dK'���:i����D����/2n���]����/4
r�V
ܵ~�4��� ȧ���`()V,k�$۱\-�����YJ�v�ؒ��qNqK
O�0m�����1�C�p�
��D�����h'��i	�`R���u�J�z�`�t��F2�ɽ���U�n|t��������鉾��-�y��U��[�~v�nz���.1ĕ�����$<�Їݻ��
mi�`�x�]���h��`�Pk{��ܑ6O,�Zt�����D�yP�E��.R�o���,��]�(;�'7WeMVjJ�ye��R��e<u0\C��ȯ\G��!��c�/��Q��Uŭ�ƞ�^��]B�x8�M��Es��j��̒�F���\��D�=�p�S�R� e���ب �_�P�a5�=�ڬ��\Y�z��tPL��4���-m�닧��C=޺F�)��E���G��_��{��������_U�~���������l:�#Gݛ6��Z�goO�]��ʖ����������3���T4�J]=�/�Tw�EsF�T��<�Im՛z��V=S0?�"6ã�\��T�Ӂ�N̧XZ�i�ګ��'�]*7_��������i��?��
ޕl��Q�L;��c�#u�7�uG	��/������f�����h81�vtt��SwM�hE�Q
�q�h��s�$f����O1*͛�u�Q
�eЦ��d�H��7j1�4��(&��d�}�2�HJ�+LQ�!��D�ղ t-Iq�s�!��Y�S�/��KF�����cz{�F��9�W{��R�n��ř�o�4$��]ӺQѤ�W//�JY[���6Z�mOn���q ��#�#u��J3����m��`[�jI�|�n9��/�	K����.����;��$�����_Bx�ղ�wq�{�&uJ���`�D痎��.Z���?,4�];��Z���.�u�;q�|
)��ݚzKo,�H�r�+�p}��ȼ,
���8����Ƙ�]�
ml�m���B?r(��c']�W�\A(l�z�|;�~��fp�:�n�4oT���烣gN��aQrPi��~�k�_�K?���R��I�����N&�����z��6Z�"7�g�����M��>Ճ�m��rI\m����М7V�ncWi�:z����F[�ٚ�f�8�V�h�����r��7�:�8Sw>4�:�~��Ŗv�%�F+��D�Y�Tv�7�0�2\L0ݓNd4�G|����qyy�8�*��A>$q���#�T$?����/���ёo��p`�Ð��7s�����P]��E�4�}�������y��}G;$㆐z#13)^�jƂȯ��-�����Tc8�,�Ϲ�[��mޓ▼t��a9�+X"%��ɜlǢ��l��?�xmй��3��l(W-;�_80Y�o��\]p݃���ԺY�4���[#Qp~�R&�J
�5��o�&ҿ������z��R�e|�_?����3�Yi�w��-�48����y(n\�n_��cۖo�l���U$��g�эy����YQ�����;1��@���,���PR�y��p�otm�D_�ˍ��P6�k+�7#Ɋ��;lK��D]J3�F���\Т�o3�=�:%x-�y�H)����FC�f��+e_���2����n��{���������!�\}jA{���q���<�����tn��g�ɤ���'�?qԻݹ�������(���s��}���������b',no�tL�F��zc�l�i+6�Nf���J�����pt��Wg~��QO�vM�rE��ިoiGe��ym�Zfx�Z�
ax��!���P.�<c'c	���7�&��n�[������8k{��@���>��s�v��7���"x�S>D
_�$���"�P?���J�ם�̿�$r��y���Z�L-)��"!�N�.0�~�Z��^�x%<Bw^_�B'����Cka]���wˌp$�b`��LG����(Ij*U|�����U�������JG����O�|���w5�t<��z=��;bD��}B�����A�Y'�^���L�[wb����ڻ��S��Fl�����k� g���h6"������!e�d���irq��x��V
���p�y�4�Q��� �װ�ʓR�`W�ɒ�`�C"��#z��|�bF��Q-�	�R���B�X'2(�_E6�!��l8�2üJ���h27�c<��;�d�r�s�[\�m�{�7aDu��+.Ҏd� ܄N��2�b|1��O�RS��R��вY׹fz1욢3����n�z�����_{��_{]��Uj�G�'�?y���]L{vgl3�(a��X��/���o��5���>__�{�%Ņq�~}[Oh��QUy�gc�i��tZ���fC�TF7끎n.���ݞ��,�U.k/S֣rK����o��v��3�
Ix�O7����m$���jc|����b\D.1��V���y!W��l��p����|yd.+�V��L������,��s�8$��o�8V�k��#�ω��)�B�)v�ȅ�(���y��7��$��XD|.)��P��r�H�L刅#,@��ՉY�`�V�1/ ��+R/nڤ({\�}�ƛ���I-����M�;�@��F7ݾ��=���	�kP��:5� ��0O�B���0r%����?~f�gP2gW�==� �������Mj"��ǁ3H��| ���ƞ������M��$��y]�t�LU��TZn�r�M���8�yȾD�1��v#�AO�cg�,�vݡ4t��v��VB����N�j�?7�/є�����mW�΍�/�����2���\�R.���A�p��h6�AD<� [��̖d���k�t�`� �2!�|���x�,�eh8�Dj����-�M����Uwn���5U��
����f��}���lK��=��N�����p>����� ����4'E�|���SՋu]�ouһ�gG���$�um�*zP�����,�|2]�������w�մ������ŪH?=�>�g'����L�:'^Y�ي���_lj�X�������F'�b4��7�':��0hV����d3�jm��֬�BH4[!I7�]�<��.���&L(�S�͍&][�j5��%cb���c�e�Mtqa�x�H�m~��!q��[ut�H6m���V2�&E3����\���3죏�R�ڂ�67+�ƌ����`���7v�����Q@:�7��� 1�6��b��Ⱦ|��yҳb���(�m�6N��f6�N�yͪy�8F���"�N��β��<��
�{�K���]_^���\�r9l��U�UN�]�,��(���E�)��N���y��@M��ܵ�+ՕV-��r��8�<�-'6�t�&��{�EB�@��3���M�|�V��T)�Li�)l5��_�1���V�@_�����_���l�$�G\��fs;�4�,tqE��L��D���ս�X���9
���X\�'�1�v�>�G\����-��l����b��L��y����X��7�����/��^�~�����o�=��Mz����C���/���o�c-�!�bv�Wq��R���~G_{�m�r%wk�/O�ԟ�_+�U�T՛���ߛ��x��G:���E��.��oכz�w��֎G͓ޅ���lp�t��dkSнbCo�v�_iɆ�(�؂�
�f�\�C�����u�_\[�\��]��kkkG�;�N��������ű>��S�����^t<7=�Uz7��W�[�S���q�HK��0O,r�� �ޝ\�O�����+�J������_uTu�n��'ʳ�	DL,8���+�!���P݂]�}�Mi���(����hOH�8$}\'zX�~�4�������þ��ך,&vW�8�y�b�<E�X*�M�-KN�]Sz�-ujYT˚D����Zr�ڎ�#�	!̮S�e��tu{y��/_
S��v�v�i�o7�*�Ѕ�*�O��Q���>���+n`�
͵��OTFK����vUWJ�UZY��p���J�.Q4*eg�X^�(��ǜ�I��|0�Z���̻Q`�E[��hh�Y�V� ������Jhzc�# &sL� j��а�*厎�6�R�7ֈ�h8U�������1����]��]�#W�:3�(����K{���쨰���v88ڏ�F�;�{�\�~�q���o?}�W_d�٤~��s'��u9�?`�\!)|г���jm}��z��[*�����C^����Ʋ����zw�������(���g��q��T��FGo?zCD]��������vM�RQ����5��.�]���@;�÷D�x�A��!�BZ䋳s�|���#6� ���ڍ�	�bYy8{|�7��胏���%"`|�4r�Y��;{n>d��|�Q*Y�Sd`޳�� =E#qqg�
��U*]Q���j��d�M4�t��t�
\N��~�qp���Gx,��n������
y��Q�pǻK�􊭦�$J����X�1���`ID2�M	`�� *wXu&��I_�jQ�VY6��ZԊʴ���Z��RNW�&􍆹&�B<�
Ǽ;9Ҩp��>�P��J����+��ν]���q%��3�ǘ>;h8!~���$�r�2���rE��zo��6�=-�z�^�3嵌no���U�CJǖ;؏���-�Yb�:v!��ou�WD�0�oT��m� �U�N��B�+��W%8B��e3�t�,��6E�EN,��ڮ 䂀���0Y����p:3�D�c�0f���1�� �����xX�d}	nK����w봕uni]�˹��s��/����J�������'��_���������A����?t>���t���9Ql���v���.n�x�-����*eK:�k;?����	�x��C}}���-u6�����^�6u5����k����������L�חjn�ԩ5���t��V��z��5{( �d|����`�l!�4�1��'���8�s���%�xN�D`\!t����V�/]�e���A���y����XY���&PF�D�%
�UJ�Z��)����`����\��[�L:E�/���BĝY����E�Ɣ��m5�O��,��`n��.�}�~��>)`�N^��"���3qݏ��p9���l9�p>��#NqC2�g�K:����ۤ��]�ϵ�����(f5���s�M��{ ^!�2�d���F���,E� �L���5�DP0L6+[�$&�YT���ܝ���\�TA�lAovv�����j����Z��z@?�FǶ�.n]�����c�	 ��e	4@&M
@�.�Q��W%O��[���Z5X�'�kV�0:	э��sc:��M'K0��p��:��g焳�]pLR�(\ȥx���[�H����p^[u�_1a��Zבat4[~u4�x�ӊ~hF.nolu~�����_��7~�|2���t��!�,O�q;{���7�zG_�������gzvq��>. ��O��˺������^�\�EP���H��O:�z���B.k?���c]^_��n������V���r�\��l�X���?��R'b.���Cu��5��Tr��s!T�5mmm����ay��P�}��P���[��9j� ��EA�CoaD4X�
(�I�ȟ'r�d�c�t�p��\0�aH�2^���<����$���A$'�J	6�=[�+>�G^��M���sb�!K:R(%.��O�\��+���"ctpV��q�15���JW7��Jz��ͫ^����q����0��.t�Kk\ʪ|o[�-��Es)-K9M��(�өo���q����6r����c�O/5%dh�V�QSc���N+���}!5D5=V12X.�.�7<�������Rñ����
%e�ý�k|�� _
�-V�K������T
o%)p�_��F@�6�`Zɵ�IdVV%�N(��֮B!�+�Dp;��Yz��`�0	��ʄ���    IDAT�
*�� �r������ [��k;�ch �Y�q8j���]��`��s������	���u<�h�Ӧ "������v���~�o������?�C���;���c��c�d�$��Zڮ���O�ѷ�{_�tIW�=?;����8^�����z�H�U���^t�����M���n @�ǥ�����t�������K�u�w:�&}��Uӗ0��Ѕ$`�Y���[~�r�5Gӑ>��ͧ!Aޜ�(�bM�:͖G).���}��'����ܶ�<��[���&
]B����N�[�դ��+�|�W�T�p���QCC�b#�����|H�ӄ8;CF+�r�q��L6��o��P,-�>5)�Sr1_���D'�?�u��^=�?�荆�:Q2��F�J2r���ե.�/D6j����ٜ�>���K�u���ӓ�D�J^�ݶ�vmQ��(�[�`�l~��6mj���ar����R��KM�nMf���j���mO8�8�ߡɍ�'�'t��z6k�ک�eB�m��H���������s�\�h��c#��ϝ�F����~0�'�ӂ��c),&( ��R��® A~���FvA6e���k޹���QXO%v�l�і����Z�x�	��%M&��\
�X�!�<
(�h�E,�"M�
�q��ܸ)p���jEi�>:-[usi��Mt8�鋫sͳa��o�~��}����|}��}���ݳa��N��'��e+v/����R�����7��
�(T4�Muty�����=s\ܻ�{�{���V8|vu�_~L	7!���-���X��Σ��n��� G���H�~O����mݫuT����n2/@��[�/��V�j
�3ONO]l�)��ku�+����y�ŲG�g������q��ݱ�<`ٔ�`���������������ǘ[�B�h6#/�c���r�_&��to�L�*�E.Q�X�n/bx��J<��o"�O�E:7~@E�"#ʯ?.���X�$#h� 1�]\���¿cLj�0r@��{kD�W��6��y�����^p��F�Fٌz빋��z�T����]���jY�k�������/��ϸn�s��I�k��.���?���~�&�>Ák�l)SB�\1`��=O�W&/��!d�"��̕�TYnTZ�l��tŔ3Y�Y�I��`b�zm�A� ��R��C��lP22��K�������[!�*9
tS�WD��Y�a�~Lt���̽��	u�U*�Nm��"{��T,lA����֋��"9u�j��,RX,d�^�X[��nH�K����Jm��j�t��[[�Y%�R/�������7���ײP�����Ϝz��Q�����H�	�G� �r%}��[��w��f�j<knNf�� ����Һ]���ő>:yxs���W�BE����Zz���J���zj7\4�\P[Œ�I��5UBFmRe��������\&\:^�L4��� �;�����5�m�Tno���}���Ӌs�i�DU���8�Q2&kp3�k� ��D*��.zQC�����Q/(���O����ȷb�㒷^�st{\J�me�-M����<*
f*�"�.ql�����Yx�r�P�(TIg��P$M)!�/�H�2��� 2�,rmE��h0T�wk�����`��x��� `;�Ԩ���bb�ԺVT�7<�����=sc�D:Ǻ�=6�m�i"i�o����i|��ʅ'�t�f]�z�txp�c[�uʃ���VN�V&��K��>�5�Ψ�ߐ<E�.ט���	Zah+�B������ �l.����fГ��*�[>�
Z]�5^t/�s�������#<O(�tmx�7r��2B��є�҂z��!�ti�sH�2�I�63f���DR˱~%uu��0�T��3������֦�Pj����ʮ ��"(�M�#ݩ�{�������,n���o����w�.#d>�ϧ4�m%˯�q��~��wlM�.f�9`U:��O��z��O���W8�R3S�v���������Z�(�٤Ɵ_]Z�D�q���n���JC%��%���r*��,���|���]�����j�R�������b��be�7~�Y�5�M��4�� ���2,-^-l�(<'��wQ��t`,)ҩ�K1�>���F¸�kyU��1ۤL���p����Sch�"J�B^u�M�.��،�ѡ"Y2����1��[D�J
���a�Qn����	ō�J�|�D�%㷥N��hҽ�������B�Q������@�|F�RN��]bI��y��j���45ɧ4!u�0o�� }C�y��Xa��8ʂM�U��oo8�S��6��r!8��8�f��݌��%�fq{å����Mם":U������㑱/˪Џ"�*�Ł�ӵ0��k������rB0K��3�������C�!ۉ:��&��#��K�dJ79��	�+SF(flK�P�"��1Y������uNݴ�H�@9��Âz��Ǔ{��L������.R{��Ɨ�i��;]ה�Z����֟}���dyě���wN���E����㾉�����$ c�Q3���v8�ꍝ����E�(s���p5����>��|6��}6�ڈr�T׻����u�I����f��Ǉ��*�����ÁQ���"!;{L��!#7*�2�`e��_�\k�Bt����ԏ�ֶo��vG�j� 4��>�P���ߺ�Ar�Q��:1Z�E�{�2$rٸy�0� �z˩Z��K+Hw��ţ���0So�-�A�0M�1�X>�����Մ{����(9���p��$E�]&�tx�;z��6
<�}�T�6v涱x��ű�x�>������Z)V	�8)h�2#�ɛfA����ω"g��@�B�ωi��涧��Z^��o��_ε��C/�;�;5��5��C��I�Tİ�s�	j�`�B��l�X>�D����g�.���/{8#�΍���8��0_�����Ԁ�ҙ�ۻ�jԔY�տ�	�;�r�k+�Y��lh����"���]�j!e|P�o���1�t�f)�ؘ"�r����eJ�f���)v��ٴr��J����l�.�� /�U�a�W
p:ez�BX.���_�US��b�/ju�kU���U&倠����'֢��Uk׏�;�'�����y�;�(��>����dy��7���9�����I���ӁW�"XN�(YY��_�����4����}ߗ�׭�����d�B`P"�	J,�$2QP��(Dٔ����xc1�e<��Q"G����鞞����Z�sϾ����<ϭ2Q4�sZ��:���9���<����R�6v�p�Ne2�d��x���zԷ'�g�Q��rp��r����S�+��:6�u�wӲ�h$}��m+_�jl��Z�'Kf26;8���N����XQ��ɠveɨ�V
E���67HH�W� ����O}&0D,>9wc�����>cIg\0��5X����V$]��Ӗ:5}�_��g$D_�Zn<O����~�	��^�7YS�(�G�247��@�#k�kM?i�Sʠ�������4�H�t2���a���3u�:�%�&�TT�`��xj3t� `���M��?Pp#��D~�i{�ݩ�l{���fncۘ�SQ�mTm���,���v�v^{h�zI|dR@��lZdpd~8�S�� #�
�j����]v;�B9c�T��0'���7�:>�b:���i⓰���۷j!(�F�����n��N�b�a�F��LY
��M	�i��W�7a� �Br-b|FA�����+V��sJ����YKf����D��5�����ʍWSF&��no`����S'$���7˼��6��2�:#��\��w������v���	�J��躕˖*U-U�����nZ?�g�����c�/pn�J�+7w���������sᖲ@������y���'��C����ዩ�(�R�؇��=h��v���4�@2.�3Y
����s�.jɨH�x0�#)�Wݲ�BY6�u�\��5��HL� ��ۖ\Ω��WAd0���'GjD�����E<��	��\(X�RB�� pqv�����;Η�w���V<P��^��,nT� �q�\+?��(�F27��z�UQ�2imlAO�� ƽ�/841"�O���`�Pv==2Ѵ��#�}��V $�3��m$��� RD����P�������Y�>+��F!�:Z��-4��3*�s<P�zx��^))��6�T��۱!�$,U���n�0�nl�J��|b��Y�Y����������2��揉_,���{��21\ s�_t�wݨݷ�uK��Z�&��*Ns�9S�G�u�n2!�0�wK�e�"\F����S���D�y4TP!��P��,�g�j�0C����+�P��4��d���Y�\�ݭ�~��{!M�#���1~��i�A[9�ͅ�S¤�I�
�����0VfKk��r������|as�T�½��ʹ��J
q��%u�P8ᾎN>˕r��Vq�<6;;�l6��سN����O�3X��XE��*�Νj��=[o������|2�o��[_��v�y6��lҗz)�(z%�\�x�U�2��d�0v@��E��9�`���-m��ˁ�M6��f2g��B�m3u��A�m�d�Uc��ʶ���>}�T�fЁ|��$Q�ղ�nGVb8\s���8�{sJq�"ΆD�nc��f5��>�&��%�2��ra�����¦fJE&��e�W�����Y���Ea����<��M�����r���X��W����W�4}p���w=��E�X7�*	n���[\�(����Q=�TJ�O�V����%p/J̾4��!j�Y�n,L{�C T=�pa#�����9X�6;?�
.*㶵u`d��\�b֏��E�eW��Y>m5��v,Y)ؚM�K���T9?�dt�`���)���/��ou��;=k]^Y��R��8hax��������rt2���/�U��+�-�B�l�� Ѐ�8�� ��̉\F�M9�� �u���8��IQ��RߪU�R̫���� w�"�`&��y7��� ޥlȌ�ED�m8YX��W���l@o�S�y��B�|���E��S��e���cM�0���eMY$W�����[)��b>����ɑ�l.�����Z{�\��~h��k�[Y�7���_<���y2��0����(���|��޷�틇��-(0��>��^[k!����$8�雌h�@fDZ_Kfm+[҄i3��x2��zi�2���h��֎�y��t�٤��N[��)(k����K���l��Д�l��D���c�o������W�j�8�$���i�Ԯ����R?*��@��'/{h��J�0Y�V	����L��E�L����}m|�P��EWf��J��ZCώ�@��A2�٠���1d� ��vvd���u�p}�?����h�d\E���g�`�C�V\�]: ��=E>�2>LH '�R]�'��X	ٌzm8�u�����&��Rي[u��4-Q�Y�\��&���� �1ML靑�ჀrG�)YV2-	����}��c���.�J�H =<&��d#�z.o�v�l��۪�w���F
&�ʅ%��Y}8�2�d�3��`r8�_'�3�7N��;#�Y&���{!��d�R	(MBJTO�b�2٬Z��M���՜ �Z%��Q������<.�g���Z�L�d�D��|^	U?���K�M�g���L�U*c�J�"���b1{1��k��׶��$D�JF�Y,_�)W���9���?��G~�b�s{��.�o�w����g��J�0���x��썭}��݇���+Z��:����3á���+�C�A�X#zzSѕNS�>5za�,���#-�҈����]�AL�Z5���Ɩ�����N�eن�X*����s��i�n��=Fؖr���]����B:::������p1� Ǎ�-g.��Cp�W�[P�ı\�ޖxv�D��l<��	48>*� �?��󿔉y��Y3�A)G0`S��-<I���4�����pL�9vo�	�aHA0�Z�"����mepH��`C�kt�� oN��SU1+|��)`n �	nj�{1�cm��LA� ɿ�P���$?�L�I����A�`��弱.?=?��C��ֶ��坦���C����Q���b2��Q4�Ԑ)Z��i���Nߎ?�u�-7�@L�RE\��S�N�z�wG�g��@���w3����,M���
C/!�Zs�%�a9�ش?�!>��W:H.�1�P��֖���~2�)AN�N/N���~����g*U�o0�A<�	9{6j+a��¹q� ρe������$��*�F�������^:��*�/[�X�E*i��ʞ��v:�K�r	�`��kJW����_|�k��W��ȿ��w<P��o���'�������T8w|�� �����r��^�:�3Dwܯ���.;������`=��㫠RL�sqD��L<aL�91gk�r�F��ի5ȄX��W��Ռ����M��f�n�8�]�����{��#�
�����������L5 -:��!}Ʊr�.�߼�$��-��+$�mOm�T\�@�Y��R��O3.,ж@Q�}�]S�

V�"��zo��2���[��J��M��z�Y����L Β�Z�R�&�%m��V(C.�NC��-�:!��`%t�7�	eo�7�s̅��T�+U�d�ָdm��*u�c�r�������
��ked�|����m��*�!H)cp�����;\̧�\�OPA .IiJF�}pݵ��u�Z�'F�PB�:����52���V �S����` h�T|��]7�֯W߃w.�pf�`GP�`��tc'֜ӨB����CB��n�3�g��u�&:pŦq����0�R�������j!�"�߶���>\�/��nJJ�[����gN[��2Zne˗���[,�*��a,jgө����I�¦�V�I��Q*]=����#_����?EP��ޏ�qp��{x>�������<t������-�Ca�~�/ڗ��ai[�����>�8�S��l�p:��OE��9����~��2&�3'��\6��BĬ8YYe����,=]�j4��vlӘ,�8OOυu������ �?5�K�s�������7������5��Jx8�Ar#��4�S����&����K>�J@�>S�D������D��(�F-X�M��ƢTs����||�������W� �%.s
���)AC�[�s�ET�(F��v87]{.����?��j�)�C�H���@�!�����&�D�ގ2�xRSm���9O�����t���t��LFmH�Q���vB6i����;-;���n��&y2���V�v���ۤ֞�l�,���'�����D�07ܯЂ#`�n�/����&��t��~.�VS�a��gҨ�t��t����wa��H���b�'�h�**9=m�����
,Zb8_�Ĭ�^v�`ހy��#aT/$��/!ɻT)�����:�/M�y��T� �ޗ�p��|a�
��*�ד⇞��g:�>�&�U����ɣm�A
��筛���|l����j���&��f�r�hw�O��_�c'��3�>88�����A����c"1sR%�6k�����{���Ν{�[j����{f�/��Űm��X��q<�����gr���E�e���s�'�R�PI��Z.���ba��¶#);�嬴�۴�Q�+v����J��Ϗu��˫�kg <q�n��D
������
pdP�>z��@��K���( �.�d�E���#���3&���w4�ہ�?܄�B�Q�|^����,N^��A$��[��?��|TC�Wq٘�W�Ρ���`�%��,��q%�+eC?���/�����sLO$Ž�H��g�|6�`S	Ǽ`��#7%E�F>A�ҋ�L���^�un?o2*��M�`�zA�-Z/�*��k���;���A:UL��G�t��b����Ώ�����_=G0eж��%2�b�>��x����f`��XA����=m%�rф�2��    IDATE�lNmvӱEo x���dl�9���OU�8<Z���u�(I���zr�mlVn��̸�A�-�+��S������P
�$�$�$9+GsT+o3�;ŧ��� �J��t"�����']?����\
��-S�$��R��ժM�C;�gǆ^d>�Mdi�R�����^��?�w>���o?~o����g�ֿu>��;�;A�l�S�Z�~��/)s�+7�����=�<�O�Nm]ix@Yz��o�jVʔ�3���Ҟ��(ZS*��s���mD��-�V��mk�{ي��Ul�Z*�1�Ҕ^7���T}�H4�$]nBH��*�4m%˒�j,mo���Q�R�~�����ٙz>�F*��XF��Sݫ�B��	��T���Ŧlϋ<�s�W`���ml>�-�k�j����F��ŦN����-h{57l�^�;,���o���y���W*>kp��`�V,޾?����{:BE�&�k�K�p)�8A� Ep��у���E T��q(��e� t��*Gc	w}}7��`���xdn���Ewj�\�36�G��B5��Lk4�D$n����wI���1=��	������O]/��"������LC���6�jۨձ�hl�t�*���bq����;=����E�b� *��P`������<M���A���=5¡�^�"�����gРl�;�		�M�]L3ɮb.x��J֩���e���������t��S�x�V//dz	z���%�ί�{l��%-���k�H�i�"��m��V�����G�v�k�p1�h"j�R�ug��_��?����E��D�~�3����wwO�_x�k���i?��E��B:V?��;����+�ܕt�n_��i�l�1��;[����VJ��f6�������qd)uI��6���,;_Xy���h�^+6�n�!h�U�Ʌ\�����~	�v��IY ˍ6	'/���E�
lp^�^�=9?sY��i�66��Ғ̍2���Gh���PI E�֌�5���5��A��%S9z�BA�Gld`;&z�4���K��/8�H�pm77�Kޫ~���2Q�E�
A�N���ß�9� !��F� ��,�������+��j ��6��ե=?>���S�9�iO���ݗf���&��-��fŢ[e[2��4����Z���3T9%�mig[�4�E{Ӂܯ���B�FS���5�Ɯ�0˝b.�����HԷ�����b2i�D�
@K�Au�6���b0tަ0衑7�	����}.F�7:��{8h9:�i �JγF^������̷�`^Pr��:���M^��E(T��r�808�������^�r4���)���y���H�E���L$��H'�g����2fɴ-�s�l�f�֥�}|uj'����}K�c�U-��i4������?~�ѣ�gZ��k�b����֏�O��q��A� ���V�=�w��ڝ�΄�q��?��g�6KFlIp[����{{�d�ړ�]�;���X����H�@ NF-Kv6�[a���d�^�n۽r����Ŵ����ܮ�a�~ry���C��&�{���0�eJZ(�ɓ'��.<#!d\�J��˾`EGXt�&5i������G@�,HD�MO�($�����R�Њ fU`�p �94CC���tb�!{
��@���9G�"$�C�r���=O��2�Ϝ�/ב�n�R����֕�������S�K��\*P�%U�ִ���n'g�������]���V@ �����ỚJ�,��鲒��NEr��T���G66Mկ�]˜����X�[mwK���r*��R�$����>�}��=3�v�tI�Nm��X�������WL$�Li�L+��5���|4�,�ܫ�*WZ�r��ʩiHM�ݴt�?`4���;��s#_�^>�T�Q���ڧs�����˗�8�(��8�����
)���]>�b���p$vˢ�J�g� ����*K�ڊ[�	n
l ��E�[&Cpk�U
���Ԟ�/���$l�V�����������7��O�_L������^��I�g���b�?�M��?���}p����$Qt3�iZ����mjn6���C���-I�堭�/���$��El-�~�������}�wD�"s㴄H���g���'�Y�.�ɉ���hø^��./.��T�&b:�ܻ�,�Ӈ))�!�UФ��=(q�����u�,��a���8��'�O�/�\�98�dn�z3�P�9��T��0]�6�[��e����'8�RE��I\p �X�Δ�r���C��w�2b�q�-�tW��f�6�uht�|�O�1d��\*[6��T6�qW�kk���a���١�9�=��_2|[3)�%�։,l�v�n��Ld&���/�U��yK}0|䈕J˴$��E.�R�v��C {�I5��9.��3A(��!a4����n�.m9��u���iej��-�	�x(#��)E��+*��\i� �[�\`*ԫB	\�˃�=�{T.�u���)��WbF���k	�/[A������j�u���E�3����.��b1q[��6�HXaȞ�(����
E��R��G�'vҹ��T*�z��٭T�ܗj�����W�߫$����R���x���F�?v9r�� �S��[4m_���
w�{�����=�:���6�Om��@$jo?|ݾt�5�ǲv5h����=~�\n���Z K�2.�Yz���%�~�n��l�\�
�m�+vrt"�U�Z���	�P�����7��k��dtϦ��F�4�L��Ө�b�T�7�)B0P�a�t�� ���j�)Љ�#GX��2
@��X�e�t&^���Y�%o��k��C&#d}�+���kP�x-���J@�g(C�=�t]�_���e^@+�	��hԭ�l*P�g2z�XrpU�`��^������j����~8T`�W����r�)S~"�5N��8��>��A���u�-��h���~���d�rI������Z|�a��m[T�ց���x&�r�H�i#U�b<e�O��u��ViT�P�2��P,��8=�%�N�{�g"@���̦2�a]�dКJ���A��/�!���´9̣�9r���1׫|���ޙI��0��)*c��J�%��{���T�����\�@租��<u*JT����Ap���\
L�/��d*��F�rE��߳Q�F+VЕ*�䢆	�xn2�5o�L�"��-�y[����ՙl��a�*�w+���ˍ��_pe�~�G/���N('-N�ˍzn���M����,��倅���|�o޷��}+$2֚�}mO	��8���T�1��SpmS�%����m���P?##���g��]j�K�����$���,(�����l�F�n_�җ���ߟ�8��pF�d���u# �,0�� 6�w�
婀�c��t&��zC��l6���Y��d)d{dq,�S�p�'�1�:Yq���dN�FCY(?#[�%h=6*�!]`��kJ0Q%�Z׳����-(�p]d_Loy�)����t恚y�ˢ]��J&d�g}#���|��3��!�#s�����ե4��1U�N��/�R�ar�x߫Y�ޞ-�$"bm	������1k����ĬzeOb��k+�*�تk�Ջ%��201�#A@0qa�l�>Pq.�wٿu}m�vO0o�!���Z�:�5�}EV �)S܅lG@^����2���0�N^⧝r�b:�Wc��*�F٩Jx��������|L�e����y8qs�wK�q�(��W��-��Y�Z�c�#� 7XD�(��^����hlY!_�������u�e�6�n죓#�v�/�g�^,�6�?�}_|�7?7�J
'��_yֿ�w.���<b�nӥ��q��G_�w����nlgг�jj������JͶr%KŒ6�N���
�KSW=7�U�.qJ�Ƕ������a�nw����/�x8P��A��̛!C|���4����EHp����-������Cׯ����:a���T���L� 0B�C��1xZԊ�i��?�	�� #������P�����0�$������̕�Ng���������xq*F �k��g�,`q������=�����O�/4�Ĳ�Mv]f�g)�ᡌ�9$�5g6W ����Ж㑂e�2�)z~N而H��΍�[��i��t2 T������XF"�_�l���f�dv�m�Fή���V�I&<�	�7��Zr����S;}v$�GTw�w��`wϚ(0��N6n�H���]�7Y	�.%`Z�gݞ�kf>u
)��$H����X�
P�e@����!��� *��|�ҕ�xCޗ���d�n=M��t{��a p�i� 
���� �q7�z�O	P���Ry�[(W^S��?�eq=�;mNdCe	,+
`�J��+֛�u�Um����bf<bW�����G�Q,��j?��[o��?��/�	��x���R2�����[
n��j�ӛ�-��ڿ��M{��C;��6P<��L�}S�� D�(�.-�ƺ����w���p��4v	�1zݾM�o,1[X#�mUda5�A��Rv|tbg/N��%�������l�7����f�j�Z�n�dE,`~��M�zX��`�H�zD`����j±�N� 	�ґwٍ(�Q�o�Y_Uv��	 <�(���FH��L��R�g�T�iR;���I<������� ��-��ŋv���>$z^�qTc�R���4X�����5tzm{��ȎON�g�
���w�	C�Sؔ�;��O��p�Ab"�9��T�sܗn��h�\�'���]�[����π�D,��H"i���Ʃ�-�9[�Tm\�۠��NteK�Zә!���o���Z�=���S���| )�v����tG�m\�,�����2?1�����P� rM]7�	ĔmXJ��#�y�<��$�2����~z���R�g��@���%$�i��h~��a�������)�L�cC�Wի��R�[ghc���T�ك� 	S0�[��O�dX��9��_E1�O[<��J�V@͚�ָϬX��fi�[o>�(Z���U��~��?ߝ�_����W]�w;������u��h��#��8����)`�Z"oo޷w�n���s��ϻ��j��#L���s�����*����ق��jKFf�RXӔ����XL9;7�����)���ڧ/����BZh`���6��%����(�I�~c1�Ak��*�L��g����Aa�C��SaB�
dr~N�c�Vdqd���L�Y��|1� W�P�ך~�}���ٱl6��Wvqq�@F��)LwC���ޅCZ���C�%�c�������������Y�B=�ة�B͉[�����B�ٺn�,�g3�8��3��%LJ��Ю�/����i�aj�L9A�����(�E1m��M�9k��6��lI�Ak0n5KZv���uߞ|�}K̖V�'��������m�k6�4`�	Ԩ��z1���[⩛r���k�\u� ���٥* ����P\W�1�QɊ3X̩�Y[��7��O�����T��k}�DҐ s��#� �OBU�z)�p���u��~��.�T("�a ��l%_�2Le~���{Qma^����WX���E�/M�)��lZ�`�2�[2 ��%V���zO�{�����ݭ��<����
l���E���s���{{G��7N7����+���r�N�����}��vj�W(��K)x�i�;m@e;�@E�G���g���l�;}�F���x�"��4�a>�ۧ�?�^�	K5�>R�����h
��F���հ��ݤ��y h�C�<�7��M�Z-7�L'��s�� \բƪ�/@�|��'�O��t��zi����J�^Oٍ�>"�L/C�zk5g�Kkb������B���w�VF��s�:h\��`�b^A�V���u$3�=���K����v<re�+S>iZ�7=$l�zCφ�>�n\y��&��Yz�6�67C���n��$��p�G>'0�b�֙���Ӷn�m\I[�����+]���IZ�R��,����O-6�H:�+o�i�4Áj�ZX-$��*M������s���i�OA�'�Q�{6t����(ŏO^X�۵�V[�A����%o���Q���Y&8A~�i'{$���?����,o{r�Ӕ���� _�/�[TJ�EC�C�p�~M8\�2=@�7��]N��_�	�DNId��$�45d�S��+%ySd�In�e3ME�M���H9Q��r�����Ӈ��o|n��>�'���7N��i-Ƒ��~MT�W�~2�5�U��ܶj���F��w�|p���ρۑ�lā��47i���B��ئ;��j#g���m�8���da(7?��6��(*զ�j�SpO�v}y�`���W�@��w����`&<��6��$�VR�p�o�6�A�Jwt&��Τ-,$2T����\斛Ҷ�rN9�ѯ��Lo�pa�J ����n:A�R��g?��qQ]�ǵqݠ�]��	��#P������������gx�L���[9�&=A4�5=�'tm���N�����`��;�'�'|����87�g47���F��n]����Q�&0n�9HȢ��u�d�jں���QC(Gmf��*n�������i�,�2z���6	k �zG�[{vq|b���;z��M��jV�n�9Nv�Z��s����x�����s;����S�`���0��#�O��*�|>�6A�|��@�j��TX��|��$s�U��.�0��m������$��eb�� �K�sCG�ww=n��z���ɾ��%P�a��RknY�Z�\�b�R֬P�5#.x������Bix�����{ۿ��Kp�Z�"����E�0�Yln��ԋe'/N�D��Mk���&�N �HU�ZY7-C5U�xl[�=�n�w�j��8�%x����>��RJ�bV�m);��J��Ln��n)��;]7$���;�w�i��z����G>_G��qC�,�ƽw��N���,e)7UYf����r
`281TR:���T��L^���h\�tB�M�"�qw0��dl7��;u}D�0 H����ce	x?��w�
lP��l�20�W�Dx�J�Z�9<xR�
��5
{FII-��>�Mݤ��?��\�}����R:4���E�[f��.elQ�۠��n>a�LD��2j����7K&vP��!ex�b�Ѹ�	�_�p��={�D���L�M��=�F��npL��4���J��׷����~1��E�wH�;lG���	U1�_e��fl���6���{
�W�U�"�:���&J�Jʗ�А�w���I仩�˾�G�rkL8<���m��M��[Ω�Z@��(�u�{dx��Uv�,W�Jl��YZg1���X2��R��4���r��޸s��kp;��~�Š��/��X/2s�$�x6"�HZ5_��FIm��jt2p���>H�њ_.e��29��K'��:��hn���V���]{��e#q�A�^-���������Ǝ�:�^��� ���H�o�L��ww���������Wp��*l�\��Q���q��`�6e��䄍ʍ��Υ=�&x�{X!Ɍ{�I^��3@9B���%�O�/L��d196ߖpf��X�'Fps H����)�7�{}/���:�MS�v��9g�L�Hp㥅�t}X�4�ᙼU�׷DD��m��CL0�k�ˡc��r��	n��LF�����E�hkJ�\�ƅ�u3��6�&l�{2��En��9�Xr8�u�;��~�f��Le��VS"�~�����l��~s�޽g{{;�)fe��w5�G�5�=�	��o�3�8?��d*�	���L�X�6���o�:#w��h}��Lg�P*�p��	��{b�[�I}��n~���	~�CG^��ԃc=C��d�{��Kk<�zkd^@S���l`J�����k��Pg���^��F�/���	i�b9�M+ժNg�^�x!'E��̮&��ΈGT�����n��ފtH    IDAT�w�/���k��������l�K�7?r1$����-�;�2��|p�|�BQQ7��lF��1Bk-���iÃ���	 T#��L�72��N��T���v��%*�$�$�p�������::S�������9�{������Fc�h��Ν}�x���N���v�F�M����p�-���:� )@ֿ[���#� r��������;4e6^���*�W��ټ{�+\�=2��ύJ�< *5-T�S*���l�TxCf@�R9�r8��7�!k�9L�0 �P�0(�}�Bo�ϱ��[@D	2ڝ=�{���ɑ�rM8Z�!��;}Eޗ��mPϛ�7�����P���Dٿ9f�%[gS6��l��['�Qp��6��-��myٱ��kˎ�Zc�޹��1�_���j��>�������u{��}��/�_{Ce*�3T� H%�Ě�l��|4�����=y�L=ڭ�]p�B��Y�Q+��'k�@��f��
D�E��C}���֎zr(`�2`p��K(���~�����\r��6�&�$�z��Z��H)�� ]��e	__��%���B=�����l�T�9����0k��ڨ[�[�Jc�6���6+iC�"�YN�z4t��F��J23�-������_�k�ߖ����w<P 
�b������=��S��Zzn��n�K5~�(�2f&;�����9t����	��E*|�R��t�$)��K�����n�h���<"1�����B���{_J��'	�ٔ���ĺ�����)C ��������v7b�24��*7R�i)X���I�g�>�/{Z�<o���ܮ>�
��:Zv^M#�l�����U��E��Щರd�V,�`5qP
�L �JZ����J��L��%�IZ�/q�*v����D��<�}O�՛C�����l�f$����6}0��Π:��^����ޙ��zn����X��<
�l1o�B�ɸMRQ��6�%��=7ݏU�fg-�][n���ܻo_y���q��e��Bm1�_�{߾����Q�7��G�v˙�kggK����Y�<��S{��MN�1�ؘ�k�!~� v�h�-m>�+���mT������i�k�6���B��\�G��_(I_-[�A(�c� �8��9��;Bp+��A�E����d� �����-�|!k{�������*G�.eֱ�zk����\���s���m�H�f)E�j*;�)������y����l�̮~�Y���N�i.���6"<��bIz�jh�%FB���}5�I(W	۬��3,�g/����ʡ�Y�%{cc�Z�$m;���> ,P�����T+Ȥn�~�q��f
n'/^81ß��&l7�NAןZ��ܸq�h�z79B8�T>8&P��]:m%zB^W�M!]x��[�l�����%8�`���	?+���bїq�̅̒�H��;��
��+��笪�5w�pNTz�+ZR�����^�?l� `2gwʛ�>*8�^ϕ�6�ͦS���tؐ�����s�'�q�ahA��u���h�e)��	�eЖ@v��I�0�O�lU�ۼ��~!m�\\e)Gm|ze��WV�o�^�~��VffӉ-���{��������Af�����Y���}�W�"Ƀ��L�6���ũ==�-G�iz`2���)���fe��������)�J�%���r��N82�4x�)��tN5�m����<��ՃJٛ����P-�A���(Z5E�+u�ʊ�?�bZ�V~�AB	H�c�0� 0IR��������_��i���<֞=2XT]6k��"��t�S���Xv��E5��J?�����/����	����}�q9k�������M�~��������l�@�˼��Ce�����R�as���Ur%-��|��}��3�h���|m���v0���l+��J*k�lN����f�裏l�s�(���C�٩����t�.�&HHON�5W������P"�/�	&�VS�����v�S��E>�P���ES�l�v2ɟ�lZ���4���&���|g��h�J!�a@�����1�P�qF/��^���h��B��#��&��t�(r����K�pz�\����O�N@�����`�?��-��Qו��is��	���z@���^���Ip?xM/����L�"��Ev�6,e���(�q_b����y�R����o����W�7�`��Ȟ�؎&o\�%l\'>�ֵ�����=�۱�Z�JY<6�N-�3�<��/����ߘ�)SQ���z]��Ǐ�gO���!�%R��q�C�<�q�p8#��A�0nz?^����sCI��=��|)X�=&�"䣃�����P��l�HA��!��ޙ Œ)����U���穐���+�������ﳽ�}[m"֛��ӵ	��hD#���'�wG��Uӹ��z�'^���K_�ϧ,%�]�o���A�O\L�Yx{dn¾�ˈؤr�N&��
��c_��K$�є�i��N�n�BE'�GOۧGO]�٬-��|<��Xڪ����
V��-�`$j��]S��\�T��Ɔ"��&�FB������B�׺���Wn�7�إx�<��̚�D�=�t�������1�Д��Z������dw(��+����#�a�x�a��{�	$[>�dC�R�(U�D!�@���|!�����,Np,f�F�6�Qj�i/��f�������
A~h����o�4����b�� ��x2;�?���b#	:�i;���[hF+=66Cn�J�6�UR6��nqn���fm[��-5���d�<|dwww�I�=;��/�s	r��
���{�}c��ؒэmWk�Ň�m���8P��%WQ�LW־l�B8=�PomN�������&���J�S�?�Ğ={.�X�%ZnN�ٙ��w�6sL�s.�K��Ȱe��!�Ttc�u}6(T��\�Bp�(��}qN=�C�ee��x�Lydp���ܓ\<�@�\�㮮����s)�7v��Cۻs ^H������6��,nb�`���$j*�dj�_)���������P��w�m<��~�h�����0C�Mp�i@p��P<E��`,�[�܄�����&n��m�klY�\ї�ѧ�ؓ���j�<ܶ�ikD3�W*K��-){DQ�I���%�-� N).ݱ����iZ�7%�c�s{�e`�ʅޕ�llF�U�v�f$H\�_(H2���sYAй��v5�y��jKi�6M�P2M�n�N	�-2�.�x����AHʏS�Uʮ��wF�l���υr2�p���^�^���]en|v2�00!�i2�t��u�`��@'�L�L2Y�"���%��>� �O8�{(H ,��)�ӔoD��[ωk2�%��3�G})��f��l�V��-����e6���,mrֲ�iK���ۻk��v����֍��m���A^Y>R網�h`3��ԛ��7�v!�^]li��B5]ڰ;���k;~qbWP�`Z$c�FJ�6����
Œ�^�}a���i2ϡ
^��$�����K	���2M��k�6���p>s����E�$	yR������Q��}_Ϸ,���xB�#�1` �OP��aP��{V���MD���s¢/&��=��ߵr�a�|�:���ш��&�V�k�ݲx��J��p�T�������������<�~�h���.��T	..L����B���t�ܸ���&'��J22p��ܖ+{�٧���XAI�y��G3�I�l/]��JM=��l�J4�&ˍ=��3m66J*��s27���5n�e%W�57�A\��#�'��B1���f��U�@\�,L˕���ä)��,���1B�L(*X� ��y8���L!0���^����zd9L՟�M��R"������R9J��FS�O���s7��l��(i�,P��Qzp4��Tw�$��V���ǹ��(��ʣ���P�K��)�:O8Oԑ�i2Psb>�ޠ�̄)$��V�ز��y5k�R��ٸ�Q�H&܆�W6;���pno4w�Ѵz�`�,Qo w*�\=**��@t��|�)�Y�~�fo?�k;Ŕ�f��_ll��4?NdNsѾ�.���ʲՒ�51��[Ph)���na7ܴa3\k��M�R��v%r�j�i�%쏡}�7dX�hVLs��W�n�E���;�ظ!����0+4\[P�%�q_Q�m�x�dmrd37��5������s���߱���Je�gR��A<�h�Ƒ� !���Q��dT5��K�����ʏ~�����{<~��ҿ��?�:��x��:�M=7en!@.��ː�]34�"  σyP��V�v���Ϟڳ�c5^���sPdv�y;,��N�&���x�&����9>��Cѯ��r%m@n,���t�e�/��2��mW^zV�}H�
P���$�w�fA��jn ��gQ�p��2��� �f�\Z╞O���{w����F!{�uh�kQ%^J�/����^��`�{��gϞ��`3)S�t�I�R@ǔ����n�� ;{���㲳���#�+��N��)�D-�p�K�a��L�ɷ|X��}�46~5sӵb$�G�x.4�ɔ���d<t��`<���M���f,V-Hf|R�ج^�>����M�6>o���-�bͶ�#\ʚ��\[ji�U���ՙu�M��B$�+5{��53Q畀��bc�����Mg+�hݸ�6���\W�Z�g$cK&��4�s �%��OJ��汋� .����RM}�$I<��3��Ø�%1C56�����	G/ύ���]��`�M����������e-�A��L�R�c�m�S)!�?|���2r����ƪ��D�&���)5��¼nֈe�*տ����_������
l*��E���s^	n�r>�v#K�W����&��6\Q����$��L�U�$$:y��k�jM��gG�����`��/�������*b-,�S�^.��l����\�贪V�j������u�eW����:O��͕��nT�=I|�^���Bp��c���A8<A��&��὜v[V=��ė
��6S��� 2,Q�������y�|27�k�\Y(�|�P�D��!��_K5ڝ��{8}6��{%K�O���(�>x:��
b�L��vO��_�s��>s�PS�W�������<�j��M�Cd�oZ.�����pՙ��	[4K
n������m�����m���j�$���
Ʒ�Ym,�Z%�@�5u�����[OgVJ��~s�޺�k�����f+Kn�[El9[Y�ӷc&���M	홴շ�\p+�o��:f��P%'A��l%����\�*�sa��Dw2i��Ӈ���s�~����՚�=�^�7�a0����%;�p�]�{_����&/��	`�dUI.s�tڽ>�7�mwܷ�	
��d/��f �q��"( �� �:��V�8�S���;��?���~���ngn�x������g�G��lǖ�I�����W�JV,��t�/� ������e3���B��o��v��&-OO�t�G��ܹq�j����.�^�l) ���U�r��ط��-��jic��۷��A�/�?&��~lo۩U�������b}j�n�a��k[@	Sj�2�0�r���tJқ���N�����d�xu��:��smxk<5*&�޹'�l �cҌGj.�����(в�o�obx��h�j䀔ay=��W#�{0����ʰH��H����@��:םN�}�F4DxE��o7aVO�;f����y���ZE��E�B�����i�e��t{}-f�m�U�
n�B�换��)�h�Hb�Ӗ��;���m�T��Ib���bey�Z3[�Z��k8>;��ֹ��7�Ϭ��Pc�4�VM.-��¬��a=c��О=?���/�sc�D�2�������#Y����s���BQ�"��<C��+GA�s��K��#�r]��g��V�UU�^u:vvu�w:w�`�����@YL�����VM��	eў����.�d�X
*�4Mw�=�mHa�.�ʶ��e�{{V��l�^�u2�)A�6�T\�iw5�� ��w�X=_��˿�Ɲ�?�'��������27
ǋ�O�n���b�oG�6&���
�2�7�j���8�	�2fҋ�m%r�W(��ƾ�V*�n��I�
aB��[#��f*o;���y�j���g+{��w��h�=�L�.Ps���4���r*:�� ��LU�A�����$A@ ��e����#����bE	?Zt��-�4��|*�YaS���\�ç9�)�lj��0��)����Z�E���7� �2>::r�
802Vk4�����#��H�KYQ������:�O�Ot��QfP���M���/\��p�S�\�Ec�,�O�^�h�)��ۀL�M���R�-�����;���h���7�,Z��$�Rp[6�6)�l��Iq&��hn�k[\v,;_Y9��/�1+Y�
����d(�\\_ؠ߱�fi�墆Z;��5�Q���j���%˦�vuֲ�>zl�=ngX��	n;x���/�L��S�'vqղ�̉5�ۃp�Z�0_P�Ɵ9(����G�8'kʧsb^KT1��&�W�-;>?�˫+iJU$@<�L��tJ�,mJCz������Fɮ5ϯmwh;� �s��؉ftg�!i$�d\����F����\���!��	��ŜE�9�6ֆ+���o�u(�esӝB�y���?��ל$��v���?������Ǐ�7����D�6$ݕ*-kKF�V��:uS����H*�W��D-��Xb���&a��5{�~`{���W��=��ϏU�R>�ᖞ̭h�C�Er��Ҩ�ԝ�Dnח������*�̟��|��N�������@F�)#�
��<h����@q�B����&JvLX���!�S���]L+�ޗC���>���P2�	$��SO|NF�>����WGL�1��OJb&o�뫖vĝ@��޾�u�9���s7�έ$�2�[��!PFr�`enїB��@���i�su}a�N�#d��%7Y��?�y�>�K��Px��D��l�������-C��K;���X1g�b�f����[nUm^��*��5U��ڛ��[m�tG������J�b	+D�VHe$k��`g���|ҷ�|b�r�v�+�W���X.�=p�8�#�~m��{����p��Jp�P���H��Z*Z���&���{3;:>����t�P�j�V���ҥJ�
��	/^���'j��G�f�j0�*U+�����/�4�����Ӄç"��Y�V�;w��hj�����u�0 {3���@O��.�p���ٕz؈UdE���"��D��&FJ���{S.#B��
LXs��%�[�26���V���3LtK�Id���R�_(�~��_�׮�W`������w�a�d:�sG��?u2�ۑ��s�bC���O�%#�)����"+='	Ek���*"(��R�ި��v�b���>x�}x~dXfs�O7�[�����^�jە���i��C@��߱��ʗR��2.r�KdS�AD�A�ߵ�&���Ʊ���z������t�&bpĂ
U.VD#�A�(�X��Y𹬌����c�I�J@���s*�����
�,�M�Wf܂��/i��DK3���d���x��o8p4.J 5�;=7]����\O ��=�%�N�	[8���1��� ������Ȕ��i媾��95��ǹ�v��o;ͦu;7vyղ�n�RՒm*�Vr�Nml�(۲�7�gԓ����Vݡͮn,=Y	$^\�U"IH�V.��}Hy���۰k���ꅴ�+Y�F����Y%����]�� ��|qn���}�;�`8W�|�L���s�o�jŦ}|X�ֺ��ӣ�R��U9�C�v$��C2�V�e�/���gOl=�8�DF/~�X)�VsG�S������%kS���)����={��@�(#Av~%W��֪�鴮�Zs���*"��hj��+�n\��G!o��{�-8������\b\�|�lN��B�bI������)D��rà�7Oc    IDAT`2\�r*m[���~�����~��>���������l�g�����ٴ_�F�6��4*p0�1�晰��fF��t@�eS�7
n�M�rˈ=(7��ځm+6�L��OۇgG⬊��\[~�4������+$3�;"���'�ڋ'�uܘ!̴��٬l8!��#�:
nLC���j�����P�Y��,�xD��5@9x^�x�`%l���N�!�p���5�cASXi����A��?�=�ks2��'�%�gđ�Q�e�p^a�R�@�؟��~��� O~�);��Ӛs�)>K�*Y��[�.~�j>�x���z��4���]Mpen�LƷ���T|o�+���!�i�t⮹Z��?i�1LX3���W�ۨ��U=o7TK6b;��E�3�\jj��V~����V�l���K�+~lԷE�c���ŴU�	K�g��nU����,�<=���~l�|��Mf��"j��{
�[��m��7���}����:-Χ��5�[v�@�TQ�Xw��]�\I���gO��Eb�J�ԏ�pSokgO�	2B�2%�N�Y�,�ϋ)��k�)�~��j��ŕ���l�ͦ&��%��+WJV���aT$�8ln���J��Ҩ���_S���G�۱��3�����g1�X&c�|ֲ�ެ:vM2)��M.c�d�z빝q("�n+&�VO�w��_y����쫟SY������������Ӌٰ�pc[ђ^m�Ɗr @�U|cs���R����E,��*��Tv�Ɓm�k6�M��O?��^i�Y,-M0��-�cSp;�6d�ֹ�R �����S�裏��ʤ�Պ\�,�t4(�Z-ѵ����ց����y����ɡ�l.(*"d8wbaӆ>��&��sٖ���`(���:��H<'�){�'�t (����n�?�Q��	���N�,��
}5��)���z�ۉn&�ԇo�����
�2L5��ޠ:��D��4%�����l�u��� ���^�	�n���� �)!s�q��Ԡ!�u$a�b�����kW�R������=�`aTz���ڦW�����ږ�m'S��J�*���4|�ߵͰo���j٘��	�F�_I��N�v�u��{��O��ob�?}n�9��S;8�#��^s˘�#z���O�ً�L�K&dPs���v�ܐ(�b��Z"�JБcb�I��Y��5�4)������ى�8;� ,� �&�7~��ݽsW?�`6K�;�>�]���T!tJR2���wM�'/����ɳ#'�P�[s{K�)�r����T�6�����z���:1ThhkR����Rn�G��_/�׶(�1Q�t4�rrX�~���O����?���_����x�n��/����z>�r.��7�cqy�[��hb� pJ1hM~�����ʶ��u`;��S�����'6�,%Yǈe8��p�2�N�n�պ��̗2x����޷������M�lx�9��W�◂"�v:����(M���9J��uR�]�ߩ�乐!��
�q���n�_���d��3B�{����\�8H���B�w��ɭ
�4H��6;�<��s�+��k6�
B����8j���-9�/��!���8=7u�I�krY���Ʃx��ʌ���CBd�3sL��p�zMJ{=��\�������s��l��ڸ��a)i�r�F��M�I����6qa��ӕ�N�l����É�F��h5pP/&S[�f���Vsk$cVME��NX)mvo�dw��P����᷿kG=�ӧ�]E5Y��LÄ;w�؝�}KD#�&8\�؇�}f/.�Ĵ�^���;*IU����'o����ե=;V�n�XY��V*9t��Zò���C{qun��-u��m�w���$�@�Mj�Z��e��,M���_~��Ւ�-��Dy0m��u[]�89Uն��m͝m˕�6���؁�
�)��_��UO�AUU6W��`]��ØY��8�؋�kqpS�cq�e��[�_x����}nP�����-���?s2����rV����+���fI7�Ht)���(K,T��	�,�ִ���
n��-m��O>���?��r.��xb���b�7m��+Y�߇}*眫n�ط{�gvf�\��oLZ�-��`ʆl���W�-�$�]�J -��6�֒Z�N��ps���N�S��|��Ӣz�;htϽ��N��9��	�)�l������_���M�S���������SW�t
�t��J��xRM�3ї2!|����IT�ʴg��&CvJ=ƽ2�T��&��[$Ϻ[S&,�M
�e��A]��g��m��_���>W+t���z�ʭ$���2	n�1�<Om9u�K} ��n0Z�RQVx��g+�	8�]V�U9��ߢ�ݒ�ib1W�p���f��&��}���ׁ��k1�{�E���<y[1�N<6-�b�c�*KBg+节��`*�d�#��,�4���p0�7�Ä]� bb�V�mv�B�t��)b�.&�\ӆ=[`�X `�Q
�p�J��#��㰖��QCl�	���7����#&�� V���2��?8���s-�n�����XWq�����K�k��6B�h�������u�&�{NĤ�V�G
�hS�Bg<B��dJ����1�O���	�!���h2E�7����˵H�H�&�=}�T�y����L�M�?$���`*][�ZE�QE*����z�{�e���AOrHYr� ��JIf�pca�6.�����#LqN�""�Y��ҏ�{��Á
W��o���o��n���j�#����0r���v�
gB�����	�+�u�
��b�K�pZn`�T)�Wo���%�+;ާ� �XJ[��AF�~%��)t%�}1��^�y��(hO'���F�y�L6�]L�J�nWtkj��@(�ـ�,��U�7H��;y?ȼ�b�$+�J��#�|�6zK�ZT57����B�P�Hy,oC�W����S�s���ƪR�м���* nP��ל������H�S�2�j,JR�w��Pɧ�mu��c���x.s5_k0�}�AY�&�@�W++7��6�ع �Y#�@�5n���c.�Eɝ w@y�QSLƐ��aF|J0��`��`�h+�
3eJ1��2V�5]<t�dK�s����L2|���l��v��d�D�T�\O�j8>ك/��y��~��CX����	������=4�MDb1t:]�_���odʪ��^{�*���T�{�J�����{�Z]�RJ'3ȤHr��e���?�����Z�$-�RF��l�����a@�P�+�Vg�:��5E�i���cd�I��)`R�Ֆ��`���i:��ViTG����3�������C�߅�X���7
��v�f����/o.�[�Ꮔ����b�~���ώN?�Bᇟ��Rǚ���5�[㵛X���f|�X����|'�V����X-Ŏ��y�N�c�|0��/�F$��b�rU@�����\����9�H�"�
�T���e�F�)m������W����LV�lK9{��Q�@$�� �@�Օm�h4�u���S����ܤ��Oޝ���G��W<�m�m���������M�)	
z�`r�o'���s�2%%B���VJ�̤&
�5���ؓq��Y@S�l*B�T�v˱����� ��(�g��_�����|~7�تVµ��x�<���U�����*�1xVH���X�Tv���[�`�5�յj�W2O�Ĵh�BN��-d�*1G!#�a#�u�zB�x|�G���|�bxu���D#��~�!f���r8v���f4��t��4�>zZ���#��	��Q���~�3ؽ)�s~�Cj)
���s�ud�Iѿ{���^~�
���W�^-��Y�V�*;��H%���[��>b4�!��#�N!�߉Y&�$� q���	�3���� *�a�h�g�X��P]�M�:�R����SÒל���r�4b̧��}�yg�Ώ~��Y���F��R+c�`O��������]�����������L2�|��8��ri� S)���%�cLH�FQȤ��J�N�{?����+F[���i��^��5���m��@X��q�K5� �wŐ�X<"�`ZS+ƨ.!
nw���b��3xV;D�P�^�^�M��D[G�hvs�����{�qu��
ܹ���K|?�����f�X	�юœIq�O?~&�?��a2Q�l�O��(�rӤO6�^;�X� �[<�E���Ubn޼A,ť̾s�P�jaU5�~�ؔ���5M�ǣ��`D%@���}J�hة+��o��HkM�fi����ñ��%o&���e��eR�-�E֕���2X�Ұr�"�=���ǒ�V]̨��r�k��y��htr�%�&"SB���7Ǳ��ce͍Oh�X���a��c[j��nF6*��xD�$!sĶ4�M�����br׆9��j�\=��ra�]ȹ�f<�f&�g�<9��v��":C�������b;��5�]˦>Q*�����6�e2�h�����.�^���(@�JFł�R+ɒ����j+������]��H��nq�G9�DnV^3�.p���!S*I�%־{5J"T�=����5�\¡!)�4�yrH9_b��
[_H�'���*p��2�X.�Z����j���ܷڸ��E�ے�����6�xF��r�LV,��o��� �F|���Ԣ��������������}7����_[[�����Y�~���͞eČd��TyR=�"ORa*)_g��M���(-i��6 ����!�GO��m`�<\���5���N�р�?Ö7lK���~��r[ӑ�/��|s�[�����yY�tJ�dV�hQ.E�yn��	hf[�gBg�׫�&'��[K"��\��e��=!8Of��1fR��|�K��s/��M,�d�N|�IT����;G������S*J���y�,���:"@��_�	8*���܊@��Q�/��jH�+Fu�j�/%�8��T"�i0`V���.�v������7ź��?�7.dKJ��mԽz�-_/37{�R�^�o'S�8������0`D VG�R&���06ܪR<��'�"}� �V���C�n�D\f�ܴK�I��)�B��m��N��a��2{5��#�.���/���b.��	�V�^��'/�٫ßN�������7�x��Ũו�A2E��<J{�5�/�$xڱW�����N�^T��-��0��;�����]o%�fLW��
!�[2i����),H^/rq%u��-|��lC%�
��dDfd���B���-��CGX7͇c5��UH�~rE����R�x2T��lJ��O��t1��baLC~�-���7f¡K%��z&���~�?�`�GJ8?����-1s7p������խ����1pƚW��|�(����D=�Ó�#ԳU,��Y���wbIM��-�~�B�ݢ����O�q��?��d&�A�<��B>���E2�A�W4�r}e��6��h�+DV[G��x�����<�(��
�� L^�<�@jV9xM*�.{����R����N�m��m^���:����rPe�F�vʐ��j���V뜁(�T��-9<feŴ&���)��R��;�� �)&<NE?Q�YM��q�qDv�T�'���tP�J�ƓFod�����=@g�J�TPc�~����r�&��+�vi��d�tD�y<�E��r2	ر���V2�M)'�:�T�;V&|ɱ܆�uG=�1�tEKE@�\P�;w��c#eۨ�W�[&�B~e���d{�"j�"8�ݷ�>����g�8�B��\,�C�h���@�V�/�z�C����W����c6�H'�� S̢v����	��"|�\/l\_\�����6��1\�D��A�f��:r��T��y2�#�@C��z[O�
��1�`�9�M��\c�d8!U�蟷+��ŜpV��S�ș�a���0cw;YT��)�0P�@�euH*û�9�{�j��b!#m5�!��),c��� ����1z�\���Xl^��胂��s[���9�����\���pc�a`�E4��q������6pyU�����;�i�+��T^$[�A��������Ybg;�6�/F�K����'�PJrH:@��A�f<	X���m)y7��ڂ������s��Gn�(�b.?o������Q,d�k̔�y�2[3 ��!݅'�^�D�*=?����~陘���x�E�P[O�<�6R��`
��3w�{qz��0�<�LF���&��)�J���5]fǲ�#�C��0�dO�����T*�"��I���v�~�n�]T�c@�S��T%$��7�z�A�2a�/ �����Vg:���%���c���l_,�0�l����hw�+���&�JE$_�'��ĭ6R��7~$`��c���l�C8E*�E�T����a�FڲPv]�9�� �r�޳�ky��yl�%��h��B����N��}$�Op���H��&��}�ޛto�M���E�)�P?=���H�� G�9.�\���5:�eso.��+�Ѩ`��HZO����nuP�C�(���'�*{5�E2����Dq���pvlk]V��\��w�@�^��s�K0g)r-V��x&�R1+��b���F��w~��:�)A?E��8ܫ	����U�Xf��Y8�E$��v�{s�������X�,g���O��o��ʇiK�P,�ߺ7G�I�2�O>n�v+	�l6H�CxR��ZG�!'���ib�Y
��4�����@:Fx듊j����aÓ|H־�b�0�ꏑ���K�O���@1�Ĵ7D��^�ٮV�G���R!�Ѹ���Ɍ�I%S���dއ�{q���J�\6-	�|^�Z��J��E̽_E	��9�m��ig]5S�{�RP�֕�T���y����T�u+�8�X:��e�ɡ��\K "�M�H�'	���Ȝ����e�\��g�E����C��^[Ma>��u{���c���'P{bj��Tg�w3=!��ӝ_�̡%����㸂�nPsER4�mi*���uD�ʚ�T�h��c� ��J���'�d��%����S����7P��Hl�H���>�}k8@(���)^ʩ��� b[H�&*�%
�9�#a</��=A��BqV3�;<�:Ǣ=k|V���A�^B��?y�d�Ds3�|6�y@����GL#�����7��=?�����bQ��p��[ܼ�@����h�M���<����g���g�"Y������Zw����2g$͉���AC���T.�s�T���r�ٜ�GRw"��[ݫ�x��ӲŪ��^�|8��jE��hׯ�9��|0L��w���|8�o��ϊQ,-�|����>`�7l�`-�!���W��U�f�᳽����-��gZl�˿{g�Ӷe�����%�;*������?A�'�r���
��+s:�I� ` �v�JbF@����s/w- ��pzC$�5>)5�����E��x$WJ��ZR�I���-RVtl�dV�;�ʒ���R�9�C%�f|�P%�t�M_O���.����ݐ�7Ot�(�tVGlG5�iՂ&��6:]�?SvG�ws7�iT�(3)O�O�Ἃ�R��a��/��\��en(���`��V:Q؊�����'+=����0൪��Ǫ���7�8���i"���_Iˢ���	7JR��ǿ�=��(�y-��ও$fI*gBUH��J�m� 䌹
���3�;��^qj��siK�Ɉ��l�	��9�98�ֱ �A��	nhB@h@��"��w}���-��1<�����n��4�t�3,T��O�|\*�ϞH�B��52�����W��-���[c�!�(����?B,W�a:I`ty���T�n��d�(5Q}q���c��M���q��\�<��%3c����8|v��/>F�� �Y��޼���뷸9��b4�]�N��8�nMȾ�i	o��a:��'�
s�MJy�dJ��,X�1�jj(p����i9�j�Z���|��~Z6/P#�ۛ�g�B�UPȤ����֏)Z��`�)�-E��f.�q�93L��b:��g���7>�������wg��e&��O�R6��T�I���)~��r�$f���T��k��b��ʕD�d��d    IDATmd'�}��)'_���	���s��<N.��D���pǙB�9]V.2�tq(�ZA�. s�B"�F2�FR��i5CJ������=����i?���#Vd���$8�!X���I��M&��^X�^�YϤ6[U��/]�iN�xhy�	��7-�"��+�#M�U��\G��R0�*-q��Ԕ����Z��[i���
h� @����� �w4IX7�OޗV/����^�-�~>�D�{���y�@ͯ��'�R�=:�r��&1P�5n<~/S�y��[[���L:p���I��+��-g�+g������S�\���_lO�vS#nK}�\[���\�lR�c�o�u�3-U��'�4�S)�3��rI�T�[#ܿ���+��8�b�]"�l���c�<�`*�}�l���k���0����[��*���	JO��?l��ˊ�����kܽ�0�C���
�N������@,�W�/p���o/`��HE�==~���=d�%�r�-[4���R�0]B�6�8l�!W�0����4�j�e��n�D�M�l�V��AC��l�n��^������Q4+%�3Id�1D��������ho�n���!2GKN9�����?��&��̭eM���z�Z��@�X��^y��n�Z"���໴��$G�*�����d��a���9\�%nв��Y~����R N�{	9d3�.�s�up�/�&��C!����4C�B3!�FIDś+-+�d:#�����"���^K%`���񀹌g��<��﷜Rq������ �[G�6�����2@��&��>�f���<.=S�le{I�#������ ��s�\��R%�VR�*���T��RY*<[R�sxU��u;�]~y����F$�r�J:��&���fWm�U�P^�ⵉ�hY��a���\�PdY�T*4�y?t�LS8��l�TD	�BkVo������%��]p�E���`571oa��X�$�����ā#���ʥ���Bz�@nj�f[���ǧ�
����XT6���6��9���5��lW[�d����>�`��z��ͫ��_����4��WA�g(�!IZ/P�5����~�����c��5������Z�ı��q��
�o.�24�c$S	�Jy|t�R��d���X�)eTCtzC��3�j�Я�QC��D&�����/)V����5�*2�JbHY����Z����fs�������sD�;�J6�Œt��_��g;`
a���[�֘��^bKR"���?��������~��k�������v̈J��2;��
�h�k{xRo�ImO,�C��Ba�vЙq���q6@?`a��"WR�sI��B�֎��4��l���D�Y!��!��!?���N������:���e��u87�:�r9������իW�I�Ғ�e$�L�q��]����=�S|3�r��.X]�:ANoP	���7��*�B|���d�dK�������e�w߬�p��3Co�~U���@�����}�<OJji�c�������BF�y1"@�L��uo|j�C��[&��b��4E��G^��� n��S��|1�6�{�{;df+f@�QX�(�d�l�ı���.Ϲf�na����B��h�|�bV*�Z���i �� 1���,Q�,|R,⳽^4ȳ�]Xx��K\�>Ǹ;@�V�z<Gu����c�=9�]l�h���������)����P>�C��T>y.�3�|�&_����9��7X���'�(�h<=F��a�4�~�GZ/�0�~����|�p*�\��Ƴdke$H����g	��;=��3�3��T�TD��P,�≄8�0ǖ��w���E��H�e�ptr(��k���`>�����hЁ1�¿Y	�U%��y$S11�\�ic�Nc��εqg[�3_!(��e)��g�}��������/Ҹ_N������m��lKiR�M�j��r�l ��|��n��#��"�(�7���o]���6��lmI�a@?)JP���3��k�;�_���O�B��~�$b�
QZ�/׈�H��B7`�#z��@ҁ��2��{F(�b� ��ъ�s7:�L��>�'��g��+�g�#ٍ$*�Y�'��z�}mv�!�nE�}�c,Oz�R�{G���W Y�{�&�"/Toa��PR�s9�tZ����
����E���o>�<��&�f�}�
Lxna%w�kEp�~�l�*�']���ˆ6��HQ#xQ~R	!1�4��J"��4-���.l�ʇ�V��W����	&�9� ��v�$�h��2QlRQ���*��a�2YY��]��`�~�ppG��A��C(�>�~z�-�ȸk$�&r���i�Y>����𢹇|,k2��?��g�������d��}�?9F�� ��$�����o0�~`��p܂1?OOP}~�ҳSD2 �-�_��sv���-���]x�h*�j����2�GЅ����/�0�}���2�����WQv�T��h&��d����rAa��;�О�	n۹x�e�R��6��~l���]Z�Ϧ(�r(�S8x����#Y⹮���h0���F�6��^�};�*�22�����h1y,��4ƽ��~��s@��e)���������7>���_��^o9���9�w:�"hl�f�@� ��?�dF� �\�T�t^ldA���1�X,�8<�=S�6>�P4&�O	��p�fIٿY��ϱ����OJ�Gl鸻�"-����=�a�^��X���A��9)��eɊ��&���U�\F�Q�Ko^�n�N��

����QY��R�̼��s���R�DUV)�~\�4��JOX	��7�F�=��<l�\/�2����9u�W�ɤ�X�rK7�������R��\1����
Vfo^��<gRM5��2�K~��FҸ��$>��J�y(䗙�mbm/��,ȟ��65ĴΙs1���e�bidp�V�"X�`C`�SP.�>?����h&�tV�II#a7S�!��c�gZ�
;���0k��2Waj k۲Xx���{��p���^���粡$_��+�*��e�i<yz" Whԁpk��˗oк��AM�҅��������G� $ˇ(0�q���2��tZbC����%pp����R�� 7��
��
��G�y^-M$*�}t�t�e���qʙ����G:�F�Ԍ-DF���[*�p$��r�Ao���;<�<`<�4f�V��6�nTU�H�8�k,�y�}��a���d �]�ry4M���H�pv.Lw���v8�I8�G�\�i��kozY�g��'O��-~��ͮ=��wF��u�Eh����1�X�a#�V�� e!;?��,�+��E��Ƞ��	n{��k���Zyj���ٗON:�ă��j���5ͅ��&�HЋ}�ia���l��1���:;	N�IE�Md��E*OvΏؚ^��U~=#��r�уJ�/�Ei�;\�����H�w��+�����Hd���]2$��ύW�uU���V�7�
z�-<& �	�����Y�`x$c-��n�X0L���ȹ���T�x��XL
��.��]���2ó�
T��A��&�+_P��E���_N�v�3�i�b����'�^^�䞌��	�`Q_�#Z+`�I*2H9b@J��]���Qo��`8�&��?&mdj e/M��(�>+W�Ǉx~p��k��������h?t`-LY>�݃r�b1��^<C�B��H+!���k��X��1��)�0N����}�	n�lMp�g_`pw/\��f� �4���v��D� �氚��]?�����x�`� ��
�����d� _:#�qk��}��D����������"$^Gb�,��7��w��)���z%�R%��~�JY
��a1ui�4�w1��Ǯ����♘(�掋�vF0�y(��f��z�>�i�Eg�n����ǧ/~�7>T����3�����kcZn��W��R
��[�Yz��H�B��ɇ�8(װ�� Ð�@![T��Xy=�i/��?��?��c��?���-<\\��$7��#K �D&Z`��� ��(����ᐛ�x��]x�����l<A�w{����!ĺɫ�x�2D��ƪPY�+�%���1W��o[2%�"�H��ȹp��w�M����բz�e������"�*����6���c��9>Z�{m�n5D�W:�Z�r�S-o��Ĵr��' �ce�X]�I����{���ڊ\���CW���Z����<3~p:��m)bֆ?(�\(|��wn���*���xD�2n�"��b؆����l��k���ᷖyV�2�Z�x��.6*0D3�-B�"s	�B�;Dzn��t�i������^��L����s!J���Wr#� ��(^|�\fQea7>��]�Wv{�(���nOE�ѧ/�
Bpds�2몃��3L[=X�1�[�L�z	��Q?�G���Jc�����|�G���P؏�A���l`�~3��
��!.�0��:�\�S�T��b	�JE쎸��9+�;n���4�]M��B��A�VD�ԕ`Ғ�^�`�QU�c�E�R���[&I�6/�=�1G �`��m�E��H�#	�V*��/�|��~��ү�|�q9���|�k]c6]u�c;���(������)�1׏\0*�vP�K�JYή��R,�Ew�#�c�VE��0Of1;?�m�p��%n^��
��"�YrE���n-aNXb��8��o[b���FגD��<E�j[�����Ź����H��9`0(rn	���Cً���j�J=sS
���[Q
�y	��RVn٬���څ�'���%������,����MD�������������#��0Y���z��K�N%����RTZ���0B��Rn7��^=���i�<�MW�J��$j|���f�RM1I^�z��M�����/jZ= ���$m�&��X@�/�y���� � 1jO��"s7r�)QsKQz.��{���q���'[i�d�."I�B�7F�\����;�^T�h��2{y}�/�x)���RG��
���G��|���Z�����_}����r�H󃨟���'�P;�G�`�L��ww��'��f�i-�ݹ��WP���������nm_�a3] �#�|\G�YAn�&9`n���ઃ��;�:��ͨ?:�T�5�kud�e��q!�W���Ad`l�iG��ֳ�A�V@��6�� ��C��G�.&�.Lc��������#Ԛ{�R���M|ss���0:�-��B3Ä'��[.��;��󃵥����L��v����9�+䫑U�senf�N:�|"�t ��j���Ar�G#WƓZ�bqnE�t
���N��7b������]�;�������9����9;�raJ�Z�PF��%g%65"��m������"m�"r:�s�)�+��	���/_��ؒJ�iX"���A}�"V:2{����OҢuCrO=p{��%��`0G�{|��15x�g�xdګM��tK*6GA����Kp�-��f�䴆���)+ts���4�|6'���\���MR��>{��Iɼ?��T�ތQ܋=�^�?M*?i=]Y(��Z����r��}4���g��<*]���\�@���_�HQ���\`����FR:d,�H��D�b�R�L>nX���a�v�l�O�5Q���&��&(�.��^�8�P�e�+`>�7/_IR���h�"7�y4�ѓI����8;;ǛoΥ�g7��
�HH��O���yr���p�F�.�\��?�\>��m�\��i����ST������py���ߠ{v	��"E�U2��i���u�B$���F���g��n=-q�ϭQC�^k�*|�� �='_�^2T���3��a�zYL1i"�kt�uz��X�3l6�T��j���ͺ�/mt�3|qq��6 #A�Cw�b�[cKC�Lz].���֏��F����w}�.���b��w�ydF&6���=^$��T
Yr�躻� �	�K��-��/��. �|R��|i���e�g�(��XD�a����"��׷x���?��x�b<�R*+�Yl�7�%37j�ș���h>ň!�k�B�u�
�IKGyOR�to߾��� O�D�հ�N��NƔV��+=���j� �u��7��p	n��R^�~�Xy�*�rC+x���n�Ҷ{���
����t���'��剜M���\u5x�6�?#�Q��� �cd��L�m�!����-eӤ�y���3������d �W��[��hM��ۮ��9k��|��e8����lS@��`&������'HW��.&����E��eT��@<*j�B�"�K��8�~~�>v �׬���r�4V�,�ܲEg�Sz�e�(�R�N&x�tqvv!x��7^��!?��%�+E<9<@�T�M���K\�_	��[bΓ3��4N�����2�Ak�7�����L�+[�"�B����}|��J<_n���K��|+ˇ/^�S1�=�G頎��X��X��]�pw~c>����w���ZU��T��!��n�>�����۵�h�7+�;i�\�H)��V�]*/����t�Y!����l��CXX6�c|~v���3��;tyQe���)�]�ҙ��t���w>T@̏_��ڛ�f����9��w�g;����&D��+�����p��*��1D�FX�w�掅�c�^��>��Y�Ц�n����#3c.&�wW���#h,�DQ�&��
~J
3TE��e���v��6�L�漉@E�B2�N.��^O�!RdS�S��liEs�N=�n�z��\ϩ��&����&S��~���x��X�l9�"�B'��xz�o�G��Ĳ��*7]jAJ�j���d	�zs���ya�ǣ�C�������d�_]]���n�y\\H[I�;{Tϒ]��Tk^���}�b��)yl�מ�$AY�+�K��h���t�p�a��^�d��.�ٚ�� �M�|x$�6[���0%�+Y���"!1P`F&�5I`�̎f{�����G׋%w���Fz�"�d����h����~"�&�.t�5l<�������E��o �l�2N�MĂQ�Y�}}�G.�%��+�pZ��5�t���>N\羍���x��[�R��l��*>��9�K�ŏ���9�XE�M�>ca�A4�`��1������u��M=z�s�8
t��ŭZUr1��<;�j�����P`'����}�(�b��n`�V<t1�,o>�Ҟ2�d�z��C�
14`(�]o��.o��G�`�ݠKL��4E�Ī�+���������}�PfZ��G�s���Ͷ���}~�l#Wl1|�6��+�GH���f�8�5P�����d�qE�p�x��d��VʺgG/(���_ڞ�C�pL�I6���o�#��"��µ>B�$H6%�ML��R����@�z���-�_ɟb'��[���������`iøE�]����S�w�&�7�w�K�<[TO,/���2���)�c	�Q,*��J�@(�U��yL�_�|?ӄ�����荨v'���u���Ǎ1�!%;cx��q����H��[t}U�I�kh���%r� ƞQrU�����E ��!���K�q&H��ͷjҁ�s,O5H��h���B�VA�ԍH@��h!���IiQ-�Ffr!ʯ����@���!usvg��8�J���`���Ep�"�b���?�"�)"����x帲�6Zd����IW��-	���~��v���c���@�7�.��J�u6F.�ē�C<9=���G@8���+�˟��.�BK�PЇx"�J5��}���L�%�����뷒��J��P?j���H�8�[�^ߣ{5��Ӈe�drN�:����z��D�.�]�aJ�x���Zvȕs�4k(��+��,:W0C���+���l�F�f�lЛLq���G���[o���!� o0fW��I�����(�zX��n1����L��PAn!��W[Y�7�E���׭�ɡFo~��j�3c{��I����"j��i    IDAT�C��.?��落�]���J.��4��W�u&�OM$w429�QI��썃a��d(Qj9�x[�:r����V0&��6lIy2__\���* ���)a}
1`z'�v����⼽�y9�Z1�r��ß���#�����T\<<�q�{���[q��ykZQ��j�x�"C�u˸�[��
��=x�r���1%��gn�JЏO�߭I�%�_匒*"����}^�F���N ��G#16pL/�j�4�JvG�ӠlJ�z�m�N@jAw߀O��ù�d]:!�x
�{���Ÿ����V���,�q+�,Z@����5VKl�����Y����"=_#ҟ қ�ov�C���<��z���V�����S�L����h��j�J��
W痸8��|nʅ���X,�T4 �����x����n}���|��7h�wT�R:���n�t&��|�����'r8?������Q:�\R�*{���(��J%L��܎0��,�;a�ͥ�R���X���,,�!�NI
^�e��&<�E��C�YA�恛�¸3���p��9�� �� Q� ר#S���L���?��Co�BJ����]/ѧ��	&ާ�V%���'����?�k�w[����k;������J{e��1�:��0#a!��P2����'[��rO�PNgP�䐌%�1���s��ctfCt�	�[>����#,ɝ��zY�&{���*[=x��K��.6�)B��T�\9k��x?��d�'x�ӕA.Txo�8bT.D#R���C�*~���<����@N���i	���c*�NW3"#y���S_���=��~���"{�w�6�^,o��� ��k/ס�?�6��I�ע�V*�J�ƽ����f*�զd�z��PPU�z�(8�����W���d'yL�v�.��C�p+(R��h<�~PLͥ�<6��b�"
Z	r�y�-�9���"Ǔ4V�c����.%�	�ޔ<7~� ʆ��J�$��!�-$+G���0l��Ê2��� �p���M$�r[ K9g���-0�,�z)���<�Cs��w.ұ��"�"6�77w��@�3ڏo�tK���X�Nq��D���s_|��/oE=��
M4wk,���lK��$��}��7�mY��)9.6G�D�j	�7�\<$����+tG»#RG���U��iM#���.�,�Ɲ��\�b�/Ԛ��HT�@8�����=A��KRo�B���(��,2�V�t$�����.SX��xm��e��T@�V5����T���
Bmi���G{��u+6��*?��R�'���s%|������!�>J�63�t[���04�X`�u�����Fx�1�!`�-'���r�P@mr���W��,���6������d}o�+љ���X���J���$�ҋ���<iy����z:�H��QfM��hsͶM�,��G�UA#���F�L�ו��܏?��ӼU�*���
����y�7�0��R]9�@_6�J���R��r�G�$���ғ��+��W\n雷U���s��Z�%�6��K���7�NP�e�"���s7m\)3��J����ٯBΟD*K��{ϭi4�J����#lJc-L&Χ,g1�.�[�qf�s4J��>Xۥ�c���Qy ����.�IY
m=�(��n���Vl���%���D�-n���z�S��Z�͚/1[ذy��c���Y���[���(g3��tm�v�+%f�Fd�!-l���A��c�`O>#����h���2&�W
����6�ңN���/��縼��
;��N�l
�d�j��� !�U4�|����r��J2":�b�$4�\��`$�%+��)���` �U��@4�C.���Q��:����1��п�bxӢ�|K���\�rN��cU���������̂��=.-ٔ�S��4-ؕd�wj��?�`���?�ӽ����ѿ�w���`�b�\��%
�(�֚���3|�<B~�g��NGx�ў�0�-,vK6����fxp%W@1��=]����V{T�~غ��'ҿp�/��Α\�P��P���	B�����$\����d*<+�X��$�72�ecH�O�,�M�^��!�f��ɫ�-B�[Uއ�̿5���]ͨ�[���,M!�OA��Ymi����*�N�����k�4�����W��6]!*ٓ2�d�-U3�p߅Ψ-����K�)#��d2R�恡�N��ja"�n�Z�8lzq�^�������(�f8�Zy.��q�H�d\d��M($|HJ�2{UDEL�B߲�6grB������W$��{���3����8�[P��P�c���(7�R�Q�`�ߝ 025�i�%����]k'���Spϋ���|D}@!�@"@��mY��p7J�F�@�}M���ר����{���q��I��?E��C>�F4�GķC.����$�Qb2���%��Z��E���8O�!�I�[/-���,���>޾�@�;����k4�G8D�\@�IϷ�����2/����j�����p�pp�r� ��oV��� ��7A粅��#��͢�it̒(#wPG�Ґ�m�n���_^ݡφ+����Ƙa��b �N ��/j��O+G����*�������c����վc����p�>_!��\p{~pױ��MG�h��q1��a�IF�biJX.��7�̍$�Ù.Dd��7cf2a��z2�]��!���q�0�J*}~D1C6{�O(I'�'�툶P|�ݥ��^�Cp�F�*��Y�|:C�%TT�
A� n]	�aU9	g�6.4���	ݞ���K��T8G�I���ŅG����jꙙ�OU��7�<ꅖ�)J�ڲjw]5Ƞ��ᖶ١
���o�[U~JȮ,g��Q/�5N{o.�Tj�A�n�����c:K:Cu�P>G��:FUn;��1x�3�/�!Z��EQ�.	��pS��0&[Sl`��Q���vy��&R��ɽ�(DqIbc. �QW�)���H�v��+�zS�:#�b��Kq�`p+��C�&Y#	Fr,B~�C>d�t�وj��6�9�%]�	@BLH�"����69r�=u�cI�_������(���|4�r.���:"!:o�����3Ͱ�`$�H,�L6��fϞ�`� �b����ί0����l&�p�Oq�X#5Qi��(�E�O��f���pK�(��?i"[� B��0�O0��c�ؿ�[s�p���
G{(7+s>�|l⛋Y&̃Q��"�x�&��?�d�D�h�J�q���>�p�G_��G��?<.ƿ�sL��.����wf�!�e����)^��(�F���nǀ��
��J8F�r&w�m�T>��PF���:� �
��Ӆ�����K>�RL))����;�c76_n��EP�Ƒc] ��ҭ�a����l9�G���[�����[Hr��}�e���b:�,��ʍ38�Ex�'V4���bH�1�D�����&��Ǜ�i� ��Е�hD�W�W�XL�B&�H��O�O�����I�|����z)���ŋ���oV[�#a0U�cA�`!�����[�	p�Z�����*�*���L�V�ԾO�+8��IȖ=��7��LX�v03a�9�� ǒ��lQ	����҅�gy5҄v~��E�����by�s��kdV~$�6=�;Fpb �\���%�S,�%vk�E�G|/X%�(��Ƣ2�'A�ձiѝ�Z\�='�%�	6��"�l�V�0O$�v	���l�|�2�3�F�Q�V�:3���h�EB4F6�ko�$�����8���KF!oi�e�p�R�F�2[� Lk)�l��0gS1�t
�������5z0����0팰/�����`�b%�ړ}��J�i�:C|sy�o���i�
%��q��R��"�)�����r\�������g������њ��hi�ON�+�%)�oJ��ӏ����κ��[��,&�6p�X��r�S��
���\$����Xr��
�%R �����I�B������	LLM�P�d
�XR����2)<���3e����Km"PpH�PZ�x"�R�(�CVp�VחW*$��U8����T*=�Z�o���/��Tt�5����Z%��^(3o�]z��L,�|9�Y%qF�J��wޯ̬��I��j֤��χ��)T	Ъ�'�;,�Jl���U}�����+ T35����U�xo�;RnB�.���5n�U%��PX��^����ن�@�Z*��$sXA���h�]e��N%"5����`@^�q�Q��(5����u↗��VU�a��1k���Ap0�0�n8C�^#���G�#���|_u�^���3�����W�B�
�|�88��^?n�i�J5ys\X��HJ��,X��J���\��w�'��4`v/j�'#���a��/��;H�I�UՖr�asܵ��`����u��#!�կTjb?��d%��;r/��0���YZ�C���(9==5����B�}i?���tv6���T=��&B�,�n[#|}y���N&�X�<Ņ1ǔ��8g�!�R	������pp�[���A��?|�/NZ�ُ���9\�Ƅ��p�������>ƧG���Cb�ܟО�в��.�a���JDhA�6t��ʛ�L���r ��g2�'��o�p��7J�Cd�4�����F����ȇ�e��EbUē%�L��5��Ż��&sg)՛�&b{�J��-��8�Ʊ�ͥ��F��׃ojIil)��hLȾ���eՕ�V ����rԼIW0�M����(��C��dn�yM�1ռ�0[�o�di��/�u!�͵��&N�BD~`\����pQx�����?|�q������"�z2Cs<T	Y��Qd '�*��M.U���~�g (j�M8�u8 ;��e$�Xg�21�ѐ�~(�ߐ�A`#ǎ6��M�^lE�RV(|��0jr��y[����
�p��p*�#7�;�k�.��R����������W��cZ�(Bz�$�)|�CQ �	Z;�K���=#�*��w��Œ�g��NrL��p1��/@��` �-�O$�W*�89x���}�3pG��q"�>�L��U�T����Y�$:���v���@��HD#8*W���JE��	�'*��DxrQ��mq�@�V���>�NŰ�l�����Z�d�g��e��i<���3���A�dz��)����{����_�+�n?��_���?��O~�kσ&)bK��l���~��_z�1��w��,�7p�w?��a���d��c��oŶ�W�VXa1�T|�BQq998T2�t󵃇��\_�3c�4�"�o��v��[p����"� j�^�Enœ�-O�v�����[��Ծk^(p ��pͽ=%�Z�A�VʞXz�2V�"�@<�L{����WF$�����H��#�G�ǜޒ����kʉn���y�*:N�_�Pe9�<n����4J->�;F���zn������7)�@^?.�m���xK��%�D�:��|}e���zt�;/]+���!PJJ�t,բ�@�y"S�W?lZ�B@*
_:)��n.7R[Q���2Z���2��{/e�'"��t
�jyA�z���'���!v^KJk{n�y&ň�7��)i�d�C��9b�*A�VM�ֽ�m)����b�ʙ�!r&�z�u��o8�X;��!׿�ʬ��K����[à����U?[�P���C>�@�P�d7����%���Rnv����b�ʛz��Z��L6���Do������c#&//)�������rFc��������X|��2���P��$u~�\�WW8���&����T�(��b�m	g��'R�f6��������?��_m8p3�?����e��DW
���ǈ>.>=x�g�}�e
�����ږ�Y6�qF��-��v2K�+��C�B=_D����͞l_���g��н�{���9�M`!c ,�I0�%��U*aP1`��H�|�*�hI���ߐ�\�*v� !0h B���S�k�����<��u�(�ݪV�ӽz�Z���>�3|���r�V���+�ҳ'�g_�+�l�e>���YM59�_�-3���%��j�h+�1�E#n�Ή�Dvފ�GR���0S'Ǒh��d�Q��{=;���ݞ�	Ȯ�ce����l�.���Hp�T�2x`�$�}�Q����>�JSZ��Ƕ^�4A����Ȗ`bH�~�A�^J=�)�;�LDx��������:R�BY�k,$'�������#X��^?u�0|_�$qz�pu�	��'�49�}����&p�f�F�
��ՂmZ�V�4��9�?g�,���[er���l4��GiϤ�r�����m����kv~m��=e�� r&ȓ㯠�6Ityp󬖬�6���7A�!����r�g��!�甩*�I%e,�ט�d�y"d���տD�gy��$�=?�lN%,j�U�u3�`�	�kKVY*H~��R`wOϤ�v|r�~��'����G���H��]����F��v�_AoͲ��]�\�M�+_U(]�Ȯ�sa���|���������_|�^���M�`��/����.s��kz��ig�V߾�����ݯ���|�\Q�����A����������_��|�[�^a��0�gx�t�],�Ó����qz_'G�T���Yϣ�g��������:�؛m;�5��n�Ȧ�pf�vi�=b_y�Ծ��M�g���
��6��p��<]�FfHՀ(�6�8vXm(E�?��)IeY�+�`}m�x�%�� ��SJ���6���\���s��t�X1-n��߼/`L0�4�;�gQL�M7��MY�~�L};Xt+�t�b��':�g1�L�3�=��2hq��X�:{����E�U�@���e�K����᳐�2�7=%(�-�aQ�PP�����it����1�h�4g�O�|�rG�e�6aW�GX�%�J�v�H�׫��`"d��!}��z9��3���@@�˂�)�������C�,���ϖ�R��P�-4u�"s �y��"�NALmZ-@u��]�!��ָ�ޮp�B�WJY�h���&P)){p�Yl�sm���
��%�Np#z�*�0�X�ժ���#�nP"��W���2#�E��������w�ٽ���˯��J����z�W6��Z,؝���?9��/�W��4����������
��|f�J�<�g���e��=������ˏ��hj�R�����m���6�� ���rR������������~����w6U;��?�?~�ӯ<��>���������~v���
�[9���恝"X�:�Y"��ە�լlSdƻ�
n�r�p@���;w�}h�"�%g[��lh��7��o�n�n��Y�ڶ�zŬ�g�:��:%2
p3[�F�9�Xu��rȝ:��s_�,jz>0"p�Eo� ��)����4�ِ��B�da�G-D|���.�T��h�z�X|4w���m��	�׬Tv�/�O}�}����q��`¿�.A< ?��˥Ґ��υP@��.1WL�����1
	)#�v&~���T7=� ׁ��&�y��PV{9���Z��[�m2z�AḘWE0�n�@X��mV��9��x�Z�U,[���[6kѫ6�@�f���2O�Pɲ׸�1�%0�����`f���*������4�=	4D֚����%�1� ����ue��I��ћ��A������"��d�ku�\p[��f0M"��^ؼ�TW��p��r53�i�'��H�KԀ�++���ʻ���=)��g��+���1�iU�vv|h/�kwv��՞���-�x2�
Jۨ^+{������4l4���K�wo����Vz�[;Ϛ�1��
2�W+��y����W�'��o�}������}��g��'�z��t:�_�ɭФZkCs2�y�+�hY�T��jU��a�f���՛V�m�Y��td(��)K��V�jj�n���jf��~����2t���s��糩d���(���	*�7��|Q�zSXI"�e��[sx�+�������L. Y��֨kAv�mH�vL/�e
MƲ��5�o    IDAT���b+��w\@2iĕ�M���Pa�L����i�+1�S�#L�@PT	u���2��<<S�ů9��U��V����E8�ň(U���<�o�c���z��jKQՂ0�?UU�Hv��q1S{�5��S���$��Y1#�A��a�vݲ���u���`���w�>�|��������@�UP"�.-?���U�� 1@οp�֜o���Z}�Q@pÉ+�ge?IYJ��kf���s�2��)'�&2�WR�O�zMd��)^�8��H���gU�5Vz���]JR��I�N�7���e�����&1l@Y�R��tf�G�eZ�Ygg/�a�#ț�߲'o=�0v�f9��f�;F�#�YԛnOkh9��ِ�iW�$ ���}{rym_||n�����ݷ~�j���9�۬��A�ʹ�Wkv���O��u?����k/$��� ��~s���g�aa�]KrF�g�*/�
֮�dCj�o��Ұ�����:
re�,gK�Rqn��`����A�F��avcϧ�^��|ԓ��t��"[�����N?Y�f4a>n�˞-nzV]g�
/�X���$�]�-�˞���$�=�!'e�6��� �K��u�i.=�p�w3E��N��E �$Pe��0#�Cm�����&�2iJf0�����&D��T>�k���x��x.��E�
�-L�SpSB����<�Q�iJ*W��D"yn,��K�	$�7e��F���5b��IN �7�����%����e4�rP����f����3���$�� ������H��qzNXH*H������s_d���h�:� �O�<�[c��e�t-�\��h��6AS���[��;�,���b�I)ׄ�AvD��-�-��J�x>��AV�0�� #���R�z))KD)�d�P6�D{��r�3?(@���N\o�,0��e=�X�V��߳�s�^_ʲ��z�Q��Î��tdN`���r��l�L� �4� ���hF}{|umO��ʶ=�X��ݔ+v�ڰg3��
YgVfP����}/��S?�-���/$�}����w<���l�O��G�Qfesj}j~p?�2Yq��M���,6
6�l��ם�l����!4	̠jk�	+���a_x��6�쭕l]/� ��c=x90r�#�]������s2��pj6��<%�1h(-6�"�.P>Y$�lg����'���M���J����	zIz�7��7��SI7;_�'���F�@�X�2��P����4��pŒO�.O&�&�:�M�/��|�@6A*I�4�}qɄW)�^�B��!GP��e�aŘkK�J�<��28�W��\��?��eI$��B ��ÌI�{<��mS+�K�OV)YV�T/�"�3�xvy�F������$^��6Ye7�m��M��P=p[�j��� �<3v�6*}V>��P	(���1��^!`�W���"�9������
n��@ځ�5��UlP�!���~�y��bM%�J��$݄�f� ׬��O��MX<����&Q�֠)�>!�Z-+࿱1��phJ̈�b�ע�1�=;9N��O{�aCkѪV󙛤���咵��>l�$�}��z�����Nl�nY�Z���/f6�.e3P�V��K��'������B���?�;�<��?�x2�^27���/0��B���G���T�{��W;)7�~�Hd�{�����ɽ�tR~����ϟ�Oۣ��6˛M�����,e�<��-Qf���*�L�Bf[��N��l�٦7�,����^O��X����CS�Pp�1㜪lBmr2�B��Zj�j���9��A�þ�+	K�g�p�,Nr;L��d�`�=�SyYp�����d��$ˁY��E�OS�r���{RGj��|rr�m��!!��M��&d�*ˋ�C�D�������)�.�-SY��$C��CK/�78%K���u��٨)�����ЊY�8�d�䁌�N�s�C�ߓ8%���/JS6������tO��4�4���[��S�Y�` 4a2���N�
|�iɜ	)��	���]NP�bH��������C���|%�$Y6��ua�]"��]�m�T;��a,��+�"���{KK�Âl,�*�nj@����U�L+)'�q��	n��|�?�^ P񾩐����:|׎TP(�i�PF�,�}���j��Ȥ�r��J��~��P�����زղa�*�����F[��ՊN�|����{O�}�>��|!���{/?�~�Ѩ���&�"g�]�TY�Y˅J��Z˚ټ���)V�^�H�V����q�>停�\�������wcO�.�rط��u7s�첦rx�h���
��XiAn's3��pj��H_W�&s��vX�[�\�M�Df��Jn����)t}s��7���FL@��V�l�F\�}�L��$���'vy~!�$�J4���X��i>���Q����>�/�́e\�Sq�9����	V�5L���21��E�㭷�;���W���b|'��M=�0�!$h���qdeLH'��������{ٖ	�MI�~�Zh�1�#�9=�
�=��5[�A�m�Q�>(z_<�x2��CV<g��g���J���A��\F�>�l
ZGL��m�곥��Q�f��1�A��P��pߒ�J*�S0�C��f�.���`�qJ����p)��a{�����f|j��puQx� S�7���@�R,p�W:�k��u�.��iLkc���9���l��B��X�&�KK)-A���Vз�/�u�
�\�{��f6���m��H�vrl�Vӆ�]��.��39<`BK��A�����O������'_z�����<ߔz*K]b�a�S�lF��޴�ZK"�w��vvرv�nEAW6�L�j���FDsіJ���tm��®�=�+��ci�A���:�l�b�T�?8x:]ֶ���a�J�$3�Y��58���Jی5�)C�g��`���0ǒR�I�``W8>q3 ��\4�ZՍG��L^WO�����FZX|%�#`@ ��Ni¡ �'��U���W����j���BI����*~���2"8���	�b
n��QI��@�qEl��� *�O�8z�<���m>���`�W��=7�Q�%w��me�ʢ_�d9UIFVN�Z�R<F!�˴�a�ʧ���P�`ks蹑Š���n����6�:%Y�e����^��W�b���֔��.lֽ�,�n���,���WK���\��䥩:�׌���Fr��I*.n_��`��g0�?�C��l��U��P#֍k8L%e����"б_�D�c�r0�ˮ�LRB��n��|�V���z��5�E[�8o�fS�U�ADh�-;�9���Ōk�c�<��n2��h��l���'w,-�Q�a�b׶�K�xPJy��������w���������S�N������7G��!��8塰� �R88�W��޶W�Ni�kP�e����ƞ��)�ܾ�t��hl�r۵��g�ך��ٿ����z��f7�f�����싌aD|5'sێf¾�ӄd?�m=�)�1�x�TVj�T���9�Aq��.�������|��g�S�������c C�1~�=3,�"@�' 1���e���J�x	E���$�DO�� Ϥ��lH�է�$$iS�>,^��ꇬ��3�_�l��X�4߄l(Q�Ȕ���{Ų���te��[��Rω,ǃ�U��]��l\7��evc��J�pC	dp�]��dU24ze`�d�ykɇ�Q)�y.{��{����P9݇@@�P�r���W}��{��Ҧ�.�֎�)�v[z_ҡK�\8"���8���Q�W��2���L�M4M��+e%��,�q5�h�$(�2�X�d���2f��y���c�� �T�6�H0$-eT��U<@������6���J���V�{0���r�k����'�:��y���Q}�O;V<A���fժ�K���\CC%=��Œ=h��{�|�_~����B�����y��b��ǣ�?}2����������X���/�{�bg��Y=[���p5�6���ƞ]^�h�P$�W������iw� d&o�LQ��{����o�/�h����(�'�.W�����o:�[~��p��g��e���� �`dN0E$3�ò����R�{wO��载������
��"�ʗ,���gV��H����MJӔ���~\K�wa���譄!��C@����0M0��.�A %��P o���l��q��v}z64~i)�a
Jl�Tn�@?u�i�"���@R�k�ۀ(�*�½M�,@eqN���V��-s~H�r[���V=hI3���7rV(x����4HWtf�rS���l�\.v%;kS�2&��rFIO�P��6k���V��6{ra��r(�T���.kY}���Mp�������pA�ԇ�G���Fpc-��@�a�a�:
(��yt�H
Y�[kI A����m��!l�38�D@,L���)�	�7��Te��R&gU�	h&�l �'��\J�0�P��B�HW-m:[xϊC��|FIڱl�c�r����u3[�Y�m�Y(h��v\*3-��o<���?�����i��?��ﻘ�?�l2�o����f�lHN~�XVv�l�?z��^}�ݫb�\d8o���.7�����<��,�u/C�BA�߳vG��{���V��mh3{�����7�ϟؓQ�VHҨc8�DzY�D�����[��b<Sp��%����r�]�1�����N����d|~q.<������,d�l�A�Pr���EmA���Ⲅ��t*��h8���ظ$I	�����q<��y"�9dÃY��l2^r���n�&�Y��o���u�=7��"XVk.��Є�:xy�c�������.�E�"ey*y58qXF��jX�I[���g���ռ�U��R�I�(�ls�`�,${4��K�?'V���o�b1�H��A�S�Ԓ?w`ǐ3��lyze˧����[a4�,jд8� �yo����^����L��,�{��;N�B
��4��=�t=(��Y:�n� ���(�&�TL��>�L�a�h�(�y��*.y�]��5/%�k��p �e��{d��TEFp�@������,��Q@E��-�����:0��!��}�S�.���r�Jg'V�sh�֡�E��s�͚����f3kWJ)�}��9��n��O~��v�����w>��y�L۸f4�;��}ӻ��}�;�mM�FΔ� �2����4�(/2��K�D��N�)g�oul�����%IJ��}�/��>�0����n B�ܸ������ʲӹTK�,��J���`l���֓��A� .n+���]{��6�г�=�̞>w�NN(��SH�n�U�X��#�H�E�\�jՊ<-�3-9�\���A��IC=�OF}.̆ͩ�$��]C9h\5�E���5}ϛ�^��HY� ق���Bا������	�n_p6��x�	����JQ2���ĢP��r��@����v9Uq@5+�oW�ЬY�Q�|������щ�{����^���-�E!RpUba�"���A�&���q^)�"���e�2[Y�7�����ז뢼�@j"?a���bV�{�3Q��$,`��L��ny��|������J`o#����n�����D�<;�w�֠���V��5�ibˁ��.S�B��P�r�pX�>Sp��9�/�BٮW:��֯3��e��q��oj���(�����4�V��ϡ�I��'�tڱ���mZ�]pf36ڬl*6�)�ݩT���/�9=��_~Q��'>��o�X���t��4�G��G�I7�a�y�{��n�A�j���y�U�H�����}�F
�h>�Ѳ��NG~�Yٓޕ�ś�ٗ�>�E)������4o���㚅e��3;�� �|�K��Ж ��c�/7ҒC��.���|Y(�a_e�6�\������$���P��LMN�%�@��y�C<�d˙���)?rqN�?���E3<Q��8�y	&(,����D.�E�^�R�`�����O'=�o���Z��eA&����I���dQ��>�`1�KS:J//���-�����V
��AJ�W�C^LO������u�<��+��R����K@�&8ty��o�p�����hSS�51]Z�?���\�z`���r��-�#]0���ڑ�Bqe�e�.�	�ה,��[����+�6^m2#���Y��C���(~�!��Ǘ�=�� �������U�6�}x�䔃3�x$�B�\��5��=�a��=@`9XU��L�� �P�F7)�2�է�YkTv�<����3�6���t(�b ��;GV8=��Aݺ����E�r��b&x���T*�?}������^������y�����F�o{:�~�:���H�hm�B��uT�er����t\�Dx�i,��L��邫��ɩٟ]����(W��)Sn��7����.��1)�4%��t�����@��#��ʿB��/49ː���*_��3�+�ֳ;�5U�Z(!Q%L=�68,b<�Ԛ�4�n�Vʬy:�E)��xU��vvr��f���'�)������#�PVӛ�L�T�6�C3��=�p�����A���� 
�JBʎi��}�ﲧ2��A��o
�)�iқܹ�sF��� �8i�p��u��?��^�b�f�zE^ ]��b�)hL�j�VC��jط�f�̏a�6eЉ�?j��P���i���Ƨ����le4�z�L8���e��p�'3ѝ2L	a�T�jCp��S"��4Y%h%7�s�S�+z�\�_sW )��5O�7�D�?�Y�OV���ٜzW�C|_�����L�5�at��]�������{�	.$]0^�>j�$P�Q�U"S��9����RTk�����]/�z~� �0r��X<�\��þ��`>Є��ݸ{�2'��v�5��ۗ��t�R/�肃-����'��һ_\p�,}<���[��w�φ�-!����9ɀ���2ApFo�:���۵��>9�++�=���d���*����n�C.��S��,p��A���s`JGC�)�76"SUz|���[enL��rZG�8Nz�D�� V'/�E��,"o0{&�ʹ����0���t���S$YDI��U<��d�2
΃�P��j'H�Պ�dH��qu}m��P�v6�8��W@4ܘg?���'H�i���G���ep�b:���.��Ѿ�+��(Nx2 �٭�[�T��oT�C��-�GPQ֕ \�":t�IK��$��yɯg]f�=I3r�'�# �U+p_��	ԚS��q������պ�]���o,;[�l?�g�� T���ز�L�C#�1�&��L(	9d
V����'��A�J��J��F=+�[�V��&RG���U��i�3� �C��Be)Mz
L�ju��YC�#丨,�N�%�5��ʶ�|UkZ��i�o���kѴ �ǔ�kG�e��foO甤܃�NBޑM;n[�������+Q��r,Z�wmsضa�d�٭��)�
�n��V+;��n������;�AA��g��]ϧݏ=���r1�������� �Ni��k�)�qSeT葐��)�n@�	h��`b�x%��.h�j϶<yixUpw��VCRr6p�a���Z��JTEd|1�	�� O&��z�����od��5`�j�:7�[����E��%,t�¿� ��t8[�X'-N� _z�u{��F��tI��;ׅS�������K�e�'��[���ɮk=��ؔ����iAv�̔�N����O6ǁ �c��x��I�ۨٲT���'�v	nd<�ʠ�a�G� (�V�J��L|^��d�"h8�"� uM��oC�	�L��x�S+��VǶo���U��ֵ�pd�4&�o7^�俇C)z��Q~R=�.�;|��s�R5䡦������W.��r�.�n:��m��	��0��0zy�R_!���Q�G�T?1P�&d�����ϙP��IA.\�����*�>�u?�����.��� �}>pc�@
L����TQ�RKpȫ��>j��Uu�V�ϖ�u�y�A�+�m%8�c-���    IDAT9�P�EU��Z��o}�{~�����/���}��UA>��?��lx�k�'��X�K��h�	�HtG���Z�!U�fʫ��p�'q���'�FΔ	��+L9�;nFK��`�$*��L�0K,��KSS�A`�'zv<n-���G�̠��Q��x��[��|��#�4D� Qd��r��a�'��	�v�}���>��CKʾ���I�s�xd���0h:Nm�ç��!��][�����rf�a���������8� ���t�}(��L����M� �(��:�����2U�v�6�e���N�ș�9eppG���XC�lf3Wu�v�,e��N�8��逅�E~���df��\���Y�?5{vm�'W����u����j���9	2v{}�ªA���^�ׁ�J��ɘ�C�����^Sp�EBy�5�	>[t(˘jb��b�hU��d|mq�&`� ��7���24�iQ|$��^�5|_�4���`��ɔ\���5�no Uq��t1uc�|F�����I�j����7��F��o�֪[����gwmV�X���.��bAgL�%�/�۽z�����?��o���>[���Ǔ���t>���K�L`SZ+xDޚͺ�	FZԑ�q��u�#=ήoq:�ݩ�W��D�������F�D(���se����f������
I`[m,�i�a�B���F�S7_�@^<T�~CYf��@�{�P`蚂?���" 9��O��֞�tlfe�X#��)�� sS�@s>pdpOS��sC�J��,�tm�X�)��i�% �3< �'J�ǧ��/�If��Pe}dRaD�����e��QR����8�J�l[a%7`�J��Fp�^�,W�!�	.F�*�(�45��W����﹬�B��Nd.\zo|��5�؁嬹4���m���J����f�L���2 �T�cz���]���DL�ᏂZx(HΝVC�i�!=ו%��с�5�,0�,+uMN�{AK6*��&;��L�KL�$�͠����Rs���r@y���M&6�u%ѕ/�fCY��qZ��;��`�;���6�d�O_g�b�d�j�7�?���j�f�㎕O�m\/�M1g�b��ł�;����y딪v�V��oy���>��/�[Jp��v�׷��{<�֮Q�o';x)�����"���N�����{��*������:0Vo*��p�4k
 ��f�VP�@�6��8x.�$���J�A�,Sl��8�����c��$���`� ��[dqh�!r	*�	,C�B���I=<�߱Forʴ�m%t�l�h]����5HT�B9�f�5�IX�[;Q�wI�:�d?ѣ4	���~�����70�`*��)`�,Q}���%)S\��fw����|���T�ʁ�$�s2;��(O�ذ��a������&��Ԑ���k���݈XO��,_���A�Z�U��RC��te�u�ʨH_�l��S[=���x)�VQ� �ȡ����Ź��xn�v�B:wP"Ѥ<gUDYMeodzW�מ����aM@��Y�}����P������rق�!(��X)#��	"	��`!��D=�f5�O��F9�Y�O�����Y(،���B*6Iu91'��TW���7A
7/�>�-z�Z���!���� �[��\{�@,&�׵6�ۑ��ۨ��n)g�]��|���u���T�{���K��������_��k.K��g�����_?����W�%�~�6�R)ѿ֨���.w�NS]4˫��7E7��b�7�M)��A�$� ��t��f6M�4��� ��!�(�sna�y,*&���b��Rٛ2�$z	�e��D�{��d�r�2�r�5e8=&�_}�`K��$((r�-iwR:����}��l$�s:���nXA��T�c��X~|��u�y��d�R2�� �f�[dF);������arB͊�xd�)�&�R�Cz:|�/|�eq`s�I!2IO��d^di�)X�h��W��dn�BI�N�9���$�eL�$X���������G)J�C�۪K�	�x�WSW)VA�t8���k�=~n��UfK�Ŕ���q�$Eӳ�l��!Ȇ�c��?G�Yo���b����K����=�kUeas��9�,�2�`M�ʲ��A��<T�p:v�(������|>�����5�����Y{�y�ӳ�v�����|��-7�����򔭣��o�w��a��I��Вj`>Ѿe�vƍ)p�c����VL���8n���sh�j�nJ9�*K�$/T6+a�h�j��~���g����w��T�}�{�������t�?<�����f�s �� C@��͚�o�`&�n�f�@qSPV�,�Ͱ�����USY8IEU�i.$pVϊԗI����LLN�NR���!��:�2<��&3����K�J����MI�z���L3����Dť��VP�W�oT�ϒVZ:b��sc_ߜ|����;ft��#�I���}�*���C���ی�;�؃*٢����)[4nxDSi�T�mr���ӽFX�b�b�ZEޣ��Yރ�a�Y'�+�ِ��
;Z�.�#�5�l�ԡ�ir��@)͡��%h&��k��-2+�t5]�,�Mm����o>�����f�������Δa����p�ۥ�9��&�zV�v[���hj�;���>USf��2�����<j4-M���3�XY�ٖ���b�0%3��41����d���H����\#A^�rY��U���'�\�+h e�Q-���H{+����nH4ׁCvO�]k耤t���+0��[�c�V�n
[�5�f��MV�D/#��=,��n��_wp�?�����}��ל�!yt5��[��?uK7�O��#��f�9emU�O��B��>���#J1*)h4y��6`@ܒ�n��:���R��Ŵ.�N)�� ��B���[�-�c�i�HNZMYJ�%)�R��i����Ց�1�`��WXo�U/�,Mk`"�� #'�2��O7%9ǧ�K�¥�@BpK=�0�I�C��������m�����~�JI��H�5�8]�]	�3=�Z�'� �`�	K٪lm��(��y��A��I(�5JR���d��(�������.�9ǆ��؉��qMt3�w�6d�� k�UKwp+�������.�]���������l%[<�@��K\m���3�b6J�nr;�֤L�	���ŵ]Fpc�9����6 �������ߗ�'t7�V�U�y�ɍL��P�b���f<s3���i�Q���م�rDɱ-Q�T��C�nq:��)��޷ZP� ��2^Al?��Q�?M�E6��Bpk�Y�����]f6vU�غU�\�m����|WJvP,��J���ux�G�;~�/$��
r�������������\��n�u��4y+��~WF�A|�-���ƣ��m�x����%ewn�+D��$����dn��=�	9�k����(>������Ta��H���PŰË2R�0?�DpI�$z�7��@�{� �ZM�����=�=8���U�F�P�^�.��S�()�Fp��J�y���|h�S���q8�饪��y��	'���E���,����W��}6��,��"���u�S�H٭>0`E]kMz�2�S����̆	��U�����ěۜ���`l��6ytn����[��*���M (��!�>�HP��E���f�)r�����vuu#@-A��m��D}�l����U���6�����u�����yX�$Z ������"6��]�����OBy��K��Bw*$���oHzp�����k��1L�^0��=3n�^P
�:���=,h�}��R�3� ��>u 	�:G2���l;�t��<��s��J��f�h����+_x�������#�B���?�;�\M��x6��Q��*�.�<���Fߍ@G�W��~\�` ��~�/Ђ��c��k��=�T�i���Y)(��E��y���"68ϊX��CXY9c�[��$;����)S� ��8h[ҏ#R�*�jLy)�AP ��7���2H���(�r��~�+%w:_���~�,Ӯ�}{�&:P��{x<��Y���h2�9��2/��"�>"��
�������ZYPG�&D>�:���y g�A�N4�4\P�z_쀘.'��^oTP�¢�Ǒ�q��PÉ�6I�o���_�z��噦�FEr�Zp\X�X�&�D:|���ͬ!� �Yn���� �&9�>���Ö7=Ӄ�՟��7�TO�̍5Jo	{T%�]���6k�ֳ�69]O�a�MC>���zJG*pa��ԗ2����&�^���"I�'����V�CZty)~L��dʋ�Ng��TI��2H
��|Ҝ=GVe�f�J��ЋeO����Z�[��V����O��?��?|!��7�蓯^.G��d6�гI�0خ���1Spc��(4j~������)��/�uR7����}D#[ӹ(SS��O��JRY���f�����TH��Y��2��ŘP� #s!B�ps�2Maԇ�N)���|MY	�@L&3?ф*G�	���C�[6`�g�YJ*��=��a�ז�a��R�K�O�^����bA�Tq��d��:F&����~L=�]g�1��!A�FŌ ��2�33����;A�� ��E�À���,�������#�9��T�ZVF_4Q����0=�t�9�D��3�9�l�{4�oBߊ@(tW][^�X�7�RY���f+M� YR�d�R�1L0@��� !dY��0��/Gֆ\��NE�q�V�st`g�
��2�~rue_��7ڌ��6c�͖�v���r
��tYM����/���)��`B~ QN
��{�P�5AAX c��$��$Tv����dj�� �Ei�B�J)\��\��N�*0���F�!����2�Z�i�c+�nE��d3�I9oVo؆uDPg|#%ރB���/|�������O�������y>��������M���v��v׈��sS�F���F��E,�.�O�TE�7YƢ%�J����#{��$����GV���ۂX*E��f;�c9!�h��@"�[=26�W�T(a�h@R��+)(]���#�#���[r2��~�6"'(=�oߥ
u�[�샒(�����ݺ�K	e����(?T�ǄU}��ߧ�dpd���̢Dܿ����Æ����Wv���S�^�����0�PY�/�*�H�M�3!�P5���(�e���c*�.������RI��f�/�h�re�����[,���]��&�\�M�Ǡ�i��I%�d��M�f�oԶ�b�����{����F��=A6��=�;�rv�Z���Y��?�/}�5ѯ�N����X���0���D�~����v���0�Iz�
n���<~�s��.9��aZ�ĳ��W�K+���mO���Tʼ(��ѭh�|�f˕�'�>#L��5�T(9 �a��S��9�r�m�B�η+{4�·��$.6�r���m���������������/(���;/��xk2�go�n
}[�3*������`b�'[և	�H�Mj�
�$`�������FѰVɦ�/������G�,J٢�|�<%�ƴ��.d\xR���$����b��f�E��t'&�����2��]��2�l�|��F�#�K��)�_%Ys2���I�.�I��{�/ é���wz�[�����c��11r��FL���馂�������DD�W6Ϥd�W�x�&ʰ5.ML��0���/�$"�ANIr��o�L��{Pp(i�����Y���n���#HH2Z�aȚ�/xWe&nV��!`ʤ��/�[�[A�3�* z��= R����֜��k�{G�Z�9�w�q(l����?@��A�f�����ݽu�̾��2��p�ҷP��f�:-��ւzV)�2������n�)\Q�k?�8"��(cCz�����B�[��j�%�,��%�(\��g�;d8���(S\O����봿B�l��C;�{�N�ݷ�ѱ�k%{�Y�듮=�Om �)e�TypnY��ڟ���/��/~�#�y!��7?��W/'�_s���G��
B���F��i��m���-��-PO���
�HpK����M��ϣ!@��e��UG���2'�ӗS?��D��F��5���A5MR#�dv�M��/JMACd|���J�W�@��썬M=92�(i	r S#��� DR�5ٜ	���Xh��-�T���� �kHs��0dW^����]������,����CD���|r ) �9]��	�ͼ20��GqJ� Á#�϶���இV�ы��J�!ƗT�Bz�CA�E�x����Y�K��;�E�R�"������y<&���w<e6����g�K[�a]�,?^h�����c�F����Ȼ17%Y.��M��D����H1ꓬ2*���K��T���JI�~���|��Y��ʲ��K���[�Α���+������Y�À�f �%-Wk�n�}��NFI�J�ddx,ā���5��^4�j���ߥ߆����6{9[ =���X4TK�.�	6�����<x`�<��ɱ�j{���k���5Xo��1�&�=���f�Ŋ�|x����=������(������\}��Q�p�����X�h��ܜc��d��$��P �:�}
^��C�;5�=�Q�e<�J7�@2�T�@�D�6B�2EY�r4�r��ϸ��&�p��x��@����9�K�J�CG�%�a�"
X0#8����)K���^�$�c ��-���o^	��I�S~-SIO���cD�, �0�`0 +z���@G�p���C��J#�� ��i
�d|��N �0Pa3���7ǐ!��hU�V�����+dw�H�)m�H�u<!'�8����3��1�j?��N�M��ӂ6ٙ>qE�O,�ۦ?ѿ������𪨖���g���'�� �2�q�J(Uܣ#��0[*�lΎ�-	MP>wC��zn�L3IR������=;99RFz~~n������BrLR�az�l��񉵡P!Ǿ\��͍]���@y�~@`�]!�����tj���2'g�`&c$��&S�<	s��Ғ���|C2�m�>�8�SD���������U�[?����=���|1�������̟��y~/����;:�y�×~�>���b2��|���r�ko�	nE��P�-�_�빵�Z�l�p��Cq� �9���j����0^���}�C��
/�Iu�#�/�X����k�e�����k
~����T:���Q��Bdd�Ѳ�n+N���uRG�z��/ԁ;�o2�ݮ�`HMk�?���x�,/�g�l�����P捃"��z��������h��,:�t=3cahV``ӳ�чK��ޏ��� a�R0�O�*&�L�f�$w/[��M��9AL$���-xB �֭3�I��>>�7���&���P9���Α~��Mwd���2��m���W�0���0��d��A��^�R���k�rCf	E��&���֮Vի&�R�[�m��"u�/K���7Z= e��<��T�5CFȄ�Ѵ��S;>�h�cC�׵>�}�� 3 [V~�AQ���:P�08�S�� ��K����0����@'NԲ�.X]V[-�޵��^����ttd�r�ΗS{6ؓi���S�Y�/1�JinknG�W��c(��]�g�Jp{<(�!)�@}p;���:������� ���OY�hF[/+�@b����Y���W;<��z/�T�$��())v�M�(�vt-ֆ�A�P�e��C${ �zn!���i�
J�C[�O�@��aL��EI.��ن��������a ���P2�=0=��x�~=,���tbs�Ѣ̕�2�8��=s�Sߚ��kk=�F����WG��~M�\�ط�c���'�4f��I���R�4Q�F�d#�\�x��D����$��'������u����dJ��c	dӅ���zL��F    IDAT`��X��Gp��H���v�"��#��%����3L��}TE☂��|%g�� �U�T�y�-�awF֚5�mȈU2^\\�u���[�	�Ea�igwN�谣�u}��i�1�WK���eEY�+x%z�PV�������Ԟ��O&�Tk���	bȃ�/�wP�P���V@Y�ӱ�{vrv��Z��%y�����'#�'������"��l�Ke{�� (@׿���ҏ������ЯnϦ�_{4���'�a�i�~p�H�hO�/N_�K�� ���9�4ߔ�ikR�*�p�����V�~�H�
P,8�)�fz&�)�����ɣ��[ʺ$%_Bc�&���4��t,`($pU#�C�D^F�[ew/�\��7g��Sf��	�ɵՎt[�r�P���	��58y���i4ޓJ��25��4��+�����W�ha>��y�r�{D� 4zdcSV�̇{	�S�̃�Rbh�)�y����F5���xj�\32���P���{��g�er8�������~��0&3[�V��l����g���򓥰oL�ד�O���` �����y��=JxϤ��32I�S�� h8Ƚ��a�}��AL���\�~�s4� ���vm4xƕͨ����֮���c�F[H�n�,�119 Yg��]���v�R��ܸL9$��z�r(�)���$6��g�ϭ{�����֦�-��(X1q%�-��}ܱ��3;<�gͣ��Z-[Vkvc+��4��q��g#�o�(f�����T����?����?������ŉ�U�|�����ӯ<���ڛ��|:킛����M�enj߉,�[�#p<ʔ����"8!<e"��&�66=����rP�A�C��0��0�����XNդ�F CxP;)�(��։���8 ��큉�@�bDPk{�RpS��$}�G�$<�18��y�TVx�IŃ�ۙ�Y^M����;�Ԫ�s+=�2c^b�qL��*=�iR�+r�pLa�Wi#C����۾nb���)� X�w'�ZSɤ ��
�Y$�܄#�End(�ЬN���O�-�Q�B����M��h��F�� Kì{Fp�زӅe�#�3��?��'(K'��ď�1:����g�$>��A��
�a	e������4�`X@EvG��|>SV'�Q8��|:�
$`���P3�ʑ9�j>Z.hJ�bϊ�5���:=�ć��\Q�!�&��Õ��J�����xBD��z�S�V�c���
n��#�.�?ۥ������.�c2tTb��&�����o���=ǧ?��/

����W��|��l����R?�������#�E�����M�N�36`��>�[��4T�*�_n"��䖠���CT·2&��g	t��}�?n�
dQ��yY�Z`^��SH��E�zr��v�+b����Q�zv%��r�0�^�M�ސ,߹�{�)�M}�o/K�/M;I뺹��~�*	*��	����0��*Ch3�⑲��#?��ߋ����E)K�A�2D`$�E�q?��	����9�ESW�M*R)�=6��|#���$o)
7&�5��l"��E��k7�]Y��,��Ta|��������K�L"�M�-I]�m��7��]��E�'s$z�L{�
I�h�,�g�M ΋��&CM@9�aE�_����-�ܰ�9"�x�B��:��Rÿ^��#en2��d4,�����L��4%��;/��[��x:��S��^V*I��,y5����ٰz�m͓;��@�-�h��reW˙=���gOg#�ZOm�y��V�d��
� _x���g~��|�S��R�*���������W�^�����DY:W:�t��6Cß7��m��ir���n���WHMYN�q;��\
!a����L}2��ঞI�����������5�T�:K�\������xRe)p3�M0���4�&*UC$9�{m�BQ�(c��~���(f��>Ѓ[� �i�l�BK.���UC<`2�c!��/��1�K'bg6���e�⇫�Ͱa["%�G !�}�64v��� �ei��S�[�Ȓn
,]N��mTv)�>֔7��^�7Я�À�H�m�d�SJB&��bX(
���l��ۺ7�md+&��KaS%�G�]&����;��rt;5#�
�p��bރ��2ޔ ,��T���w;_JVH~FVG��S�)O��5�{���J��mIc �P�0� ��늲�x�~[��SI�k�)�A�pv��2i-��������JJ�b�=��I�ri�RQ�4�[�^��ё�[��c�:W��Od��|6�g+(�2k)*ӗ<���\Cf�/�:�������-���?���G�ޯ�9���n�Trߡ��Z��o��s��T���dr�ҍM��۔q����$�T��x�!������O�F*�U#�$�K)�s�"�ȧi*Mէ�X�LAP��!k$��7\�nI_>�]*y�9F�*�H0p>Jl��I��5����_wR�H�k7,��,��$e:�R>�{Ġ 靥�F	��~�82��� �F I�V��A[�r���m4_��qܙ��1Ō�Ab�(���E�JYI�� �8�H�>��.�n^�*�	�6�r��	^��r�M粞]�܂���=�(N�#1��^�M? !#���P��ɻ��[�"��3<
���$,a�o������g�s����'h����\��	�����q���U2n��EP���t�@����|I�O@�</��ڰ׷^��&dn�dvx2@�*x'0Ը��Ppc��\ �s{�7�d�Z��p�sh���Vm���|=]��rf�2����n0��.l�Y��>�V��Pp{���ً��O��������Ëi�W���i�$���.��-����~��d#���E�F�%zE���x
B��+c��I�׳�T��hJ���>�,Nv%/��JM��T~
��7 $i��gQj
C}9���kK,4Up]즭~���0z��JT,�8S
V��{������2��}�� ��$LT��s6a6��C�U�[�T�z�l㛞��S�G��.W���n�l�v���34�.][��㣦�NHx7�^�X<�yL��<�����D"�@�wԳ��y^pt�� 4�߻\+�����%]_5�j��f2���M�{ܠb�`�8S9+!UI�ϝ[��5�������:��A;��{��`bZ�ս�>�����]扽 X�C�V�9)�9�A� ��^���+�1!B���K�Ddٸn�6��1Vv�z_G�ݖ/A.ABFӱ]����C98q[uk7�R!�$St��U�:ֹ���R��|i��=�m���8����j9��z�!��A�b��m��l���j�������*	��G_sY������'�����#OF��(�QpK
	�CYJ=��m�~�pQdr\Ь ��2�
:���ښ{����B�!M�H���*NW?eCH
���Tj� ����� R�Ie[Z�*-�L".�^�
�������~�{``�y<��4L�,�׬׸���=&�v���-25zx�tB��a%!D���	�nO���֮�*�1Ӧ�vm�S9�?�Xg�R�}�_g�æ��|ص�vc��̃[���ߢWSM���~�a�B@3�����PB�Hel�x*�^��d�B�J��Lsyk���;�����۔�|�������f݁�)K	�;�3�ZH$q�90�͞�{2�Z�{��i(� K�j��%a��͢��o����	'���1 \'��q��]�>��IՖ�C�*h	A�>���l��.���J�[m�z��Q��m6��{ջ�Nk�>�2�Z�ڈ#(AS�g�j�'�89�e6cד����v9�,���������d�V�u05�%;���A���W����o���-%�=�����COǽ��p�,�* ᝋ&�<AL����t���I=��փ[��i2�_~�[
h�i}Z��d75��n�zg�kx��㱪]#�2��6�oʦR�K�\|��2�·a��!)�iZ�T5d�yF�5t�����օ���	�*{/c��!��qz��j쥶^g�X
��{���+O��f}j��D�Ѳ:ÄMƮ��ۼ��އR�!:Wf־�N^y`�;
n��º˩M9gd�R�^kL	`�oJ}Np�5�K�䧑�"�r�ا�! D�t�_��y��x&�ۚ5e�p�ؘ)�Mz}[Ƕ��6����3M%��Wy�������:��;0v��NÜ���=Ā��$q �2ة�h �t5N(�F_U�И��R�gq���MS�f�a��*����/	v�2%�@���4�n���Y����[?�P�O��Ԇە�Xd���U�Vi5�ztl�F�F�݌�v3�Xo>��0���va��ږ��!J�J�sk4>�j��'~����EAA~畧��y<����7���
� A�W�R�IF�%���5Q&Ɖ��%��d��H2i�:\B*/��8%L�܉9N,�K����dS�nR�
�"��E�}7p�Ϣ,�d �-�P��`3 �+��s���+�������G�9{�/e\)�'K�JV<��*�e���҈甅�� "��;�}�M额v��o��g�?���94�[*y ���[u{����W^�gî]���[�T�
�/�M ���A[&&�׀�DpSi��};h`-�̞ W
^��J6�f���Fl�029�xpb�Pɸ�q���?c-�j8� �@���i%n$܀
Iՙ���w��4tJ�-	$4@�2�uJ��V�ϱs���������[j�x���&��9!�L#r�=��z�L�*>� Cb�t�]0$�>
�({��hZ� �r�9
�2-��P�m�R����B)�@��eq-+l���K&o���&�� ��m��H�����A��5kf���f?�r��c?�-��b���],��x���g�~�G�b�����E��[Men,<���wҼw����7��>��UHنP�܈��5G0�}����[E�ԫ�j�%
h�^�R�,������/9ky�J%�"
<
���hW>�Po�	2r8E�I�
�L��TS0ڕ�އ�r*���)�y�+�y�%���;������[���7ްg1��sx�)�l0����+��N-�DJ=��`JCY �bƬZ�w~���޻�aO7j_��6��������x�fn�Ep�7e�E5���6�26̰Ke�
�NBG��B�^5�+.{76��-�'��\
J�e9��4��RwA�rz�W��>`��'��%]E�)����^�G! *�	��W���.kۓ�O�i��A�U4�ZG/O�<����C�8Ӵ<��1��@M7���$�b��j��X�_��&[Ԥ  �V�\���
ʋ�Mfc�OFn.����R��f�"�u���l7-S-)����[�ٲ�vm��º��)y�Qi���ɱ�ZVYe,?��n��?�?�bd��s��M������^��F�6�IB?�b�l���m�u<T�D(��L=͗$P�{�H/� f�����'=��
H=*Np�jᵰ���V]�2=1I�$��$.=N��H�|����`,8�b3����1L^�M��Ty������{�l�[#CM���x���Lտ�y�pPye"�'/���M��˯��[�
@�t%���2���㛾A������|:����F���fD�������RM�[�Ӝ��}Dm�(�)�����r	rx���@�G
n���U��	n$4������uW��Փ1-�v�j+`�~��6���2���uS�T�����u� �ϝ��&g3t���o|�F��t�%�cQ6�1H
x�Jo�n�w��t�%P<�������:�L��VRx�
���G��,G�^�[�y���v�pk��E8ܔ*^�f�,[�Y��A�օ�]ͦv��ëR�����bbS���l�٪��ɩ���M>�R��џ��|12���O��b���Ǔ��=��sdnhrQ�y	��P������_n�
N�(�^��(m��)��B��WIF���?�Ʉ��Ʀ� #Y��)hi��4e'���̉�WC�O;&t+7�������	iiJ?��r&�Nl1�)�'l^*w�4MִyR�&6�A��,�^[�:z�hP��ƓPg�����*�,�N�@�ψ�GOlxy))ut�(3��	۫X������y徕Z��'v���w2�nm�����)�ݲn^:9)^m9׉s}0�j*{A�U��k੟9�{P(�X��G��l�H̡F/�=���#??=:RpcZz���M.���2	���t.��t�PYN�A �RP���^�hX!��H��g
X�.���!֩�����!�W!G'��[���q�	C�8�7���c	mϯ�'���7�2��jN�"�����}�̍���nWU��2�f�d%�0����u��W��T?2���Zm�u:�b��ZhŴ}�3���Rk>n�,͢4�\��+G�~���C�����k�����|��t��'��w?���fQJ���Ά�	�̋�
��tv<������x܅�<�qs勉�J(�J�(���֌O735g�i��#�����N��\V��)=�N]� ބs��>̇(G�4���ޔ��v�-��{z�{��
h{f2B;)�F����6̓�t�-��u�:F���ʦ�GP�4N��\kT% �V29�?�����+�zͥ{Tq*�[�����mTm�^؟�����k�2��,m�����
�n��B��� �!�����$t�j`k� �1��0�~L�)M��&In�݀����-@���{��g�#��Ս=���/�%)�:!�-�S]��~F�^��Ñ�сA�W�R%;�r��?HJ���#�r1�N�BE��iT&�jd5	иX�>�a�=��&�̮�ۋV�����/��$��d�!�~�%���x�ڣy24�����T�f�-/��YP�`����ʝ+�,�l����F��e��C�������*U,7_Y�P����?�/�����B
�������?����'�^��Ȱ��&3~���hօ��p7J�@n#G��{�FE5����J#�D�ִt��������H.g�$�)~귥SQ��]��L�x��H�(���$���,e]���T@��̌~�9��o���B4�JB�I�b�����X}�R@S�>a�$}[(m��t�o3֩7��PFӣT�m>�$ �����N_�ow��P��'7�v1�[�PpKe邀_D�l���J٢��/�*��-|+e���u�t����pu~)��K=*�5\-1��erOƕ�
'���	e�SE�
[>��{��*C��]�~zn�~���� ��kB�c�xC�.�ے	w�Qq�b�>�#c��k���g���4ݩ�DT���^����N#5?�<$�K=�[N��7�zB�Zv�*����)�K��$1.Ր��H�s��%��ALv��Nk��h(�"?_��"��Hнb��m�%�2@e` �&r�y7eF֪�/��F��yt���m�/m��ci���=7�X�ҭ\չ'��,���Z��D�暆m�-3ˤl@0d�h�$�)���_�P�,j��@n��ӱr�7�l<�9���ޡ��htw�[�}�s~�������dnn���6�
n%U#;N��kn7�c��n�:��4a�i�I�YeF�Rѯ�����Og��1���]���ݛ��؟sS��i�-��|����ćQ>Ǫ��� 7��~7�aXN��#��5��nJrn�z���� ��B��Z���������є=X½;�%�i�rfTB�[^+K�d4�l$.?i���,������TI�N<�`]h��B����nW��߷׃x<�,,��/��47�Es�G�]3`������A� ��4�q>�܄�9�l��J�F��.��ں/�6'3*d��T0";�f��z��~�0��<Up����1�s�'����4*�A�kXf�\{��w�e+���g"sr�t����@õm����S    IDATu����V����m�m����e���T�N7תpC�=!�2��Zo���;@5�����j#�n5J�� �1�Zi{�mX)Nb�bVghc&8Fբ`&��i�%��1Ml��-��o~��?��W�uZ�w�(�գF�[��?b�8�V��UARt2���HQ#���� Es�ce��T�����a��θ��Z���<	����љ�z�ne��Ȍ�43�k�������I^��6����9�@�fN�W�hvp�b��.ke�.���쳘7�g>C�, f���j���zMLxJ�JZ�g85���Ws8B&�Р��E1R^7{[d&�nդYI��	9]�9$8����+�I���s3���E.�����L����vg(��z�]���G��Ե���Ԕ&���A�g� ��
Z����z6�&xk��i�
l=�L<��t�xi���p��2���r53
����a����ʬ7�Z��px�P0f��c�o�7Nފ�E��0��i�8�G��p�q�Ѥs,el��O5}��'�5�zy� cpS/Ӫ�8��37�bq�=4��Ng*��H���2�)C��@�<31�\��L��H }�Ӏ9�C/�Rae���$��N4�Qoݔ�DD��1��-��������)K�����I������_;��(����nx��r�ǒQIR3�	E�udt��Nd�qb���B�s����LG�pm#u2s���M73P0��27��?8��vJ�R?n�/��it�<��1�uC��Qj�@�m�K�H�#n4-`��X�������}�U�}��1nO�S^I����y�⣸e91f�i���JT�!���"X�_���"V�E�>�8�	[Ĺ�<(��
pa޿s�������#琐�����!��Y���JHf�T�}�����c.ԣsRo�9�f����0�*�:�*2v�qpq�멒��aƐj�Ny��E��Y�yҒjG��nO�/�39B=d����j���j#�#l�g�V�ku�ԑ��u�b �
N�uuk\� ��֕m�;��R��nܣu����pT&Ƚ��q������8��֟1���ﱛ�OVNZ�V�NL:�.!�N�_�C;�N�#ax�a���+��C>c!�cAD���|�:)r܇H����xj����/�~��'_�|����d`����
���76N[��W�����W!ZR�"�,��h�V�	K��`D����6�S��5��tL�f.�y=�)�ص;*���ocf�9�\p��vp�Y~i
g�����8��ր����;�6�T��I7jbq��3a"H96�t���eb��v�W�ݬ�8'Γ��J�1y�5��4M�� !S�hW,������7n����������#<�|�ݣ�h�W�7�b5����G��_� ������ZkkkX[[��Ң|+y�1��
���q���{x���`G�Nꖦ�:����Y-~^�(HVq�H�R���������ݦ��b��&��NmVYvG�g�"|�֧��{H�xI��$�떂�֑J�M�Z���)�*�YN o����Q�����LVu���\TAXe� �]�v�I58J�Ś��������u�;�3)��_�e��DB��b���rf��t�v@b~��z�{n��x�Ԍ�I�J�����6��D0�ԋ#F1I�>]0�^)9�7?��
��|<ux{>�������Y����ܨ
r9l��;�˟>�\�ʜ�t�w�~�=�x2� ���x'0���<Ỷa��Lps���ƛ��fu�;���(�ܿ��މ����dCU�-	��o��Z��0!��\�����++͂�\AG��=,7%����SX��D�fhܮ���4�k��Y�!FE�<>�^���ept�2]1,,o�#�����)�b}qo߽�w�z���x��9��|�
I�T1��f6��O���2=�R��ǏQ<����{ｇ����x�ݞ�I��B-~�/�0z���Ϸ_`�`_�^���;X��G&�4�4�?%U�>\H�����x�_<�a���g���:� <"K��h��B�5"��z�J��l�A_|Kfx� H�cp�|��X�8��D��ϑ~7ܴ�&��F��7�gs�����.��+
�D����}��X.���3њ�u"s�#lt�j�3��n�3�-�M]��  ��c� �>s����G��Ǩ.�#��epQXa$TE*�4��^������� �������_�5��|���
~���_>���E��;;�˟�/_F����o��l�n�-K��$�܈OkS�M�܌|x���N������J?ʞ�����{��b�����p<�p@Z��+�6�p<��)�p@��P3��/nqO0+�I�bv��	����Y�B���B�u(�j��&(aԩJ��a������}���xR�����8�)�Ǐ�`#n-��ޭ;x��q|z�gۛx��)l�[�={c���_�q,��y��dST��/��|�3���;�S�(��M#�8��f�AK�"������M�pgm�x
�~O���ZU��G�p�S9#g���o���Ml_��U����mb�M�9����N�ҩ6�`�VwL����E�R�0�P*���3�9�ǤP�[:h�����!
6j\�\�7�P�����!��E{x�{y�[�;tݞp��5c��mš6�N.C�ai�������1���M�h�5$��K�p�h�X�x����a<PU��<�W��hL��oBw$��d`��߯ඐJܚ[����Ƃ�e���+W��[�'0��q�@�K2����8�u9����L�z���R�����5ї�p��)8ܜ��d �|�I��}����zeN`���ǲ�*����	B�9&�O�|,9���.��6v
.����{������dO���F=�Qʴ����dx��3S��qoeC����}'g*K?|�
.�A_pn�?��쬂���eB���߿���e���c��j��$m���cX�XW3�(��/�X7W���g���>�W�jT%��EE��������#�ℾ��K��X.L��8��F`ꖙXSR�-ܜ�%���rU�p���s�-���\�䂝*@w�'@'\)�Ke��*]9)�)u]W���i�:�I��+�'׹�Z�0��L?�|����a�j�H����j�wz�U�Z�3�DB��	*�I����<���n�}z���y�~PIJN��x�H��ȧ�{w�W~�s���җ�����dp�wY�/{�Y������ՊQfn�J��&���z��2	Er����6����d�7#k��=%ո1>Z�3� >�˵o���JVW�1����LНTZ�Nr��K;��`��q�zǎFi�D�5&�4�@�^�Q��7*n�����!̯7�48����pM��ND�WV��e��:L���1D�}����<L��d�#�<D�v7�����?��;�e�ɋgx��ʭ���Bͯ\"�Ͼ���!Ev�n
=���C~q�^GW���Gb��D��$�-@�w~~���4�J�8���n��k�����|��JU�?�ហc��̴6�����x���sM�4���@�3$l�sY�]�ڑ֌c��?�vk�<C@D��"�t=�QN}&������̙m��(Z�e�Xf�d�!��0�#l�Sp�0�q�c2s3��P�Ȋ{c̠�Ƹ)Ks�U�^&HP��"�5CA�� ���h������"�1�1s�&"
l�0͂�s��54��ό� ahR��&�45�����[�����7"V��<����v���+�?w\/��s�[ĸ��e)�8375�%Zi
�,epsP��{g�e�Q�M(��Mq�9��uٞ+��z�=���O�j*Wl�T�`�\L����YR1����S�Yj
]㒤	Ԅ�_�-L�פ�Ƅ��Ny�����{t}�!{��F��@��@��)-�S:�X�H��a��$���t�������{�n�F�\��-<|������2)ٯM'����|w����;O6EUʤ2��R��x��<�{�3�MM��#�Z���Q�N��W�9�YY�[�uty��}��Q��|�сc_L� :3�}�]^]��N�?k�֏�Zݚ�Y%NK�l��M��^��?�5�nX��8�˪M�z�NHV2���Zq��n蠃O��3 ��>\W�Z���� ���a��C֖�nR�CB�њ�[����5��6	$v|m~�Nr� jl|�԰�{�k���j��g�F�n8�Q�`� |Q���(�N~)��o��m$���L�R��I�L�<�9��w����ʷ?%Q��O}ߙ�����g����S��/��x��6�}��e�#3-MF��2s�Ӽh�~���Czl4����O�1���� ��>����ZX�g'�rڴ�e]���(��tSI-..���t6��IMv}>=*S(��_%�I��b �	븟*-��ev�_� �G��I����Mt�Z��	UWȩ�O{,n�����:ˀ�ЋHX�����zoݾ/������}��/���p�/~�sX�]B|��������8Vnn�6���1���w�[�T�bC�(��&)�;=��ǝ�e��~wo���;���7>����#�	?ⴇ84��aƾ���`=Nݺ���el�JC�;)�0��6087+H�������E���PMb]#�>�3���m�L?�\�;�Q��2�٫>��3���긥"$���yMŠ�N3#�L���pu�[n� �@�Vq�-{r߫�V����|�:�|񈙐��R�Q���3ȱ
�СO���	?�+>�I� ��1��������_����?�����N��V/��Q��,%މ=-e7C�C�s#z��.����cIS�p��q��eT�ҁ`πs|��0�ܒa6hjey4��0���k��+'�=A�湮�n�[<����i�;�ܩ�Ǝo�j��,l�.�~��N��&&���A�n��b�*(
�F�c�Ĺr�~��?a��<˭>Dh��)����w��ݷ5���%���!*��zf��yF�Ke����n�-#?ζ�,���omH���������~�,Q�a����Az<v�Hz|�5��;�k��qC��R·�>R`<��P��u7談�Jr����ٍ���!'+B���8\pp[��_��8�1�1�&�sS��k �n�mH�G]4�/\�Ck��cu����f�)��*��ǵh�����Dn�3[B�C���FL6iA�6�������>��jv]����g[B��ʘ�@J�y�(d��(Ti��%X�5Ì-H/}���cCp��xM1L�z�#����?��T����7�o|�F�3��F���
��i���	�fn��)h�[4Z�72��$H�G&�qK�gA��_��iw��X,݄^1^�*�O/J��;Ь߀'Ǵ�	�N>"�]&����0=6'�uN�������zꝍ{w��'7'5d� �|��k�o{z�KlW�ڛ��WNm��;9(�W{B;�~9n$�z"�j/ ����@o��W��ͻx��=e���{���C\U+z�N� �7|�s?�;�� ��n��J073�b���ǻ��'��@�?��nN��@��Al�E����n-���;�tOO�W��㏰[��9}-��e�ݽ���}Yǻ��t�_N�N"�}��Ϝx��������/co룠[{?��a����S�0���={���������Wz�t-�k�P�l��w���;�,�ϭ;D�D�'���d�$ߏ�^(�.�
��&-6�9H�+���p��q�3�G�xI���U���ƞ���"NI)�"O"O@т�Ef���^7J�����������}�������?��oF����e�z�_���17)��N5.Fϻ�m2��M�Ր5�Dp�<�\��iN��ȕe)Og�+�?)/�J��ӑ׉h�)���nd.�R鯙r��Mu����9-;W�^8����ZD���M��M9|M�r�	P�bǋq2X
�b6���i��f63��m'xƳ���f�݁����Kx��=�w�-����5�4�& 75�Յ%����iqA�_�
�C'����Z��է���E'�R%$K�>�@�> :!�	`cfN���zWW|rq��~�-��QAM9k��F���\����tDs�?bݐiVc�ܺbc�G�+Q����n�,�(ee��I�e�u-Mam6g��Tu=S�'U~�qA9�@����3��{ߥȤ���p7��q�T����w%��UI��E4���K��\�z�r@F_p���'��F�V�26VK��sC.v��[�hP � �(�W��CU>3��H33s���a���P)��j(���ͦ���P�@�1�n�W����?�fzn���/�j���W+��n칑8Ͻ�2$7-�g�J�Eo�S�&)h�(Hȿ�3��-}}cN=wB�Ū�5�D�*@����-���;�{�������^�u"'p2Ⱦ�3���il낙�&���g{fщ����TA��&����X�3nnwO�\	��(�X3�����GA&�nN��7L�F����9?{���s�'c1�^����Ul��!��[o�x{_ާ�H��s8.�xo��c��E���xk��Ã�:o��@g��lwV7�#ｏ�׏��s|����A�M��1��6�0�Q�ϡ2,qp�$�"�<�0�O��cX��F�x���>'s$���)�v9\��t�MY����$C�*9���4�7NE�I������,kf����(�U�qkV�P�Sv�����=c��p�M0��$�F�@�a�f�d��>F4Ͷ�ٔ��Ma������5��-C4���i�J����� ��h$�����ssy���#9;�B����S\������{nӱ8fB1���On�-��nG���:bp�4b���X]����~�lJ�+�N`��Gi����B��I��r��mrń	�x�e����fr3�a+�ZP�d�t]��z{�AcYb����<���r�ؼ���(�s�����^�k&[m57g�<A���k�5�)w��O-�;$oc�����1�q��c�
���`7<�|�ffpoq�Wo �)�<99���)
�W2 �X]��ħs
�J[O^h���`~q�Z[G���qٮ��1{.�����;��~���I�Z^�۷�J���p��~�8�:G�7�K�x(�I�����'�KaܸI5�&��cZ&�Ym8����v0�p������$O5�	iy��60볒G�I��~�>2ofp���`Ь1r�L��&��,��|�`0��J�O�F��+�0�k���4W<7F��df(�bK����������!��BQj�L�K�U�A��DA˨��\�d�ك%v��Š�xT��*�J!'�����4��s�B��Vq|q�B�
д�o�+D'�z}��&��F"�7f�~�����f���ou�[���V��&sk3h8bf_x��2����j�I1�1	we��V��
�.۲�W�W67w�|��pCgv��;W�!�+=u�-��5v��F�M~m���I�c���^��iw�6��x���WH�&�2�M:I`�(M�&"��2�f���7r�g2>�@T���{���븯�:��!8Ԓ�	<�G������i������:n�.	)>�uP8�@�P� �K#5=�z����c�)s#u���t�}�����+E�;M�������7ـϏ�����lV��T4���=�/��qY���ƐŰ���X.o2��{ؿ:;���A��iA�su=-��fC�� �0�i�kYe��l�'�G��2v<�t��v��>�%����L:��כ
�Z[�X��7�
�Lp4��y�T�&�D�q<��~IIџD��jU�a�FPu$�^�fx����B�P�4������A
���N6�v�:�鷒�����	�(��2Li/�����}�)�cQ$�2
n�a�|>1�4\�EQ�Pl�Q�Ք�y���5i}	��F�>Y�������_�� ���C    IDAT3���k�}ܬ��a���<h�M^�q�����L�4�9�R:x"�D�77�O&-�QnE��Z��Q���c]��Ԕ@�\6�-vG:Z��G�s  �^'2�n{\��)�z�񹀬A����`�=&���A� V*���� _��:��o|����O��׽C3�5����Y��*Q5淧����I�A���V0{�����|XHM���*�-�b}*��/$��V�(���\U '@ؿ�8)������+��yun�oݑ����gg*Cj��2�H(�T6��D>���w��j�$Ú����4�M����˃]�.�
�#qu�����xxt��'���>9�jt��!
Z`��n��*��&���Y�ç�2t� y�m�4I��+�d-�@RJVR���aP�:O��@�Z3��}��A��I��} ط"^���v�/�v��C��Х��5{k�i�-U?���#iOg6͝w)3~C{4��0�(�XLXS��&�v���<
v�m!�M�Y�@eXNWa0+eB�
����Wl��s�lZ����
�^K�{����@b��� �pȠ+x�x<R��Ɠ𴚈�<H�}O6rs���A�o���{����I�����V-VBb�.���xB�'�	c�F��G�^.s���ƾ�QV}%�	"d�a�`e�,m����]{z��E��˻�45�дb�R�$1Ϳ�.��^W����'�g��8�n=x���5�:F�S},�aޏ	B��.ss�����=Yc_.(@��E�J�r,�h� ���{]� m�u�j�"v��@`��̣7@��G�F>����<n�,cij�@X�pNL�^��:v��u�����ܴ$��,� �g�h�u�{�Ⱦ�w$EkЕ�Ь��>��~��YI*�L}Q��E��5%�X���QA�<�C��ώ��2����{�b�0#a�Mz�e(H��i��sV�k2�1X(����LY�͹�q�YZ�����VHb"u���t=���A�f<|}^'36�@$S)��9��t�����ۢ�5秒�`��tW�����V�4m	�>2׍���S�x&� �l�Qi6����۩���v`B��I�v�G�P�Ϩ~�5j���xM�$�6V��Fi�c���~?*�=j/K`<�I:~�W)#��#<�3��K�?>���<��}c�S��G��Ϟ���p�(��B�nD�3��$\��
e_�,��%Vi<�����[��5�dMnx:ܸ�Ͷ��Q�7�S�|Be��d�#k��}��LL�'��5P�	21z�`�����P�9�O^�	`��.G�c����*�p�Df6���D�q-'�ᦹcr���n�eO�qiQ��~��T����	��1Ka=����e,M�"�K �e���1��p\:G�Q�k:���S�|fV�hʌ+� `�����q^����)��x�M��oci����M+8R]���'f7�h�͢T@�mb��@��LJ�}L(��}�����<̴8�� x���s6s\Tez�K̒�b�Ɣ)��1�0p���5`��o�PTY��I�o�|�x@�rYL�rʠZ�"���,��=-��8����w�g��h ���0y��@*&ʐ���~��$ܧSD�It=�j5�DqX�5�QN��+����b�I93��=e���^�.Հ^̮-#���N�+�=�l�����k���j�A��?�� ��D��]^�ۍ���o���O���9nU~�Y���r���D�O�M�H
���(3�Lc�a���讧|�%�&�� ���ds��WP��&�6~Iz0�2���=��0H�|���izn��cl�-�^n�S��^~�ei
�f�`�f� 	�k��8+t��l��ۡk���W%�a!/NY�&�\Vfb{���Y�z��\f(����X��{#�KH����X+�y���S�yG�::��y���װ����`��46��6�����bi���(1l Z�uZ�=>T��r$N/3���y�^]W�cp�]���0�tL"�~�h�v�}v��fU�4��pj�gJL�k+���H�?35�H`�ӤT"�VA���;}5�ō��V��IƳlで��(k�P-��G��
��K��m�'�5(�MT>�������B^���h��F���y�� 1�9�AUr��F��	��V�I�� |>�Mz�R���X񩴔��
�J��LV�@�e��ϒ�!�J(���J��K����Џ3�e��� ���ߺ�A<����YG#@�=F�#����փl��A���?D��'��V�7~짾�i�����W4e>�V��q��S��Z�:����fn,K��'
��2���[��prv00�`1C��u�*p�D��2��@X��)_��Υ�B�����>N���	�e|��Th�NK_�a:��0������a�(���+G�Ӗ	�n��3�V.�)Of��9i%~#�6�9+86��taqV��&��q�jy�*���������Y8`x�93R�Ng�W���q�
�g'��z�q�ډE�7�L<����SY�'s���$w�����E��m�~\���m�Z��Pm���:6�KRP�4Z��F��?
�����Lj:�x��������>hcD�&��R���R�WC�H��T�r>��-:��V�q]�P3�` � �V[4ŋK��>D�Ĵ{�6!�^�/-bvauz|Vk�wZ
h,I;���=Y��<�x�)64��02D��+Z�>��Y~)9���p��)�8a.T�(7�h���Þ���tp+�Ʉ�������R�A��K��}�u�W���XC?D���UG��\��l;��>JN�)9E��H�8��w�V��o|�o|�����76�;�t�*�M���+9翬�F�?sp���ۈ�h�U������K�I�K=W.NH���Aӓ��±n��*s�b�H����Š��=x˱�i�p:pn2'a�rL��D+-r\�'�3������i��	"��ǌ�I�Og3=M�$XіX6�Pvh�o��\p��kN����G�?��4
���(+���S��5NT� ��K�!fN<��a꣎>G��6oo(Hɔ?�\ ��hFx�T$&:A�R�N�FU~
ln�o(|�Ǉ��9,�,�Ԍ��d@�}��E���RW�
��"I;ԠK�5�IN�{���_�-)s�ka�C��EU2����s�be�l��J�C����̏��Zs�:(]�scP7 b��L�Tk��>�Von 3=#ɦ�rI=���;�:0T9�#�zG���Ϙ�){a!b�:}�Z]�9��A�á�Y��( :��G<�A�U�e��,�i!4<T��)k� ��T��-�`ʁI�QW ���Q�vK�Vև6DC�Z_Blao�n�~J�E�F����2�öu�t�u�<^�ƒ�'��]Z�������o�C���a��;'���7�!܈��jZj�R�]ύ��&A�?%A�R 5����6��i�+KUJ���8�B�{X�N'���oM�ݤ�/����<88�Y�/r�J>ı��U9e*��d�b'�����U�5�j�#�����L�L60	j���H\���D��L����ף���K*��S�P��h�hP�I5{"t#��s��4��t��<��P� ՙ��|D�K

Z`�|�f�z��R���z�"8A��G��o�M�@�;D��7��`��@��f��/`�)*J�!!�e0��3��̬�Uo������EG�����̨
͍䋅%�Ĭ�O̕���zo<HXQ��̭�U�ff�
E�Kbv�~+�;M\'3zM ۝18؁z���C�%i0�����>Z�:zVb���N�������C���p��]$�S�FϊW�4��Y��Mã �\+��3� �üʊ��"<����ǵ"ж�аX��ZM,��`qm�T��8��Є�I
�1�q�� �u���I�"���+e��Ѹ�(����:���S��ـ/��Q���zU���(�	�۸��l4�iQ�r�Q�����8qn�����K��O��������W�ڍ�9�~�U����&dc� �><�!�Ѱ� !�v�����f�Lp3���y&?�����5ev�E6]'���]�Po�N
���A��U���J�Iܗ뵩e'C�\�~�����J=*f��p�%����73^+���^	��Zed꙰�jpM�T:MbߔLy�CN#� b}���2�
��bO����sc��n�^��r^�R��_�v�'���2��ZW�a���U�ZS�D���0V~}*?�Bh��RXDC:h�1��d�d|a�=��tkm]�7b��վ`�k���R�h���){Un�����d�����ƴ&�S��Fft���&`���ҟ���� 3�vW��dV��� ��0�/>SN7[�A��J�9
W�D����#N��IJ[!:'o�ה�/���kwqvx��I����/bznV��F��b��R�X��M���g��053�Z��Ó#�]�K�D#
�<X�!���hf60+���A��}na���F8S\n6Qn�������;92��O)�`$�h��r��z` g��k4�3����LJא]Y@�lNqV����`!D�y/[&��Z��ø�n!��[>�x�����n�MMK��?_=i���^��3g�z�:���Li:5�H�"�hZ��7�(�3>c@��Q�����k7'�勨gd!#*�/�Y�P�v��pN��������L���j����U�	�4�<�qg5�xmA>~/��!���2���yiKE� `��Bׁ�c���'@�m��yu"���{�aL����h�Hf5-�'�
n,f	.�1K`i:9q�5��a��f�YIQm��q�D�{��C�%����W�,�LH`�h�FHIw�xߧnTkaPmb��Y�pP<d6�U.���P�F�/2`�U��t	a���PD�TB�A�ߑP���0��oev�6��+SE837ra	?h��֚*�U���uד�de~����Q�XN������|�c@�^Ҕ�_��1أ"d���vWA[��� �W�����K%�)A�Q���N��$
�`��v��y�El�l	[�v��y�8(��6@���Ť�)R4��/�aiy�pDX�v���n�J��$i��Y��D��y��F�H�:~��M�����-1=�A�U���Z�^[����
�����v�fM���
*L���'_����_짿�Fpn����6/���Z��:�Pmx�����7���@�,5���z�T��(I��%K0v��J

F�I�=
6|������bIe%�i^A�}7[ۻߩ��"��ԝ��f��~�F�ሰV�f5<�I�G�o�!OpL�=�ٟ�)�t<�B��R�d�=��ya:!���d�N	�d_I�`N+�#Ľ�;t�5m��A,D�Ȅcڄ�v[�D�\��%�E�9&f��Rce��P'݅j��'����_qe*���8�d:A���F\��^-��>�g��ƕ��"A�� ���*u�
5��@��>�Ʉ�/3���2�10g�i@(�w���L��I��;�����e)�f8�6yI�Jf�H�R���O���Pe���E���ʥm�{��i��\{��gX,<0�BR�����V/���N���҉�🎷I,b~v�xR���4�9��-�!��Vp�=:ĳ��qrr����w>�{���R����prvf�`�Rq&��RvF���U�BQ;/�H"��!cf6�p4j�����Z$���wt���S��_��k�+��G�{҃t:�u���^#�-�fM?�Q�}>\v�8kTQv� ���^�W����{��QoՕ����x����^�����ҟ�����7�j��W+��g�F�7C�7����37����c3k���&	c<A�,���R��K{��q�:�2]��'�%qR��=�O&EK$v�n|]7�f����;����d�L�}���B���f0B6�d��r���bъt%�̓KR/v�TK�cc9J��7��/ ��eճK��Ć>�gg�������8�1�`[��G�V��	�S=q/�'��$����}$��ɅH-NzF���2@.�����L%�-���*k�V�]�.T�Z���a�8<8x 4��|�|V��s%��fy���tg߈�-ɾ��/FJ���FA� !Dɧ�i������Jin��Y��V*�f�pB߻��֒�#t�/~�����P���iTV0�gnl8�e�זW�x�T^ǳi,n�"H�m6�j�����8�;T%q�������k%���'�Q,����'1��­�5Ap�g8;>�����f��v:-���J�r�MO.��C4"����	����,���}���i#�8�r"���jn�]U;>?*��k��m1H�k�:�	��?Kx�p���"�E�fܦ"q,�[�.l��\|�O�Hp���uk�U�'{��O�w��On,K�\P�����KQ�ޘ��� ��˙�L�_�u��,m��}�zYc �E��48�	1.�4�fe�d�%9c�W��I�x�,Y/�`oKg$֢�8'f]1�PX���cl54]�|h�me��K����<Hx���$0�F�Ї�;(��[������l*c�cv`P-WT���[]^A�RA��J��e�0hz���R<~Y�����,�777ǁ���$	�͎2��D�w0���g�XE3q5�#��f�3�R��Z����R��f
;e>7�t!��jקdp`a�\������	�q� ��c�/�)�a��fIJ��
yM<9�`�Ȁ&�N�FK�s�2Y��l�R.��f�Y-��,��
a�a��sv٤�v7�b�zt�~�o666��BQ�X*)!���4�#O�������H;���Օ%H�51���a�:0�sy�^^Í�e�����C�_Z�R��Npxx�B�d�뤊��"��fg��qtq���:z��|�3���D�N��1�)��=�A�խA_�m�(�@�?��Z�3�\�շ$sH�h�^`$��Xb����/ߝ���7�~��|��I��O���������E�ABD�W37�o���h졠E'�RfOײޮ\ �rK5��p
'}<9���Z�.q85�5n�� }+nl���!#nk�f�t�X��DvʨbaX���b�6���5H����'�����et0Ppc�D�Q�^�,��2y��Lx���$��૶�����_h�8Oc&��;y��~� .N�T�R�a>���,�A���I� ��A��M������)���=B�X��Xi"�9Qe	�Ǵ��"a�A-k�'3)��?�� R��]�������.RA�0Γ�'�ZV�ө��=�9D�D��2�T���xR�t�x�%��D�#�ӄ!Х��<!ӫcvʉ"/�X�. Ą���2:��BH&
�̪*����Ѱ%�����Ѐ��1��@���}S�n��*��°�ѠL���d��i#�������
dL���{�垠1wn����wx�s2,���6��t�7��qsqE��U�GG���	jR<���O����Z�� Cy)f����	�g�ܶpp~�J�n�0 �0��Td#g�I�g���Lb�#���a#�A���(t�����[m�����m!���`q�oN���7�~�����߫��A��Kg�&j$�����5-�,K�0]p�_��f(@���.��B��B����enn����� x�@������{D,	5�4��q��2c���z�
^���	��FΓRN�d��g�H-4ꍯk�Lɟcpk��-Q���Y� >�^gf���x�/��)ֱ��Mc#r�$B�l��=���
ES����707�k�3�)������Q}��m�.-#��ŋ�e0i7Zf�Kd;3%�l����nJ-ҀWA2�M���\f�h7�c_:6��T�p���bp\�tBA��p���2�5_W�'~ U�����1f�����tA��5Qf�&������RY*a)l�YI��j۩��>,7Y)DX��U:��4鶞�ϫg@� ��,��e1.xk�
 �I �ˍe���L6+��栋J�#8�?]\    IDAT�uv�=�..�΍���#��n&r����'�:?�j~��n���MԊeGVO�KHOO��|w{{;q/��@<���*nݺ��TN�Z���+�Ѽ�j1� �����]��	h���BaN�M����1��-π�eND�*|�_��a�-��t����_�l>�'?y�'������f(��G_��[���Z���:�
2	Ѵ���!��\�,=�s�tmH�.Q���ˆ��4:k�>�zhV�����j|\�m:*�S���?�(�1kb���.�f�٩��������/b�T=3�����G�����0�d����&(N����G�㗱1_���S��L.���]�51����&p�~����{��j��#� 6�#����l����w�A�ZF�X�I(.��'��i9Ƞ������%������X����!./��
���Japc|�dH^������Trl�"�NW����������:
�XN���r%D���jt��P�x�*��;�5P��'ׇ�T�=Q�S���S��3� �k�Bg�~O��v#�h����*W������}���g*i*�y/n��zuNA(�t0sҘa��v&�d�G /A���[����Ю�%����ܨ�"�:�!D^�x�g/_`��Kd�)ܻuW�[-��wx �"����l��ᶆ"U�n��ծӿ��]Le�qzu���[����RSܠ���o+�6���0ݬ�(
jKSfol]�j��)`��x���IP�fߕk�U���Q�����7~����~#��w?��=��~�Y���VU�.�Zk4��[���5�B�ېY�27�����h�A�4�x�иx�&������a��^U0���LZr����)�pL�M�$r.�'����4��3"��Cm�������Y�))��d�Y}-�
���wTF���$I:����m������[}������)W�v��T�eq$�\��9��T^����+�p�r��d�>�G>D�4U1�9-��e42��'��he��+%a��Y8QA���q�rC��E�n��L	�P�,�}��`E���1Cb�Y��%��L��Ϧ�2`b�L�,tz�d����)�k[=82&B:d���癹0��a�|F�����w��ra�F���:z6��Ig]�O�X�4�031"�	˰*4V�03r^ܸ^3@�`���{�@˴.�5r\{}ӷ0����<\f��ԻF��LO!�N*�eB�a�;�o���[zН��k#�L
��R������,/�w�A�P��с��ydg��d���ob�`� 3�A�]�f��t�J/v��h�J��_�e�T��(�`�e3��5dd̹��U�h�~AtH�d2������f�{dY�![8�fp��XI���ϯ��ʭ�?�o־���gn��џ��A��������^��ϫ�-�x<"�!}K��&ʒ1R�F��\���4�(l�au�"����E�cw�i��e��/���s�X�D�DF��ܰ'BH�m֫���h���/�ꝳc\6�c�_%S�!�b1�CQ��꠵nU�$y�*ݫ��E��$�0��F&y�3���i�MZM�\��	U��*��з�L���������bs��SD�]��>d=A��^�Dc�G�0���2�ഋ����墲n&�f��'�8?Q�Li�R]�2r#Ca�':�W�UA6rӳ
����Nt~psI�KɎA�+���F;�Q������E�O�"�l��V��%!�<I�CR�l0D��l�N��o <�,y-��`[N��C�f� ��(��2vV��,ǉY8{���d]k22��))>JP�(k�i����9�1 XZ"j��WwtbQ���"�I����4��p��
y��[/^j��ֽ������s4�U��y5�yؼ|�\A�Y�;wpuYTpc�9��n��{xy�-X��#�=ݽq�������p�϶7�`�.�9Z�����p�B!M#P���z�^�1/a�B�����a���%�!&�@H�2�}�=�;I�bp[Me���/��{w��՗�>o��?Ȳ��}�?8jU��A���I��7���9�?`6Q�3�*��n2��BU��u�[R;$i� �ĵ�<Vg������[�{�j�vcʘ��Y�/,am:�$��������g��en�wl�2-.��8,_J�����NS��,f���ĕ�q�P(���T�e��r�t���,6V�8���3{�̍���P���e����#���A��B�7B7���A�$�~]��@���U�;�(��:��),�s���t�V�kq�czfƸE���SR���4��h��p��p�M���OrN�պ�)3�S��}x|�����ɥ){��-AJم���Od�[e��t���T6� �L�V�j�Dc1�P��3KJ�38*�S����K��Z��9�ｴ�8�����Gz�̇x-~�YjuX�SX,Uǔ�7��G�p4n%�M��J�b~�S`�����3���r�ԣ��[(�I.K�t:#��x:�x:�tn
Ssfj�������������T|gg�'�t3kO%����}��E���cgO�yy��O�_����Er��|xw6n�ޝ;X�/���O67�p�9*�����,Mc��p���ZC���}g�36����o��:�|����,�^�ʐ���!I��`+���[󫿱����?���G#o��o���v�4�o1��H�����A�1e�GT���(Q9����9�̴����T��1�t8.���Y�Es�Z�(W��U^����6�Z4=,�,cei��<�l��\����յ�0vb��9)�5KFh�hW��.%}Vf�qgy	OXM�z�1r*E���JQ��p���U�Z���DoH�[7N��qj���G���|OvwT7<��}��'H7K�� �.TP><Ai���2RC?ֲ�X�ɣ[k�Z,�m=��2��Nÿ9L`�"�RK4����/��h��!�?2��F�`�Z=ee-j����"H�jt�8�8S_�A�7ș�ƽ�X*'�Ò��6Í4���:Ii��l���1K�7��6��Ph��`����:���+7��.�9G�#6+���X�� R�9�yܓdi�>�������3�k�Ϥ"�@	�Gf������ngw�����W^S�K�p#�+	��$AL�L+��#QcP�W������2�S����������n�n��=��g�����uMI�����v������f����e���}��G�O�|kSW}OЇ֣����oɥ�8�Gϟk��F��X�G���z'��>�2b�x���9�`� ���>��eMP�=b �PL��j�V�n�@��V�S[��-�Z&��o�8��|�+��3��:l����f�6�[� O��#�G�fl���@����n.�9��w$�I�->0*�X�Ss�9���X	_��)������Ԭ��ܽ8�q�R&��b	��u.���T�`�~W��J�.�)�e�%S�8Qd��Q���閥�!e�j]��u8���q�Gg'r[b3xmi��n!Ok��F?a,�|A�l��@rzH<>f�����W8�A�
�aK^�0�Uou0h�Ы6�*��<�BXXN尔�	�OC2��Uh��?��a��4L 05F6��T6��}4ZM�_�Y4��p嫒���N_�'77��TV=�b��G
j�n6���߲�� b��X���mw%'j��\���W������,6n�aeuUϋ�\�^����Qk�li��1�87�7ql�F˔�v�"�˨0[%F�V�4��[:N�:V�ˍF%���JP/%ٌ��h<n��DH]�(�&\�X���+�Zt�Ji.)���]�*��P�n,�%	��/��`���N���X1���[
p�jC�ܣGt}�9h�wO��4F���CGJ�K��/b��?�g��um�Ff���w���ￏ��<O����<��B�;D�<r����k训�g��e��R�a��bY�zx�Y��� J%'h�3�ZE-
��p�F8�r*��~n�W>�c�~��kj�_R�~_��?���/�|Ԯ��a��~ܨ�J��tB��ƍ�q*�׸��ۮ{n��$ �uz(C��У(}{f7f�o����������Pel����ÀW��a����1	NѬf4o��ڈ��^\v�����<��ae~��y���Y��3Ǟ%a�je����\d���*޹s�pZ��˳s���{���� ,`s
�y"�P�5�u|��<y��l"�+��>��A�͎�*��
��%�����G�D�\R�ׯ�T�R��6��`$j�N�l;n����1����:�G�%9O]N�Zm�V�h+@0���_XY���N���K|��_���!�..M�F�l ��̆���ш-�������,O�Y�|�V�� r�)т�gsȲA�l��r�d��|�Ͷz���)�����
,�����5^�����~�~��T�S�5h�B���cpY<���,��Leǥ=��H$��C��`5�%�ym#)�*c�s׽�*�e��`�L�	���*�Vn���{�[Z�����x��}�.n޼�v���O���ÏT���r��m,/-
��u����L�RrD�K���������|�g[/��ʨ�<��m���{��̊~���3<|��nN��#�O%��$��t���*�� ��U���?��\4}O�j�X���j�,@�o8gn���˷g��G>���xp���oF��ÿuܮ�O��ʲn]&���A(�ϣ��3�$>�4�%�h
.�����Eէ!�Ӂ0nM/��5,Ħ��N��+;%�(U�&�P�CU/��t/O4�Z��Cgp|k�&��zh�FU����#��%��TLX��ǭ�%�L�a:�@MK'g�U�f����^D��i�g'(7*����훷�'P�V������mԚ5t�u6�#73�U;b���h:8/��k}_� �~��$B�?[�1I��*蝗���E�ᶊ]/�
$V*�����3�,��L3~�A�}"҆�a "��5�t�bE ����y�I����C`���c��&NO�����i��F��x�l�������bN!�M3� iN~dRi7�g�D�3@��)ezD�
�zidKK5\��&�)@��$����sxD;d`�r�U�aW\a���?<�s���(�A�ו�eMp����fP��'�L-;ԨU�KEN�k(�*:|ܴ���σ�33?����P��cR�jY�Xtcko[;;�f7n���Ҳ��'O����b[�0[]Y�ﾧ
D��
WEj*��T~��p�Ock[�:��81���o����*ҹi�����K<�z�b��QdП�h	7*gK*��#�^��/nZ�`�?�Z�z7���>�̠���Aª��� ���{3�_�b?��?p��>y?��S�{��r���e)��x�3@Nfn(0{}�nD�k����n 9�0��.0��3�7q?���7o�/����CI��(#����TN�x.�j����>�~�`��vDg!�<��ݛw���DQhV��s��;2�e���3'��VpoyK�",G���.qzp$n����Y��%:�^�Y�
�����rab$�������e�4?;���2�ݺ��?&������#|{�)J���I�A[�����x���"�CfBqD^�k-1 �8��8��t�(g���s���(-8�Ō%{<�7D�M��)gݳ̎��~���N!��Q��?�����ى~6����C�[ q��e2
;[�ꅱw&hIؔ��d2�H�\�@ȉ�2F�
T�Z�}Q��mԚ��	&��0�8n&����ycX6�5y]�/)��az�V@��U���Y�q�E-�ʸ���,�\���Mg�L��A�I�A��NO�p||*m3B}\pS�]�PP@ޙ��֘��"�-'��ܔ�1�0�q�Tg0�w?�}�����2�4޽���X�/�*K�YU�5,,-j�P�qtz�ÓCe�*��]���&��^O��6_����D��B�6Uf覿fX<���
ǙE���=s=!V�u���lw��]���:I�P(��Hb��t�W�����?p��n7u����a��뇭��9�S���4�z	��N7�ٝn��S�^y̩n��}M9�B�@�-m�ś��E�V�����
��NO!�������a�">���^�\j�T�`p��E����5m��c�hT����I��˛Ͼ�o/o`!����������)JW� |0,KhEG��;D�]���|�<ɂ!���"���Q�3 ��|O�X�Y�o�������񭧏���gh�<�|��B�k<?)���ux�-�O/�s�zCȅ�h����*�6Nn�����s��
n"\��^��X6��r��=��A��Y��ݞ2�Ľ#&X=8;���啚��dZ%ԣ�ի��
�"N��!n��Rpѫ�J)C:�?����	jT�E՛��I8�,Nس�@��8LS
�ev,f�;Q�W��p~q���=���#��F]��U�`0Ѝ�2�O�I4����E Ȯ�o6;b�Dc���>��Rc�p���9H(���"����卥����eHd��F6��$�EӼ��.���Ln
�d\��dz����@���u����|��x����~PIemi��,���q�4-�����0�P(DRw
��ܦ���J�g���K�<����).���J!p��ב�5�2X��T$6j}����g791���S����pY.j���"�b1��wy���3��>-�=�P���V�W���[�Mb[����l@JQ�ˌ���>J�����N{
nܰ9O��8�]����u����3#�X��s�jd�S^�W2��">�}���J��hv�zB��{X�- ��QŃ�x���0��u���[�e��_��]��=���7		P�B�<yr�����N[{� �!?F����B���c�	��rg6��j.�l0�n�+��l>�Ã-���!�M��]MLG�6��6ZG�vF��V�*	
�F9�1MhQd)A��w&�[��6��N���f�$�v�K&����H��9!M�����'O���l���$��o�pq�ʠ���R�(;N��L�dg���7�F>)�&�9����E�;??+ƄhS$�ǣ��*��x)Wj�����F>�d��\&�2�Ns�@�k�x�A��Qϵ��L,��3��"?р���H�6�@��ܜNr՘g�t��bo� /�w����j@�lL�:EB���M �	>�Á*�x���W1����&`������<�9��SU=3������FC����(�&���9� x��o�\���Ac�(4��X�t��}]�wC����U�H���Mw�9�|{�{���5:L����=L�x��}&W�T�VXGp _��>���n�K���4Z�&�1Ǚ�p�X�<�:����&��A}R
��C��㑠ũ&Gm�kF�34�D$\��M!MN�'�E�L�C���$�P�R�B%3M����G6������:����Q�����7��P�Q�5�� f�_k��n���ɞ���Ȉ�/B�0��CT�-Z�.�SF����12X�Vj�e$6����P��Ϥ�����Ѯ�Iv�al/������?���L���\�M��y��ݷ�;��r@}��Y��2LO���5�Y�����z���@b��d5�ӧ=��Q��*��F}�h�n�������9��7��/���z��i��ͣ}�Y�w�����ՈI�<uNƌ�>+�*=��F��g(�D���+Ȃ��D�L�����nP��t��#�>��i��\+E|��+4^�b>��sP3�"Ræ}h���}����:��t� n&qp`P>��&��t�;���3��v���0��H����)B8�+%���#���2�2YN+!	׵ڻw?�Q� �~�"Ŏ��\2	�Xs����}�BVD���*5[    IDATkc>4���Y�W%@<_���ؤ��Q*8b�q2#�kU5i��ôs�n�羟1�k� ߇��57+j52Ӗh����n���j�\�0s�Wʤ��p\:43C��E�3��H>���O�� �禦9*�����0U L�X���)VFA�j�ʨ'B*j�٠3L�ut�z�> �5:N9����,��r*Kâ�n1�=_an��(�.0yd褦,VO^�u��4	�) �M�6�JM�2��M )@ֿk��{����w,��&�����������1Mp�Ps�3w�
n�\�:�K��6�e��|�NZC�C�h`�\��]4�9_g�,1�����"ݹk;�\����#�q?��b2�T��~��޻wQbR��u�A�<���WG(-��+Y�m�Z�����ٱ$J(���5��/�����i�n��\s�-ކ�=�ؓi@�R�shog����=ph?�U��e4�Pü]@����6��m�ퟦ�/Ӡ�ap��4�0&�z	6�����ۜ��>s�xHY �ͥ��0�Շ�h�'��`�#0(�����q
���!����t�R��cWq]
����8
�-1���I����Ɔ,f5�gԩ���PL]�0�2�WE�N7"�c��H�J�	��ap�օ��㱈#�����O�^�1�x|���[�L ,��_N�k��
HK���S����]���29:FyMI,�#Ti��?�x�h��V�T�����o��яi���Ȩ\)�~�fh!/nX� #�<j&�T]�SA׭0T�|�ȥ�v��t�G��N7D���e��O����V���P-���/������:D=��'���#9��f�P�|��!5|W�Q���!:��p��$��	Pdx��QB<�>�!��x�*��Y�� e+%���m�=3E]��@��r	⛩�����j�X�;G�n�uoeε�v������R��R̍rMF��Y=S&�3Y�7ϯ�{����6��YO�����Ct��8�e*�}�v:B�f<-NFѨ���KDS��k�vڽ0AK^�4�K�!k�=}��<L�l�{=��N�g�.�tD��6^���Q�o�=l��,W��Њ�x�@&�&'��yڽk�4kRR)�Ӈh��]dKb�'Y�JӺ�=o�3h@�Q۵iOk��ط�~�/�[K	xJr/�Mb�1X�-vȝ���H��jq��iw��jP��A�87/�A�H�oL���W2�DӬ��MG+�#���S��i do��i��s�驙Yz�����[BS����yUoƔ�r�	��(����gDIHYy���uEg��ivKרR,R}h�Ny�S��ςP�U!�	'��� ޛo���m�4�����q����
��\H ;�#��n�|��ypp�����%"�LF��b^��{ĳ�j��N�Ӟ�4��!}F�fY��I�R43��͛n�6�޷��	���H��
+����g5�V�D�\��|9�Qi�FC�$�Mv�:�l���ѸBe`�
đ�0�Q=1�����*˂/��Pkz�Z3�\ !�`}��Y:����)����N�ڡ+�*��]���(q_�8�N�l�jV������~�O���u�E(d�K��T];J�e���8�rZ�{��Rɴ�p���u�o>�5��o���;�_{��T���GfKpCA��H ��.z\sc�]���� 7:����%1stR�N���P�DQ����8����Q�����U��A���ݳ{;텠��f�ktZ@ACam�Fiͤ�N��߷��ڽ��@���0�
n���T��@����ؿ�CpIx(���ӵ#�4`e)��h��;H3,v.��;s��!z���B��F��Neh]e����T�r������H���N��}��jH%$W�@�����wIk;$/t�����d�Iv�<7��� ��H�*R�,��ӣ�7:��ST*8�e��Y{���) �jHǸv�`xtlڹk}��ߠ��I�s�\E�/7��EWL̓2�L���@p&�H�Y!����G�����
�Wj46:B�|�3���1%D�h޸�#c>m�A���۸�����0�B���{!����g���I��R��#c�����V�sdT�� �%H��Q����=�y<É��<�#M��M�v����=����`\6������z 7p !�M�'Dި�q���-Y�<��_C�j�����D4e�0*��h]p,���cV�x$����Esk��in���x~�]Ԡ��V��G�L��u�J���4ow9���_�NA;OL`� �a�BtA�I�J��c����NߦV����le��7�%�V���Si���$�
 735�yl��6���uU��=|���o�k�i�w���%�� pK�A_P`i�����WƬk��<n�wbv̲C2�t�� �J��CZg&hǞ�l9��58�Gj�t̚�T��C2�Z����t�|%m���v`��m�`���N����Mw�~��|KD�Y5R�q�N��l��|�Z��A\�C��K Eְ��{��:�G�w�û�f�2�ُ����<��G���]�T�i]m��~�S�l��T:�o���Ow�}��j �M���e�g:]2I!��x�ҽ�F�,Y=���#ݕ�熨u��-7QP]6�2A���ߠ�F�e�T-��7F/z��\.������Iب
����������o'#��6�I�߉.`&�f0M��$�yx��Ħ� }���)"PU�4Ժt�֏���7m�Ӟ�L���[�>j�A>ꑚɼ���	��7���57��#U��a"�I�0 �r3]��z]�IR%�;�H���Cj��<������kuKS%Őhh�F/zыh�T����7(����	��3�s�o��Iߺ��,
[>怩B��P,r��v���,��Y��e5-gRm|���A
,������") ���K�!�I
D���b�z�}��!Z�s�h�	C��
��T����>ni�M�-���<"E��{����1��&oZT/V(�,�.�I�}�J
e$MW��N�Qiw&M����Hq��M5��󜒕�����<����J�ƣ��od���;�^}���L9]����8�- ���b����<B���聡9��>a���PUO�q�c�ax��i�K���fh��},��s!+��Fc�q��y�	ԋ��C�Y�ܴ��7��-�3�=�F�2o��v�>���޳�Z��ĉ5`���Ik7R-?@�%~ϟ�|��؁J�����`�D'mD��F�@����9z`v?��qH�kr?M7�˅�4T�њ�(���x*XY��:К��w�O��y��jDM8Juݞ�:����9�̻�Y�`�7�$�ѥ�v�{�G�-��fJQX�r\�A���
��u�b��4G����追��L? �3wB؍�.�؈^��w�K?����w��9 7�s�����?��:>�)`eL0$�������)Hq8_A�8�>���锓7���<J�sD����������R����_o�7NQ=_lT�J�o���i`@����,,pD�>&��z!$H�b:�i�5��SȂ�&pR*���������k�l���C��t�u*���顇w�?�����?�Nj�"ҵ2��@m����	�6�s!��5�@5Z��406B�a�\���d�� �a����	��ޏ85̪�\2��]��{���ER�K,DZ��9{���j�����Z�f�.-�g8�{�D�j�P���ʔ�B��d�����*�b����u�=n��c�f�Z��K34�Z�i �� �)[��G�ߺy�~�K�"�_����h���;<�7�^}����v�Ԋ�A	�;��WQD&��t�O:p�8\&ʲ_ �A}3dpK�e쫜b:��uT6KLd� ���ãN������ ��&_�z�Tc�v����Yjy=
Qc����n��t�U��M�K?;�������������	c���Lj��3}�~��!�1�h]Ȍ��Cr��z�(ȴ4=˭t�Đb��ʩ$���Ȇ8*�P&S4j�!��? �'������������#ؚlJ�Tߣ�Tre&&��L���A̍���̶�+�'FX#&K���1w��n�hE&*f�E����q�C�9���^��#��WU��l��Oo�����λ�D�TL ����B��@���]9VU�U:t��\Pw�b�NN�DO}�����=���g0W� z�-X��)\�@��ٽ����tם����p�����(����R�>L�n�f&��F�0aehQ.a���H�L��-&/�$���n����@��� n��n +���V����I��m���=�)��x���e3)2S+��Y��u�{�t����^���v���-��mp�8��<�]\�%ϣ�g�d=�Y���
J��E��
�U��K�I�OS��S��"����hb?!څ�������'�5T�iH����¤�4�p�	D�%&Mc�蠕%��y�&�[��/Q�H��%�����y���֝x�jeN��7�i��@��.7Srf���Ɓ�O�����R�����9���;�_�K����ۣf(�5(H� ����0H�0��c��sG�AF��B_f��X�c��Q�,��v�3��P�n9���ô�>N�#�^���K�ԁx�&S�0h<[�gs����V�ҽ��{�!_GA�����6L)�d�~���LН;���H� n9ՠcFƹX�֜���&�`��C�P� eB60iqd0@���w��ٿ�v�N�X�g�ԗn���PwbpT*8�s�L��Y��}VQEj
�&�#��hc��0n�,d��&"
Q� ��.�@�Hk֌�0���-�Mt�c�T_@�%�v�����~��[��;�l"��a���AǴ\�{B-#�f>�� ǆ!�Rׇ5b� �q��|������>����g�1��!��0���$�tm��ޟ��������g1�%CZHc�\y���[b��m�b
B�E4	R%�o�^c�f��8�ei̗��tڰae>�#�yC5�tڷ�0}�71����Q,t�uCf�#�P��i��"f��?�¹Q�ӦSN"���9�G�v�";���"��v���h`�g%��:f������Q��*RnD��_��{�B��m>�R1��@	��	�ʞ"d�?N���@�%�h��$��;d؞0Ǵ��A�A��&{�n~��8RtL�vL����Ys^浨�3����02�������
n߼��ڤ�|�a�u�Ag)3���HG����LE�;��*�(b�D�
�,�����F�CO��bк�0mĠ{�� �@Dvp?�:�����5.z�����o�ɥY�3u�&�s�ň�*��"�36��D��
K���� ���^�2�P5�۱cki���d��%j�H��Lc�)ep���n�����BjH�t�#4��!_^F��ڃG��Y�����~�C|x�Jȵ�XP� F��d�\*b�lAvΑF�B�Bԓ �6u���v�!%��	 �(�1�����{%E��.��6��b����gK6PpB�;F��*�f�����n��N���i��K�Cw��Wcb+����\C*�n�br�����f3���&���g���O=�T7�b�`��� z�^���{�cp��{������@y�i�ДCʎ������H�
D�A]a�� nL��5f�i�������t��J���_���	N$��ݮK{��Y���O�o�x>�n0ꄹ�f�M���<2�6�ll��FZ.M�����=�ɴ;�&hڵ����i)H���%�@�T��hDm�܌H���,�g�muY̆�QJ�PoX��)�<�x����+��}C�>4�b{ ��K���M��Z�T�;�r�Oa�C��P�@�#�hfa����y�O;��|���=xx?���n ��Y2��Ɓڇ7��� �V����?�N{��L:�8K�Y�OM����%�Y��e�[�t���Wn�������!��]��� �T���.���+�η� �m@A�V(р��Ej�m�\r;�k](Yae�5�4R��)T0#�on�xM!�D-`|`��=�Z�]�p�ˑH���!5>ۚ���Y�D�#�YH� n�� ���@��j Ԩ@M����}3�t�n��"[��.�
Ea$���Pk躔꺔u%*y2O]��BP
i�Yj���nw)t�Q5А�k�@�7ņ�u���!�]�g����I'�D�}*F�p��D"7(	7�:t��ӏo�	Gn�M�um�l�<���7b_t����"�c�����ՁE�7ӯY;��; 8P-pp ��B����y������~��A��2��2��,EL� أ���B���6����&���,�k��<0����7m�@�/fs�b���&�2d�����l�i��}��3��owP��e�u��&���Y�	\ZX��!|��Ad�(�Mц㏥��7Qa�B�'�}{vQ[����6��-�
��ұt=�-��(l��=3K��%&��K�G�	%�z=�SHͧ��t`q��:K���":�T���� &8��2P�.&4}�.�[���K�&}L5����B�G{g'��C��\��
^�� �l��.;�>��s�y�э��s[���Mx��K)NK���c�|��U�^ظ �ƪ�Ѝ����O ���A}
�R�Ų��L\�p�Q��h)���<����ɨ�<�w�����`~��?����u��(��q��S���Q��44�p�`X���xXd��l� ��3R��� �w�����f92D٣��@��4�!��R/�VG>��o��Sץ�R9P�iT�2�u�<V�8;CKaV��h�a(����
���֩>:B'�p�� 7 >Z��3"#�[�ѥ���n��/`pxu8L	�,8Ʀ/���BVp�X���Y��a��I�)Fd�J<L뻧?�����e��N�ǯ!�B���1����{��{�B:��5��ryD�B\���Gl�8��.�#T��|36���#bܐ)ܞ��r��2�bBDQ)_(q�%�v�K{�`*��X�k�Rv ��5�g(ɸ}1I�g&Y ��f��CU����˾�ir4��h"�>5�_	� � t�U
c�z8�nh4`f�iIo&F�Rb�*��:5}�&�t�9Oסn�������!s��V��F��`��7ZTʄ
)���#;4�PN���LA=�N��b_ Bl���n��Y��1����}��㞹pT#7�[#t�����-�@Y��,��!jtZ��� ܠ��mj�M�x%ܭ�
N�t}��eN��a�C! �p8p��z����s(��˱�87�h��x-��F��!��A��XX߳�� BS��� `�4s���f_F����E8u�^ȡCw�Ue9byā<� �h�X%� �����P[�M��{ ֐��t�f�N��8-�J:�%C [ߧ��#J���\�g�Bv�
�C�cp::���0��z]�P��T�;r
j����'m>�N;�4�j�: ����P[�;.A���l��<H;w���N�ↀ.����Y�ud BZ
��蒁�x����Q
����kC}5�Ye�ŧ=�T^4�M%�5�t�5ZB\����O{�d
�y+"]E=�K���2��q〹��P�eB2Go�� lEZ�(�t�f�Titd�6n\O���,>��B��w&���"@�>45ó��?�SCn�(�Ӝ-究�N�B�3���4�S=�H@�@�mϡ\���v�QTΜ� Q@Mf3��&aj�ό��� .�TF�%<�>e���R��uN�Ģ��:�B�MS�%��uy�J���Q�������l�"|1r�)v�*i�k/��$�=��L�Yy.�5i�Ӥ�~�&K��k3h�z��*�T瘁�-    IDAT�e��F��죝�~g׽�))x���>_gΚ�Cf<$�B��q�\sCH�]�`�ŏݯX�g�<�-�4� ���h7���c�j.��1/a(L��>>���=�k'�#�Pv�4AKM>�q��P#�XH3�Q�`�YN+�0� �� j�A�{,s�$'Jr<X���Z.��gH���bP�3¹I�������,*���gL��eU]�
�i{�a �!�6`S��Е����;�,�<����C��Ӟ�57�Ȱh �HT$����M��A{��c�H�Dj[3�n(}�&- lvtK��	�a�=.�Ǿ��h�N �=D�+��bq�Ӟ���i DF�B�/PIX3m�I���f��� �	0�ẒauD%��@/���x���),_
S_���O8�Hs�Y��iú�t챛��ͧp=���B� ��z @��&�]l��C,��id�̘T�Qi�ʶy>�)��P��cW+~�Yǆ���@V8m�x�Q��2���x�N`aJ����!�����j���T��S�J 8�?�4��Б�d�� ��t湳�K��CO/�Q6�P@����HU�4�!f����8�1	�ua�2e��d ǡ
pC��bY�c+Տ��n�g�^{��Q�� n�r��)�s��ά5��'���l��LN��p�C�/Ո�5�� ��T��a��1��/u���k8�-4X9��Ɩz\�)#Ȫ�N r�9��Kȅ��*�D�xf�G�s�8̻	����`|��"�� 7x� <�w�QI��zL�#�l`'��;��[�a�8eqB��G�,y��"2]�'��e<�Զ�nXn��t`o����d�V���p��gITf�}�`�s�Π��u�x��\תժ|=7�7����YM�	h��]t��$G���P�:HM@��f3񸓈� ��QKֈk��`;�J9�A�:�"Q������È� 955��0@�czs^c��ӄR-T/pLVEtp�C4ߏ:��H!Rg�7��q}�|���{�T4"ʤ,ڸa-m>���o�ʵ։�I���en�;�el҅f�f����G�HGQo+��4�v�R�"ua5��9�Taڃq3�fPD=tna���ɺ��*�v�{u�x�-��/Uϭ��l�	�C#�7s@��g�� 6<����0�l��L�:p��ؘ߯\�c��������Q���ԡ,�E�{qG[��@�m4��q�� C�f���Tkל4��?����G�nڱc��u�7e�/�ߚMO�۴�h��-���]���"���/C'��s��G6#>ҩ�����8��nӭDK�0�1x䏅Y?
`�� �NT���9�GB��hN�d
��X5��x|"
z�ٱl2GDp$��tx@E��JL��8r�k�2����Ʀ���k*2w� ���⺂��m��'�-��̎C���1��v��R\�B�
\�xnpyo�l:`���BF;�^<����#dhP�W��@���Ƙ~>�G��V�e_̙����T[Ã�X���<�L䅒")p��� ۅ<� �lڢ�r���s<��a����p:&_�s�(BL�7Hs;�ЕkC��H_���Q�%��J��f�N���<���N�r�(���O}������uk�M��ӟ�4nv`�B�3�s493�ׁ� ��^���SP@�EG��~��7m��H�f;�j�35dp�*x�06��Q�Ğ��TLgp]�;n�v���^���o��Ĵ��U��r�%@��A �2�5�O��E\�+�xE�G�[x��Y����"1�Ƣ��"%<:���t���g_=x^�W(cV)�0�/����������;X�򜵧�?����={����i����s���65d�l�"(2�����B��P��OP��c�DQT�oN qj(BMB�����ح:�$ 7N�b�%���a\����Er;x8��b<^?���}�[��:YP3V9��Dظ���Y!A��8>{ "V�����Ih�' �(d�yZ����=Y���"=��IЏ��s�%�Pk�1�V�L/�10���e��bg�\&��`��$�?x�7<:���8�'Q�\�n�0EFW ��� �����D��"��{�-.1�e�Vc�P��D!]8�c������9��k]�[3N�t ��<��rA�R��m5439A�SS<Q�v�{`��� �<�Gj�2�o�c��%�q�_� �q���p����#:[�^�U�'Ky�W�&B�nn~�S[�'ܱPD���"^��S��� mZ��N9�dN�!8��C���71=�T�{>-.5hjn�"��ajdp|�;�F1G��y��4X�;҅�'���"��]��?p0�
���$�'b�@�7Vs��Lf&D�/�~Q����މf��T���4���i."5�����m��`�9@���,�؜A?w��`�/*�CȺ��QW��m��c��p���q�J5�8�_���j�C����=G�n;tȚ�[���[�:�]��;Ԕ"�+#� ;"���Bk_�s�ƹ?O) �("B$1T
q� ��4�� �H��Ŕ����Nd���
I$_�C�w��ش���1�N4�+$�|bAv���	7`��� �DnlylN�Ҹ`��p<����\��&���X'B�L-CD,(��DB,����]�Ĝ$��p�r2�A��A��*e(�
�=���/�3����p���-ƉPA}�3<<�\-� "`lN��Y�������`*m;�㇛�;�����=,��TjB�(6F]
�w��gY��Mi��ť����&��ժ�f|����B��\\`J���
�pԤ �v@n�>i��3��2>KJ��ƀ� ��}���u~x=���`�44=$���T$*�s\�<����(ds�̪��MNqF��#m��M��D��u*�۠&�.eY_p��DM���#�D$S��E�tT���A?c��gq
q�sS�k�EqQ����k�?F���9h��W�|��k����y�x��������/D�#|"D��S�Ĉg'ؿ
��(��I&<�m��c�-�
��fH��ttl��O�W��}�1�~���[E���<pڢ�~|�m�2k�L��	P`�)�p]�ܵ�eX��wS:Ǯ� 7�)2�����!��A@c���9z,e�������f��ՎS���>��n$�k���w�Vx]���R�Iׇk`<c	�A1^U��ч���P��E�"�mL�E�'),ݠgj"��7�"���/{r����p�nذ��[h�(VN39jC�����l�ݣ
�\|���''�^��Z���L�a�����P�ذaG2��D�'�=t_�@���&�;��<�.jX�~�M�C�Nw����k#�2,4�,�� �X�N1�M ������:^��������yK�6���q�8�N���Kܵ�D��� �i�uUj5�>D�f�Z��8<��<��6����nx�K�<�`Zf�*�,���N"��.�_D��<�9pQ�74�[�4�����J�0`q16kj\�b[H�P���G�q�'���5��V�=�Zs����b�`@o�C#x��=��uR�8N�q���+�&��>�. �1�c�X�O,���dn(+ r�h1Z��C�q)oXT�Dn�i`�{������=���
nx��>������/����7ޖ���<+���I	�c7�.�z�C�|	�I�F2��O��`�'7"�~�N�4�BI�{p���8��	�~�4�8Q�@��������"P��4�'\_�
�j�8%����D���}�7�W�%��1���
`r$�C���k��ro��遀��HOḍ	�"�p	�b���p��IA�4��b���/�l6�/6�T�/"|�|Z�
���� ��@ �$����:��?���Iw�^E��ވ��K8t�B� ���NO��lb�*��Bm�J��!�� �8��\"��p�y1��{�iG��ڊ�D���dCV)(�
�v������닚`�(㢾7<�C�9iצb>+D֭��o���pQ��Z�
�t�uP
L�%��ݥ�ӧE��B��h�z�k ����GN�NA������p�J,p��l�g�|�1�QT\�fH����q�O
 ܒ��-�z9����T�5"�ľ��_�}�_�����P���܄����/p ��[�E�Yi�T��h���[_}�s�;������w�m�n[
^�J�M�s�p_��@J�MFq�n�_�8g-v�!^'>��kq1��3Q�K�;�����Pb�:���V��Ϩ�ŴN'�v�x"����e.p"c�t4�]�A�H���& I�T 4���'#���|o,\cb*�a?�d��P���S��	����<$�	�h�A��La9���1�,�Q�	��e����"���Lg��9����j��ֈr<P�$:� 7�����;@�'"�N���� ����b�x�  �DP1��'\���e�T6\��	�t)�A�#�� �"Jvuo6(0�������+<Hq��}�T�/�j��X�d�c�Ls�!8lF�쐢�]���+:�I���xx�x׌��� ��L�9}�$6��3��#��I�:9~@��?|����*�l�4��p���'�~�!�/�p��t�J��<�b6"R�^�:O\*���s�T1I�EY(���T��e���q�F<�&�f�^jl���%�0,c�� =n,h��� �"��
	�df��X�eM���sO��_,��E���'C������F�ɉ�J���L)�M�49p���(
dO�d�k���\���:3�������'�"�Ʃ��/DDH��ua��	�g�C�x�;F�T���:
��h����",Ce D�
��1�V"��8����p�Psc���Դ��r���"��S1�#���$B����Q:-��ŏ��n�LF�6�=�����q2�x
�1�w	�)���:A�(HW�fÐ�cכ�Cˬ@��
φ�}=�8�u��?:sX�TZ��I����8�C�  $n�Ğ�\���_��T�">�$�~=��B���UT��,�YN*P��dP�t	l��������rBl���m�ݎ#MD�
���L.���-�����O����)��9u�;1��J��̢����)��ध-R�ƣ&�)���9@(G ��@I6�(�hi���X\�{B�;x#!�Fq�Q�ǒ)�ԅ^߿�6�g�`��
תqء��&xo�떨Y�,2"���T$O4�pL��a��)'����B�
���AH��f�"�������"�=�B"2"����˖�?Z̼��N{h��/|�����`9���Z?
(�0�}?/�a.p�|$�i/
�F{A ��$EA�Da$G�/KR$K�SR�(R� g���9�� �P�$	߇?s�U�|A��i�dhj�HRER�G6��ˋ9��T,䇠�O	D@��x3��;�`�sp���"%����h�3O��8G�$�`����T�ൄ$�@u&�2eEaQE�'?��c�ҡ!���kp��#�? ��
u�H�E$�c�x#���P,��"3���i0�� �UЁG(</�]��u
v����czL�K	�H*��4;8��PK�'?���8���w y�C=B7���yʁ��4�d������������>`L�Ad��XByW8I�>��/�$҄2p�<�.��������?l1'��������8D
��p�2�x]��5E���+���t2�2PC�$<�tX��9!��������`,��2��gB��H�~$eD=�)�l�@8JԘm r�#�MAWRU5����n�^�L�Z>2H��� ,�=��LF��oH�qo���,��>��mV�q�q���P33_����y�3�-+�=�ŷn�*�^�b��hh��$��"��L���&���E�H��a�	R� �DA�+
ô$�iI�@�Rjbb'ᓪ � ��Z��l�J�˪�i�,Ɂ�ㆶcG��I�(]�W�0L���k��*2��X�v�ʒ�a�^��پ�9�"��/T�TUU4MSE#��"�{��E��ya�ы$EQYR�>�5���Q\;�Dx��Q<	 1@��*�H$�
8 �e��� P�#��-��'�Ma�#���K�*+V� �]��1�;���Fj��d|J��g'D`�+%�-[�!�°���aů/Zύ�qQ�����ʍS�ޜv#�øX\�\��"D|��������K�g�Ѥ>�"Ɇ\7�g  ���iq�5�����n� =ˣ�1�e�H��AR��""A�@�U��N���+<d��D��f=\�7t2�I<� X �b�����جQ<�A�ф� 7$�� ���E�ɑ����&uj�a�s�1�@�Ah� Fm�zqGTdC<��*&�']ͤ.�1c\��,�%ymű�� i�!����&�$*��D*�Ϟ<����B:�����s��_q�gK)����k륗��Y(��qT��M���1M)e�R�Pt$�5�g�Ty�43���K�2�.�a^�I��yn��8�5�0���V���iYiE�R$QJ�|h��8c ��繮���۲=�`.�KYSCWU�#�D�P�$Y5�P��-*E�燡�wG."+J�2�,�rR$E~�y��@�I��6� ����BY�d�)�*I�UՔd�B���6�} ��|)�TI2�0�d$I�R�1�*��RT��d��0���	�0�Y�x�t ;�)*\��0�S�	��x,�@�;�{NS�(�"�M>�،�����@EUU�PQ��
��%�8�BE����l
��`�p�8PTt�А $�\.�Ʀ��%5YE1��i:#��+���ZR��DH�ٸ�'�A|^�Bt�Q.�J	�I��pim�@��@@
	k�D(<�PB� �YP��\�/E�$#:�����S�eهXJ���<
��/�M�5Ufw�XNJ4�b~�#X&�c<����v�̃�	�\LĄk�WR�͇��?������x���Q<���X&��Ч��S���bN* ����*���:�/i�#�JG�hB��[3��5��s�-�����)�<���[A���i�J$o���������Tk���l6�u�����`�֭���޺U޾}�477�k�޴IZ����[,Fٝ;�J���+��<�N�Y]��\Z����Ț��2��'|�^��# �V��[o��:�NG��j���JYӔ�fS���׺����c۲$���)a *��@1$U�K�T�iHU�Y�j���5Y�I�d�ZQ�-]�j����x� G���B�)���>�?h���_Q��(�p�D�,)��*����v׵HK��AЉ°��j�Ȫ&ˑ�(z��]�=;��U����EM��"���u]��1b��b���I3H���	���呩��T�4ͮe�|YUd�U"��+��מBX˃&I�w4SVQ�G܈1,�A�z1WY�T5�d9�%92YSU�ʦSפИbQN���0���בj� �Џ�i����p:�?�%]�eK�e]��n�4DUJ��(�C)d=H�PLMC-F�A�*r�y�|X��(�.�(wSE��"�6b�d= `��J��ʎ&���+%�BsV�#�eI 0�._�0��y~WY�BY�U��� 9N�%�_\׉� 䄵�T$>P�w$I�Y��J�iJ;��yYR)��S��]�����O8A��>�ד�ka~���\`lQ`�)ЍP1�B+R��D�`6c=�2�?*��O��)���ԥ�<n���*��n���q�g;$�W	�92�@CU�%3#�u}!*�ё�H������iQ��$�<�?\�>�È�mSN�{���ZF��Q�a8���SӖyF�2��tMIa��16��%sƒ4���N�!G������z��<�w=�\�,�Bѳ�hZ)��HuM�U��5UAN�    IDAT�E�zv�v"
]D�<�'��H�A"�Җ��M�:�R.?U��N1��1�A�J0�����'K�Lϵ����7�m��%��@�����W�(G�=!��_ �����<���z$Ij�Ry,�&�n�_�X��)!��E�I�K(.D�P:�ˆ�R5v�&9� p#�q]_6�H�(A�E�7�@�+E��*��+��7�:���6~WY�4C�̔��iEU-E�o�a �{�"��<�(J����f����<וy�+]��~]PK�l�~�P��</x-z�_S��7�!� �t��SR�SJj
�0FwHI	�����1�1J���}������s���u��G,j���,��0�s*�xu|gS�ת�V���;nM�^,s�5�m�b�����|�,�c]��hD8R-�8����Y���n��Nd�f闽ve( �v�HU���.[ �[S�Sa��[o>��;��x�}�G\��a8p4iʀǾx�s�"�q��$�s���h�y�\R�O��AI1h�њp�n�_2p���Av��[Wb�f��~�o��M?��V|�ʅ��>�j�Y�hӽp�1�Ǥ�11��f���C^�Y��@��s�\K徼G/�F�o9A��۱� jT܌�TpkDxlĠ<����V4i�if�`�ns|=�J��A~�x�ߦy���p�S8SM�qշ�Zxr�յ˖QFƜb�@g�;S�E���̬���&0p���[���x��Ϥ��z2�����m���Ŕ���LL��`�~����������m��{��|p��ЅZ޽��
Z������0�T�X!���~f%g���p/����,K��ܒ�s��uW�Y����$@D�����M�\���xeOV�Ȏ��~xX��;6r7��C J1-�j\�����h�G��l!�O�����uF�^�����_�������a��5*��.�H�LOW�����3=Ehx{�EL���M���(n��8sIQx��p���W۫pm2m��-��H�Σ�K�L�WbD�A���J��r��t�O� 0�~X��p������j�� ���ŏ�,�L���y!�vw�oH[)��_���~B��J��&bgͫ]�uMzQ��5�t�[�(��|K�jY��"�\v�Ԉ��:�N�:�Ԫ&!#���}5��K�E�v�ư܈o*���9�1p�o����7�J��ppm:i�;�%�-M��l�荹6�/if*�{�F�P��	jqZ@y#�η���p��_1���oNo���8�}��Օa$}}�I�d�e�����㶟����6��a�Bݝ���e*�my��m�.�hf�<�G]���c�l�Mݨ�K��M��x�a�.�������N�|��L���]	L�1�t55���p5�r�A^��/�F(}�~����9�� �zp��=��G,��T��cy�}~�}��0�پIz=�&�)CI ̸�Ύ�ZhBG]�@D6�KPҨ`@��$nx(t���C}��E~����;t�2�u�Q+���#O�ё�l�ێ��؁�ۛ��|Ӄ��n�d��E��Ǳ�k��
u}��V���_bK)��~�Ch/6�U;��{���]�j:���a�p��1�!^	[��`������M䑾��FS�Q�Z��R��G���j���+��`i������`z*�̥���>/��rd�����J���k�4:�S��^�����C<ih=���U��S�;�X�o��-�����~Բ�������әM��r�&T����b��=ot�����[�3��˥:]Qhݨ�W���IMMM�d*�
.��n��3*%���!,�K[�疇��������T>�Y]��^�З���=���/Bs8�fE�NR�a�'��-�J��L(�^�D�J?ޝ�;d����A	����oS7}������Q��u��?v��7p�'�7�HN������BE��k :DMZo?�������O�oDз�T��"�+�!ӃN瘫������:�=�H{g����������a5���$�-@�7�^K�� �Q�G��n�:��R��`E��N#L��B�İ/%൐2�t}=��fn�6?���{}�"{�N���k��"����ֺ�Ia�[�U��NU6��&K����2�Hy��AS���}U��
�"9��Ma
��rKo^�]O�����m���i�e��%�m &����A<À��o�N�D�n��-����6�
�&����£F&�)	����O�A�
�Pn��w|/=�N���ϑ�E���{��{ա������'���3����2��sgђ�=B�ϛ�ϽQ�����S��~���}��I�B*�I?>�a��Z��a�Y����'�U`��)]*�J&���V�J�(	�E�]bbnn����gV�ˊ@�U�M�1�U0W�O	�V��/���~C<Wҽ���.��J���^�����Ó�.'1gR�q�U��%K����.��߀˿��Kϕvg6N���T׹��Sja���D�fs6�\�e]`�����
M�h���k��#i��^����}��vv�R4Q�$ҟbz���f��,��~��)���K�*��Zn���m�>+ra�]ȯ�K,���s�hYB�Ȉ%L��WbB^�-�j�GN���駦�����/���7���F\�+�P�p���j.����[�1�����{~e��Hأm���Aa43��ك��^F^.�.z %�[u�)���5UJa�W`t:}ʹ�E���[0Y�OCK�A��G�&���R��\�Q�<�=���Kxș����'��Tm�X��؄ �F����Шa4,p�,8�{YF�^/u��T�����tmQc�&lF�8�������b>ʪ���^�ҺQz���n��s���!�{]�UE�e�1�^�9f�Y��R�Ix��6.@��56t_K>��Z��jX<Y*�ϩ�5)E�*����ϐ�w�9<#�e�푇�����x����:�s��N���Ҩ�蟷:�x%Ug�>��Gǔ�ߣ��Y�?���"i]p0=�ј�erM�L��tyD�V,p�4�pP_�y�K�$8Z����7���-�� �pT�P��t�?7{�,]��(�`��(���F�Z����ڀU ҈�"#��i#""��isl��<G�+��^���l�8T]�,^���=ޡuh�pE�90�[I�Y�:�]9M�/7�m+�!�s��=N�<�~��j��v����Y����iYM���D4ӿ��7�C�*|�}8FM�}�ڒ�8ٶz���R�S59d(#5�9T0�ye|j�p�����r�$	(]��>���}c��$M2�� �xR�r!c����-�����}@����;|x��}�s	�lŏ{	l`�w�ͼj�C��s.�*M!����`<�K�W%�o��6/W�MPe��>�LN2>�6���e#6�N޽v�����@.�gc��A
�3AdMU?E�k�-���jXB�rXK�\Z�U��S�n�dt�>ޮ79��I���Y�EN����Uڅ��5��7n�r-�W��B뗡�N�'1�R�NR���/�(V�/�;PO��=��^*�tT\�)�4�׽��V�������$��uz�^E��遽e��u��N���;^ۤ�]�^��w�>\h�ԉ� �D���ʰi�`�-�fx���š�h�����_/ÿ2�UT��*��pClXW�(�4����γ��i[u���AN>�WR���������oi��|I�mR�^�F�}4ǣ)FP�[?4�&�zOm=B���������̆O�rH���T��ж����:��?/�뇻�G	�0��(��y�VA,d�/]��IW��5�Vm�t�ͤ�r#%2�r�٣|~�l^�˘�J'Â'y�6��� wh�D�͛@�ϟ���=��US���6Ԩ��GC�[�����ڼf|C"8���}f���ޠيװ���Ӡs鎣9�ޓ�}'g5�SJ��e��6S�QR\�����$=���L�j�]�K��Bij��å������ګ�!�6���B�������fɹeKt7��:���Z�
MN�b�͓|$\��҈i���|�2��h<?ڰ�����o+4W��-C��Դ�#�1�滉�͹�C�D4�.�����T��~��_c ���>��nl$ x>ؠ�8@8�(q��s=�GӾ�����5si����|$��lYn;��3]���}ގ-�<·H��t�Rq� ��"�Ns�;	7;�'6e9ˇ��`5{�Js�VQ�n�:�c3OU���p�z�Rjr*��;�)
��J*�r�?�� ZQQč,s���v��6`݂�Q��9���.���_����r���;>d��t����*瑺V)(���>!�<w
��k]������|��)O��<���:���O��wL�.��f*�DE����^2U�'1TP�Pxa�[�����ɧ鸈�^|4�n�9��5��?�^=D�8.��j���Jem�5�n���dA��އˍ�����? �{9@�x��	/�oj���ϖ0Y��>5�^y���<u��p��Z�sU��0��U����冃}es>�jx	/6�������/��=�I�Q�V�<]��:
���!~���m�\�����fj�b�\��ي�s�����|^(����!�"���K�k����K8�5{����z�1
��!�ɠ`��3� �;�q>�̉S�8�d���L`��i������k֟�&��m/x�<�¥���i:����44��b��n�fK2�4��c�7NbM� �S���	�h�ʍ;t�Ē���B+����n�W
����h�S�r�kXf��a蟀h(�kN7�U�y�^���'ߒ&�m�]d�O�0P��������gu~��uP�zfH�O���{��`>�Ɏc�`���=��if�u_��*�	$�d�7t�Σ�9-���h-�h',�N�QZ*yc/�3�lqO�x�	bTX$%��s@V���j7��Ƥ��1*��6D���:KO��ϫH��HX���d>�i���J�r:���T����Zlƚ�M<[%�瘾�t�Ӎt�S�j��!fI��wY����d:4���رi�E�A���T9�L>����9�f	6y��W� ��2z�I<�Z�3E��ɢ�0�<����Q;�PClTNoL�5j�l�o˕9̣�5�j=�~�� .���4� �c>��<h���b���乄<H�Iw#��������|��MD�ݵ�Q9���7���?YذB��P�{D��6=Z�8�a�C��Ѕ�ӧͤ�r�y��
�)q�� &B�ܫ�7�+�tX ��j�3�j*����/������'��u(|AT�g��n�)��Uz�<�|m7��f�v6��~�1�nnQ
<� #���M[���C�����D �:�.'��k�c~ƛ?��==p����i[��A�RF�7�v���j$�fO�NR!%À�e�_��[�DD�����4�R�u܄5N��ځ=)���̔�&3��b��|6��#�y���{w&ȶ7'���s: ����M�V#��������u��âV�Ť��:8���YԚЄ�����!��"��o��qTS7�@��?ة���B\�	Y�c�,�Uyقk��ZV5�S���gm��=��i�bY���n�ng�C��T.fsߝ�������	�>�n���>��\��b��)�"h�q�{�w�ׁ4#�,d��%�
�	L���������B�6��b����
e��JYÖ�%��k�7T/�����(����*.@6z�@Gk��#v�U4�����n"r��%j���u���״���tP�pxu �KE2�[����z�'�j+��Du
a�j��??��q���oxz��e�u���H6��Q�wk3��Q�$ySVR!�����*�&x���:JEQ�~co��x �
zA7*L�\�x]RX��t-�լ�yGF�������5O�𓣡#	�ƾ�S<*D�tp�Q�	��|�;�91��b��ixBx�]VGڝ7d<�9�J�J����D��T���k��ۡ�n��%��I*z��#h"�R�SV]z�E�xu5�m|�@�2YL���	�,�7Iv#kĩ�ޭ ݔ�9�`K2�"��'X��'	�$ �����leV)R��J~	 ��_q��_\�9�F�)���7�
�xd�r,��&&n�ɫ�+d�U�Ѧ"k�eғ��x��<���;�����5��
�UN�Wc:D���g�#����I�R�Y����ɑVMZ��Ú����)L��}�&;4|{���|r��f�YW��������g������k��\����LLI�����¬����,�U��I~����+c"06��XF��,���ǹ�r�}�
"9���^��ۈP���V2&�P�y9;�R��ة�̚�9?ȳW'���g/���_��P�<���� i�1@��U�T��ONq�7��_%a�z�ϳE)RF�j�:B�lE`��j+�jځ}k�3�����,��ł�9�$N�q�|4j�Mۄj�c��\q=�.1f>�p6��Z��_�} U�b��
+���uMv�Z�4��w0daM^0W�}@J�1 @�lw[�-]�[��k������_ب�K�a��m9�[������56����*-�bFw4v���@5x��O�7+���jl�'����7Ȣt]���c��kQa:5�4 ��xE��P:����������N\�̚B� ����{^
�x�+�&
 p��b��-T��+�i|K
�&Si�԰
bsL����1�pmw/]��1y��u#�����IN{�*�R����H�%]V���8�0�^�Д��Ua�c�1����&Ŷ�>ϗ8�E�|��2��d��:�� ���Uf��J����=�4��k�� ���Y}�E��tMk^�C�uL����x|���
��Z�>zS����mI$F�@~�`MQn�?AS�2�vؕ%���IZ�e����R)^&�?l5"E[$۾�v����ɿ�J�]B�2�z5�hl��aԕ� �	�l���	/�	y�(p��@�޼a9ҿ9D^��M��$�z��
V{w�Ϛ�2�����	M!�En��,x!���H����`�=��1�������M#��bŅ�Q���b���/yY^�!diA�2c_jQ�'�6��R:������RA6�T�/#�9�:�a^���B�RO[u��>6�SP����T\����l\>�@ w��\�������p���?��yFoZJd�"W���25�؞M>���8����546�Ae�����%Q'k�}�]�+��n&%����2�W�Տ�XO����j�-Я���i}"E���H�J��U<�֣���<�m�g�D�R�����W��j�Kȃhu��~��������u54�w.���/nhHY�, 3���Kڂ��bGX(ňH�D�E��%�9y�5'-[����a���xw���T�	��|]ڊЙ�dE�;U\[��(�.�]��?���Uf3�{����a˨�W�Z��ja�ɊJ$o�\�C3�D�I_��'>��!���o�zA\#���?cN�Õ�����u�,.�%�X��l��r�r+)�V�JT��ґ��<#�<��b�������b��߷i��ӯd�I��M�����~��-xAP�����mK�@�h1b���W��L}@����v3����̵ږ��&�?���鑶ӂDEO,)�+�V�ßQ����sx��7�W��ْ~��T�N�~��v��;݋ޫf�+xAyg�:�+���C�H_����\ˍ,��!���ka��V�į'����O�b0�Q*��V�%|y��]K�R>��=���۽E~���6Z�w���0__���&z8C?yC�o�v*����x��������U�N�L�U���+���&2&'�����|�&�<av	��_{��Ƌ��PNN����@*�j︭D�j*␪L�-�`��&�8{{{���W����������R��4���\H&\�(�D>�Uu/O��Ė+DM�������pDX�!
����M=��!�I=�jA'^ճ�>:.~�9^��{�1�-4�^.K�m�'��cb���0Q9w�Q|o�X�76]G(K�L��e~d�10�B����f�9�b�!:Jv[pq� F��!��B7<�d�����X(�b��'��b�(�rF)�
4��)��㣉�7j%2�J�S�\�߿yH�B^�L��kM�RsY����o�gUW�ҫ�2���߸#�,d˼)3���(c�@\���F�!^��˴�=N"�}��`� ͗��T�����0L}Օ������៾�ޚ�_��3����e56i��A�=�Ns���v�mo�f��{��<����ĉQ9�i������@2cޚ�)�@�ZU����\5 h�t�sݬ�6�cӻ_�T���d�+]��F�R��<E���[^4Ӄ�8aڮ�Q�;;���,cbU)���@+�EҼ�x�9��>��ۿ9��g��ZW�N�ռ���!���O����$�!�3:�M��:lT(�Pw�F�>�~��ο���ݫTъ���`��+d<�ĵ5���w����l˸AQ|z����^il�ջ>t���I�]:^+f�/��)΄D�Wi+����wj=��(W7�,ͻ[Ӓ8Ʃ	kfW~�y]�/�Us�o��{�%���>�Ԥ�L�]RjШ⊢����6"�@ �
�<���2t�c;��s�˻VlP$�RS����=���NP.���J'wfm��oAԋ��0޷��?6f�Eϵ���@�i[��{ݲ���ɭSNI���N����\1��q]��(����}�
1�|k�'0�d���&�X	��}7��,kٮ~�2w�L/����f��?�cߘ������`�c��9���2�N�ϊ/X��^�I��l�)G�����%��`��f��׍��1�u�S% D}4���қ}�Bq�E��9�<*�PB���v������>����-4�1Z���p��-rQt���Q, ����O�O����ؿ�͑�/pO��$Q|3ߚOi �+Pݡ����s�*���?W{��\�ț%����ǊO��RF�rF7�z���n۪We��YY�խ�\)��������}��cva u��bOSo�Uoo3�H�=�V�x	E��$������&�jf���13����{����,��VO���L��T,�LWk��r���*wy!JW��YF�b��;�ؚ�������+ז�Y���ɏs����~ŭe�s��OU��z�w�����֯-a]�*t�M����˺HA;'��Π���̃�M��/6K=c�}��;c�5�|||89�cX-vnUU4x�������S�ڤ&�ٌ��Uƙ�W��&\�b�:�£4��V���I�Q#�o}N,�%��jA�ߐД�'���,b7�N�h*+2V	��쐵TN:�֬ˈ��"LH����]�|��eNig)3��}�S,۠�����P,.n�J�!�b5%��XB�a]����*�'ņM�jAZY�����3��_A�j,ろ������1�1����MG�"�C�ȷ��B��c��!a��x��ٌi�_n�U�O544�CYG���9+o���U�;��]�^(��K�@���t�1�u�3��~�4F�X\l�5un����׮ȼ��+"<]j"�gf29wц�H�t	���Mu�"���,���\5<��H��݃!�+Md �0<�{N�l�4��m�t���[,]@���uE�C����Hu_��Q���Ï*w�F��R9����W��ƞ������wKS�?�^t4Yչ>��.��5��9�.��z�
����K�p�"� S����4����2��1��Xt�"y$O]����#�c�K�>}�e0@{Z�-��gJ������Nfu�Qʅ�����]/��\9<��m�ǉCc�*T֬'��i���2O!&�?q�)&��z�f��8)`Э�9t�b�_wF�:d���d�<�!�6�� �=p�j,�e!R��v�&�l���l���1�w��3Wo��k	+\�U��(�	p���s*�7?~�;7����`�� D��������@��n��Pb�{�<����f�3����5�/�u��7�ty'�U���G��-ł�D�<��<�QC�B>dU��E:`2�%ޠ2=;���yȞn} �=;�P�Z�>��@x�Q�[w��t��,�J
���@�=_|�׺����kl����7Ղ9�D�֧WT(��UTYa�ŜM8�R�����]�����G��57�'�n�M�V��򨉪*-j2(� BNM$8'I�C��hK6�(G�BǤ;�lޘ�"��t"��ւ��T�aUL�D峈��;�~Ef�<��}:�+L#9��������%��2�G��hЎf�Gw1s;}�i�p��2�/+��z�(����]g|�� U'_�"�v� '����������B���1�����ƃiz�	0\����,k���w�&�;҅�e����n��(iA�~ʫLM��E�pw�
uJJ����a��y�</�)���E�6� ������ۦ�$䪁��ȟY�򍭎;��l���	�Fw���M���e��3￥*��}(�L/�������1��������O\�k&&��c�QPoѶ	�4V�W{�Z�8W�{N����̎���CH&� �|_O���v{�L�����c��:�w���	�D;��Ֆ�36Ζ��Q�N��l.���%�7������ۈ��3��8�����-m�çO�r�j�bl"A&�%��J�M��<IK�'�7P��D�KCp���@��t	�$)Q3'ׁs��e��͕��*��:(M�l&�7�"Ν�06u�խj�_�A:,-*"�����6����/���Τ��w���������%��+�
�\�Y�$nc�����ޗ~~tB�P2)�R��TY�����N��Ĝ�3�Ɋ"j�K��d�v83��u����b�F����dzc��M~���7U�\�'s}��]��4,�3&tA^"Ť�=E�_Fo�����d��>�r%�wS��p�l�.ʷ�T�h����!;go3_��Pnǲ�D�X'Y]�Ş�'26Z-<�FD��{�x@������)�<m���Q�V4�9)]3r�wŪNw?n���w�ǊhÙMh�jg����/��Ou��B�������E[[i#���E���^�q`=~����-�;��rbiI��[�K�Wy�a\��CZ�BZj��k����y�����'����U�j�0����#L���=��E�eD� ��r���4���݈�d��`�B]�E��s����M��������!�d"N==�Bm�4g��Բi� �Q�]wc�����a;���U�9g��6A�s�R?|o��q'��g*6t����� ���x�^p�ҿts-�����n���q�b�B����~5	j�{;A�3�^q\�R�������ҏ��e����;�z7��m"���
��Uwu1�M�m�����??5ܽ�s	����� �^���%"{\T�k������K:N��kN����^ɿ;}7�g�t�
��NWlh����
����]�}��2��N���}��n$�[���z�����{jd��F�e���O�ӟo����l��� ��SO�^� <_�$�e�W����)���&���h�ɹ�oN*]s��,�e�uMθ-UG��@k[JZ�!��r�a�K���?���%� ;o�\�@�0-M?77��^���I��CDoƄ?�}d��|�x:F1�����sPf�m�v�L�W�ȓ��D#J�>����8���D���q*�ʂ���p*+��c�J�r|���1��>���W9�8L?�H�؞����^�St��M�~��
�u&9s�I$�y�G��X�	n%W�� ��N��Ɔ�?m��̌$ =��&]Z}:����o���4�@	^u�����+H�WG�ظ,e����!KB��FR��㑑Fb����0��U+� S���{ޭ��$�>9��t��G����|����63�s�$`��	Q8e���ػF}�k��aw(��F�YB�����ҿ�|��[������&�/T�vg%�S��
\�Lv?���^��:0��t�q�7.�Jf #];���-6¯(��ǯ���V}-�|^8��!���cP�E[�!l"��0�3��MLDp~N:&:�q���+\ ��r����c���텅��C4��
kZ]^��k�>�����Դ�V{�u!�aR��q�E����!��=!j�M���ے��Z����<�W;��b(�
33�I<�i�m�݅O�n�d����.�C��+�BV7*��/����F;y]ԊVR]�A]�d/?�_/8{ѝ����~W���(B%��~D{A��6@C���dN}��!���C�f�m*��Q�k�C���o	ݯE�A��r�\��}�VC�@�<�D����]E"hI�(	pR�kh�C6E<�2#?���ܐ�x0�_���
ڻ��jf<�	��ڊ��N�u�P$�l+JQN�Js�c4��� ��0�ǶzBH����x99��}���i	��#_��w_Rb<?�+���_���i�pr�:;�D?��:C �5/o�:�%΃���<�H!��x͆O���as���C�9�O�N���^JÖ5���vN �3|ꀜQ���l�p���:qr�w�BO�b���kf�Z��Z ���(�: ��X�.��ZIHw���y���"#W|�e�B^w@ɓ�yk�t��DK�T�Ik#6��z����s�W���OL�*��)I�z^7�>�~p_f����t=���LV���A?W~�gV#堎��Vkw(����mq����Io�8>��_nx�r�3�Eh��.
�ښ[m&l�}F��r���^���u/�������ƛ���GM6$GBJ,Cc,ώ�Bg�tţQ��FuZ`{N�-��unKQ)���M��+�������|Ce�����J9�)Z�Ş��L	���vc#���m��ɥ�LO�]|O�b�2У���D�ʒ���%#B5"b�+���Nݛ������Ҫ��+�$]l��5[�¡�Tٖ��,rxm�������3j�/�/	F�b�b*1�@�J�]F]��D��]N��doT���@��T(��ǔt��{�O���m���)��U����ݒ e���N����$��9I��`vh#�b7��0�QU����ڽ�A]<Iw%]�0f�; ��(h�W�~
�PK   F�X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   '��X�l=�o  �o  /   images/2c21fad4-931a-4469-89eb-1a483abbb87a.png @鿉PNG

   IHDR   �   �   ��o�   	pHYs  �  ��+  ohIDATx���e�u��>���^O�n�1� � i��VDɢLSN,F�+�TJ�@R��/��|H�JR�S*9��R�.�lI�̐�$�i�bc$Sݯ�7w��{gM��� �F��}}߽g�{�~뷆ûǻ���@�{9��w�#ǻ��q�xW �=��
ĻǑ��W���v�L:)���5`'Ʊ�Y�P�C�t u_3�C2XM�y,�����J���K�j��zY�������������h9ϲ�wE:��|�E�@��46�c�s�I�>ߩ�[;��������mԇ)�&�v:��62���ߢ�o�@��g[��lu�y{��K���{G�޽�x�b\�4u����`0X(�Iӗ.��E����~����:ơd�Iڜ4���A���j�w�zk?+�aZK��_�}�߮ۨyج���w�1~��k��7�7�;W���p��s_?=�>P�����=��>>�,���j	WNjy�%e�����ޑJ�zl8��7��¨���D�Ag&J2��I�ԇsK˛�[�_�^�7澳t��u��o���9��~�K��}mak�`��g��\2��Hg�Ƈ�7n�����l� ��"_�
py��� ��C��F�'�~�ѐ���@�&��@�i<��ȃm����8(c�l���/�7;����W��p���O/,���~�����,�����1:~��s�+���k��ăׯ~fp��Xo��ɚu��4i5��V|���X
?��f�R&��A	P��;"n�8�@B�J����3�`�L�����B�J�>���,�����v1Ɏ��u��_�da�ͅ�c�?s��]��߸�v���i���G�������`��������������Q�}������JZF�) �8�9NT>�	� B)HP@ꆴ�c!p���x[�, ?��@��w�ma>��dBȚ���T�#�QBVN`ܛ��):"�\��?�ˉ;>,�g���n\z�k�������v���q��_�7�?���#-�oo������|����˿8����Z�=���"
.�!�I�C	1N`���8�8a����\��p���<��GsC?_�}�(B��C���Y	�+�\(A�@A�,^������1r���(�v#�Ql�Q>X�\[{׍Q�'v����v���W�~���������?��/\H��<����u�֕W~;?���׊�Z�f��!�2��ĉAP�R\�1�bP[��~|?�QHX
�5M�ŕOf����'r�h�ٰ���:�@j�8 ��p�c��@&���E��Ƴ��x�?;As����`|�x�9>��u������_����y�~����|~��9���ܟ,���_9{�?�y�՟i���u���MVk�Ԋ��f�(P;P�Kq�"\՞x%�o�8�{T�dO���w%�ZPIf��O��wQ�b2	�D|�?
[���н�5HF1JF�C3è��!��K��|��;�{�ڇv�_���{�r�k��Bzϙ���~�� 2长�;����������w�?r,v'����'�U(��j'�����]��/�#՟���L�f ���4�HPn AplY�ӈh��T� ��jt>�1��'�!>�A@�X��*���8�;�k�OT7��ؗfg�D�7x$�������~�����+��oF~$b�ٯ��������w�~s����=sv�O�f.D�R���6�
�)`�G�t.� W6
�>�����u,4,/�	��$���U(�4�Z�,3F4�`��!�B��P�#��$�9(�c�b���o���0�i��w�.��97�wܿ������]��S�*��t��������k���ƫ�~��y��I޽;��f:M�эL�<X��p�=�v^�1<O$c@�k|�HC��r4������ �Jp�i� -�HPJ�4H�"��H����;~�=Z=�g��
dQ�i��CLdh� �,�7l'��l�=����w�'����o��啿�.���@��o�?����g���`���A��-?:�H\�@��o�vHȃ�+�"MD�-N��4���!ZhB�aK^� ��)7$��\����5��V���mT ��2�t�?l��7��)ٴ9h��EL(�oY
Q�$�õQw��z'��o�g���/_��?�����G��>~(A��?��w�x�O��������>�A�ȼU#�1V��� ��30A�{�0�(,�:�K��sī�>C.�a�!K7�i����3\M�g*��D �4ť��T���&V�Y!�4B~�P:�9�'�͞�C4�)H��>5t��z�ܴ����a�=t��T���/��w��{~��\ <>��������������U�m��R����h_�T�$F����o06�c[	�ER��'qj&<���٦h7�#Z�p�*ܙ��y��Z�EX�Wb<����Lx!��_�����$�4�{ɋ	kK����_���L��n�8y���č�^v~��?�����_�\�A�Y?P��_�R������������_XL��I�r���Z5R�9�sr-c���+60ӕ�4�nH*>��MHe�(\���HA��	�z���>�Q9���@�g#/.��D[XoU(���J�y�.H�%FH2r��'mS"��g����S�4�xn����}`o=o��|�3|ߟ��n��w<�&�������|��X�]���w_�ߖ�_ƃ��`�T��B�Ѿ��,�sO���	g�R��55	�l�i��p �� E��A|�6鰬a�^�e��U�O�{�yf5#V���(��y#�F9������p��At���:7����^��k���y���Bq���@x�E���pߵ�����~�����f&}Hh�P ��1E�r��0�Z����"}QAyZ��d/De;��,Hhn�H�h�\z���a�R��5��@�k0�� ���E�y
�2�����DtqqT�W^l�@`&�NS��(�дu�qE�莺�ﭿ�+��i^���/]z���g��\�@⥯�ή_�֧:7.���'Fg��\�-,s1��X��a��@pdJ��8�P!��<T O�cD��@���,�8�&G���3��.ʵزx��53n����3��Q�H��&>�}��q	yO�0�h&�J��	JH?��k�F��׽��y���ƿ��^~�q�q�x���S�>��g:7/�WM;~tn.n���Ř�o��� ���<F&�'8^�4	֪�&A�6�}�����Z��C��d�8�$+��J�D�hbE���Do<c)�����&݁ރ^Ո)�w�a�H��wJ�&���L�4Q��@0���<�۾򟏲|����72�މ�zG�ҟ���K���ý��ER�m�E��sW4�ʍ$V�G&�H�ѻ^V�lU��~��>�U�A�葜�!@���*��̩�+!��4�\�^Ka���� �r=�=�����&�p�0�Ť%�^���MQ��%�#�Y�	�)j�J��@�ժw��Y�=w���_��?}������=g�@\�_Z~�[������:��[��\T�p<������T����I� �����N4P���P�Q�8Ti�Kj��x��?�8[ݥQ2�T�:| �r u%)�W��fI��ގ�X�%%S�F�t9� ΋�`lB�:!�����'��B2
���Α�I���޿ws��/?�s�ۿ���a�wD ��_m=���<�۹�+ロ�\o���@VC�"��>���~�x�
q5��`:�C>Xk�O�[�\k��)0�$� �2B�Pc�`Wi��@H�,x%��W��b�Yy��
�r�[$,`��P7�3�Ƙ"\�E�&+��&mA	`�4�q��F�(���f���k5n����_zf�m���A�˗���ܵs��?����Mk����s�`B���2I�3��ޙn�,�@H�N@�C��)��Va-���
�zj���{S�������Bt9�JD���ɣ����=�)E�+5�BH%�TxŤq�+q�!�H+7BW�Ok@��Z��r���ĕWL�L������S�}�mI�}�b�/���[W�����k?W�)��L$Z I�ɐ�B�F��$���0J4) �l������ ��xPK� ���5��� ��d�{S�R&�k��X���T�pdU<�NEehDT��S^��"v�5	Eb�M.$�+X)�uS���ǰ�j������y'R�N僝����=�o���x�혿�U �����ן���]��Z�wO
��]��&Jgs�c/�4�u)�p����w@�Q��`>�EUˁ&� ����Q��>j�
��OxrhB�ac3��J�: �V�BPI���<�d��aY��D:��B��[�6W�8a��0�o4,��"�Pfh2�8)���
���A޻ˏw>}�����u���p�N��m��_��'�n���>P��vT��N�d�D "�N�������SP�[�Ahh�(38�Q�H"rh2��4a哙p�0:3G0�	^G�8�����K�'N�r�U�9��3`5&������hjPm�=���1H��s�O"�)=R��<�G���@?S�2������?�}y���7����O�7�;�ǷM �����ׯ|�����f9\�i�?�	NY�Ǽ�9�@W'3�ڍ"��[�`X���K~�Wn �M<����T�
VC�!�9J�V��t��L)�^SpDdM�r��A ��R�P��3��X]#_	�
���TlN^r�g���� ��|�I�xN�2��:esdp�(-���߸��ڧ���_��@��"{�<��_��`���MN���MD;!,S��\$?Ҥ/@2R��wM5�A���a嚐� �b4B�K+�{s�)��Ձ���rt-N-�����`ˀ�z'r�,��C�.3su��׸
k(dUN*@˹����܇��M�S0n$чr-J	��bm�=���˗�{�k9ķ޲�x[���U��������z���P�NB�vrL[;e�(4���#�MC9,���
� R��A���z��u�[ate[���-Ѐ�%��-h�
vJ03x�s�X���3���7�q�{���}�wWV5�,/Dh��ը1�ڒ,�P�F��j)�>��Z=�ə��+�KZk���������[ʸ�c�8|�O�.>���'�<f��ˑB-)�n�h&J,�3DT����(
�[�$����a)�I<;��P��8��/	��R��ʌH��'���"�7�a�� ���ԺXy�ª�|.9'�_(�55[Jh�@�����K����H��
j�1 ��磻@�ڍ�q���[�o�`�*~�/�9���?9������~r:�<���:eHSb�e~@0B�v������Z���:�'T�eY%ŊMU�Pg��m��b��*Xt!h�������"{#�Th*��(�����jT0�	q	N�)#5A��d(�e͑Ƚ���,��g-0)A�k-��� War	�xvO�a�{t���w~rs��_�B�^|u�w$������x��}�#m?^j&��T��&�
��V�]"���*�|!��**)19|p���+�M�/\��252��8��L�/����:n�� }O�9�e8P\#��E!(F�D�� ��QŦ�+cU֖R+���f�;���\8�*�KA���ʘ���Q-���ߺ��ݍ͋���@P�˫�~�`��g[�8�c�D̐�����q�X�>�t^]D�J�/R� /}�k0�����s3���((e4�C7�[�,7��.�t���ߓg7�t"�	�'��(
�Ẍ(�{-�Ҏ��ߋc� T�c")U`Ƹ
(3EIf�e�1��b�5�$�ߨ�Y�!(G.*>��Ҭ-��r���(����
4��r�������=��čŻ?y[B��5��������ýǬ,&�"JL�*�r"4����V�����,PL���(Z_���]%�~I/�@�s!BBd� ��*����,$�&=6���D���}�{@a6���F#�2ϙx�*��B��@�$Ϛr��"��c@��$�`�����(��$��Kݑ�EP�`D�\��
>Ӑ��$��I14y��`w��֟���oY &�`y���������1g>٪���D&�̖!T���H�%Jv���K��I�(���d��>R	`Q����vV2���c���d"�R�QhD��/�n��2S"�s'ʂ�'��4gD�Su�y�VqR���xҼ� gj���*� �!��a���nv���𳀊�D��e�L�k25��A�QU�4�VO���'��Aw��7���/?�e�}���H}g��S����/���T�K��";Lif^Q:?�<7���,��D��!@PR��[�ohղ'��#g�%)?K���X�ۜ��6��<�ް 8��������Pl���Q�\&��e3���
Y;͠*����ޏM��qkz�V�0�#u�:�)��څ�$����`�A�!�KD{ʹx��8���N	�	;O!�����a�wV  �o�����Y܅��M;�N�A�tTf_���q�Z�f
�4DL"�ҶrhX߯�R���$��8�1OFI�����y��d�E�����j�G+pyM�'�ǂ��!��՜�Uo*y�	��L�# �ؠ��z!j*Bf$j@a���r,�
+�Q�1�(:H�j�*�ʴ�K��#�`8�tJ�!LA�*MSNF��0� c����c���`��{7/h�{�.�������9�('K;7�~8��Ϸ"��='�r�+ 	H(�<:�AN���3���Q�O	��s��u<OX����V��؅)c��@��Im8hP�pӨ��n���Q��/��s&��:�����om���.M��a*��' v}R�$-�k�"�@��Q	��NUᑸ�$ Fc�(,��/��B"F�W�Ad"�:�JV�2x�l�&����cQ��U9��������O��K��wF �\o^\��ݻ�a�7D�##�>�lg)a���Ϙ+��k�+����0�b�p���L�;@;9��0M�Y��4������W�s��P��=*���$�a������}���rh�X^���B�)
H5ޘ�$wA��]^�Q�iR��0�,�����8Wǉ�K�Дs�
22��D*���G��ܘ`���y�|�e��֋�о&��Knm �i��C���9���d0�����n[ ������|��X�V���2�ĉ!�2�`�oJK��F����F���)��E��3jo����y�y�#�=x��&\�~=�T�(pb��{V��3�������Qh|2T��I}����}X�r�����#��U�D4v|������C���]k��6�&��
kcJ�i�*�Q�l�y^�r /]�
�{��E�G�[���]�t��n,�1����@��j�E�L,ǿ�{H4�Gf5s;���R�L�=�$�� �"LRǓ�Ҩ��u����4�^6'>�Z�b��\��~��h�� ��t�P�zZRy�R��5r�^#�I乌(ND� ʧ�g)����l�Zn�v���C�.\܄��]��K� �6N����9�.��f"�2*k0vM��N�;�߀��v�e��ӆD�;�!7z��[p�����j���ZL�u���GA���0g�� +ᕝ>�_߅K78D/�u��0�8N)�uʄ��F�93�LfQ�	�>�����լ���2���1K�����.�'�ȋP�tvT�v-�����[��ݿ�,܂ٸ-����7/~s��9�&M.����j]�O���%AQ.1_o�h (aC�3�7#�$���{���P��K�\�օ펇K7P� #'y�1�����W�"��
i�QC�0d��k����:$Hx;���N��Ѥ������@9hE|+'���a�Z�騁�C�Ʊ�z	�&�ҵ��݅�.~�u�2�@Z4o�q
{7NL���NX)�h4�N�g���P:��ϬWR-<��NjD��R���8S��(YfK�p�X9�|�V����?�k;��dyo%�c��	W[qޒ�{���H^��@���I0e�$iF�e։���	���^5�6�|i{#�]<��E���M2M@,�
�Z�0C�07v���+peX[-����}��>�1���9�p��%CK�xyVW�P_�!borc��+�k�t��%ַHP�ь��0�%�ߠ�Q�X#��,vť�ʼ�`��\����p��h
��U4�
����t�7=��r�+Z�hxn��.P���
|nK ��택���`1�Q���'�H���K�@GF�=�a��gS���.@q��WW�X??�F�&�Ga��	��-h%�zt:�l��%j���],p����3�8�P�,H-��O�=��g�9����vqb��v�������	,�5�QO�b;6)<�����:~�K����焞�zi����Z�����{�U�){$Nb!a�E(}�cxu�����˰�*5�!Y�ڃ"&�DjSrb���F�����Ω���|?��U�,�"w��'�PC�KL�Lm�Ax &��e�	��Y�b�IH&5�N<*�\�RJ7��hkB�.C���Z��3�d��}�=��%�D�E,�Z�ڦ�簏��?|�2�����"zx�l⎝����<�����  � ��<xf� j��C,A=���Ao/#�|����j-F��	
n�o��Ed���"�sҽN"���șN�j�H=�|:����ZQ���5�+�#���@�@�4,�n��{��6���Qs�N�bt��	�e%�f�p�9$��ͅ����5K)t�5��,��W�߈t��S�8m����D�����A�8���:>0�B8IF����ǷSN]����z�Q� ���sm�&����^[J��$	�-�G�BK������$ps{^��;4W��.�!6A7x���/����QyF�H\K��]�҇p6�h��Ho#�1�L�.�f�(i%��s9�� M��O���F�Hc�Ǒ��g�Q3t��Ǔ��M�-Ġ�7�~�ASc� �(}-��8F"6��JI�g�g��6F����� 63J�r�-��;��=����Zg��^�Fn�'��7�y�T3Ը+-1��S
�9P�"�$���넌h�Jn�JXL��8z�������-B�Q>ɠ��C�6���p��o൛�.ބ�;�8)8q�YD���jwp��%^�B]�fN�gb**%��"m' �]ªZ'Q���rg��t@�m�8cad7ɭMB��rZk^b6��5����^�m���~�w�|�29����� �U��M	$�	�/UՉ�(م����$5�"Y	��	"N�!��00_�!G�P�N�}�U9�Z`��E�G��ג:��	N&���j���W��%Z
�P��倘�tx%|�5Lӂ @��b<���tm��-�u�a�ۃ��l���fy��x���!x4h:&����a3��e�J�z4��Ϣ�G����;���3F����&������%D����9u���Q�en��IŌFd����]�nY ��Ak��-'�z�f��^�gL�R\!�c���ǣ��p2,��� J"��\�*Z�.����yj:�8O�
~���p2'�&}.��F&��&�s�4rj30�+�Cg���_pN�,�\���9	��!4�桎>|�pwh��hJ�+Lz�F��+$�z�&l��jq��������yɅ�5T3I�".p��qe�:�CuŘ�&(�4�c
̅���U��� \C����i��g�U�DR	�ۺ�E]Is'$-������͕�I�ם��x�v��?n�|r,Ƨ�U�%��"����]�b8"�ڱ�m����d�N8��k~(5J��ߥ~�Y��#���d�j��(�2��z+1wl��B�Q$�i�\	��v��h�j�Ȩj�� tzyϿ�|��+pu�Z�	w?x��i8q�$���Z�,���^V�:!X"���&m.���գ:J����-�6�Sʞ5g)�3�hi�5�V�:Vp�a��.��1�hn4�;n���ߗ��5���*g����\L) &�PwL��3.k������Z��8x�7e�����ϗj��;�h����La�W���P�7a���)Q���*ɢ���3c��FW��9ne�BB�YZÕ���k��q�LH&2�̱�z�����`���:��O�����6�l�`���t�p�:��n��h>�S�8���DLB�/�	r�H��$�c�j�k�Rp�G��ǡn5N�ډ&��Ĵ߆c�/a	7���`0zC`yk1I�<G��Ez ՚NM���r�Stӹ�n^���=��	�9ǀ}l�0�,Ꙩ'�g�#�J�盐 X�)���2j'QCs� ��D�̽�r���?G����U�:?ø��J��6q+q��`�MB��iϰ0F������أ�l��B�{�נ�/����[{@�W��0�\��M��	�1J�Z�b��Uò��n��'�!QO�u(���ېt�ʫ+5��AgO����w�D>L�lp�qC.`B��)�#:�r~�eH|@�y�K�Ω���UK�jM?M��Zr��f�a9���I0J��z�LD)k��̌c	���V+hj3<�('YnB�����C_J,W�ՠ^kr�e�ۇl�C�����	��.~&�L�Π�_0�c�cs����[�=���u�rV�q}&���M_d�.��^��B#��Sa����j��2ѩ&e-�bei���kn}�ˬ�ar�1�w�l2^C뛲zR�E+�-<�FLp��!�DB���͉- C��(�c�6X{	�F�%p<��\)%�s�Ω�ԋ!����;RJ�+Ku�b�|f�Ǡ��9�ۡA���GS���\�3�X	��|V�Z��`����k	�wQ�I�$!mE��F����!~���ML���a�r�T�҅�p-]����M�Q�R4D}��bz�=�H\~-���#��B��П3�n|�s~K1)FQ���,A?�eetx�)�ҋ�rh��8��f�?]
��@N����� �˿�]5,ζJ��1"t�@"*ỹOA�#���
���ڕ��X]AO�6;����~g�!G���`�p��qHhH�,/�C5��p�y�gW���@�Q���q�E�ZB�	�-�@-��ŵcvх�;D�&����b�lR+�q)��hc2i�4�4��h����ԥr�]�^�0�$�;���R��Qw\�c�Ȇ��Y'*��;�L�w ఐ�0�~6�l�@k����)����8cH�3�l�\W��0�l�C����jx������dʁ�h�(���	-5�pb�	-2����6wa�F�W�����vz�=�9�3'[pr��BևF��{�� .N��[0#�.)��E5Gl���k�a����
�<x�nx���p�x�N�`�j���ǖ&k�i��c���4s4�����1���I��h
�A	M��1��,
T�>�Gu*�0��3��6�{��7)S�����K\���R�IY;T�@��,�:��|$���!E�����Hʄ�0���~
���Ŕr�>}�E� ���(%M-�����F�Q�Π���C��싇�	������`4i�`P��k>}��J��[���	��!��>5.`�:�Q��P ".J�K(`1�r	`g'��B�q�n���<��I8��A��B��B	�)E�M�ێ�r�fV��k����!�������ZM�g^��m���u�J<rҺ�D�M�62����q��ز�e������:5-����Y��b�v�������3�^�Ĵ`5T�e�G��H�/-��-�����!��m��@��6WI��)_+�XQAZew-/�{<t+/ma�������r�v(Sp5<|O8;+�8��	~R:���`�"	�7��;��4�!,�rXk	��kP��8=N����3�8��#�>R -QM�N�w�;#0�bP�jQZ+i����LM8aZ����֘���go8����$�)q�\�$��.�t-��ʽ�<M��vZ�#�\�?yv�
�"�lzI<��XU���T1��9�1�����9�p�ʒ�1"��qu��j�y���5nX7nB|�#`t��ġfX8�f��O�C�V����(��0�%�8�`���R�����:��Y�r�ڱ0��q���=�{��t}�Uo��P@�>�D�9�F3�JN����8L3g������3ǫĚA���E0+LY|O�p{�1P�P	͂`^�N]H�$I�ɔ�Bm�	�6����	h��e��-��������=�0��
�(-�t��p�=sh�	`YE=��&T]��j|	���	8yj�z�����tܿ����+X��li\�E�S�9G�0I���j==]��Z+ލv��w��?�S��5S���b}��c��$���h�W����RU&��c����3�*��'��5{=o��������sR8<�rI�p+�7I��z"�%��+�����e���nfV��>R:�h<��l��O��.��h|�l�Oxd͏-�`e��zj�ܚ@�:ݹ!��u"иe���T��d��:,4;�9����6($���Q�Ӟ�q�'q)3�=�B�PCR�4�1�*j訞���qBXb�.f�5ZL���dU�&3*��j�&�xo*���La�|�y�}:��"�@ �3���"w�{YȨ�(p9Lz߷�̭�`���7�Rx���hjv.B�(�&'9�c�V��b�A���a_ˉ���/4� ݉��L �I�	�T
3�:҂��1P-GMj^B���6\�$ȩ��G����EA�!�q�5B�b��PȡNI�(LT�I{{%	!?���	�͗� ײ�S�m��L��yr�8�������P2�;v��d�c��hi'�:��=��ی�Ly�]�;�l\Ȯ� Y~�V�s�;�k:�7�#���[�4���c��8�� W��`��� Ց�����j՜��T�rG������,�6���	�7il��s���w&��)"����ZqQ-�d�!N^F� �"�8q-J�"&�\,���.<�%�h.G��RIN%{��g��&���l^j�</��b.�4L XUQr)�]N���}9��u�W-�	���(�0.1��y���sS#�ϨV$�z?�5�w�6e�#�G��W��&��w�!��n���7C��l���u+�H�s)Ŝ6du���V̅�1���:�9P��:5�D5=��λ���
�,\��X 3�j\�D����Z@��ߗnp��w�&���&���L���C��-�I<A�"ۂ�M��̈́'��Q���r>A��������UTYy[Dh�q��\M�tO0)�
��W%q��@)��+�-�s�E>I���N���h�oI �z=���>JE9)hUQ�H�I�Q��p,�^��o���6��lz��a�Z�KI,��@�!��#��@UȜ=�?��6pTCapr���-��PJ:y��+�K�de�Wpy?�T7�p�
nWD2Č(n�aW?�4DS���҄�%k���
8/{�G��؃�)' +n��ku�l!)1禠<,���TXպ�9@�Ƨ��h��J	��[�=Sezd�4N�IT߱@�$�MuM��F�N�o8V�#Uk\�̾�[RB�[7�2UR�m�@t��$��������)�6]���	�
+�Ɠ�&�SP>e;!��zh��8.��e1����Ij!r���6V#���܄>G��t��aPP�%��KE�B�i���ƶ�3����=39d�/�6Le	 �P�R<m_�}�h�+���
�������Sَ��7�|�b��Pv��a��I��j�m|)>�����V;��eYE��p��k�J���xb����N2��Oe�9x�j�"J�R���J�M$��D��x�&^:��4j
�F��s��*i���q�+����0� ��=1C\�h�d"��d4yM��Y<b�锽MMT9��kn�~b��^z`��0g;Q�<WpA�P5%�Z�)y���p�
\rx���(��
/LI��*�(A������n�tK���y�ټ1��$�["�M�E7�>M����l&���qJ�p��*)F��iI�X	�R �C��Q����C�f�\d m��8���&�X�|C�3�4E�D��Ny��	?�q�I����2�k1�✪��9F1�H�S	^�"e~8eV�JL�F]t4���}�ԽgOF+m Tf�1�TZe��?�LLd��� �����G��$�q2�՛����L�i\��7a�G?�����4JVE�`Wqf �Y�sl�&�7RW�TmJ�CJ�S:��W7�Rsf�p`���1���Z�<���h�]�j�.M?��=jc��+4�)���&"㈠�4�Ȱ���r�&�r0b���KAN)��!(�I�:��s���X�c���͙ng��U(x�]��eO��T"D�RҐ
�UO�U���� '��b���������M�b-����]EC�ۧ��H&�&� ���!�w���4�P{&�*'�Ą����n�*>U;#�r}�o`L<@-⠚��(,����ĳ��e}U�,����	���Z[�f+��`{{�\IM�����V:�v4�g�S�)��Q��\�AЄ��k�58}r֖[��e���xX�/Ey���D�2�W"���(��UZ� ��� S2�	S^J'^"��zmgniyǜz�mn-c�d;K��Ei��L	�H�n�D��F���De���ꮲ*,�-T*�`�+���Y8��ps�
h�O��=�2�T&	2�M�/��x�S�|.x��6O��ɨ�wc��]�^�ft���ɤ�Ę�����r�������@����7��5�ZBO�'�V���������d"㴳�\���|�F@��h'��P-*�Ҟ^&��Zc�9�����o��0�*6����=���gDe�E�X��L��ܰ�k�����tx�&a�xL-�8�w�M8q��X�P�O���}�fZ�q2bm>*.��~�a#�$LQfR�E������ۭ,,��E)!ހ&���R+�d�.��Rs�l��5>a+ך�G�&�h���. 0os��<�����q��W���Y��ЧR]Y����o�Vy��*�H!�d�kz%���`j��ּ�n�ߐ��e�`�h�����~w��$A7��%�f�d%�l����Z5ƭ=T*�M7^c�^j��}�[���\ZI�f��C	�S@���`:;)T�j{���h"���S��{X�K�����[�\����`a�P�}�\�\�v������'U���[C5�jP�����F�C�	 c )[J9i]�6V�Iv���1�)�GR&Jysꂂ��0�-�������r�%QԚ����~\�¶���+iտ�W�!�Γ�L��K�1���������75��cT��jQc�D*����R�6ϡ��S�B��C(�G�z ���X�l���A�}��-t��I0�Iכ�vv�Օjx2��7���~���R2F�x���МY�o�{��5��U\�F-+�O�Y�v*Ci#j�Q��v}aec��}"M�'��֋6���̯H��Z4U�3Z�7L	�j�c醄r���wU�=��j��?S���H���s.�
�P�2��a���]�l��"�ln�C0B�i�aSXX7��B�S�>G$j=`'c4|��Ӊ���v��M��)�	Fau�@��87�`^���ԫ7����G/�) �x����F�z���o�������b1ݠ9w�&���t�P��P�q
�9T�T���(/�������v�����V�-j�C�qF:�}͝،�iEǅ���aS��l���t)��6�1��>W�}6�VfG� �p ^�O��@��7�5�V��/_�I���dB)�"��e���r� ��&�� �����@s�E�U��`>�^���Lu�E����W�s+��s߭���c���~\ol��d��ibeRi�*QL�6���H3o�B�N����Q���j�2�t�*�\�����c�+�ne+&���L#�2(f��|%�n"+�4�� UD π�h ���!v4����Kԉ�YNc(*a�K��z������Rv��R]g��Ʃ"��B�8"j^�(�M�B3��n7c��v{w~q������ۖ���~��j��.N?��b��]�@�� |പK�*�`���U�����B�g��k���hr?� L�0�"�N��R�ILMC��^u�ftU��	�0�U��{+��A$i����4^��;#���<k̙b��j��h�$oX��T��,�i�$w���9�3��Q���5M[��k38�f�I>��v���|�oi���j)Ԩ�����7�z��x����fn\ԨX� �<�u�+�}"��[I�!5kU�H��$�څH�ӕ�1�K�A�"�P���2<UA(c� ~Ai8�ӊk$���v�W�$��@<��8:W	6�ZZa����^��9;���"�!̀`v�x_�����8",^�Ċb�%׹�t��LG�t��/4w�_��	�Amnᚩ5��q�Ӵ��U���&J�^�ts��:F]"b�A&LZ��v�	W����U�h�$����r��0���<��v�7��������,)w���H8���D��T��}8������"b�Z���ם��*T��D6~	�DG �U\È�
G0!<ƹ�9H�8u鍸��v���-��oyw���د�[��B��H��|�_�(c���0�+��L,��U�4/�S^t�u���8�u�4�֩�tAv4����t%�i*��?<p��<B�P6ȄD0[��G3���-L�G�TS��E(�+��@�󈙜I�j�%#�u�w�����B�p��Ƌ�B��hv�819�*y7�8G��?�����;#<�sk���ڋ�q��mҬلwH���2Ѓh���m�J��H��Ia+U(6P*���o�%kz\��rņ��V�;��0���R�>(� [,T�j��R�*�2��Z��vv���v��n�(��!0�b�"͚�j��ddf��b��{ҹ`�&L����|�����ʉ�҅�����a�s��m�Xk���g�������5�\��x;��9	F��(a����V���
������̪t��\�7;����P�@TV瓙��cF^�NJ�-���iE����LkH@�����y���MRH�Հ��σ@p
���<b萍���]p�$��aE�"`�CEK.��O&&m�v�=|��v������k�G?������Q�J�� �7 ���x���f�>�E��e 
�,����a a7�{s
E-�a~f`+���+�܏�6����&�>qzٻcF8�>�pD�W�۫���nD�S�"��*��Y��;s��upJ�!��a�<WoR�8�0���������{ٜz�6�K�#��s�6�{9�w>V3q��R���h
˭sf�]��2� 44%	'o!b��;�w�j���δm���z����	�Tw�T ���,^��Rل#��M�ċ���U�^.//gr0�΀Q��@���b�0f�}�"hX�{md�!���]�(�l}~��v�/�w�ؽݹ}KѨ�u���tv~.��V2�;�c	�<�R���2��I�q�x�) U���|�Y>���`U󵂐��
��MV��qĮ�,�&4�A��9���Jk�訩���� �����8*�D�gjNF��c�$�ߨ������sͱO��6��$����n~�7_q[/����`Z� ��b��%�k��8w�3�J�XSh�ޜ`b��3☂b��d�"��!prw��Ty���Z����Y5}��_fLD������u��+р�&:x!��	�5�4�A$����0�ޘ��6O7ְ��	+�Zc�^xu��]_;���oen��&l�S����'F���ҝx#9\�5� ���A�~V��x\����ί�h�檾<�b�nQ$��I�kG^&=��8����5�	�
�^MT�����F3A3L���`uA�����\ �Uq�׷W�G]N�6�;S>�ZhBCD�;QD}�ɻ����6����œ/��>}K���oY �q��r�����UW�N8?L9ZH��r�b��#'/^T�q�5ԝ㭗À���_��J�J\�<U͘���,;�,��Y$N���ghй1��\���'��A�%�Ϋ�f/EE�q�3�O*)!�_�(y/l�4��(�z-�)5�B朙�s�I�AK��Z�8��hf.��w�$]�p�ܣ_y胟xKځ��,�md7��\�/�~'�?��5I�(�G5���Q�A�h�P�@^4�	8v�V��D{*��$K��P���Fs
C5�U�Q1�G���:?��. �k�׻�:
S*y���i��n�ѯԹVZ/Z|F!ָێn���d��E2sr�S�?Ukޜ;~ח�V��f�|�M���qG[=��V�����t�w�$`e9`�y���=���dcN���ʦ�,Kyh�2���B�f�����H�e#����'V�P����Vg}��" ��9�u2/���T ؔ0s���`���j�~��|��xH���R�7�\�@�H��X>�-��&.̻����3�?�s'szG���_��7_]7��K�0}  ����[�P^���m�X���^(ZV��V���ӿc�&��Ю�G������4 �+S^)�g~?�Zis�;�S)������7q?g�A��L)���'f�w�e���:��dF�����g�Y���z��?s�U�ح����#��A�;���z��q�~��z�[*V�!��S�^.�~9%fB�G�H(�,(:63���s�3�����$Uv��o��a�-�'��|&c|���3OW*��3z*�`��h2\���!tV3�zY��"�SAB4��~@$��}z�4��\9s�����=����O���Z�%g�.��+��e�i�5���8�Y+�IG��c������MY����
A��r�(`gN���
�G����#B�"�>���]��Ui���?B�x���Xw��$fˬ+X�lR�{b����o?s�-���"O[b��\���Pr#����U��ШT��bU�^~�t��QMnJ/�UV��W�s�֋V?���<�o
'!
�N�4A�o
MޔF'�|�5h:a���'��aQg�T����J09L�pLJrC����굹��7������������ ��)�"X�=*�u���/ɪ��i�S'J�� W��W�z��^w������f�aVC�� A���;+��Hq/�孆�KM���m�T�<V�o�6겒Pq�B�6K5{���.Nw mu�냷�c���G�x�[0E֠j%I����4���Q�Tι���ka2˲ԜJ+��pSR��`˞E,����[��&4�j�pD�W��u�º*��(�!���6l�������X��h��-�f�����|�dZ���v��/rN��t<��,���Q�7�o�M}��D��;����Z��'2��x�ұ�y�Q*7G/�rߛͯR�SP���3���!xT�3��z�*A#�C
|�
�]S�% Z��{��8����m5�}�Mq�.q!���>�jVP��1w���1��vxF'T]wpܑ@l>��[W����f��P勉- F�A�-�Y�׶���0مL�]h�P��D����A����ӌ(Se.�l�C2W���^u����;��]�	�̪K�&�L��X�k�ޟ�{ 5B+ �t8���^I,��MeJ�ˠ�[*���!!7�>Ί|�E�/�p�щ�\9�������j�I3�̝՗��]�P�q�g���%�JY�JZ��p;���V*��/�t�B��		����HfEZ����A�kZ��6�V���U��ܝ
�D�c�,(_���(�s�XH�fSF��4�!Si� .�H��Y�Ծ�TpɄ��ݣ�l�߰���oY ���K�{�}~���؍Ϥԃ�	mMh��5���X�i���)#������j!��a3.��2� �V�n��.T��Rmm�\O����-LR�֑�@X�%�[��N�τ�s1���Z�:*_5�4�a*VQ�E��f��d����Fb��'s����NI):ޒ@�k_j����~�p��/'���C����e��K������% 3P���B�j��^��1���r=��y��w-E嗕��/��q+#Y-�1��Q gD���|HeS�3�Ӱ��l��	Znf凍�=�e�A�~�9�J�}�BƏ��˩�C��:W���iXئ��~8qu���ݭ+���'��/7b��2��:$�idS4͓dU��IT�V�dҤ8Ii�������i�&N��e�D���p3F!ͦ�w���U7��}0�k�
�H1�N�A)+& ���gl����M8�K��&�
.
�[x1=�
����ly�<�v߻���u��-gW���{��V/�x�����϶lvW��R�ơ�Tu���M���
�h����m�J��?N����8PW��e�eVW?�*���LMʌ9�5�����E�f��UV��n���*x�/�)N�D{A�B���rqA���s�]k�k:7�r|�D�j.�zD�<ƎKsr���������
~���q[�ѫ�x���6_{�W�ϙ{�?�$ky�+:&�(%��	W@G�e�������T���@��^��:V���.���5�AI��LQ�d�wZ�1*�fzCT�5%�"_�6 ���>��"T����\O�b�c�@x�!/��w:�g��_���Ehp���h3Gli�#�4�����\��N�i��<�Z���m3�t�~�y}.���r�{�?����~�j8�X �������'[�������b��� ��@���xfuSWNuҾ�P<��3!["Pkbc89)���L8G�7_)' }�SޜvV�F�h&�^�rJ�S����o)	Ĕ�8/y�m�t��l�襕�L�S�ȱ:ٻJ�3`*f�VW�?��B,&B�Z!S�-'��$��fM��l��v�v�z��ݖ�]P۵�p��N��N�w�ן�7ؓ�m�ޓ.o]{⣇��?�pũ�A:WGA����j�E�ﶓ�x����(88C�%8S�:�s�7��(|��ה~��!�~�qhW_�u� �ϋ�j�'m߬�����dZXHU܂�	�_ D��|ĵ-ecu���ԺH4S�����=Q&^�!'&)R�z7ks������{:i�Z\�z쎖�ɭ�U,�m�BUq��f�����1��>��1�G�ݽ�Olo�~�_~|ߜ�ԛv��#����_x��n���lԽ�^��j*MQ�u����yT)�"�Rfm��+��9���e�]W�[sͅMh����HF��j��
��/��F'd7Ie�~[�k�k�X\���b�$�R�W��nl^�Yﴏg��B�QЇP��ń=��Tip<�qZ,,I8�i�1W�Hˁa6��,q�FčȩSm:?&��k�\�K̥/��u/#�y��%���Lz����}��u�>غ�Hk��:^��M�[__?�u����{?�4e;F��n�`P�����T&�'ڥ�i�u`!i����E���\x:J��"i�^�I��F�dXv��b|�(���=���L���Dn<O�ڰ�O�G���8��K��p�%"%��f ^ܶ���%����R3�W� �����R�L���k�t������b�=���o�r�������#M�?���	��	juD��	p����ޣ"�k�C�|�juY�?��u���c������UN�M�_���x��=����8O� �zJ*.�	��dC��S W�(������n�0<_[��_.�y���3�g�.��� ��?����������l����%�1�wN��d�g��[bp<��3�aG]R�@���Ȫ0�w48���T�T��Ӆ"!uW���J:�}2-���$P�p%9m�H՛�1�A�������m7�]�HK�ʕ��s���$sK5']�k�����ޭn��v�M'�RKԄu�"?�����vv�>�?y�
��[J�{S�غ������������Lk��m N���k� &�.e�g�y�T�è��}R��o/��_:�;�<��}�����i*����>�ǿ�Ql^y�{��ݨ��x�������n��iT��%۱��q������F�_�������ACp��w"a(��>6�3���y��6&�Y����k��I`A�8�M4*�x��ͯ��K+O�-/�8�vl�9�:*�5g���ΥG]o��yw�cnxx�TB-�M"i�|"�(8+tĚ��u�6�G��D���ӽ���x���y|����}[�_x���g��l68��&�Ԡ��m�&E�Ԟ��%lߘ�$0���Ȧ����Ǿ��мY�V�j~��?[:��3�~���������SM"�l]��7&�ݧG��c�߿w��?�'����M]yi�m31���V�q�h�����'�WQ�J!49/�� ���ڱ�3�@��$Av�(P��E�{g8a#��ަ[`�]Tj��է�+k�����-$��?���D���_k}}:[/�n�>���όƝ����gOne�]w�q:E�U;Q[g���'��Q{'���Qg�}�흇�/|u/q[��o*7z7w6~:5�݉���gB��.��}���3Ji��|-��`��w�S�:
Cm���=�<���|�#O��ԯ�v�ᣟ�"�������u	.]���k|������n~���h�O�( �K7n��RG�H=���ۄ6mO��8%���Id�W@�����Dr�����>����E�'���Cԓ�x�=�k7������ˍ��F�\�O>�9��_�A��}����l��/|�pk����/�xi�����/Ǽ�z\Y�}$(ᄺ���)�������L��f-���`��O��/�N� �}a�����G�b�%q��@K�JD��y�R�ʢG�$e �&�I�t��������C|���a>�mq:�ss�q�����Y��R1��][ldGZ�˹���n�=3���̊d ;+�P�E��-�eY�	���}�w^yB
��	Ă@
D�U$�]HP.�Մ��s��3����s�*�:����}�>^R��=��8]��_��l�W�[����T���1�0gu���D����LQ�b˫��1� F��w�3/�M�2J�D� ����ےn�o��Y�+�e�6s׫�6+v�k5[��j�W[�>�������Nw������<^�U���%���*QqPu��8�T3�GU��U��5H:Y3�[�]^�*�`y��#b{j��}���po�7c�@���{H�9.��p%�4Ւ�P���'c
�&��%6}�ܼt�g��x����:�!�a����e1�4�Zgs��=��}��Q��'�,K�9�9��4c5nŞ�2T�2�UY�|��P(&�򆆊R(}JYV�ڶ� ֎�b{ġ�Z�T�\�x~�_��3�˿�;������tnnvW�n����tl�P�sԖZ��  ���f�-h��9���l���}i���{��7�=�ؒO���EWp򅔯ˆ�n��E^��))�4u�����������\���e�;��p�@d��8u�m��v���+o�H�%D�>�|�Z��ܡ�f��GL<^�C�?e �#R�v�b��d��"���)`v��󿽽��_�B�?�} -���J���Q���DF��TŸ*� �t=�e�����ƽ�&q�A��Z��ݼ^��v�p4Uq�j0�cȡ����Q����:5����|Q�U�?:��������=��~�v��!�p��2�zR8��_ۻ�Ɵ���_�~����_�6_#�b��8�H�:,��hd{���(��%��GKΊ�o��ry�A�ۯ�|�N��yJeP�ȪX2��S�H��F�"٦n�r�/�U��#o�v��3w������x�g�_�V����c�ο�Y��a��e�Ȭ�u��`헁�َ�\�D�d���#����m�@3��Al�؉�N�'�4g�S�Ht�0P��@!��l�)%c�X���$�;��9�{�����7�~��_������� ��w��3{��/:Q�B�FӫZMdQ�{Wi��Q1�����v�J��C���0���(�p�(>h0����j.H�fQE2��#�B�KȜ�k�f�k����o�]y�
��~cg�?x7�����zq�s��^ ҊÎ�W��	��ϕA����)��4&hj�OH�G6PA���"����8P�ݐM�\L�Y;}�;�S�ϫ�篽6�����a^7ȇş�W������t������$�^�!q =6�UK�D�e�ok�w�qli#�(��!�A�#��␮G2V �����Z 2Δ�j�@|+=Ebmz��[��K?��Q18�3����Lϭ��v��\Dv�wI�����k����1�P�5����F��Qu�	�*����@/��V��g#���@>�L+�'b�=;����++����XE�?X��_߼����__�0��_�`��U� �W�n���)*譋*��O�6�s�!��زݞ�|�b�b�X�X����v�|\l&���Tgn�.>�N��o�@rBh��>��������/T-i8II_���V�M�"-�P�Ѷ�5�����e�>ô/]B�1����RF�;�p�@c.�VL������,\��x��A>̼����������w����9J��a	3�B	�1D�Pz�nŵF�j�P�{��G]�z;I�G�<�ya����D�T{�۰�Z��^�zK����>�sW�Z�.}?|�|!��G^	�eR��YompX����zd�қ��5����N�`Ro@�Ƹ@� ��bN�]�^n�/�>5}�0{�������/]{�Ng����%��U'R^J��ب�:�n�ܑ�#�2��ԧg����F��0��)�;D1J�>�7+͹NO���2�8`4�s�oܿ]����2��S59�TK\��8&6ݲ�3�O���i�o���ËuזVP���]ǃ>|ͫ��ba�2ϭ���g���3�?�N���h,,l5δ?�
��Xbי��Zl�뇈x-�V�^>�xq���#��|�/����GI?�.��K,2�iE��huz��:�?��M;�$;{����^{���Z�`�c�Q�j=�T�4[͑��'NL���:{ờ��+��gc�=إ�]�jҭ����͹++�Vi���"0��p��+aou��a���tlgA���j�o��./���_�������x�~5`ȅٱ�[M�[o�]|��Xh
�`<�[g:������� �&d
;��2tV��g���WF�� |�A@M�{��V7����f��lWQz��&x�:w�A�]B���:�.u[�+�����j� d�[��?l_��c<����1���������#���׆!U��bJ��Jc�x���Cǝ^q*gT�d�´>�s�s�9sfq2{2�HӳAB��x	�(�x[��{�Р �
�Tg��ٽ��d�*e��� ����̳��5��o��6ū�\�q�f�v�{�Z.C��)S���ŉی���2�k"۱P%�a?d��\X���� �]�Yg�E �%5ڡU���F[2�Ku�(^*�Jej�՞9�Ȑ�C0lN<��
&�lc:������6e�'��)���ƞ/��K��0��X�S+ӭJ׽�he��<�b�:���N����e��g�RN����R���څnP �D�Q1�%G-O,���	M���ejӝ���Vߥ.���eaN~<�8�[Z$Fd�C,#��#��`2dM��5�$ؠ�1	5Q66�|�r�!0Q�Zj
�8�GjA|:򥝂��we��@��16Ae��ן�T��F���d������!�P�� �"R)ť��ANA���f�H���x��@fe��"@��Ȳ�,,R�"r����8c�U"b���Di�Aj�]���<4�x���;�П>�s�a%vPB�g�LZ�<�&V/=��LCLih�1f�p�=%�&	�� Nx�Ї� 0��@��5�"K/2qr`�2WFYhɷd��x��.<մG��2xvK��l���d�D�+e��y��T�$��b����Gb��D�T�iPP��\�<��z1�'a���-�L�P4�>]0�U���c��f��`#�J4�bR_2����NJ!��8�J�F1�(�� ��fҖ��Lr�e�5���4nj%b��|\�z4��T6FUCV���f���n(v$�*�b���1�ĩ���h����^w&4�
�Q^��fP�\ĩ�� �L�DcniQj�=Yգ6��@�C�{*F��އ\W��i�@�!d�!���T�	�����5>Y�$����I��J�6�MQ*�0Δ_��!�SZl�9_��m���@C�1�4�T�e_گ��
x�|A%T�Ru^�23�l���(\^�<Q���#�N:?�,#�OC-=������|�况ʃߙ���!�e���(0���wC)&? ��Z��4Ԧ7Q8!8Q%L�)�(���s�s�r����/���(��&���
&ze���q�C����F�0ۦ�!*c��\W�e)�^ŧL���:X��"���8*W��*�4<=���	2� �	(K?L���G��%�<��5:8��R_=��{z+C�3Š�	4�h�?5YM
r.K[���O�5�'0S	8hTT��(�Y��$@�/5���?���c�n�ip�$�v��2��h�)]x�Z >��2ʇ���T�Ui���_.�F0�,�B��j0�o<Eɀ�V�<�	^<�˷���� xC���!���6�n=
�1�v'� �ӝ�8� ��f6�T��ߏ<�o�SP�Rľĳ��t�BC�Ups�����@�]d_�I�`��G�HG Lqj0�IQ�h��~&}e`���2CМ��t"%9����Ƞ\(���\�D*��21(G�f��Qc�'C)D02R�@��x*j��(�&eh���z�&�<�(�R�g��ӧ�����O�XJ/�;�d�2�Â'�� `<+�C L���`�iV������8�%�Z��%c#yc��2&�(���7f�I��<�?Đ!�BD�`i�p��1��!(Uw�`=�|�Y�)Y`H�ɶ���)4�2Ɓ��Cɰt�8C��aE>�"];��Ν&(�Fv �s��yy���A�{S�(�ړ��lig�i���t���*6�|%#;��8��9a��3��2�P/Ci%�ĉ��,�A;�C�|�o멨�CPsEe�K�����"�2�x��Pb�I�d�N���(M��B�st)�>D/@�ɕ&F	��hQ�/�b��%��L|���=8��*��w��na���M-���#�T�1�[���*����}�3� �PFXa�\K�BCidJ���g���+N���Q�`\�PU�tC�\�v}�@=��,�R�s�P�5�/�'�cp��U:h=�}u�
��Ե��!�$�4�F9��M���˄�C�L^s)���#�Vt��R}a�2@��'@Y�$Ȳ�)=B�dSBXh�_<�f�:��g���/CZ�S�%��vB��lp-�<���B�5Qd@���6�<��-�
��B~�0�Sc�a\��XV�j�li�Aj���dP
,k����A�t��y�.*��Uq����эA��TYy���`6Y�<�+I��)��P��U*`��H&xe@P���"J��c�CNX�PȐA�7(��H��^>��L���g!�-�R�lKB)�Ɛ�>F9��o3ԓ~[������	ed�W�|j�0��O����̠j~�x�r����ݸ&8G��4���X�?[eO���o    IEND�B`�PK   F�X�0��^  �  /   images/3cc6de24-d07c-4ad6-96a2-959384ef4fe5.png��w0^��u+�.V_e�(��m�UV[}�.A�.Z�.Voщ��%�H�Zt!zId�r�3�������=3��̜9s��9�<���PN{�����:��7�	���?��p܀�G�ҏ����_A�顉��"�_������?��ׅ(((����~N>.w�}�r?`%"b�VW5	����=��7������x��vӚo�5��t�[?{g[ؖ�RIP�.Z��2�m+��<��6~�3��q?�/���54�!��K�͖���*�3嗺����F�[��
Se�۽����E
6!d����uH��PM���I%�_j g H�yх���Y�zy��s��+jՂ����D^�)(~)��j�W9��)q���[��}�~
lpy��k�mnj����1-�rc�V �߬��g{�G�lw��JZV��������aQ\||U�6�ڋ庌=�LLL��9���*��6�%E�1�*������� ���K^x�� ����/7Q:���a�����(��$��'U�U[�������y��ohE����n�5Pi鷸�.�kKG��l�������k�
i@���p�.0�m�T�;�4����*%xϴ��J!�:ٺI����F��Ip�R�0��@2j���Z�s�D[e��i�~�L�m&&�$���]DC�G/�4@i��.�.�o�?��=zj>uv��ڰ�@1�r�py;NǚKXT������*�� �a�{xx��wץ�'�0X�aFpA�c�z���А����e�V����5�+l�hw^�!AE��"��d&*˰ |j$_�D1��sg�l/�K��#���e��8azj*���%K$��U69--�X\\�Z�[�k��I7[4���&1����f �IKK�#�=�".{�t�R�PI:{�5i�(�уm��QhlVMFFƤ��4�q�v1�2�*�g������A���ji�c�(Z��F� ���C�nH��<=2P������LL�m�F���KOMM5�!���3E� �V>�%�'m������$H4�-I����.�Z1��-�#^�4ො��°�2MP����F�)�y�D��ߣ]�Fא�7ƒB���2ee%�Q��tg����=-���9��uI����EļW+� ��A���\q��Jx�$�k��T�HS/+��6g����sO���mFm�tρ�G	tx�����SX��c�;�<�r�
��J��p��Ȼi�7��?{ßS�g�f8J=��Y��3��&?*��x;6u�og�N��~Dh�nI}�v4J��r�9HF�n��/9��`�;��c������i�v?��7���8*`Oz�H�i`�*���v|�w硱?�<?�7�'7 ��k
���<�ù��sM�6."�w>������v�C�' {[���i+�YYq��O�q��(Ȍ��?.c�(`�l���P�v��2�HW�����Q�iVf&]�p��]��M�Jt���-��B`����sû��UH�G<ȫyԟ�8�t�Q�=�ň�ڳA^V�=���:EǴ��B�"���aB�F!$�R�N�&�e��x4쏱.C��
�����%9����U��;x����h�2��`;�����^�;���;L�J*H�p�� �!�iޤ��#��%c$�z���G��^;2�fi�Ċ�<��q=���0�ݕ�p�3P&���&���[�gc�2���.j*.�5�瑶zZ����ظ�Z���M4��y%�&z��e)�ґ�"��&-�1��CT{����f $�a�wĉ2�M�F�E�lXlR�Ձ��H�p��r�C2��AO�X��u��r5J`�F�y:F�G�WJ&���R����7�4xYٖ+��A�D��ˈL�������s���Ι�+��?�kф��5l{�3v��F�!�ee7�e����{e�3���T���-Ǌ���ս�q�r���~�ڢ՚w ����֌\ݮ� =7)�#�ꬦZ��3V�6�����GR�I>y��3��B`��g%�;
��Vɫ����]Wg"{+Sӂ �O�����LML֛zz�Si���+kkg�a���R=����E|7Wd���!U���	%"�]Ώ�a1˧ߧ�g�.WC��8.ȥ����د�����9U@�n<�CU켭O��5��M�4؋/��y�t3"����Z{�֨�u*D%����R�:Eo�N��|`���g1X[��O�c�����
�ە�	}c8G@�c���}��e�qR�_���r�(���Mj�*]�8C�6��N��7{B����_��Ϗ��윉/O�2ۅ=����e(ۅ2����C���j������\�����M�TD%���+^��=Zh8w7��(M�z_+�C�,7?h)�U-�ۊ�Lj��Rgni�^�uydE����^,�^u���U�\k��,�13enW�(��B�]��I��k�eFV�N���&h!���P6�8J���m֙��Y�
��>��LN�X��a��@��`��������ǔ~X�>��w��b���X�F�uU��?x�����AV ����s��?+�V�HE��_i��ߖ�����qq�����:%M�P�֭]�T���F����%�;}���x!G�Z�%F\�=���+I��Yқ���I&��t��n1�
̴��92o��>�����
�ͧ�ي.x'���sa~Pc�ܿ��[A?���,�B�1b��<$�ۭi�dF<��j M��X-��]ĩ��ѬӜ~(oc��ka�囋x]�J%���G�����:��F���_sW��Z-C���w2E<�)��`�~F0��f$��"/��\x��J4+e��/WAgB��^H����pKqR�۷f���yP�JA�f�����i>����vH�m�C���yy�T��C�U��x��, �����Qw�e�vGP^ >  `W<�o����Կ�ͳl����dO�d9�o��(�A?��]������X�%��S��׻0�(;��)MB��w] �r|�B7+o�M~��@N0� =�3�y��8�p�S[�2���G6�q[`s�HO�Z�_��D���p�/�td�O�.�/,�O7%��O�N���z !�C��d��f����l���%�Ko�������)��N��
)?����J��B�BL��5�<c�B�6���j��[�tu�+������0b�ud2zӇ�JJ�:ƹ�(PZĤC3�4(���k��ӫ��Ψ�G��QET�/��.B�d_"��}_@�*�/V��ƎO��MP��o��Ca���⮷^Nca�N9@�W>�Τ�>�RT��ɫ�4�w�, ?�5� �W�6	H��I�o�n��]L��í7K-�{#��L �'JF̝T�ًdn�HR�K͋;�x�Y�B :Ї6y|s
���%)��ԮD/h��5�w������_��2J3H��$�Y�ti�����W�(^y:�.5)|3ũN�G��}�+J41}���QZ[YNbo���4��S<A�%"���y%�'M��*�]�R�.�0���K���$	�/iw��Z6fO8�q�����.��N��,�q3�`}�*G�D6�T�,�*-���M�������RU)H�f����\׶W�T��F̷�d ��+  ����~"�R���ַ@����-����@��7�"���	�o='>�+�&^'��pqc��"1�Eb�����w��w۵��W'%�6��;�O�nGY��O�4�KOm�yw��YN�f�B�ͻݞ󨝲�q'�Dp�\G3ۺ��I(��>O!bm����z�ANtd��{;�+��}fw���w�E��DW�m�.P��(��8=A�t��tJ����-�W�!-O��u����!��Ќ��%`>���8�;�c�ߔ�8�t����b?�7~9���z]��0�K��b @�?zv��m���iQ6ң>1��%�!=������c���FJ�$�#��SJ��,��%����;j�,�_�g�7z�7��(	لw� S�>�Te͋��=��3��
wSG�WVm�h��w������2��[)�b NtG�E��4�����[�u����ik��nʒ�wC���O)b���-�:�F=d��A���t���O�'��	�6Z����7���K���k����%��@�I�ws�9��%��@�f�	=���P!�������1U�@�?=�0I�?�����+�%*�x�!T�����Y�1{6`�c��y�Ҋ���k�X��?�Ӣ)�x��#�[��E�I��uY����T��H�R�<)����,=�����30���)a��g�KB��dnzG�A�R��WF����x<���O���~	�z�/�C�m���4�y���>�ঞ[��7�?�|�_�~=Y��|BsR��1�1c��v8�poz�59׻�����6��I5 dM����,���vf�����x���J��gz��{-[A���7--2�=�_i���y��~~~/5#�eaw�M���33�Ĺ�z"b���>��XT��[��~E|v*h��b�߲Ō@����1��{��Z|��������������NڧG�a�U�\���!.����9��n����+V8��|���[�S�|���ff
9���Ʋ�@�F��4Ð�D���#�����❒3r;*����a�[�)I�U���u��f�ٺfm�u�����ް2+k�K\�؍j����xhq�ޮ�<��3�}|�Y����smy��d11t(>�x#[���J�*����h�D�3gѸjNO�����J�g��n
�d����b���{�
y+�Dʣj��R��=�����]��
�	���Z�Q���:�XMv]$�$�dW?�%�1)��?\(��dk���n�����[�}�PK   ��X�}�R��  ��  /   images/3fe24426-b06c-40dd-b590-a579c31a1c4f.png 2@Ϳ�PNG

   IHDR   j     ���   	pHYs  �  ��+  �EIDATx��W�eW�&���>��Ȍ�d&��E�XlV��R;@#��G��yI���� A�z-��R������e�2��dz����������7�LF��&�C#�c��k�oyW����\:q����=���z95i�O�u����cuk���W��0��C�/����С����}��P�J�k4Q��ğEe�CEG=#Gy�6V�V�JY��}e��^�G�	���ۖeգ(Rqg��~*W���[U���&�0�2��܈\�ҋ��9���J��DW5��9�r&��%��
�m��r���\����o��>zN("N@� ��ժ*W�#ʲ�[_��ވ���7�#n���,Ie�^6�~3	E��@���Hg��͍�g��U�k�qU(|���GGG{"�{N(Z�6�e�11�ń�_�z��F3���P.�mҭ�����sB��6* �d6q����F��~���WgG��8l[e�hq/��Rj�~2���*�� [쯨g���b��$��[*➙=')���y���N�sY����GV!
��`��^�K�	5<����*�&,t����Q���#*0a��@������J�Fd�N/��KƊ�UV=GE�D�,��m�ێ��W�3@(�[�~���> ��(��#j�E���}�&����Qǈ�.��0d����<?(�g���`��+����6�c��ս<�Ra6�[oG��u�aֱ�A�!�6O�%iL�(�}�3���@��T�['[%�U�N�ٴ�|�Q��D�(!��tT�}�	��dۮ�d�f��\����Ê�<|��{�ҝ����g�P���l�Z�F��L��`]��9#>�8����!�,
NY8?���X�z&�+���[�u�����|��F�(+�BR�>/qٻN�z�^bC��-�˛y�Dv�o�Q@�S��w���=]s8D��(��/�A���f�B9v+"m`�Yq�D����L������
��������<���8
�q�bR������Լ Kp
U*Wrv��������P&�[y=�+�|�����"�ϱ��eY�U�7��ؽ�FC岅�-���vIEq� 	���>41����~zN�(*����cǞgٽ��0���8�!���J��!m�W��sB��;�{�j�]�1Ic9�(r�{}_�y<2r�L.�`���m�a������<�V!��ka�|B�=�R��Qພ��N��j�^o�ӟB�Qi),m�!��睻ʍIۈ���Gz�I�س��g�Pd�g�C6�~52Y����ɸ-"���|�s�W���Z���Y �[�|�HJ<����y�@��8A⮘3@�X(�=��W��L��Kz���7��y�XЬ=G&C�3Z��s]�6:Z�&Gx�O��3��^B~ٸ瞉����6�0T�zwE&Dг�z�؏r�яL$�`�NOEq����O=p8D2tы�����L(~��k��o�PV�����B,�c�X�@N���n4�(�1)ێ����3A���z�/�.�7�P��Y�٨�D�b{�8�%��Ǿ�;�Y) GY��E�I%߃���yͬ4`G�\�Ŷ����T��k��5��N/��
�z��h�G�;�>��ޥe�(�D�8�8���w�{n�6��j6��z�ӆ������ކぽ��$�L�<����sB�Q�_�V�|���PZw~����s�ް]��d�,�8PD�S�c�	E +G��A(��X(\�i�X=
P	_���i�=i[ ǳ@(�F -�hA2{}G*
rae\2�� ��4{��"�qm��drP���=ݹ8��AB�G :qD_Ocd='m�����TD���!E~�Ѩ��z�y����:��l�A�]ő���yt7����z����>�D� �7�Pa3"=`���Ђ���=99�*2��C�V�����zN(�se��n?��O;���FG��]�>�k��g�o6G������h����fz.��\&��[���~����l�"n�*+bn
� �m�焲ju+
ђ.b��c�egz����"�{Ȕm6����>��ݗ'NY�qˎ�����sBَ[�f�&�C`�B��tf۲�<�]8h��z�l;*����&
�ȸ�� {~Oq�|p^bz���Y,
G�	g�ny��*�Ej��E4��~�e;�V6�s9
��g��͚������w8���F���T��	��v��M樅|&�=��.��	im���	ϏrQ�kv��l�`Y;��x�ʊ�Oh�D����*�韍��3o��#������T������Ξ*�C������۪\.���r�z*bp�Q�N��%�����0�S��SB��;X�6�j���ߪ��#4�T=>�fs�tTV�=��㸷�]O	�l�'	HdQ{����f{.���?�h6=��}�[���z���G�H����@u߉��A
�P��KK��^4���=��P��<h[�
Hl!�Ps���,{�vQQ^4Tt,kzbb�kGц]��� �@�'�e�����e��%��G\�j)�A/[�������pg�B��z������}E
Y�� �W�6z}O=%T�\���X"�P$P �>Lom�u���,�H�t��B)���ȋ\'�-(�N��xQ#��B޳��R��Q�� �l+ �{�C ���n�`�d2����z���˥�n�i���r����x�x�:��kw������������:U---�w������?|������h4�ʵ���7���@����� �*�J��7=�[���7#���rvL�����c�^��(h����@_3��։s6����B!��7PZ���_������;���ѯQ�:U����7���/����i�nll��vx�ʕ�E\���;88�.]�t�����@���Z�CRf��`6� ��c �QM���иyp�\q�c\b�J;�L��8��\7����;<y����fNz"9��C�v���7�^�����V������0�,�/[7��\��h����V�}c}�c;^c�r����[׮^���흃����D�Z=��J�D#��a=(!qc���
]��K�!\��R��x%�Pb7H^��r>-v�H�q
�7xD��4UD��kW&o޼=��뱱�?�������Թ+����'�N�_�<���������WCժ7�������o��_����4I�4G���Vk�����3�<��˸\��9qscK���R�*���M8�&/?��@�1��\���Kއ��f �{g�������M2z`,R��M8�c����W_}�l�U������p�������g�6���g&�쓫_��v���>�[�OE(�)���9�����Wn���c[�776ǯ\�:x��̈́:t�;��*z EJ[�p/���رcjttT���3������ڪ� �
���\^Lᶾ��d�&��J< �&L���;�0��kjcs��#��@X<~/--���-ڔ��Eu��A584���pOChl���x�����Α.������t��ӓ�O��oB=x������_ܹ{�Ϣ8>��~���裏���,�R��P#C�jrrR<8ɄYYY�_R��E��ׇ����gZ
@��*,>/My�J�h��p.�; 8�O����V������Bth���d",,�)�E��tC-]�{����k�}��y��Q�c��s���|/���}wrj�wn��#W������k������+W���>�ş��7����߾}[]�|��x��{�/_����� s���8?(\FM"��!�pp'i��x��a {���'���d!�=!8O3ga��~��u��>&��@��<8����y�l��_~�����AD�P��3�92/�ݻw������?~\8t����︕��[[��샇����W/��C/\��q��Z���E�kw�������[��i��x�$�E�/��Ļ�����n^< 8	�����޽ǻ=��!��ϋ�(X^^�ED���x&ԐM�~;�Y�Z5�
Ko=|^��#���̀9s����⒚8@���H�U��V>�'Y��J:m�3J�r��	��7n�R$���6���E���v�*K��G�3[I�0R[~p|g{�����[gW��jag���{rq�ĄڮV߾~��_�"�{��:w�E�kY9C|@ǜ:q�9J? n~nnN����B1�.WL(A&Ù3\�t��b���ݿІ[�+���b��p�эTNp��Q�2���ApẐ�8p�l��)ұ}�oHp#8�5�\7n��!5�76��i�K��8I��_ax����y��髿B�g׶7�������r��a�"5H����#�K���+�̙3�3��p[������qc�]�8/��ax����h�E����!HL_��JHB߳Ş�4�	�I�B�!��=�5y��F�1A��-u�����2�;�U*5�'��W$�I��0q@�H�F^`k�aJ���v�����l��_]���^x���<�`�ޞ~�_6��~qe����/��֦���e��!���=���!���E"����X,��J&
!��W�5��Eù��C�p5�!�C�s/H�Rv��8Y,�*�f�ek�X0��T��k t�炘�ٮ�w^�L���B���ł:D����f�Ty���e�f3*���p�s�j~q�;��o����W'�N��7��ξKr���;�w�q�fff�gF����M|��'�浫�\+�m5P�S�|!1>�Hn�B�5�_7b�Ħ���&P��L*�5�l�Q"dHXD�D<S]t�WdD#E�:��U0.�NB��-�r���!���KO-(8�oݼC6Y����o���u�Д�|�<��Ŝ�+x|�F����f��z��n�A�]	uccp�έs�֭}���f�J��whQPUWV��zg����SDv%�71y�9��2/ޛ��g.c22�:Ds��'E�-����0ZE�iN���8u^�u�骜������m��"%]��6	�7�f~�ZVWh�>��e���\��6�*h��ɽjE�LG����S�N������O����	��_\X|�ٟW��Eehae�I��g�-�� �.%ѥ�nԊI��m��w�v+DT.g%���1�������{k���������7�-w-��8j4Q��p '�SC��e;k��!�0��3���s������M��3g�WSG�,I�
<,�������C��`}�o����o��޾U��IΎ�f���h@;
���آ���m�������U�ʣ�6}~P�odl�v�6��Y<�W7X�'6���0lAv!>ǪJD,��M�PsM�z�.;[A���߀M����,`�h�5�k*I����x�*mTӚ��W�d��#��s�ՙ^ �q@M���s`�d������
����_x83��r����[�;t%T�V;A7� U hh�;G���i�$��|����믱����e�X����D���s��Ő�!�f�[��qՆ���b�<'��8�yeY/a��a�B�����+���������9��hw�#��퓸�씁'U&�E}���l�5	��+�wY��t~��'o���z� ��������"��D��6	)C�C�?xx��j�p",�_��	�G�~:$�;�o�x�E�G�����,0�1v`B:t��W������,�8P���k��ɜ_K�q}r�Fы��E{ѣ�3�b9fI�p�e�%��R��N���*���
x�����a{�d�;�,�e2�㦲�����5������+���ϝU��c��f�xc�^��b	Ql50<�F't����������V������q���N� �k��H�u����h���E|�w��]Q��%b����`����=��� m2�l!�D���:?8��h&NT2��g�\MЦ@|�3��6���CWs�O� �E%���k�?����X�g�0BǎW�^<�N�yNy�q Η��R� }df�y�HM@�ɦ���'�q���%���48p�D�e�ߵ~��Ф��B|g8����,v ~V3ˬk ���.-�A�F�N;?��ZHAm��d��:�Lp"�a�8�~]���F¥b��w�.sIo��y��á��M��Hԑxκd����A�7���u��HRL�B�������0�����'0qo桺v�:{mN��1m�E����蹧?��쿐Ε�I:�>�\>���5w���Bo�4B��V}�Tq��*�"�B��a��`}L[�%v'�nm�.ih�)�-��SM�5 
DX���bD$B�j����=3���I���P7ݤ_ :�.T�5i�����(�MPtNp]�!R�y����/k���a	9to>��$
r�LϝQ}�O���mu����uWI筭���k���Y��Ͽ��z�uu`d�A�*׍P1��PPT*c4Q�"�hi϶ev3�׈.����n��\$�C�#G؆�xDas{����-؝@�a��}��7w���=p�Av��^�o��I�q#L�ok�W,�1��%΀�p��u��	����F}��|���a��Hӿ!aJ`sTh�D�)����	���Ç�p�J�. ��¢BF���p��(�6u&��"��5	�}4V���8 n��x_Ėx�����g\M�q��; J���)�m��<�q�C��S&n���]�z�	n���.��$0���$�KB(�Z(A���̨�V��\s�������j|b��3@ܺ}G?�����LԳϟc������>�1�sP�vc�\Ӣ~Ko������Ј���~��}�E5�p�1<�5�#��ʸx�u���������������z״^�!>7ǲSW��Ɂ���AH
烛
�����Ͽt����w��S�O��(��\@$q�����q�:�� j���� 3�,���f��3d��l��F��"���׮]c�r嚺K��o>f�~�{�Sg��0�n@:�4�@��8@�+&�&h�Yo�Hu� �3�٧~�Z�T��
G�ͬ"���f�h�E���L�N!�X��L6 �DfE�I����`T/,-�=-p�����C� (
��.��|@2�֭[l4������'O�K_^�H�vz�\a�}mcC=���� *�&D�n���f�����^V^y�Dڐ�r�=�K��eB����/� qa�Zc���{�Y��������)�?ٚ��F�M��H��:�I�d3�{e�v%��y�!5:iQ8Et��b���]3�VnJBx�4Gb�y�q����â���y�]|�GO��c��G������꧅�̢��Ԋ�d��΁ ��q=��{��"D�_���q�:uJ�;wN���?�◾�	�����jxlT=�?�>��oP��z�L@I$� ���� N�w�>��\6w]�qt�(۞'W��,Jn�p�p�0X�e����6D� ���2�q8?$Y�<?���'5*"��0�as�@8���/#I'̑�v�l��/�HGT���/���YK�M؋�U�����{�Ν;��O?E(m�q� �o��o��a �^x��'�'���?gn��~1G:gC��o~�D>E�ݾyS}���L ��jYg<�����3��:P ��\�Dn!���(�j_��^-�
�����I�<�= ��;�Ƨ��4�RVY�Y�b�}��/���$���9 �Xf���C��l|�@"R��h��u02�I����G@m0b�-�%8�6�����#�3`�g�X�bs\�rE!z��������^�$���L�M��`T��&P�!zޣ�O0��V(�@f&w3wc��b'r�P�2���E(4�-�.�r��T�bb�
�3�MGJ�[�>��g�)]��j�C�1��)cN�X -t�\������^
���X-���go\�0ǳx6b���W_e"� ��~�Z&}έ}�su��֩��X�:4��7JFn��yY��b�Й{�lH%C,
�����L��|�yaz7�|�Uկҳ���l.�<.U�+��&+����(���ϑ�/�$=��,��x%��%y/�iM?A~Xh8De�I�KbAM�%�{"2$��?���g��ay���� ��Q�l[A����/^d1���������������0r��E�v6��@����x=v�(��0��78��P�~��p�:�ts��L)�~�s����+~N�F2�IO��K��T�'aH8�?�	
�5[�!
�)�dWl�Z�1����Ֆ���˧B�9_&�h`�P��//]�����S+k�|}D�(�RS[�#�c�"�s9R�!� Ȕ��)�bro XQaK����Fh�}�d���O�����"�[p�����Nh��M�0�.�b��Y�I��������o�y&V���Ky=}^ܗ$[JDB'Y���4ͧأB�s���3 ������CɎǀ8��lN	��%����s��R���bo���r�b�Q���0�N��g��i}���J��|rز۹lOBM�&V�ǫ? ��Z&G��M��s�T��D����ɢ��&�š<N�^�{,[,��rmw����N��xmx U�a��.�8j]�8����7���H�LO�[6�k�"HH ������ܪ�"��	"бc'8�������/���tN%���1�8�V�d��s�k�	�=	����?�N��iGI/Fפ�z�d���NG>�>G� �t�=�0ViT����MM2�=[J��t��|�8�����vvݫ�?�|��������qn̾�L�C�Nc�gn�l��S��W�����0�ח��&_!�4�g�"�ŸM;k�ôR�ډ�^(i��..ۿ�Z��=ٺ��ѝ""�ϒ�
�A���O_[ϒ��<,*[����3�ׄ�6:2�F�9�^�E{ˍ��ʯ{^��'j��XB�
����R�g�p�8�8SKbR�"�(!�,dz�;�jh%����οb��'�{�j�s�{j�=��i �2ɝ*L� #�ޑ$�(�ŤGb�X�c��+55�����k!뉛���ɼ:�c�9IJ|��XB�E�nܘ����3�Lb�,�,\��:-l�E��]w׏����:ǝ"��V��:�9�?���~vs,���D^r������gH�qBi>��	��u��j�Bi�(����&iQ�z���'8�(���}����_���[�^�xG��vp����m����)ݑ�ND��t]?�\D�ٜ<�g��̚+�Q>B}��6�v�я��pq��PLu3�B�*F"�N����P��A+w�������gA�:�J&����,kw�d����R-}��i�)ߑ��tK��')J��+�1�}�m��Mƺu����J���*()P��D�τi%�J�QL�ضkq_���p<�HNGiB�Ŕ .��ҋ�N\ym��ܖ��"\7ni+�k�ŝD��g��X�d�(q�""�4G�r!rjd|�9H���k9�\�%�M#��є�xM�R�OB�'/���JɃ�)�[����󨳘ڋ�v�Ƹ�������
ג�g��%�,�\��zُ�����,46 |~[�NL	�k<v��ń�Ԛ�	�8�{-�jW��I�T���(F0�4���f����*��l{�����F��Ig2ɱ��J����J��#)�?����U+��3�"ɤ<�f��]�/	��/�i4#��U&�a��-��$RC\M���l�g�P�) �ڑYPo��#�ϫ'8��>���ʕ�t!JZ�	a���M��T���-b���ծ��"�jC~�(h���[�	�
;�yv�خ�M"��%��yN�uS0��ix��{�4�XJ�l?����	-B�ttOhR�VV����:qB{�]:/G,�)6��N5���P}��?�+�8�9i�J�@�#�]���x�a�Z-ŏ�F|��Sg���;����vy}��� �$��s��S��8��<�c��Na�<��ĵ��m�������L�<��F���+Ľ�j�����'8K�F#���"���&�ҋ�~�ݖ�?����;�99:BuC��p�t���0d�L������~�#�����w�]&��;��|u؀��0�%�C��1%������BK�l��:���o���Mv��黵��676�8��"�M�u-5���
��k[ߦN�<�h�<i�ۋ�҈�a�M��&�~n7��<h���B����2������:����{�ҥ/�]"��1 ���չZ�&b�~W�"� A�8a�g��9UADd�~�*ǭ�~ k�t�F���z�cOB���ܛ��Sܬ�����J/v7�����{j7H��;)!H�=X(pPl�}�X���0J3d��"}uL5Q��C.��tϋ���
�}���4k�?�M���/SC;]m�;	�n�g=<��dp�w��-N�F�e7�8��W���P;՝��;�oH�4�@�64��t;�4��p�Kʲ�G�q{�N����k�?�����:.b�����k�#�2�~�}����.3H��'����0�s����Y�әsH˦���dPA܋�ٝ[�����A~�H�vL�bΘȀ���T�͒<T�#=����_�i#��y�	9$Qk��ђ���~B0)�R��O/->��M�r��NdDƭm*
�@i��v������<��q4k��ՋNR��Y'}1;7�v����$�+���E�[��P��ב-46q@�k�,�]u�'8t�m��N�����z�'��X�NyC�F���Ї�I���7����z�Re�L(Y��<F��/Bݻw�T���n��(@ki��#��t�Q,6�. �kE�=�FTm�ƤT�����zC 8p���~;�Gr	�7ZP��+#�><4J��O�?^%]��m�)f�~�+.2c<����\%HHm#Ψ"����wWy��ݓM��A��A�t��Fp�a�{g��?���S�����qi{Jz9��thG{�"P>+edt��Ah��݈����� .�!�q�5B�@w`5�Ğ�pm�x��B=��s�߀ti  �����3T�g�E�x��֮M�8X�Z�pܮ��t�;$K����/����%�B$u���kr���|�B^��%�kY"����P�`A�\�E�	��hG��Q�h)}�@2yq�Y@d!A�C�`ǲş�iX1�b����U��i�]��D�X˴8���i�tėP�����`�=F�����X'�}��M���EZ����o����m���I(n�,���gI$}饗�=��7���ӫJ���k���	�Q�!�䶋�vCW8"��K�4TOsR�4��[�V���A���~��j�\e�y�뫜���Sf���>�8����@ON�kts��¼��/�\�
 �8Qdp"�7���U�%���;�}/�s*з�@i2������z<.��ɀ�@(l�F�g�ͪz��YK�*��YZ3�NZ���R���q�%h��4���!{ӻ*)*k��ڎ�B�W�t�͇��@�юFi��ϩSgN�N�}뎺C�h���JE��ydð'`CZ=�T�q&N��:$ γC�R�(e��kg3�N���Ç���55G\���Ρ�c#�D ݍ���z�.C�&
bv�@!�������H�>v�X:��bu���	e�6)�Ӏ ��k�7-�q�_��H��.�l�B�Ǟ)h�`}�������3�,�䄣 ��7��t���E�wY�`sT�a�42���v|m����L ��cǎp[ 	�\p;ٞΨE-/��c�ܸI����I��uk[mml���lH	���)C#LD��:q/82�@�͇�m0�]G�;��aN�qt%T�Dnl����@��DI������m�w�&{	jY�i�H2���P��K���jxl�A �|�8�8>�&N���ja�����X[a�jV+*gR��T"\K���I�Ǐ��!�q�u�Ψe7�gӢ����悙-��A������{U*�A,QذE�~�ƛ)������{�24q|
d��&�_+�5�Ъ�݅#]��kC������7@�K���<T�}��*�pe�-
�.��2�^]F��5����{�c�fY#=G�s5j��8��QR��\�൹;[w*��<�.� ��"���_f�gԋ/����l_;�J�Ǐ|uR�[������C�_C�� qj�kٍ��w2�z�#��LٴW�=E�p �
�3��;8� XH@o�qum�w{�t����&�||��k����T�ϜT�#��"������@ݺvC�2�t3�dq��>�捶i��(k�Ӛΐ���_�K����O��ӧ�/~�3W�f�#v����p;ӆɣGA�l�&ط����+��s�(�P��>J��|�r�Gwτ^ɨ�H����P���msvu�L�$a�.���Q�+�L.��+�D�a��p������y8�puu9�7�M�,�?4M�gl\�^ׅ�Љ(�p;T�gXGIḘ$ܚ.�]�6i���	z
�6����RC���n�	é���� L+��{�7FD&	q������J���L�ι�:n 7��i�F����N ��Cp��Yu��Q��@Y(��pz���
�����nݼN6V���RGg�R���Gu%g=ݼ�]Q�菝8N`�('��u�/d�>�G��������d{�=n�z�2��u��8�&�kqN��(/�Hp:E�R ��F�#��7���2n��P����q��&���,0\�3	�w�	�L� 5P�����gN�9�� ��6��w��f�{w��̼�������=p���E6
�*tc��G��<�^zE���k\MQ1�i�R���(?{����/����d��=p]�&��$ez���ZE9�=��ɺ�J����`����5�!�]؉�KWq�Xөb*iq�$ai@%�HO�	���
�P �M��WbyuEݹw�헍�5���B�n�&����$�����MB��� �i��;�z��ak.��kH�8@�� �Ңބd��޸�쑭'��~`4�\��P=�9�`}��ܘ����T�;�1���nHb�%G�T5F��W�û�B�K�)	����Ђ ������H���?�][hq')X�A��s�����+�{������p�B���J�n�4����d�������=ml��1��G��~֣	;y�ys~-Z����
�����	�/\�F�~���X��I�G��籖wq�X���C	�a���]�)�y���t@Ow��U�z!�y�}����9��Y��-��CPe������3$�$�Y�d�\9�9�p�8_�#�-"��n#4:ԅ&��@f�r�t��K�M=��)�i��&�|���N+du�\�Td�oaa�7�.(�$Bc�S²\%φC���'%T�<�H&���ѕ�l��-��n^�MEJۣ��dD7Sl$� 9^kDZ�ɰ����'/��ې�}�=-�A�;��+1i �r%�7�� ����	�(#��_������ك����F��8�9�Şc� L�C6!8����<��%��̏��C�]�%7��b����`7k��(�f;)a���0=VOg����������Fs�$��L�R�ĠƖ�"e�eR���P�L$��xF��D�:��I�v�>�@?'�(�6]�ŬXA��ŕ���L�	��n
2�%?ϊ�%l��b�z���ͱ��Y�f�iGi�J5M��2[��vh��M���BͥD��	��p⚂[(��f��-�S���Z���F2��s�$��MSlJP�6>7�K�}�`!q��j���-n��@�	�C,Gi�m��hw�~nq�� �b[�|�9:Tl�A�,�Svȉ�� ��ݰM.��N����v�ʿ!^��pB�g�J�숨�L�k����x"�������ѓ�w�D�ko|K�9���ƣ�!
����y��ǈ�Q/��9+5���#�#ݬ���Ֆ�������>[��lhn�&�ur�#��U*��;qG�x���DJo ��3&�u���. g@�h"0ᤚ0��xrޕ2N�r�-��#����d���ܽ��^�y�]w��i3�4��H!C���s�����ŋ_h�	�f}�*c��:0l���56#�	��JՏ�i�
Y�(ܧ�c����H�\,IX�@�v1��^J����D2�AmD|����c��� �?��#����qs��f�X����x�9����P#&��<F�'O��
:�d��c]��nb�7W����(.�\|K�J1��}������$��.��4w_CYI rhd���m�����5���/�f�{N��넦�ؒ.���-�S=dc�}t��ް�G�+M�@|x�e2��[�����b�"��k������X�3j���`K$A���8�����#��M#���qD�ݘ+�8�����f]��h݆nRưƿnXZ^P�/}�Y��A�JR�j6�>������6�M�8��[�gY������2+
1�{wn���6�u�'LZ���}-��+bY)w�(�����Y"��e��۾��bM�Ҩ'}Ӓ�'��`k|�7��!�<3s�
[�8��c�o��m��/��^y�e����j�>�+*t2gю��f�]�������֝��fȆv!�b����y����9Ҍ�bH���^�;uey�m׉9��a���8��-����1󳊉�m��?E�Ý�G�S�#!v2|�}��N{�Z�O�'�|Bp<�ؔ��{�!��29y���K/���6h�1՗�)	t���@K�? �:B�;��߈�J�VU}���ru���w��m5;7�]S�9��6�j�<Pro�� ��~��=߲��8RO�&���G�sP�a�Vb��_ҷ�.�`gB���7���l�k�v�_���z\��쬚S��]HĿ���d�FeM�L��-�L�����S�E���d��^��f	@bHe�} RL�cR�E�
�1�"������1��,_��/0|��ibaB`:���Qu���Hol�]����9R�G�>�5�)�w��=c����┡�C�J"%�0��TȆһ��F��M�i��H�!¦�w��ٸ�B���9GS�t�ֹ4���C��j��x��.���jG���i��2�����v���}�;��4�˛!���C�ح�7��G���?�N�_\��"k{G��F����HO!�;3����x�0a�)4p-!�]������w��r��jq�E6M����0fO�g�*�5���� A+���-c8����E��S�������X�E�{��6���\m�������������8�8z�8��#�[�
����.���:G^9H��g�h��p'i��w+�`�bq���=&��B5��HE`�_��7�d3Y�LM��ҝk��.N E�v�R��bq�9
�9\����Ƨ"�2юv�Q�#�I�D�n�Kǳ�t����L��S�y�N�҉ ��lr����77�9���͛<�A�;��,�נ������~>��(�&�����n�%2�6�&�ӫg�E�QY��D��ۜ9�>u�h�B�>L��g��cE�P|]���K����OP����N�'9XN;��y��<����y�2�BGf� �$q?2�[%��#���.�n@�Z��N=I6�UE'e� j�gz̾��K�4P�\��n��N���XP<�)N�ośf�EzS&khŜO���c̹�?���ܒ��~��8���7	5�KPj'�G�Br"�w��O���ruK���	WR�^�g�X[Ovq�� ;g駐�9	�OY������Y56:�N�z��؂����;b�5�;vL�����0����>��7�_��Z'�aV@�@cr�	$����|�^��8����!�_��N ���� 'Έg�W6�癐�OvI�nQ��N�N�$}}W4ز� @��H�7���X��iB'� ]Z�Dm��$$Q���Q��烓u�}��Un��֨�B��j/n�����7�őW�3��S�:¼��&^|���H�h��總���2&�9��}>�1-����A���	�psKb=ϳvO��Z�j�����kCm���3_	��m��k�Q[�%��@{&L�L���H��6
������1��� ߃{ ���cA�Fo���̧��A��?�>�Ն��gt�+����.>?��q����&~?�c��{��뾅�y1Iw�}�h6���J���{���`y��S���}��WT�.��3Ӵ��@�� ���@kX.[��Xt�@pd2����B�f���4O���^{�U9������B}y�3�F�8E���d�����sϫ������$���7�ɰ�@�j];��`�����d%����J�d�t�XPn!�Ȏ�}zϣf�{����鬿�먘sPf��Lz�K�K���ϩɩCj�8NP��G�hI"�	�f��.��R�n߹���HX(�u!yz�e$j"�ٯ�~��Z^\�vd���m�uBNh��j�Y3Y�I�s��߫�J���y�2r6��`�!�eqeY����"߫ǎڳ�bw�'}7��I�����>=0�}�M~�x���/ �_"NC���"��)O7x�s>a����:�� �e����ʢ�䓏����B�^T�c�3�!L�"����]_Y�q؇M�������j�sHjbC�F�U#��ᾀN!� @4��}��?=7;�R� �$r-���8���Y�u���:髽���h�_�(�Y@p.!Ė�����v�U_|�%s�q�a,��s_~���h ����Ϝ
{Sl~���O�`.e�Aׂ/SjW��"�<�,߾qS�"��ib��\�AQ­�Q6���T��-"ȘP B���y����I_����+g��Y_�̄���{��~�V�{�t�N��M�I-�$e"��I~ @�_&x�:���	qWD�
���}���;�v6��wr���h���
ܲ�y�҇�1��b��Qe9\���!f��D��mEq5�������/�bQX /Ov3����[�"�Rީ�����2]���I���k��k����؋@i��p8-,�� �@ 4"�qQ���h
�����0jh��}����Q��̜��ӡ~ I4��3�w���š�-���ąL��hcm�6N9��
ad�|v�yNܙ�陎腔e��AN�#N�h�f��#Gս;�%�;�����y'��Q��'��c���ҥKZ�;�I�N���ex�91?�Y(e,��1�y�z�lN\�����P�S珞dOD�������_dor+?�9����o�E���>��/[�.�y9��j�/]����H��t�V�a]��Q�Ց������_݈���o�Cl�O?��kk�pL�rځÃ�̩�j��T�O�T�O�T�ü8�z�+<d�%�%|t�o�N�x9u� �;��MC0��[�9�3�z�ӓI7b�$����#�S�+-Y�zM�)sl�a�@�, ��W�Wt#`��%��A/��" �����{�#T��W$w�ﴇGv}?FF���߽}�E��$v�9G�n�r�e<����
�
M���/L�Y\��S�܈b�9ǪHQ�������3A*�;�8��T��_z�ꙙ9��ո�H��H[C:t���a=�ml�C%��T�9��>��:��`
�O2l�bc
���:=���y�a�����M���8��^G{Qr�(E�'�4���b����Y5?7�C��+�;�����/?d;mP��\n�;�SJ?�#t��A4����Ou���fC������z�[���HM?�Q��,�͊��e3�(�N�Y7`L��Е��ͻ�����aɇ���m:�`O����zjw!��� �+9�_�P���U�&B'�ޞ/�X�DR�(���(}(`�4׀�z���7�=\����؜�� �����Y=E���ڪ���I/ˋ+�-2H��<����܆��c�)�fӥ��l�$/�5{�9�5@7��+�F)�y�����q���S������;�RJ��+��l���A�d@l�fŐ�7�j��	��T�{'�9Bq�����_t�zcs��M����[�\c��ya��짫׮��ȓ�z]!��9��h��6)o������V p1�!��{�~DB	�"];�K��j�=���L�i��'�x��Ǌ�n���YyCd�v��H�_##�3-�3ԲU����a��-kZ�a�%;D�8v�kq���;�K���K�P�49�Q	j<�n`A��!C�jtd�ŤT� }��'�i=6P�ů.��Mݓ�����q\��f&2������������r�ȍ���(^d��E�A���t����Hv�
�#�鈧�?Z"@�{��z%+!�|��tp����� z\G+sĲ 2��1����m;�/?'�XR���Ν=�~��$>�H��q�E���eu��-����ν�z��o��5x�k�PU�`Ͳ��B������|_�:����@0�F�(8��d��a��s���H=^&���Ҋ�&�,Ǽ���������n�k//}�:�n?:�[������%��/~��� �C��V�27�,����aޯ,-�VVى�W,��֬W�no�����6u�g����0� gcX�J���=nI�Xlm��#���(˶w�@�0�^���X��"�4؁؏#^�܎��pI2#���o3�A2Y��B/$x��Ra��hѤ��H�3�#���B��	��,̀����K���[g�ؼ��ﺗ��ΎjGz����s�Q��Չ����h�u)�{�D�����$1};���R�$��Х�I� �7����,�$�{��Y.�RD�]�a:�xn�����٠��I?F�o���z�v��iџƧ���-OFi}_������~Y��L��ح��rMFu���Ju��+`�0�W�w4�<u���"�,���y��p�C/�j �z�t�5>_3���.�d��آ�x���u�X{]���^E��9�J_S2�Ѓ�{
��p��vW���~`ϡ�Z�y��J%Tx� ~��^[�}y߶���4�G��Æe�w��,��B�G7��M$v�{q�.����/����ifL����-�I|q�7<��_�9P�J0tޞF��&C���r�}��X�ýpm㉀3c�Jj��Z�
�ㄣ�8ܿg{���0;Uu�N�Ծ����������p��L�[���J.x�Mp�s�,�(5�K�6L����*�f�ܤ�x���A�9=א�Tjҏ8�H�}Z'b�=�����8q{#�4�Hj�2]#%���Hn�vsQu��]fB�/1Y��zt��9KbF���|B;uY2,��f�xRAe��B�C�!+����ʆ.Z���N�=x���栿�G>�ը��ػ}�bNo=�'��w��������u"bG0�R�i�.!.����.u�:��Z��&M�AW��p֘x��g��~���Q�d�������T�`��a�󦏽l�]�i�߽�~�5+~$%�t��d�IM�1���'�Z��R�]x��dV3zJ��#_���%]����N�w[��gWb�G	�p�GJ''����LI���I�g��]n�`�����I��x���O�Q�(��Z�nvP�H{���vr!��n�A�s�\�>P���nI���I�|��ۜ[��N�tju�m�V�/������37F�B�8�SH=��#:K���k{�vLvib����|��G�˦����ڿ��^�÷��şC��R�0�n���6��!�:]'��ҩ�V���MFv]헣KX��-�X�?�<�EN�q�����:��i���&�ef J}O%E_�{�摆v�LU�E�Ȍu�QG8���ޢ �A�:T��)���2� e�D��?��(��1m�ǋ���rS��G:�L��>W:��n۔���Z��`²3���E8>�gۮs)�y���̰���j�%��]�^6w]�u���]][fO<��U��_Ҩ��P���5�~E��Zv�I��X)��>�+���t�>f}T�[vF�2� S���8"Z��Z��PQ�.�q@;��5P;K��\x"�l
�@������B�g���ѩi�
��h�c�X�a��͆oF���F��%��{�g&!rxj�E���y�n�����`���k��[��~R��N��}�u<��]CƸ_D��$
Ӑ����h��/A�wy__I���r������"9Do��`�9:�l��d�8� G��Ԣ��V�kj~iI]��"����/ ���\embV1�#T���]G'��;���i都ږ\H@K�a�8���	��X���@U_ vP{%=�������sh�~���p�\�0Q"�"!�<+}P+H�*L��͘�˸�����n�ߓa*Ȥŏn��qЄ�kO�,����~�v��;�����fI��+y?�J��S��h1	�|��K_�(���B ̄�g:��;���o���@��'��"lr�J�#Ʃ�Z�q_A��R��-GWs@\�P �YI��A�!F&*�����|?�����ǰ��,��\Z̵t`�OJ̙Ik=�$����*�^������آE\[�dNì�,�:,��Bal;[`ɖr����ɺj��*��غ+'����z�x�h���vp� v8Ļg�Ǟ��V�cE'C����ͺ�Z��'84�Մj��V��t�8��� 	�L�)�tǒP��܇��R��0ՊwYmau�(�&< Jj��ڠ*=lfi╶��o����0G��bl�g;(}t3�#cHp�&M$����v����)�j����C`w�P�E����"�.��('E\�,%/���9nh�������Y@b:��Mk�;<�E�� �ѕ>�<g�%,�az�i�,��?G����o'��8��o�H�>�0��/�bs��p+JsطF U </����v9r�q���YN�F~�������`"l�P6w�l����:i.j[�ز���	訴;��X��eH;c�N�e6&��MD�Y"�X�����ǐe�x�pf�6�x  ��s~�`���$g�㓓��LSa�./��/��{�{�� �<�������V�b1k�H�l���gC�#��<�I5��c�ݐ[�Ʊ�f��QRȶ���8����.�y���Pc]P��������>�tI��E舸��'[6z<`�޿�N�9˺btt��� P�d�Bdޢ�r���0D�.�9:�l�(�G�ѫ�kSs�u��k��K�o$�<<o_�v�^�M�����Hw]�ױ㐳}U�33z����_��N(����/�q�A3�>�X�E�canN��?�����~���d�������^����g�XE��J��;���{����`���GTtrf�fdIo�ݙ���?tu�,�S������n\��N�QX�B�#ǎ���y�M�lT]�����2µ��I�8��:=����=�[,���0*ȏ�����b�Md���c�Tl_'.g�F=ic�ӳ���&�cwk ��N�����c//yW�kOD;1���n߾�lz �� ��g�'Qu@���h�Q�E_���d�z�g�&T]���6�DR��4��5C��I�6�NDa���d
D!
��"V�w�w(I1��k� ����#�"�4!ypK
T�q�kz��E�]^��ӿ����}msC��'Os���F����C�>,z�Q�a�.���G�i���fak&.��I'��s�Q��>nmP�Vb��ej5Ҽn^��Er�_ᆽ��۱��\lq4�\O2DY&���.]]����Q��J����gĦ����g:�V�� H耍�-���'�|�&�@���λ��G����;j��u��5u��=.jr�!qӘW�ǌ';4
������g�|(r�${g�Q�Gs�8�a��]7i�\����$�0U<ц�����Oa�ڬi,���N���ڻ�임��!B�C��"��ὀE'?_��3�b [�ݙ�+Q ��l_]��vБ�����	�����έ����+���S��nEf�ݠF$��Iya����0���!���yp�DL�獌�m���j=���.��msi����н�����%о�
���nGO��b�%�&T�<�L� �HG3m�ډ$��=�����f#�z۝�
.��^�꿥Ŭ��
�ÏLV��>WQ`߾yC�I���f8�K^]�����8�֬��sU8� �n�#�8�1��믲~�&�� �B��s�Ë�R�����W������#�<�1C��(����~�O�n=n!��tN�t-����ݙ�&�^�݄�"
���#TR}��L�b����{CÃ���i@D��c4��u/�����Ut�i6+Z�l�܈-�(�mӶgD����I�#��YV#Y��;��Bl���窅��='�`̟�\�3�\��2��5Sp1��i�����G9���#M�ǁ��,U�N�a�5��B4��,�c�TR��� o�!�E���SD�Yќ��\3g
��:8�g���`���h����#��O/�Qh �`v}�mL�H?� 	�.:��|ҕ���v����vT�xT��Оd�������K/�����'�m҂�c���֧�S07������hL�����,�)AmOW�=�-F�r��I�ê������qq�]�w�Q�uO�qQM]�~��P��54���@c��p{e����0O��:b&�%
N7�?�xң��y�����|yyI}�ѯ���ayi�!5�HH��(��!�-�;�9K�"rܖ1)�K`�q���&ۨ�ۑb�{��R��y��.����w�pu"1�gX�l���.R���#V�,�2:�MH$Z�D(�����í���T�6t*f�{��I�tߊ��t讣�zU�Q�.�mWL�{
X�!����{؃�l�@Wȣ7s�gB��-�yވt���h�?��`�J�L�c�P��#���B�M���CD<�/InWkɸZK��x�S3J	�p.�U9���� Qgx|v����~�gÐ��].���n��݉��뤯��7o�$�����
2pL,g�ƚ@����C$���F:���, \�i��΋��j~q5Q�;�H	�H��j�)l���I�i�ϳ5��m2��=*�syz�����^��gXB��?t���D�NfD��Z!�)P���v�j'�pigl�#͉�sI|�7-?m�8�vd�pG���#�I�76M�z�̡�E��xe��Ô�ƢK�q��*�g,7�/�#� ���qq��s��	�8�פ|�0�/8yem���:xx*��$́����q��sȮ����D���]���i�����ЈK�~L�cKg -�kȊ�$T..��$���9�����Į��������R^Oɶ��(��NBR��ֆ��d����Ď�k0��L>�N[gؖ㑲��_K�*~��ooB��Q;Xh�n�M��9�;����!7AF\��kG,��Qi�؞���VR!ч&#�J����E���j�T�'��'R�@_L|����F"뱡j-�!8A�e����Ɂ�lI�pk��~^+]h��	E7���vw2j�	�Io�,$ '� 1�vM�А�2[���Y����$�5�!��a����g�!�ͫ69`�'�
B---���!�.\��7���2Ľ�ɫ�W&@
��or&-G�Ø99<.�T]����S�cr�lX�'�*:�ku�N�S'@����Jg��SB<��o���bf� �P�)�1��*���8�G*��ՙ�ΪW^{�r��Ok{L:��#�	�ʃ@[��Q��B�7���� :M�`SGl�`p�n� ��R���#2�d�t=|B��{d,Qz�g�+Ml���Ń���ʬpz;L@�zU�:��\g�����w�<v\H��:X(x�F'�����o~�a�!�w�[s!D�c��+^�T�U�:`%"+L=�k�$_�Ir9�h���0l��Ңl�����IOL(�0{�����F����8hM��o}K�Ew.�sQ��$E���4�� $�0��O&Q����ߘ��	\/|z/��ym�zS�upfp�T圮YN=��1Kq��+6�M� ��h B��S�I��D±g�C�Q{Ǣ$���h/�"��������Wo��������626��.�eN�y1����s+6�`yv���]�w�	�ġB����>P��	4���Xp�wET����WΟS���k}e5��d5-3�׈�tb����h��Y�l��d�uh%�Lh=*;�ӆ����ϡ��A�!�
��Xч~��Kǌ  k��7��[̰��C���2}oR]����u�
�h�M-]�����;:u��3���j}s3�Ԙ��A��v����_�>��S4u�?'�a:%L�e�Ԉ%^��L��3r�X��aq�i����@��=��	:S��;j�M�,v�@+p�&%ʍ�?~��f���{D7���*ു�����s�E
�ʘІo�#����>n��G�}u��a�l}��~x��JCw,<���Wձ�Ձ�	}�B �T]YYfW��ʚz�ྚ��c��,*e�^�@�!���l`�����2eްHo�)�+�W#«\�
��*W'ʊ�P�#�p!�f���o�h*W�'��@C�p,z���F_��1�e�ðk؍�} u�r)����/�xXd��h2��V]�<�V+˫ܲ.�J���	1zcll��F����༁�~�%dPऺ�HY��q���J��
18I�vZ��H��ņ�kj�Lt�*�5�{����?��o;o���7�i!�s�c�� 7o��e��q�����_M������@_��Uv�taˈ$�A,K�h�奋I��rĖj�,V,\>���ۑ'^��u��l��f���bY�k|�fT��WE��,'Ru����H��I+����ߝs�x��vv��|����A^�cE�̳xi��HG!�
�n�3Q��t�q��-0\�>��.��8*Z�7݇|��A����Zޡ�2�%��;~�&h�Rl���$t����6��,q+L��紾0x
;J�}��m#Ƭ�:��>���U�f���B-�.�'N%Ę:4�G� QY��[��y�ʥ�_��R�+��H\�=4F�	67L��`<$���
�=�" 9�E:~�z��wԇ�q�]���.���r���,x`죐E>cA�r�$��F�!q*`�Ls+}޽���I���}])�5ӯ}�;QZ�#LX_�PC��Ȩ-�lS����h|���6�%�
�D,�a��p�:x�o$��2<�� �L�OC�.�����f:6��qz��n�Q-ƭZ:�P����%��IR�`�a�%̄����u-�u(����?��^E�1�?��(�%�M��v��!�����[���͟�H* l�c�b�T��}�9���7�PgΞe�s���픣Mq��)u��Q��|p% �V�����C&���b�k�s:���1m"�
�pk,�?��ݽ{���x�����N�I	��Q�����V��u
�J����~z!�41$�	��Q�!1#]٧ �\�D�$1t��<���i~���>a��eŸ�w�yG���k:nĥ3��-�9�m���F��=Z0���fף�hZ,��W�6>·ȭT�yvb��>��<E� 8ʶZ�7ivO#]R¯�7y�/��H�6V�s�Fص�Ȧ/�����]Yl\�u��2g�n�E���EQK\�V��Pe4I��(4�C��S�`������'?��@Ѡ-��~膠M�M�cˁ-ʋ*Y������e�{o�w���s�r��H�M���pf�����쨫E���I������U�TpQ%���f �֡t��ڰY��T$�hvzF��λ�έ���g��N�$�S��|��(ӐE��*��r3�W��[�
=�!��z�� �P���n������vu��i�.}��9����{�N��_J��y�lZ�X��qP�h�	�[^����r�#$8-�Z"��&��yr>|�U���Z�0}��h�_��5��?�W�ۦL���[���P.���G}�j�M� �z"�<���)�8���k��YDMU����]B�Ԇ}�ǜ�s��ҁk߭6ح��_P�O�hb���B�qc�7�)&pO�?<���� ����{D��BPP#�T!��ۣ���������0��;��2�w&wn�����m�a�5�e�!�v�B/2����	���e!��/��'�0�\$����-�`���L��I{�pܶ	�G�6���z�_O���^Zd ��H��1:&�$
Q���'Dgw&j�U{@N�?Pٍk�ʤQ����b��_�p��a�`�WV��) G�b���D�O>���F���ZY�Ĩ��u�P��j:��{9ЦD�d�� ��ۂ�C>M�i��r�qٶV5P
;]ٙE7d0<u�z��M$\�o�B8�롂��S�P��>�C���i�W�^�遅/�Mk�^�8�����j�!��x��}�6s॑/8Ekmu�]Mܔ�0da�gq}��[l�ւ�A��%=���Bw S`�A�9��9���LD�!�8��^ ����Q���Gq9)1��6�
��A�������&�{���a�67(�oɴʹ�$�ϝ;���3oA�~���;�bmu9G����Y���f��	Fm�Z��ߐ�#N������s���6����¢�s R�����F�R�"s	���]&�=�O]� p��{0u��G:�F��B���S�T�F�zӞ���c$����з����kŒ�'��#.(���U���r�[��F:�bejrs���*�+<�u��]Pk+��L ��7	���i������Dy�u�Au���g�s�CYe�B�P��|�Dٿ�(餬jDb��k쒂�e-/şit��dȰ}0aɆ	
L�y֖$�&T��A�z�%ԄV4���smn_x�(g�5��M�w��>ڋ*9 �8�"XsK��{�I7h^��"<hoS����L�l����sq �"�n���ҍ��H�m���a{���s}���K�<�aѬG�ZV���P\c����Y��m�,���&[���t�-�Q#��D��ste�������]ny��j������hCӬ|�����[d���2���sS���%13>y�sd�y ���f�[YGtЦA�$���9S��֭11;3�i�1��Ј�����7���*�J܄QN(S:]���D:��-�g���Þ>|�k��'�o��(F���8�Æ�����Hj��+���KސPtl�|�����j$Þ���"L����f�LLN���#�$�׈X��/bc?m������N\6��g\��=8�0��2'�?��3b��1�	�)t�����d�^��B�U�&�`4��.��,ä���6��ϖW�l����>�I�	6����c�A�9B��;��W�q=���,���+�*��s�c1��pǖ0���abh8$8���	�M�,�2�Z�@�d3�&�����~�l䢸v�:���씋\��1����ʏ����Sb���x���#CC���26��+_q�x@��2QqrC�B�2:t��^|�q@�ӧOsJ5l(D�5aT�:��=�d\��0rw)�F���aoB=��	$d���� �#O�"�@��ݑ��,��nzܽ}G��?�3��Γ�_�1SlG�Rry(��k�H�`�� ;)Bbs~�	��p�Ϝ9C"2#.]��u��`n9�iӶS���	�T���q�l9�N�Z{���'ѪG���0���>�pw��)�i�b;
��	����&D��j�ɶi(�4m��8�`�}P�����c��C&WV��w"���"Q�E��pG/�ƨ/A����+�W��#����S�4�bB;ѲJ�f�×�t&�B�em��	�ԋ�:���!�̊*v G�\.�фWÿL��.0".6]	U����� ��Q9�*
>����/�ز}��ܐ
{�\V�r8<���ڣ���x��U7�^!O�����2I�8 ��[�#�.���i�V:^�!��"Y���s@y��{��02D�&@���a�u�[0�C�5�
H���*�q��~ћ^P��\=�VCd@d�b�3'�Gdw�t�s�뭳��pi2q��-y�����0#~b��7���{��"�9C:᭷��ĕ<�,����-���#��ƛ=���!;���Io�,c�!Q��$��;���'�di���2
m(�gTu=s��E1��
�~ч"�cҿ�cn$����
�A>�6��L9�Q�(�,�t7&I��$������r� ��.A�"�����sp��G#��)�)b���|��y1�`�= �_1u�Ó�5(Lq��䄘��d~��1��[m�qT:���s'0�%>*O���;z�]��tF�ᚨ0$o&���<���)�Ce�^%B\����"aY�����!��*�3?;#���?�e�q�&
 I�$=��V�I�7�EnaQ����\�I�;�)a����BԍOM�_c�
t��BT�,"�1Cfߺt�5���nS�kc_�������wlw��V�w�s:�[g79*T|��q.?D��^����6)�v^���i%?�[��Ns�(�8n�H<)�;:���A���Tj�iTgFi0�.Չ�3,ݝ�/�<4���66[���D�Ͻ�������L�B}SБ*'���*������E�X�4�;;U�Nt%�{��q��b���-=LUp�{f |�wS的t�a��MQbmPl����A5"P���hinү�V����@��1���P�jڗ.�DD�Ϯ�0���t�?6j���_%Czמ�qsHt��9�9J��ɬ{�����Wcx�L�z\U�X;�j^^�s���?�+�����-TB��Gq	 ��]��,u�/���_��uQ�����g�8p���ςm-|sd9���(2��1j�l޻�z(����TW5�6�L���ح�]�*�낺���JAC2(�bRO��^o���.�,(��fZNY,�$��3��m��^���|@ &��'�tȮ�GM� j8QM����k�th=�dF�j�D�z]6�� b���Mz� ļ�zEރdkV�3]93֐@"�ٚP,ZM3���P�}�RI� ����ȜzD�h=���!��&��/�T1��$�}�A���Zg�g���Pp�����k��zo� �fB�)^����ʶy�:�:�f�lp����k����l�Pt-b{8A��`(
���J�OYYoNЖ
��
�gz�0�����kzn�Q"*Ǝ]Y$��˞�4�%%z�
�ޟm�`��.v!	4�rE<�z2|���_m1'�� �֔~J����-3�*,��:[:эu�米��D��.����\�w9*| ��^CI7��]�+���F��wՔ׭�s�������S!<$}�4�� +��Iݤz%��@��[R�%��"���kqj���Ϸ"mET?+|qg�5hb3�q��<����`������z ��ZB��~��.�:UY�qk8ٮ�C$N��϶����]F�J�$�VV��I��;��D����z ��h�.t��|�:a��&NČ��z�2�n�pZ5o�������s�]�����+�+۫Emr�`�#T��������BB�M��:@;��L�,��Ujڔ�*T7l=|�p�z�7�#���"r%� .�,:��G�˞J��J�IW��:�w=��R��\K�>����^ĨX7y�:��W��U�6�]ɜ2m��̊S挱�����2�H��l#���f����O�9��oD� '�W]>���H��Y��J4�aBۃ�����,K6��b��9r��Fn �>.n���8������h4^�<�����R�9̸G䦈-��/�$�۲�jm���������H��?G�I�0P�j�B��nNC&J6˕���P.�?W�M�eI����G*Mn�Sf�Ok+��,md3+!f�e�w_L<ӳ3�� mN%)B�!ďX�feG��.�k�e�Eʾz�X���&y>	���].*gp���O�x�I�PB�U�9�.$�`3!��!2�@�����m>p��(�A�[DƧ*��(�"N�ԜL�Ņq��r}p:N�k"��$��-����8��,����(�B�Q;�5���Zth#Q�%!�2:�%�K�� $�������v�X�Dpg��O]��X�G,,�ʾ�6���W��&J�K����� �8�ey����"�Е�rπ�,��F\��$��VR~(��s��p�w�����ݻ�;���������m"�_e[ʒ���
��m�P(�����Jw��ꉼ��6�W���[��~���f���#��� <�ٴ��稄G}��?����@:*�!.c�$�e��,�	�ۈ��<6h�~B��=��2B���W���Q�h��={���� �}y�,��%�z���,�Ų7��ېPX�L�'�d�^�P�3M�z�^�5����aT�f 锭z��9 Bz���U�]B����F&,�xmJ5��*��Ŝ�FU�X6�������T <���t�,����<��i�	�z��Aq��A�O��YG�B��`��HinJ��~�^��G�������1]dP�L7[q�MQYi������0���-���w��������ҽ�36�sX�Lpt�ΰmJ��t��#��V���)k~<N8ը�'��q:��06�����E�J5��P�s�<!�j6%�G5�X��4�ySBg�+}���'羿�X�?kE���}m$V�I�o�z��k�&b�����QD�=���u�����nJ��B�W+/%fg�� e������y�;JYWg@J?�7{���	`0=�@N.��)��
��:��/ȁ��&ϲ���j]�K(�T"�a"���J����^zJf=K뇰�Ҡ�е�Z�0�&��V�{!q�fWiUGՑ���1�Ι���޾}����$�ĸ�fL$�������� ����f	����dB���FDH\"gH�$�U!6�� �!�	\�j��h9O�����ǏO���_[XZ�Gx�_��a���	� a����?���FP��<��gꮔ\�g)W|o��($c?���k "����v���"2-�2M�އ�[虲J3�&��'³��t^��lK�;~�H����� M˥��u�n[X[��c�u�X���0/�͝$Bq� D�ί�_(̓�饟�D4�OC�#|f<��N27���q\�RO��>@/�\~�`�S.[�ް1�K����ؓ��e�K�5�L�1��A��4�g�x|6�<�0��p�s�`v��H��@�~*��X���5C�� "�`�B?e��Mfe��]�/2��?�{d�:s���?��Ϯ]���O����[���v�s3�t�+|�Cd���#��V"D9:!{�'S���1�2H�R�����wH�_��MjW�=Bz�B
x���#>��#�C�ufq,!��T��ݖЊ[U���=n_��������hN�X�A��cq�� z�c��A�O��9��,�-+�1�%�b҉ؿ�����3��w��Cu{�O�����_�/.�dyr��mm}�R�L�L�UP�\�$�&�nB?csP����s���G��'O�.�!]x��7���<��B�GI̡K��	ls�eH7R��^~Uz#���+��˘P����_�ϑ?1$�a��S�H�#�1-;����x�L!Á3����d]�j�N0��p�|$����ή�s������Ж��Є�z�F���7�|��L=�~�����6{�M��� yqg-�p=����
F�Ai�ǉ�.|$f�z�1�RN�t7�f���Ԑ�k$ZP���Қ��mX�����v��<����d*ɳ10*��8�UbT�	��N�Zޱ�7���s\�@����Q�/ax����2g�������@\�Ez����r��������w'���$�vD(�?=M��{v�~�����������f����?H��e�e<�JP�5�#����䕽��1/^��w��fk>��-�;F�f/���[\��4��uɷI����@���� �uuf� ��b��H�n8�j��g Q��ׁ>!��܇��ʃh���ȓ}�X  �<��P�_$�����方����~��o���������^z��o�����\����\��ح��tcC�(��&d�OTN� ��4���7B\���A���s�+�N��"b8p@����2����f�-��4��zAǁ
HU.����(�*�㎁a�-��0�9{��90�q^D���|��6Ў����,���y.q��f~��+:���v�w����~���w��;�u��Y��+x��������O���?�8�æahJ�;#�����`8�"�bnEvq!�k�AYd0��߻�����H�8q�=���CFk��l2|^5�Y��!Aq�o.\��PY@&7\�O��ǟxB��!�G�#�~�&� �Ӟ�nvE͐X���!�.��|ANe���.a�wv�_jmk�Ş���9qbV<��cB�+��2F?�^��7��r������wr���B����LmN�6 Χ�6-N��NF�с#L�R��RK�:Ć�9l(zF@aOL<��Z��zC�d�F(����.բJ�ŤSu&sy�i��%�$�pmm��z��� ��؋�9&+��PC�^��dƳ]�_f�������spp�����x��J�^xn�;x���k��o�{w�gjj����������0:i#S�x,���h�7%R�):��A�����E����ΈE}1��x��6'_b��ioc��u���	��"��	��6PAHn$��-�#Q�����s��LK�e*ٔ�ߞI��;�}��-9AfLA|C�!Tp��⋀O��1B:���^j�?7ז���'�$�|rfvz���u=��6>%<3J�d'Dh�,�H�����@#G�����WU�$$�C4�'��e}!�+z���X��d.
�d"�iIϷd2��'���lWW�]2�G�������sϝؒC�Q�o�P�tڲz��~M��gf
MS��:�V{k��=�B��Np+�^�Sv�{��WF�T,�2�H�KX��l˳툧�Qxr^�T,����]Dw�J��Q)��%k�P������b��x�i���T���&ى3{���e�����vB�[�!��}q���N�36O8���Eʳ��B�-�	�9�Ѽ��<� �K˶]��Ŵ,��J��.r�����a�K���$��J��L���#DY�����[A�͖�[���_]�+��K���t�`��6�    IEND�B`�PK   Ŧ�X���j_  `_  /   images/43e0edf9-5f24-49a3-b78d-83485af402b6.png [@���PNG

   IHDR   J   �   q�   sRGB ���    IDATx^�wx��7~g���^��m��^\��$����$��-	��o�|!		-T�)6��n������}���{��^�W��}��_���ciwv4�S>��s�ߗ"EG�� �_�
���/P
Px�%�������\.W�^-j\�{P�rϹ\���`p:�Z�ˢ�h�N���ʡ҉:ѭu��N���	q��ΐ���`p̏�G����^�5.�[��B*�Jp�T�(�A�V+�"�?�NE��t:Մ� �QԉZ���k�n7����o!��������)��,9�%�+�(]�v�6�T��Tj�Q�p8\�cF��[BBB����'�V�6��w�ѸL�&�J�r�/�ifg�����`
0���wt��Wxh�S��;4Z�j~nN�t�Tn�[-�.!*�R	D�ֈD�":����]�FT��*��Ѩ��F$D AN��h_XXp�Lơ�ʪ����>�y.��3P�ox7>.v:&6�ob|4��L�J����r���� ���Z-�7;;K�v;��V�TD
�t:��fs�N�K�պ��Z��p*�J%j4�V����H����A܂�h�jA�ӊz�^��'���p��zT���.��.
�h�������:t����8""¼�@��h -��_����z�N����Qj�Z�r; .^z=wb0��Ą<�I ���@���yx��v�po�Z������ ��A�v�J�H�=�#22�8�vz=a�!�I�I/��������y�`��D��/���Ё#WE�Z%�������A)@ H�
���<@��V�=R �{����w,0z�*��\��RQi��-,�Q����$d|bt^P����s���1�+
���h��1�����njh�l��դ���tvv�'���������<7�  �KJ�*���F��=���M��^�Fg�.������I�{:m�A�{�{�FW��ٱ�3�Q[�>�UT���a���K�Z�(�(x  �7���z�j��K�b>�N�" ��TZ��t�,<<�$%%���b���j��m�o���{r3�!ˮ���^�_SS�M����ܹ3��@���������@��E`Py P��j�_$�(�=��Y �M�4�O�n�t�{N����d������:�Ѩ>_����M�ٝ��B@��f�����T�®ήo��ϗ�@�����Y��<6% CB/�OA��y[��S�����ޑ����=�(���O�L��ד5kS@�{���+~���� D-(�&v���D񨶧�t�[%d454����^�^MZ[[���	�a��`�7��@�T���Z������d�s0�T��>h��Inn6IO_C�&C_Ey���ܨ�DT��@�Y��\��g;Qw�=��di�:���L�vbw�����:/Q�/c̃��H����Nn�x�AiB'���F���@ge�?��.����
���3afa.���������� ���N���_$N���N�<��-<H�=[N�x�$^��=��R�ז��Krss���?X^^�pvv�k� ����Ewuu��8fz��}��7n���������AP���(�zH�(�*��
ԙ<"����UjF�G�Y����/����׮��X��V���ڞ����ݏ>�u�J�Q��G���,Y\����!�pq��B��%W'� ��%�[b��w��y铫��j[�t�����]���l�ɬ��dff��z��FEJ�1�.^U[�w�s�ӳsiikHgk7���!�[��� r�&gپ�R����o��	Hx���tJ8��v�����_�tM�Ʒ!dT�"c.�%<��}��;{6���&�'���Y�X<L]>�Jot�裄ɥ�W�r��xPѠ��C�9���a��@���[�ܞ�UP�$z>������~��=rmNvill%C�a237CO�O�5��
]�rj� �R�,��r�ץ�3�����deeA���l��m�ُBCC����� �}��?��[�ޒ��G��?H&'��(�<�D���3��<y��y�ǳq�J��̛?�/��:�DP����۽�G�6�?l�| ����y��}��HZ[۩D-Z���Z��/x��/���?9�Q�q*��}�HEE�(�F��������/�wŁ����?�ӿ>����5�������Ä́�W9��u1�Nh�����Of�`��ǃ��U/55�����DY,˱�}�-i	i����^cc�nll���_�Mkk{EFz��3���J|d^���ST#�s���a��Er;%WK���>Đ��z055�h�ۏ|�_z�Ƙ�W,{ l�޽������?y`��KM�@usK����Rv�pS� �?�帔8_ �@��!X<E�も(�INN$���$,,d$77��ioDF�w(&&J����l�'>�裫C4�ݤ����y����Qrc͟�+��;�+��V�A��ˡ<��v\q���ee�(��e+x)JEUWWK�ɓ'�����i�I_� E�@2��⍽�Fy{şo��R�&�������H\T�A�
�պ���=�c�s�(����N���+�ݠ��u�M�da�Bff�<@�Ҁ?�]�/c�ߓ{�3�(�k�@3������"z�v��������W<�Ž�����G����������H]��2>>I��(P˽x��1H�&��r�̓$'�,:�D�]��������ྜ��'��S^��9Z��F�{�j&�&��jm���^��h4�::�H� �G�nV~�o�/����>�3�r;���_6
%St���ei�N"�K�eeeP�U]S�`vv�NA	T�Rj�4��IG�<y�����F??]gG/-0`.J��"x�*�a�JN,y{�p9O��-1�R
��~_Ra�^K��gVV��h�k߰n��̜�]� X`t%�ꮮ���Ύ�_��w�Z	H��1�S���Ln�y��?��|���B�����$��񜼺���Mdaa����ʜ�A�e�����ql�(v�6}���a??��������%?-_�O\n����7����'U9��UU���uj!AAAd͚4����2��[_swnn�W=������Gܻ����j4:C_�2���H^5xіmx�+B�P}��3�{N�KJ��[EF:��?.���L&���D	gPp�9>!�����wCO���(�S�l\����y��?��Y�EGǒɉ���O��fOSs�xp0�ؠ'H�'��c���CP5*Vq��������Nk[[k�w���߿����2��N)jnn.��'�����͉��BwO?�(�Ԙ�K�<<�x(Y&T�||L�D�D���������y4_/� � (��3��R�92:d����r�=�gg4)U?�@AG�s�=���o︲����������D�=Q>W���{��� @|�G�o7a-D ƍ�X�J�H<K��]WIQ!)**"=�]����O<��m��I �ʔԽ^f,�w�{�_��jbB����AK�v+��7S�s�j�CG��x�Uxp,J �R	@�zB� ��1p���R�(����S��{P�+(��z�}||����|�δ��c� 0#y�׹H�z��}�.+((�N6����0�%�|x������7l���ru��Ҏ"R@ ���R��y�{�p0	(��JtLL�bY������ӛc���v�)
b��顸?�ṿ8xtsQQ��T}"V���%_���Sp�p��ox	D��*I{�B���R@ �l�)�X��OV�{���FJ�덎;�mW_}�*+��R�������~V��ϛ[:֧��V��h�6z�v����TU���EON3()� P �s,��cA_��n�Pi�*�6�e�f��ZW�|ƚ�SSS�Z%��ft�?����ڷ�~����i������'�ԕ�s9�AJ���A;��d���vy�9�6Ƈ��ǂ|�J��IA�JOO'a���e[R��|"(��\�͈IR!��w�>u���w�~�.B�@�0���m?��z�?#���y�ÎP1hoDc*����%��  p~���6�Jק��.j�!��Tp`��m���MOφ�:#q
^J�RMN���:�����x�&��O���C{�,֥ޕ�®8^"�<���S[��qx
���g�a�
zE|�0�;4�wҥ4KPP@gIIٶ����+�%I�zx�cmGk׏_{�͛A���� ���0|8���O��w�@�G�� �z|:�	m$��@��nRb<)//��***y8**��d8��z�477����~<?��"���da�J��<\A�xu����$��"��>s
��P�@�����p��?�z555$88����x{^^޻�#͢2��W��C����ߣV��<`dMddi{3z;��c���̝��h��-�޴�j�R�۲�z �gee��h�k[��z[zz���%�233�t�x�u��x�~�S�Cfzf����Q���7�Rg�(_1!/M<PrG!��'M�b9s`敕�.�VӲ~}������·D	#��I����������̛:;{��������"�M�xy�����X�GPxI���GҶ����N�i���~��� R��#�ٜb�9.��o~�k??�qxh�ttt�{����V����z-����灒S *,,��dgg�������*����ޯ4s@�
A��>97��Xt}��7ߺ�bqG�����8�����O�L�WET�z����/r{��:>F�C�%��BCc=��0  pgIE����V���ݻ?�~�O�>=7�P��[H&'�ICC#�9g��������v���9_�k�S:��.O����z,���-��x���K�v��*�+�(����#���7���T����LLL��E�@I��}�1�$
��׍/���$�I?���9���AG)@���Q���t��-w߶fMV�Rϧ(�p������Oj�YZZNZ[�I[[;1�h4kNx")�Q�I�&r��3�V��A���Ͽ'��*(�#999��=�G�l��qq݂ �v����'�z���w}|EAA	�7�������^��tʯ���3ly��Ր�����z��^d@�ff��f��~���OIIoS�P��m}{��K�!��(�z��b9�Z�w_��7*Wk�d��`�@Ch$�J��i���O4������D����ju�ɞ�ԯ~���PeNN�����(4�&�Ln|��"^�������E�xlT~~>����t�t���+)��0""b�ljGϧ䠣G�����o�۷ykyRb�jpp������ �����z�o��v�l��P|!��>H�/��FML���"�_��򥢢򷕮ZW\���lx__��x��'�gCFF�HwO�{CÃ��>����y/M����}����L6��r�|TZZ
�p��7]p��׮�ܳ�.lx�'���|�k��v��.�`acSK3�Z�4{p&[�ˆ!PhOPbx־e�����Wm�Fi5*�e URRB��������ͅfewp�����;{���c�u��*��0&�3�(�%�a̙�;�9���Й��<|�����"P�INN&�����j��,ߖ�I�4���(Q��������{�~����&���Q20`��K�|�^��x��E+�C-����ӛi���Po��(,�f|�CB�zJK˷�:��]]!���pzSC�O>���f��4���Y��X^�1��K�|˫"���M^-���ߗv�iT*륭��-=��E��q>�R��mki�ɧ�~��ؤ���Hf�-�Q�&r��̙W/�t�L��r'p�7�L���M�yb��K���Q^U��0�����sQ=�3��6���?�~zzVj7<4�d���y����0*J^<��o���9R�BRr��,w�������m��E`��gQD�R9󱑱�_~�??��Z菂���$�?��<O�I%��K�䡍/�� c�ܞ���;=c�p�Ɔ��=����@Q�w.����Y3;;}�o��ea�����#��r	���'�_����������J��FQp��_fV:�u���5TW�l��M�vzs�2OV�D�w���ݻ���T*�axh���������g�zr~����A�c��'o�P��[.�.�t'�JM�EC�����]�k�UTT퉊�J1Puu_f��������sCFz���p���zI����r�|q�%��=��T�ȾX������G6o��tww�OL��_��k~v�P�7W�Y}����er�j��f��d���j�<IJ$���u\�.����/��^OK�|��j�o`��G9�������z�k�fC#�"�~.@����~��K/�ZPP�3��'N��[��U�/��o��9_A-��~��Z���FALF�Z��i�٬�#G�o{�������9��*=PE�SO=�;�]VV���Yff���,��x �s�Sn{xi������������JES�����[�{����RO��U��x��^[{evv��~@��u�g�b�B^�%g���KU�D:q�~�a����`�K�i���Z�'�[�����'7+�H����v�\ҟ�}֎uQQ1�!����iFC�1��S˽ ��Og�^�����w�X���o��'&6�lذ���fKKkC�E^��W�z���^��h�"�� �����Ç߹`����4���F2a��$O���m����xIC��E�z8��R���x$*44�����F��1�*:|皵��I�Iݟ��w QaaI#�#?y��������?�N�j$��3�蓖��/�+
A�K/�yE^��F����ǭ^�Jǎ7VV�ݓ���w��,��8??3���g�˯�z�¼���Γ��f��7��i��9v��7��:��	���!�P/f��)I�`���m�99Y���o��P�`Ia9t�(���J�[j������~����	���Of������Sȥ�l���\�x���<><���LLL��Ln����ks!�[q�Tfso�������x���c��bq��SMd�a|�v%����4 sr��c��E�R�p��թ��.$4����t[ff��(Z�p.�2����N�<��o^����Er��)▬����������.�OޝM�x�)���i�b@��y]M����RH��t*x�fh(>����}�_|sb|Z ��ob�-N�ž��Ao�����9���zSy6����
��qq0r�V?4mذ~{vv�{�A��j��V��ut>���ګ���ԝ�ݴ}��`�\�C	:S�Mn��(����1n7[J�'��Jk��nb0��H�K/�:����������hv�9��^�ٜ�:::z���?����� Z��������� 6i �r6�K�|99sG���yg�1	��{x�V���Қ��鴷�_��g��Q�
B�w��f��ᑫ?�h׽��&0�'�N�����K��n�1f����9r�����&��z*���qka��cɺu눿�_Wqq���̜����0J\�K=�356�����Oԝ��444\?;��<_�K�(-�<���_��n!P|��P=�;8���6>��A�%%E�Ok���7_��6���l�N���ɿ:t���ZX<^WWG\"�-~y��c�pp����UHp�?��<��I�wb,[u���	)* 
�b�Ͷ�������ޓ�_rT)EP,Q@:��׿>����q~^����inn����Ş*o�Q�+�"������E����	��X �L�W�|޵�𻟞5�A�����,.����Ǝo�z�mII���
PQ�s��m���37l
eN7H�*9Px���yiA������y�|�4z?[���š�����"����0���	��������!99��<���gϮ+�灿l�pA������Pz|����}�8<�>R��ǅ���
�ǎ?xP�r� W�    IDAT���o@*���z�upp���m?�9!!�RԨq.����+/���������B��梫ԧg��x=9��Y�p#8�D�?�9�����>D�a���x~u�Px��A3� ������{���]ii�JKV��������{>ٳ���/7���QC�Ta`.��$�WG95�Y5�����!��� ]i�I�^���#M~$66�TUU��!��Ȩ��_�ڳ6\�sE�jll4�v����컷��u�V��.,���cu��|�(����T��Bi�
��ދP� ����9�4(�}-�\3��{ �����e�]Ke�#��_(.,x)3�`e��b�nd$p�������ޏ��s����K�v�	'o��F�FQExW�^��R=J���e���㝆F�%3J#$��3�ʅ��r�g�w�[W�5/���ƍ��VBK��gl�=wpt�O>��FsS�zq�I��ۉ�9���s�n���Y@�7��w�
t� �5��������I���w��Se�' Q U���tυ��2�]VU�����YV�?jl�#opp⑏?��jsS��;�׳��Kt,Ym�/X8�%�,7�@2��B4���PH,��r.
���\�	�f
%�����INJ %e��h
�-�.y����|�n�C��桱_|��˚;�m�E:Z;�[����;��h[x5 b#I��*�l�@��@���](`q����&	O�N���V��?#�d+�z�����ёG>����-͝�iq��f(��-���%
n�o������F�?�D!�|���#���G7qK�'5v(K��^k�$-9�S�������EE��9�wT;4d���|x�G�|������n�
��ܞ5�K�xf�x�ī��Ѷ8h�q+&��d��B� �ۢ��x�4��
[X�S��INJ"ťE$ ��SUU�pqq��hM�B���Ƕ}�ᮯuP�;�@l`d�~}�Hx֎j$�� *�uCh���g�� �����5a����&�쐗b!ӝ��L�+Ja�AgEE��K��u�Uott0kbbl��;?������v79��H���e�B�,��(M�˵�`�@!�h�S���N�ZVW�'ÿ� �+-%�TVV���ť��H_��x��9у��쉉�?|w��]����`e(��ڈ�bc?�����
�	U
�����w�#=�����eA�%n�I�T2lKT0��͙������2��iz�rҟ���zkժ�N%��\�R�wvf|���O}���W$����"1��\8H�?���v��F�j5���;��H�����<F�J@U�n�&�r�>-�؝N�*Ņdafz�i_<���]����M�H�rA1΁Y�w�{?��~RUQA\v9y�$�-,.).����n
?n�8�_a�w��XRqA$ ��E��!Z���m��W^QB�NM���'����RSSa~���3���Dԟj���[n��������F2�^�Y��?q��Fw�7���/��c���^U��6*�R׌Jt�B� qs�&�CUj�3���z0�fbttVC�����;�"#{W<54713:��~���s�s������&�Ņ���rNŧZ���@�ǩ?0t�b��$2�',p�Q�T��p� �tz��3�n����vV����Ķ�wŧ�B>JQ%FQ�5??�����[�_��`�3��75���-hx�p��r۲�2�<ú0s���v!s�i����[ q�$�[�@����S�Ewr�@A�fjJq-Z��;Z۞x����;�Vb6�j�&�zg睏��ѻ7\���NN�,n]b��� ��,�Jz3����ÀY9�+�	0
 ��%* �_ J-h������K�&��a$55���EbwLu�4����k��.(ؓ���h�
E@������ګ�����C��ܴ&+��L����Nb] �Z:!�'��T�.�G]��f9(�?#���d�wA� H$�v���4p��	(�D���VQB�*���2�sqa����RS\��_�����̕\*{Tk2��F�����ޫ�����z9z��,�h����9F�]�D��Il����&j7c�ni4�`*]�J��<��n��0�gNiM���A�ճ�Hqb�AM3	���,:�$*&��F�"��D%�:�W��&3=飨�$󊖫�����������ko�x�d��Z�G����H���u8��@�j-�ON�����8a���A�rjԔ�E7шrh��2��)�A!at����4���%&#�[�Ġ��6 L���&.����=��.�`�&�\�Z�TV���_��de��ئ�[���}�9���"C~.�S541�vlh�]�|~mk{����"ihj!��.�#�[TDBU�9>I�μFG9���H��N� 1�������b�C?K���������zp"D���.'-�A���f;����۹DB�� *��1u�� ��g ��1����8��Tee��S��w)�|.@�����Z�۶�;p��޾A�yd���O����A�0IC�"��Ut��kz��=�7-��U�LTtn7�	��	�_\ �1��$8 �,�/���iH좋���(�Z�@�;qX	�� N�m��FR5��R�-ml��ШHښBj�*�űВ�����䗲�����!�Ql�M���'~�����a���)219I���n#��9��DA�-�����v�L@�A���r�D�����t���9j�"BB�9����8A�T,3@ǰA��� nh Z����i�T� �3�?�������R�Sp��PRT�l��a��%�@�������-��r�X�ƞ�23�J���z
�(u@5�j(�Hܦ "�.✙�mU�h8R���̆hDo ��H`���h���"8$�5�-Z�R��$�w	�.,R)3���حj�U-86~7��H�)�@Da0�T�Tm���R�+ۚx��I���y`p���S�==�&�>r�8�HZ��A�CK��A�-��'�	gj�8C�j�g�vԇ�s���p,V�����ề� �X)�����T��@#�&���U�����P����\� T1	�x삒�WWܘ8��
�����<]�!���� ����F��V��71��/�VP�"���Pzs���5W=�CS���}C�1�[����ggg���*��� Lq8�a�D�i_����":=_EV�(�͠� �/�D��		%�E$(<���������_�*�^��䶵v��ԩS��Z�₍t��ЭN`๩)�D��R�R�X�/�F[��@JT����:OU# (�J�"Z �j��Z��� �r�K�ń�HlNQ�b ���5��I����퀭q�Ep�{��S��HvV1�+*+���&�j��Xr���;E�fki�8|��G�[;.ѻ]]S<==K/Db�f�8 ���4�8��N�Zq]BD�^\�o"�V�`��[��.�k���q�&PM���N�Y���3��1�v&�N6�R�:]@�hfTA���EF�թ��H"##[�c^���� *̯A�6�J�Rw�>�����]=))�QC����-W��
3�ƖUn���(�$0P�E����p�?�HTn�h�[>HX8d.�Vh�\��.'���zV`��T��j ��� Rε&!�N�_�۬��';���_\aͿ�Vrڏ�P?���~�UU�N=3�@��h6HE���E-���	b`�G�`Q�J  7��Y�M���[�w�n6��S�C�N T�݄8�RA,5����M�h�0VE�Htz-I���ö�Vptuw6>�u���9iG��P+�(	(��?����۷?SZRi�_���'OQ�M�kt�:����u�.�
j;�%J���}D.-��w;`�
3�n�L�S{w�6O�h�p�Do�)𺠢 ���F˲�NH��D�������nJKKlUZ�9����}ս������J?��M�����@ᦩD�R�TvVJwK@Q��DpI����B�j���
��{ ��E ��r����4Z+9�|��@��w� �\N��<�w���6�|��DR^RJ좃t�u�m�r�M��ٰ�l�jJ��(�[o�|��O=���r�~jj���w���I�;K�sQKD�HD��E�����UPvw�[�>���� 7�n� �@�6�3�fp�5(�
�VH��`�4E�t��J���	�FEO���fgA�!���?���k����@�����3�{��G�y��˳��u6�HZ�;�ua��mE���[K\� ؙmrk��V�^�`�Y�T�Ŕ
p�����R���W���w��W��!m�*:�����d���S��"�HQA��������[oy<7�����xE�"���]���ǎ�mkhj�6��uz���JKr����j��č+��RO�z lS{:PT���� ����w�<%m�e�h�����	� P�t;�ƭ"`�v��ӓ��hRVZ
��pڏ�?W���3"=]�{����,��ӷ~�w���=�p�����=`��.ǲ� ܼ��ҁlJ����C���a�'GoTZ�a3�@@!�$[(�j�����O�.���EIRBm�V�sUu��5���+��\��Do����=�}�ŷ�9 �lXj�3��e$̉c�h���ϰ�E���eD��LTGL)��cok�*�'�g.k=1SI� �n;M�[_I��=�5��*J3��H6�V�K�D�yFF�s����۷o�7�;�@��b��w�Z 
g��a]�J
�>�j<U�E�Gp���0��6Jڡ���&J��1��G�a�����ƒ���`�fy��4�����hw�����}���v��	�W Q�uI/��u=�Z|%{h��Vy�g(��b�2
��º!KC�L��X)��cwؠ�����=�!!A}�5����8/@��v�ON�޳��}�:��1?�{������/+'؏ ��Q�=|����rJA-����P���ëz�F�EUWr
��!�@A�thH`oeE��;A��z�yFGr��&���}W=R�@�NCts
n��LS����f�y��4O$��qڤ�d=ؐ���PX�cR��܅EQ�(f�X�+UG��H���tK�kʡH1XZR�����*{N@������T��7=R ����Ff�fe��e����U{��� x�ao9��໨zhgQ�(��uR�f��(o���`�YȪU���7�ѯ�������W΋������/N_�žw9r,�j�H]<�%�� �.���%�f$�6���G�`�û�.�3�kIz�����L<���u�n����
�ZPu��>�n]��+��<��Is�����8�����J��'�N5�Ͳ�!�n:8(�N�����C	
��U^'�b�0 T;l���9�$����f���eꏶ6I�5�q����8��L��\z�OccjW\� ��޶��k��������ёq:��.u̡T��ƦU�AA~@���J��B�Ǡ]�����'�����*n8�Y����D��j�����55?[�xrr2��������Ʒss������nd�̐��,��Q�z�@z�u`�,M86��w(T=8 ���.)����Cj!�����XL�*:W�,�}��W�����򯾥���p��?���{����� #m$�28M�xz��G�J@p���c�	;T�(����tP�Ӆ�'OD)����(ޣ��1���Ј�#q1�$/?�M�斆�-w�ukna�I�������v�[�<���`���5.7NEՂ�9�(��v��X�xB�F�W��t��7��A��h�&��u�x��:KMR��Inn&	�uu��=p��'��A#���޹ �ߵ��>��C���-
��P���aY
����u	�ý>af/�2uJt��T/�+z0�(�h�0<M� 
�R5`#;m�����l�Ã����u�)�~A�W�pH1P0���7������ܒ��l4�ȉ'ɂ�y0sL(Q�9 j���`�w1���A��cCޘ�t�ĵ��L�92�;��H� Cl�v�z`�E��2>>�p�M�ݕ��������G�j'&�s�����X_�y]ll��d�Cl�F���W=�!h��5.��!%T�����po�i���|�x��(,�e��`.(}`"��Ҍ!Q���E���b�&�#C��^r�KYk��*��6�u��Id8�Ğ>��s[{ۥ���p�JG�O6���yGc�.T�	n�f�M�����4XeA� ,l�ƖEx^�;~��oTl�#:PJ�8��,��u��8���M}_VV��e/����WtK&���ŉ������v}�ľ}_�Í�@I}�%���ax.@ ��Wrb� Cl���ѽ�ic��������,GdHTuu%��������ZQ���R��TZ��l�J\�Z�����=r<�G�#j�3���!�;m��@a�'��5�"P =|�9p8�8#_:�;����2>��TLS~Q�#�հte�G�ō���L������>������1uu��{(����x��%�r�aL�F��:�gĵ�x.�ЎE���	�����z��c�1�o�/�{t}�o*��%
�,��]�.�������O,�� s�Kw�����a�#��j�@�{��H��4�6
� �w�E���.�C8%˲2JC'�GEEu�?RV\	�Q+�é��i[m�X��D�����/���2���Q^�)�'��	V@k�7�"~4޼$"P45��fx��N���K���'C�.tD���J ��[X\�DeyͿ���s�(���`����7���b˗���B⮩��z=|ɟ( 6
��c���p"P�$�dHm�R�	����ׂ-�@x����p������r����8@	���).���O�|����V�n�^ofn���:@21e��)�*���Q����>釱";S[^���̘�sP�Ņ$<<�����W55@�VV��u'���o:z��/>�����#'O��N9�1袙��VEХ#�Df�|>q1#J! `���:�wO���C�ו�*�����܃��bgdddS^^�/��ׯ�1�4��	��(۽���w�� 10 �455�T0���zc>������`��N����u�Ui-��c6P*�:��x�Y.����U�z��������'7l�S��c@|���G����{睝�<�|���)dnv���Q���1�X�����'�U��
@ 7Ți54
�BƎ}SP���'�<I���S��v�1��� �n?�a|lt�qӅ��|��+%���E��O��=�ӟ�-�/	���5qlb�u�Jq/Q��E�-7��>�m�0+lx��g��+(�Л�?(ګ%$22���v����M]7�|�S_|PE��\�
ؽ���?�٣/��͎0�Hm�~O�<�f�h�����-��.`\�!����U5f��&AO^����Up���(:IC���{����ߝ����W<���^���ǟ�uQaY�N�'Ǐ���r�1gZ�H�� ���� ��ю��<�N3	*֜~n��Z��FE����\�uֆ���-[���y�s�(Ë/�㾧���֊�# U_�@&�'<��(�z(!|ЌO��q��ta��e^*Q��3x_�e���m����ƍ��q���$�:8��x���ܵ*.�>""b��~���#���_y�׬]� ���NҺ��ȣ<�q�9c�7���>��Ǡ�ϹC��K�ډ3�C�7�yT,�J�:�6�S'�~t��X]]�ΪU)#gqxLZ���l�?���{�F�k��!᤹���ͳ� �����||�vn���xgo��=,�:@��� P�c��"����
1)**"V��LoOOwZj��o}�?��T5(�@P�H��ߑ4<<|��:x0�fu���&�vA�K�  IDAT�R{�@����B�����9PH\Q�>�p��llr~N��&!!!$$8�N�_�UV^<�� �+���R<;;�ս��>X[[J�<@��.ߧ
��or��8:;E�����7�<h<-A������q;X/iRb<����B�[
�ذaL�Qd��811簹~�����{��H?C ��d�/ɃR��L@���[^�=�דy�&�\.}��@d2R�&���b|\lgFzƯ/؜���>m6w&�,��<|��ݻC ��֖%%�u�(qx �6fiy�?c<f���#zGz^X��s������T��@��Ą�����kjj^[���ᩩ�����[�;v���Ga'������*Q�� 2�«,oԽR���v	��K���ԇ-?���uÆĠ�����>s�9?/�,cc�kgffn8x�Ѝ���Ch�Ag��x���L�w�Tb[4�)y�B~�4��`/
(�����Q-2<���Z�۴y��կ���C����\X�|w�n�ݷ?w$P�淈�9�4�$ϥx�x���m;�R���c�˶����T�"�B�e�]&���޲���+J_V�P��k�������~���W��ɑ��Y>\Z��{/�N�G���Ͼ��(���X�E�"8v	��4[�bÄ�r��*���L�ݕW|���f�r���������ＳJդ��I������%�
���������9�/;�)��FU��1&�����ꮪ�|��,�%A��;��~WD8������]� Q�8������N6��w9M@ �$s�1Gu��	�c����߾7CcΤ�M���d���{3''�����A1P���!}����^z��:�!<<<�?q�7���nS��%��x��NX��u�����zrIB>����oܸ�,��.tnܸ��/��oqqq�6�P�(���ڽ_����ϚL�ё�Q������z�B�x WTO
�|˫���?x��$ƻ�OPeV�z�䢋.�es�޾ޮ믿��͛/v���Q���SU�_{ӋiikB������o�� 9�6/���{��4zՓU[x�F���nY�%�А RYY	}����������-�������GAkbGGG���^�#>>1�~�ם �W�PZxZ��Fɍ����vr⾀���У���{Q��e�1jI�\0�-ͭw�y�}%�k���sP����ơ�o�����Ā� r���3��	om�����y��B`�s��� &�n��^���{0?q��F���,hzu�����������r[[��4w&����/��ϟ��%D��T}#�����y�cɧ����p9�U�;х��M�L��N���)���&�N��P���K.��?������ZI4�54����/o���]��j�BB"<{W�!/M��^J�������Y޸��	k��(gZ5kن�TEe	,�����-'#���kSު��|PI�APpif�9�f�+oi�x��ߎ#DC�?N�2ܼD�Z�q�rR���0�T)�Z<�VRU���4t���udUD�pqq�3�����dW�б������8��G}�h4�cǎ��YoI����f}�K���J.Q��I'2�`;�!9�$!.ޜ���M�J�G�f�<*�J�����������/޻wo�ۭ"mmmdxd���A�/��K�/�+�Ug�>�z0i�Z%���(�����$'&�Y���E}�YAV����x���ãG�~��g���\�qWG��Y��r�%�Q�19)��T�0VD��M�1}��1*BbbbH~A6����+��˦�%�9/9s��qá_ޱ{��P�Ο����+}%7ؾl�ټ�� õ58��[ps�rB�_aQ.���/.-����E�����������ٵkW�������>]>�t&�B/'�2^e���tUd)bX쁪G%\2�z���K�IRB��ڌ��m�/��vl4��������[kkkW����H6=Æ�-w��$��Wt ��b��`����b��{���/-0��`9Yy�����x���~'ʪ��d�a��Z�������;vD�1�=@Q����f�&����#�@^v��f~@8P@hTQq	4��K�a����>����u���󒖖�'�{��0�Q�����4rD������m�/�(g��I�o��� �� �K+Fa�) 	cGj�U���sII�o��s��j�*E��s�������ƺ�������������������ȁ���[�w}��yS9�'Y�o)P���ڂ�HuM%�X���4���Y/����Cl���������O��_�����s8ј�f���g˗�y��H�rBY�P0{��f�Ҳb~c��h�쒋���+��G����(������7�x�)))q Q@f�X$^����UЗ=����M�FCǟ	(�(���;h$���56��暫����+^8�;���.�?���5k�$P�>(�i\jOXnI����
8����=����^$-$$���eC�g��;1p��7>��"Z�l��9ITK˩��}����'���%�C���(_ގ�zri�BF�ǣ4y�����<S]�Fy��Qc��0�RG=�^��H[��c���|��Y��GF*������Ѩ�{���O�������АH�����������Z�"0�k�]���?�'g�x��$��a�ebb<�,544����m���+�.//� ::�_ɖ'������~���w�y�/l���Q�����40�!J �}(e4������|�(_l�W��;ƻ	>�%SSt�y��c4�Y�<��Dye��l��ƚ��a�Y7�Q�n��h�d�kff����9@P���� �+7�x�x� ��(����w:`ɹ��͌�J[�9����`���;������=..�DRRz�ʩ(����VT?jmi���_	Pkt�TH��5/Q(q�ұ�.��rf�#��.N�<���ӆ�Rl4��-���ssr���g�K3>ޓaYt�^_���w��b�3���&2h�d-��A7��+r0����������L��NU��f-�@**ʈޠ������͗�*((H��D�@��3:ڿ�j��z�x�u{�|��aЖyh�����i����������ۼ3yT��|Q�0�깥�zLL�&�Xܱ���^���_��X�4A�α�'��ڵ;����V����/,K�@�b9��k�i�\����y���q(s �����2����Byy�S�E����b,����'w�|?ya�B�[��n�] /��1~���$C�/瀪��P���x�3��zP)�<���3����*Y_�d�1B��9�zCCC.�b���߾�Ύ5��&r����'��]B������(��%��J�����~�J;�`ΰ��&��Q���K�y��\�i��G�������[���O��hX�N�Q\�O:QϦFH*坾�񐛡��<�oz�b�1��p������ 44x*;;�Ś����d���b��fs�(:
Z[Z��;;2a&r}C�`s��A|�:�Q�l��k��;O+���$�*��RP=S�?jժ�ɼ���>�4spN�����h�[�P���'{�f��������z��B\��K���_n�y�?#QE�/���ǣ������H�jU�Tdd�7n�}RR�)%U�sJ���\��g~����DjiQ)�ol �!��Y4���+����	nH>���c�8S
���F��`�TE���� �{`4�Y�fs�w��?��⫫�'�w���w��s�H���d����Ϝ�NΑx�w𞜰"X�+�J�/Jb��[�y.�����D��doii��[ݴi�nS�W�b%]��[߸���5?-9�4�����!Oo��'��hr�P-qI,Ox�F�4�����,�2Y��%���<b��
�i���@��l���[����}�t=̹e��5?�;11]�:mM����p�|��\B|o�۳�m���$A����8��r���U�_��| 
��&�u�a�������n�VZZ�x��b�`�^RR����.?�V�r�hffn��������c��?|�R�S�p�F ?�K`��ha�"lh)�]ֹ���J����܋��q���NB������F�ux��s�M7m������"(
@"�$�l�{�}��͑����466���i�RU( n�>� J>q8G����O���%�9Y X�	����1y�	(���dS�`p*�U,�+���/��9�&&���;�JuE@5v7Fu�7_��������7���&'�&MMMd|�u��<>a������*�������R
)-�@�(Ps������s9<ll��@#���!&������PNNΗ���/UWoأdoE@uwwG-.Ζ�l�M�������0�ם�����w＋�8;�M�݀�	�%�C�a�X8�)�5�:�Z��ԏ�]���,ˊ@9lv�w(s�͒�7����f~~�#���^P
�A�%�*��ͮ_}�?t"lw�?`>-q'�K<���A����HZZ9���y��7�$�����A�1���d7�m��f�EC&�?ac������_,+����d����Y_����@�������������|�GA��r^��k�j7�3X`Xn�2Ж��ԨK3�qRx@pK���x��?C�nV/��'P)		J�X��6>c2E�!� �@�G���TC�3;w��v�����qcܖ{yK�,�$hL�����?�3�7��� �N~�|���>�flNdEEK�U���2��:�_�k.|"88��8q�5:�hZt�r;Z���޻;�a�e{[7M܁�C�Ğn�+�k�(Hx ���ZB(q�9R��e�p/tw4���CR?�3t{4i��o��B^~IMM�X�����5��L�I*1~~���ށ�_��aE����B�ٻC�ܘ�,��C��JP��s��6a� �=_/DI���,��q8��K�&Ⱥ���B\\�Tff�/����|$�K�"M�'�|vǻ;��p�����0@o����X�F-�Cq2�碠p1���g�%wIȤ��v��`A�
xx�������ת�+���[q@���G���ϮZXX�O6�fW
����	\��(H���� ��{*�c�wp�%�4�.��
웚�Y``iTT�TNN���5�����҇�QP=�V�28�w��;w�41>�����sޣ�M��,_�u��
��d$�AR	<��i��z�(p��Ġ� 煺^eU9����}gs������9'�@���.��b�����:�N��A6o-'I��8M�$��i��K�e؈�����*����0	 JĊ�g�Y�FE�
�h5��W~���22>]��0?�X����=��o6��0==����N_@Ɂ��1���t�4��@�E�/P�%/�(�*I�fi$/��-**��0���6������_��5k2a���.l��Iu�7���������������%�N<X>m7X��)�(t���ݦn�L8^�N䆭���Xր͕r;Yvb�@��2992��η�����S���1������Ȏ����iii��O���V\�E���>��v�岜b���e���
WMI�/g�\:�����Mcׁ�*��b=P���U6�^w�o�			 �w���bc�G�?����:|YJr�����LOO3�q�m'�A:h<&5��s�ԶP 0�==��ɣ熥�N�w�Y��M����Za䈖J�
���������뮏���Yq�kn>�t��7�87�X�������%��,m��v�3c�DC�D�μ�I$�+������y����L*�eh� �GX�.{�׿����z�S���\\\t�mSgE�`x�?����7_�ǿ�����*�����I��+_�@Q������.�Eۅ�C��v�	YV��.a��	�ˑ������@��f髪�ةRk��k^����u{g�]VPcc-�N�W�45}grr����!M��i���Ą��x���
%��&�����2�|N5�� j�t�L��u؛>g�E��z M�EF�����啥�2��b�S>�&+H�ݾ������W^��M�ӳ���A208�s�
�{_l��~�1w8ρ�!P�}��ɘ-�c���;ײ���@�
z���l�qQlذ񞨨����M\\��l}��$
z8;;;���tG�<���w\�r�A]t�\��1��Y9c�=�\��d$=�	8&�n����a $8'lti>�f��ρu{�����/���;���zzz����g�(��XO��!Dwuu_�ګ���aw�����4˒2���xă�n����-��F0{ÑJ�nb�?Ý���w��L�ဂ�}H����XKbR��6m�_�h�s�Q����:	����ƞO>����T� �-�|�aز��~O��t�����t�� H��w�+%��@� �A1�Tpll�-1)�͋/�������3P����!����l��_x�)��kaff�N�#x> �ri@[�=	�f�l�=L��3�)ߒ
��9~އm�,�*yo���m���VGmliPP�G��R�q�o^z�ƻ��9'�jllԍ�����olmi��fuD@*x~q���� 
����D �aU�IP�D���>�U��
����:e�j�6�F{H��\:��P�.���@���It�*�ZC�U�U�zMfΞ��(E3��(	 ���ڒ{��"��׮�����&��Q�|v�3�^Z2�6� ;��l�4N�Ap@�p�.<��HY�@������>����&�� 
���v�?M��CI�U�hU��V�"bՓk�$(�$^�ɳ����x��(^
z�Z��A����4�b����|��4U�-�E��,&��͛��|��<la��8Xw=�9759�r6s�aO��HYw��j�e��\x%|258x�DUY,�%g�R�db��'x�큒'j��mY�����=�,%&�\�F�)mU �oA(`�r8�&�C�#5��@%����ڇܥ+�d27��I�P3׮����??4�� Rn�KˏB�MnR���F Q���>����#��(��2�G:�y� �`��	�G.��n�B�ŽH8wܵ�\'����t:��I��������''V��j?����OWޯ^J%6664�X<_�KIzD%@&��DT�9�R����i�T���%��pha&�O���<>����r qP=.t]wJ��27w������_�J=������7���ҽ���=��ƹ'8�}
#��I&Rp����E)���q��s.TU�\�s]�3�8������TQo�U۶��i�Z�2J�p]��:�,��A������[�nxg�N����G�M�=�uٶ}Y=)Q�o�G�/.�:�ۛ,����m�D��@���Th��F%T`��(1#Fj�:�-����P�T(>H_a��N�0�UF1$+�Jʕ��6\�0��w���|Ϭ7\�)Qf�p�0�'��!<A�T���2�2���'l�K�+���'ݰ��ӧ�EU�-/�զ{��8�Z�iB��eY��
�١]��ٻ�0��/�0��<�'Նs���q��h/����y�T�c��)u���U�a�'�o�}ȃ! Ÿg�OL��0ٗ��/��S�P{�T��Dl֑��@� ��߷û6�    IEND�B`�PK   ���X��Y9-  �-  /   images/4fde46ef-4620-45fe-a6b4-d27a85e18129.png�wUW�-�.��]�3�ˠ���w�P��ݝ�"�ݵ�S��a��y�9Y+ٹIr�����*��B��� /�M�_�_TM�b��]���AAa�ϡ�Y0H�����%�|�.Q���ӏ�!�W�����XH��d��P�p�|la�!Ss����ۄ���:^ۥf=/��;�?>_�i��FK�CC�EA>��J�Y��$��׷?	>ia#��ix>Q����z����	1q�������Z�� ����Ӷrð�dy��'
Q�j&��	�*�Y�L�ⵤ�E_A�(�٣��ELz�F��h@ڹ>ʻ�\*ʅ��P�5�-�/�j\~i�-�vu�mrq1Qۢɨ#��&��̆Ɠ�G�9����mty�y�x�Ϯ����e:���U��.�2���P��a~-*��X��r�yTi����!�T�#���7C�^Uh�;r�� ������e���n��0&-c�"�5�y�_ /�P����6�j�ڸ,�]}$���)�����" �"p+�%ұ��<���}Uh�a�ĩ���C�t��'����#7Õ�Z�1!O���U�S���z��J�b��~q�:���Y)��;w��y����,�J��h_�m'W{�E�+�Y}�]8>�,p|7�+�"z�õ��#����-�����M�ԫa���Ph{Ji�s	�\ޤE�/V��	��y#F�]O��c���}-�s�.\�{�&k�?]���0A��4�J0!~����C�X	`x8��c��Ĥ�r�"e������G�^2����ێ��+�vʫZ���j��ɀ�	8�������m�L��{C2ء�I�9ɖh�m��е��`RBI�,J�|��4�Uc�jX�jJ*�Jo�LB��o����	?9q��"�X*T��;+*���=}�5��td����ͅPl4��=��sM�b �L�j�~���VT�����~y�F���1U��M�դ<��#ZaHQ�&9☞�f�g&�ܰ��Lx@�]�$_'G=Q��Y
EEe.�h�pΝ�P�业>-]8?��T5:琺l�k�0�{O��X�P�?��'�݈�)�1����������߇/�_bR;I2ӳԭ ���W8�,�,&���B�ܬ�r���̯��H��j��d��n!jIn�������c�g�o�N2<%^��5C�L��l�m�N�OB�ۮ��<j��?��Q�I��f�!��R ٤�,���8ɻ�Z��yHa~����4˿R2��խ�$��!�a�Bevq�_,ʁ�_=o&/�gqK�A-~�����'�D��'�s׃��bR�M�D6ß��t�>���� ��i&����UN�lʺ�[��7���.Ջt��w9s"s���:Q[`�-��xR���M��	��ǘ��U>1�d���8��R
�ާl�4j`�eW���6x�����(qV䩄#|�����q�gu|�ñ�w��[�N2����IWќN5̮>�+~N7-Wm��jr�m��˱���[���mX1�F��S��d�/�{ss�G�k9���ZF��Х)%h������~V�*��L*����~QV�����	V�,�9H�c�x�~üG�Ϗ:=,���;��ٸ�KСs���5�+�4����ԑ=j�2+2=r�ur�VTZx�������Ĩ�_��%����2�X[l���Fto�]��ZE�*O$��X8<h�r��l��G� �w���Y���`�hQ% �u��E�*b�Ճ����F�2�� ���.l�%�]C�4��1�Ha��M��%6��AEE�Hv�!��NS��tz�u�?�s�7-D�2ųYHǥŌW�E���ٶ����E�~��x�� a�Y"�����v~?�Z"Y�%�!h��<0?Ϧ�iJz-��}GD�d5�؁=B��\C0�	���]��-������d	��#=R����>G{kIM�2�A�R9@"�1̠�$�UbA�AZ�H:SF
�q{%�*}��Lx�%S b�㿍S ��II�,��'��h���ٙT��J{�v0{��2$(�7(����4���GJU<w�� ��{#�	�NDH7�9_΋��n�Pr�6/R�> 
+N�t&����s�n`�0Z���^ٕ4D�AWm]8��7=*�>�t������u�Q�^
Q�2[�"F��1Y���#6Y3&���&+����/)���tFU��y�?_��X��La�.���R��^����Z���2�by��"���.�xj�����^�~��f��F��lW�e�2`�3_.�Z*f\��ifn��Xu���R�?�v�P+���]_0E�.:/���Phe)4a��W���þ���ıh�e��=-� �Oha�2Z]Hr*HB����{���OF����[lQ���1����j���|>m�֘��ۢ���_�p8��xnn�A}�/X�&�Z	�CRG�uV%�!/@\.u�d�Z:�Ϙр-gH:g�8N�3��Ÿ_��A���OF��bj[Կ��i��I�[۪(2F�@����`����O{�ķa��/7��p��s����x�����%���'Pg��
&���W���<A��ij���'z'��9���bN@�Z����y#®M��iW[Ţ���7�6T����4��ȁM�g~)1�Wb�W�Y�))b�J ����k�p>Viϵ�όC�~P��ԌW0�����`��V���Q�����!b��L$����Z3������+�}F��Ǫjʃe'a���o�����W�-XtJ��~�``��73	E���ٲ/ϣ�����)pv��K���	����,�H�h!Ҧ>�c!�v�R�b�n������2�Ş��2�~���v-��5�HX;�]�%ΔG������ǃ�!�gB:��r,�`HRI�����Jr��G��� ��Ĝ!
.�b��� �zT�����4[E0���)�<�5�H]xᰏ��,�1bz"�ˇ������T�v�qH���4q-� �V�J4�BS�:GE�\Ƙ�m���0m(
.0g�<�"V�o����;�����Sj%��QZ��?q��?�ȞԁDlU��\��W���X��b��~y��̲�-���&�U�貵�fǅu��g���}�!Z�����TwRn��('0�7�K>�J�R�BRw��k2�:���Yi�B{5�������OI�x��p�h�ſF����$�S�f���a���X嶈0��x8烵�^����;�7�������Y� u��<��9F[�zo�Y!��l*�Z���9t:���%���^~�J��W�1s\B.�6�
���4��\&�K�=+&H��I&B��bu�s�y�g���ݓfi�X%xIۭ�m{n�� w$y�3PH�;�UnD CJr��:g�C�IS3�L�@�ʃN����)����t�<��Θ�����A����
)�sʖ�=�KӭU���k��u��w�o�q�`�N�Έ�:�`!�<U^�1�˨�����+�2��`�QE-�>��$�z<��}�7{�
V����e��xsz�!':@� �������Q��!�믔�3�5����U�ӥ<���Z6�aۥ�!�/M��[]�	-W@U�2�Y��>����U�rЉB�4��5J����uq5�n�_�Xn�ܝ���[��Oa:��7n*S�>`��:���2�����x.��u�񹠠n�1��m�-1�b,t`5Y*3H�i�O�wҐ��y_Wf���[<�\�$�������;�����Q�C!E�58JC��|3�PL�E�F�ٳ�.��R��h��ħ+<W�A�i�<��FyH*���%�j�'�r��Oib��=S��\���_T �w�'��dP-H�(IhO�ݼu��С��.�Ө[��k��x6؟���vK��?���axebu�/�{`;@r��5n3���8�ea�p�.�4�N+n��P���E�ܩ���́�4%�2�&��0q؛�\z��u#GČ��`FW6��G�>�a�W/�ga�)oq�e9��Ѩ�*��Psm�s��~��@V^۱.��q�� �IYa�?�\���v��A{ؤ0�������L�c���[��ٕ~9xm>�g؉n�$�&�&������- ��ʟ�uć���8�t�\����Ǧ؋`&v [��'ۛ�Tk��dJ}��P�Pd�zi�R��+e@CIZ�wmN�J�5��NFꍚ3v�}]��r8=W����5#�b&~�`�oM�Oh�G�G%br@�B+z~��Mp�� }! 甖G*Y�wh5�JĘ�X��Z��E�9J͏Ө6�x�d?�RÒ�7f�xv��"i�1dTW�Ƙ�6� � 2k�:zi��u��@�)r�gT������Pp8.V�׽0:N˯B��N1��-��W�ߕ�&�Ò%�@A�KB+	H�~�_WX�S*�ػ��l��t�M�X�*c���N���{�u���Ky����^�f���T�e�R1u�#Q�呬�YŤEo��Mg���W���5��3*��2>�s�R\'y��FW��Ra-�Smf�������	�����g`E��E��o�m:.<K�Nz|su� q��꘱�MXy�^_�B��G��)��z��g9��m�z��������T���5�&a��3J�E��3�V�d灪�x��{?���o@|w��G�{0j_�����☍Bfb�_�2�@������)��Oo�'�Ik�oR�5�@$]�i��,�K�l��L��r�E�Dp8��UQ��(��Y�,e��'`ן���׺�^?�e0ต:�TZ��(���]�iK���N-��¿I8������z�S��'��H�y��&\8�"N���ft#�2H$ Э�({�Om�OY�Ciξ3q�Ӥ��	C�(����}�M/�v���G�8�p�"X���׶�������=�Ҧ���m�R��p+�|���qu�}{(�(S[��m��J��Ɠ9�~9�н��3>�{e��CkQx��t�n��F��n�'�h��
 ��l�W��.��|jE�I�8��"��d}F��K�K�ʗ:L�K#>`��{'����n�j�Y,��2~��.fL��[K�|q�m�&a�����!�7�ؿYzq��w���u�XFfFw�-��	�����<l�z�#=Ô)W�#*�.F�M�5��ؽ�.R��������{���1H�]�t��m�d�
| O�����*�s�tWp�	b�����9D��f�a[�M��[����wg�|D	�9L��\�ՙO���xRqGFF��0DC|� �|ۭ�Ծ��s�j�QI֖��o�Ԫ�ѥ�".J��7��J��76������Hǂ��/E��֎���O-2��C��EH�\��[gҿ�cB���Չ�����5gn��8{B��������kFn���ių�0�<;�y�HBT!n���7i�����f�����g�b��3���s�԰������{��6�짵��A����w^6]�v�MD���w�W��h/u��ϝ�0���I����yblrL�!-���f?�}H�w�M
ѿ\�yt�1[|w��}�C��c(,��%p�꼣h�ԕ�׈��a���!�?E�Ijmʗ+�}��+V^�kiC�����Xϟ95(�O�\���񏉎Y_}l��,,��9; �̇�Z��Q�&(-��{ ��
H`J׿��:˧-~�>gׁ�ǯV4�Vy�e�k�����F�SN������5(���yS��v9�x9Y�\#�y��!��OU ,а����8����-�W�Hm�<�t�k��.'+�m��ZM䫯F+�W���E)'P�%�t�*��1�
E�m��͍���a�:T�������O�Нd�-����V�\j<�u�{�˦	�G�b���ZǷ���zI������4�ط����K3�����.��]���P�?g��'��O O�l~<��_6���;"�~S�*��礷� �-8[j��.��j���L�ǘ'4Q��x&A(���|�W*ɰH�K(r�!-��"'�qghTO=sݜ����D��J��jȮMR@�Fc�!h
�<5wKyI�i�\���>�QoQ���RB㥠7��[��k��iX
O��iʪ�G57E��ת{W��c�G�C�����L��\nUX"�k���0U%��sS(�2�
*!̌%nz��O�b²�>x,��!F�$f����İM�sl��qH��C��3,ˌW��I��w���ÔoW�L�ȓ�~�t��/	b���)�&��Xe�P��.y�l-��W3��Ldb�R��#g���`3i�Qh��<�o� )���+1&�
���F��V�&�='�S�c����j��g���h��1��-E���=��D�7ʍHDG� c3�)���OL���$�G%�C/)�v�4nK�9U�j�kL��Sp�9|�P��Ԭ�t�qB=n.����=�s��q�T,?�;�Q�F֘��,�Ց���.Ocvn�4[I^�K�u��>���vev�<H� ;���z�DuUu��-;���F�Cgu�����йlr�J�o`0�6ט�=�-�+�:+7���1.�����A��i��^����:m�ݏ;S�5���,+S2�ደ��;���ݛ�0?Ȕ�|�r�I�:�ϩ��~�jɼ�Sai!z���auקY�Ff��p
yq��R,��=�^� U�tNb� i���N��p�bs��r�"�	��5�b����V��|�T]l��No.���LIEOf/b(����ZVظ,.�9�4ξ�_ 7=I���1{��l�j�޿���z�E��ՄE�eO-t�OaP�u���7|�ǚ皚Kؖ)��n���	Ǽ���t���?�̓D�������dg�:�ꪓE���t,��B�&���^�U��n��\��9
Ѝ2(�-��S�2Xښ��y���'���⢵~�y��[�����lb�Lo�5��;�~4�����N�(�ŝ�`i��+��J#��K/<�VZ�@�vV���GG$�</E�����x����ZY���M= rъ�E��y5"s9��?=�T�P`̥�
�� i�1�$�,�َ��$ ���ӐG�ɪr���)8
��=k���rM�O�����Ϗ�s�=��a��6���g�LS���b|����]�$|��a��l��O�58�Vf���4�A���B�[X�`5����f3٠_ZU!�P���ETo���&�'y��a�a���o+=�qb��zd��*N�񥊕%�MP��޴Vf��V�n	-�'�Q�N���g���9�s��[F�{��C9p�{�s�����cZ��8�H�ֈ)�*>HTx����EXԺ]s�i�����i�27�~�����[���O�c�c����[��X���� ����W�8��b6Ig��������W<+j�A&ZY�8Ã)��^�`�ּ8aD4��[���c�c������ՏX7s�O<����9�K��=[��3p�ǺJ���^[*aT���[���-���-U�.�f�1��A��`(�G�o �%�@t���J�H�A�+���5>��G/��]l R���ɖ ��<-��[��%���Q�͢Mi�h�����~��D\�
� Ϫl�	�1�K���yA��ɋu�Yg�:�~6ө 4�tY�" �C���"8,/�|)���q6��PJ������F�����K#���f��>g��C1�-�W�y���۷��*2[o�~��z��t���t��,��;�kc%5]�xI�E�,��9��e��!r�$��|������r�G'Y���}�� 4��a�J�Gȹ�(5�zK/�Ƿ�v�G:f{�K(�Y1��O�F���U����yp�`�;^��K�j�mn��P8��-����r0��Vc�E"���K������{�U �
�|��[8  ���+l
:�&�
?KU�����֭�,C�9���,��tH�4Yf���T�gYụ�ݳ�8^�68�O+�Q�����ѳ��D�D��*�`�k�Bl�X����G'�&�|�R�Z��ʧ7 �!Ȧ4"
��D�+ͺH`�����l��(��W�?�yAB�)^���)DJ�����h��놌�T��d<B�%���OhL������w�ɞ%� �g��c��[>:��je��՚���(�[�<�b3�`��ʆ���G'��pJO�o>f�u�E�h���Pu��������ʏ6z[<�#��mh��c��� =rd�F��ڌ��<�"�!�_�n��Wl��Lt���4F����]�W�&�q��̉��}���n�����^<�3��S��2��-�~{�mENƻ�^_�����t\-<]l/�k��
"4�}���J�=��Q9i���fw���X<��ivpe��m�Og�a ����@�<}�#]F����������ʼ�觕��N�W{� ݆~���7oǅޅ�8[L��`�Ȼ���L
�+��P)$�����a�e��٬���R���[��8�|i)�SȒ�I]�<r0�=�K]�aM��{�N��v{l"�N��T���9T�ZG�l8z
jZL�\�}��" 1�.=O�]+�r��/)-����Pvm����\y!rc�?�>�w��$1�vx�yxq��t��u4ǚc�U�l->5�1�(U�o6�ah���rn���]d�|�}KǱ8o���*TN���&�G�_�k�{��vhkQEQ��*ThRA�/�@�dx0��RR��=�[.�Om��G�.<��.������C5�ݛ�hJ�Я�vl���x@��b�D���,�5٤�Y��,�� ������tR�Z#\�:2��=e���W�:�+�kצ 3hS3557*#���� "t�k���"Ȣ~=����Y"�\��xdV4�7� �o���|�#f�𞎢묂�c*�r��DUN�,���eI��l�P6�s@oҨ�?� +F�	�`�n븓����P���Iq�PwQ]DP�����U.��Ұ)9/�q���y��ׅ{35��00#�N(x��aM��"1pKk�/��w��m7~��HY�/v��#����T3��9�1���>�K+��V7ü�g%
K
��Kob���ve6Y�61��!��h�ĉ�ￂ�a7�(�/Ev�5�XfP�d��^�_��>R�Yt����y�&v|,�_V
+�?D��(o.����3;}�J^4�1P�7Z�\̄��46�J9i�Q8K�D9�E�%�qBܰ���x�m���RY%���'j��W�`%�$OƝj�}	7��:_�v��L�*���]3�Ơ�
)˾�	jz���*#(VT(�\�GQ�!�n�G�d�p�5�vMH����L�Óh�1�V�K�HWd>�V�'���Y��c��q�Wdj��D�
���jD7�p�>J�?�#���P�i��f��ވѢ��g²kꑺL�%4v=ѵ�)@���O�]2��,i�OJ�����nkSCL�������H.7�?�����G坯�u�_�O<���9���G�럋
O})��k8�Ş��^w�����Թ�\*޶��-S����V��*���mČ��ʲ+���qIy-S�����9z׍���	�󯔴���4}�]�╶����R	R�4T
�rf\7�7��U]TU�����w=���"��T�~�t��lQX��0j���Df�$�q�4�re��j����Jx�U��a�*t��b:����Ȩ�ݑ|�>w��3<٭�Z^+#�Sp,�!4��H��[�
�q����n}�X�`��z�n����m/;'g���~ٴ�+2_�u��M�X(�0��6泷>�_����k-��+[:������Y�n@���ʓf,QY<��7SS�t�^����2�<k��wmh<�	T4&2�v!�7��#�&\�f�"��\4�FM�������g�h�Ŀ_|�|�u��5B�9�Zz�_Ἲ���D��m����� ���_Wt��Kw;JF "��]���/�-�ÐE{Y��~
�}�-PV=�W{@ЮA쮸�a�Eas���*R���T�0?!m�HK�_�A�x@�L�uKdFA��˼ �Y[i����ׅ��Ӭ8ɽ�)|���M��P&�'�����7+p,s�m�[���[�h)�˿�����합{߹�z� 90�A%�wQ+*���b����K8�y���~@�O,=�9�`9@$�	����
f[�[��H�-3G����,bof+E��}�E;m"!�G�/���##�J)���N�U�Y�E	�m�ZǓi/�q�B�?U���Q6��rї�#�sd�����@G������S�Lx2����U����f	��_ń���z�����T�.P3i
�R|g�^�n���휦iJ�AN6�*5����� : +��j-)]uݜ4=C�c�� �l�*��Z8�`0t|ų�C�A��=&z�� ���}�O4�3�{����ׅQf_�'�������e��u����r�Ң(1�2��F���\&~H����O�E��5~���8Z���%�~���~��ǒ�zBV\��Gj��~��ڛ4���V���*Tv��Ҽ˒��(��ڬcC^�"���r���O��"���;�l�&Us���$��uV�0��WVe�ف��^ܟ4&���H�~)H+���\�ׅ���`��H���{:��\�
����^�)kC:M�Va�I2/�X�+/�.6�#����z8����]sj����|�����6D�cZ��Ǹ�T�i�a:�+E5����d^����a�|�a�bVzI�����*�o�}��_DA0n�j[�`�\&�4ę��|Kn�q�ș��I� ]X{&�7��a����/�?����s=�M>g	,����#������T��*���cRV�Yn�$eQי��(�C��RS��i���C��~m¸.�r@�s��-z?�g���v�A���sܾe{|�Y�����-���wV���!��^a�T�K��������+��Ɍݔ>lP0�.��%z��M���B3��|B��@��r��A�������Z��b}��=��#�����1����5������_�R����/�ߍG���41���Q����Ѐ��h�}.���t	Mޱ"_.�����Wg�Am|�-,F��_��]�|,gg����/��ecÍw��D���J��3U�78����s��P� f�p�̴U�T�EY�va����U����s�r�;�fR�M@2��:}�d��/:�4�DM�T�����gz��
�t�e����#�I}U�}b�<������bV���cdf��$u��j��Z.���/�7��|/l&�-k���d�gwm�:�6Lv��5s8+G#&qm�4�*+�K�;^�2EKB���������,Am <�[���	���	����=�����Ox�;�J�[�42c$��ݱ��~3��{�qѠBia��b��)ȨJ7H���PK   F�X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ���X�j*�o5  �5  /   images/5ca6391a-909f-49c6-8bb0-8f0a302a1c0d.png͚�S\M��qw]��!�,����X\�����w'X����l�Źy��'��0gNW�3�S�===5_�U�1�1����e4�������P�����\�^�^�rRp��pp4p
2�ڟM��SL��!o����0S7��fAk�����&5�!�Bj�p?�r�e�2���nm��5OJ�D�u:-�4O>�����$ܚߌ��Nt�^�{��o����H�9����2��Wݺ`=�狷�Y��d�@k�q�s*���і��4-p|��4-m���>����U�"�aZC'F���-ð�זwgJ�������\��2����Z����w����G滟�_k���&��E�C��K�bg��o��8c��������v�W�?X�5��J4��3�.
r�O�t�����m����=_�"J3vV(���~�E�q"��6��%`�Vd�P����d�-L. �ju:���a�଺������~^���O�E�s�rN��Hξ@�"ܧ��G,`��������L�{娎�Z�@���z���'XclLL��7BiZ,*$�;CG� Q�k0^U�/ku�y�e�Ke�]{y�˃�m%k<��>9�%���ai�Q=鶁���a�IY��m9S\���4#QAl�ǜ�.䢄~R��*�x��z�W��4��7�T8�!�gk�W��퀡ϣ�Pt�H�t���}�3u	���a�`����@�+!9P�I
� �#o��E�qf/WS���V��C)>�A̖i7��0�&!�?��|7P���u$��G�&�<[`h4��*�qp�|���a����m��>�f����b 5�7L��&KPJ��a<ܥ�>�����k��o�������jv���Qs�ba�����!����ߧ�.c��6b����)���p̏fRo�.h(�����u�&� 7���_bYYf2�-���%G���F�U�8G}`��1&������0Q�z;�x���G�&�8����o/�HيH�r���Ch�����8[�G����� �״��iH�ȣGo$t6������B�3��5>���Oo�T��z%孯�W�}��|��-���_g�=�4Q���M��>�Y�?��o���4q2���d U3����rS��� r�����!�)�z��/�K�m�J�c�j*7C�y�S"��V�n�x��dH��2>�M�9_����'r�����<~���/�c��T���C&��R�,���H#�1F�}�Z�O ��^�&���6�HT�d���g�v!Q2�޺SnE�!�g5��վ��m��䃠q�˞]��Q���W|]\���ye;�E�#ީR:bv���P�6F�T8TZ�XR����/Z�ON�!�6h�+�CR�LI�юb�'��,	r����z'Y�^��WI��O��a��g����`g���zo��-Gⲻ����>�ĳ������T˽Om����@:��ob�Ƃ�����\����<��T�G]o|(���'ݤh�:��CYJ�t���2��mH�Jk�<���I	M�|8�G#�t���k�:.��m(X��r�?�z*��C�/[\M�q�x���W��Tt�q�"����>zCY���5��9v�5B��j����>�%eS#5"�f�\����:1<��QG}w&m�k�s�7�FƢ"_p���D�9��>(p��७�W'��,x"���Bo�I:/_(��փ�t�UUo{��N�'�?�����x���U lz��Fڛ�r'��`lqjTz�?�%��A�CG�5��T���B���_���Qf�"Pw7��*fL����]�V�� ���WM����y^���,���o��=m&7_n_㚸\��Y�љ�_��1ݰ�P����ƤF���o���$�Z��J;��X�4���R�V?� 6'�����]R��a���m�݂R?PtPH�N�����Y����g�D6�/| �++͍��=��5k��=�/�����m./�n0�YM�6`ؘ��F����x��kk�|��{PN��B�����ָ9'����Z��
IL��h7}����~�� -�(|���sθ���4+�B5�/ͳ�I4v%,\��d�m��6�ш���7���)�(�&b�4����_*��H��e�������4"�uz�4��0��M��85a2���Q$�����|!�)���ǯ����w�ȏ�qy�Oy��� WF���]ii�2�ϱ�r�r��[7��k��!�i�s�/jmؔb7.�e�6(P�dE�����Kj�P}��$��`I,������,��:g�B�d�ꕾ?�,X�W�F��P��,��f�pNf�V���(��%f��=z-�MJ�8|r�j%a"A�i�z%˾�P��>�Md�ͭ.��7�=��r`��f~��c!��P��ג����k�\òԕ[�����O-�S���;u�2_ .�1��!W��]~Wf����:�J��}8"Ӱ��O��y7�<Ab�b(9�7�G-�H�ͬ9����!~B(˿1BP�M�iL�E���ЦjA����a9{e��up�ޯ���#g�z�^Gj9���}���I���5s�����Eݥb��?�y�����4nʈ�q0���חs�>!NV�_���Q��&�DXJ����O�g�Y��m��ѡX�*�o��At��u�������s�:���a���J��AVN��^S��m|�fu>��I~#ɂ�����-Z���B�$K�jZ�QC�ֺj��H�G8Ͷl
 ���4�d%	�g�Zb���~�B��������ƍ'�̱*�BzɴY[(�?����%�z�}OKK�B~QQ�ÊE2����n~�B������g��V9X�,�i��8��:Fx �k1Ti(�7@=���͵�_��;���xo��/}M��{���_�n���=9w�YwV��� �|�]�yh�}Y�����7,P�c)���!���13�w�--���o^̲)X�ܽ�6:#,G9W��$���`��@����U�{S"�]i�}�aݿry���?V�L[��>������aV�n3��8��ޕx��i*�@8ܿ�g�������lE�8#=C.�DRX�F ��K�C�_KK��.L�ڛ����ҥ`N�f_	z���S�����˸�>��!�y���	%-5x�);�O�6H����m�O�!���6�c�ZdR��Tߝi�.�;{	ȓ���4��i��}��pr�ۓvgm�KN�4�2�E~��'��`��W���|��L,Z���}GD�dV;{�)7��j��`�ȭ3�ώ�T�K$�Ɣ$>��ӷ�RFo�*	�\��)���=�j�O��L�b��˻f�3��{�\SP���}!(WH�d���Za��Q�- j��i�c"K��R)�x�TׁP���?;�J�|	؈�x'��]�X�B+�"'-w�ǄSU:-���"dڋCy��m2���U֢��R���;���|b�Q����ǘ�Q��W~I�һ^0'F$ˏR�H�D�����O�j�R�q�64��STe`T��%Ak�WM���{��$�η=�����nM�eX�@mc��X����w��c�����+MI�A���G���pv�4OL�B��DM�.oH��&���B)�f��i"�`�ؿ��+d_��?�ϒz�z���=̨�YB�=7c���~��_����$F"K�KbԷ����닔��y"$�P��3>�����e�"w��:Ӗ���'�Q4ƽQ������1�
��	���g�W��u#0�� :�{0+>�"-	4�_ns)��f����߸V�fsq_�D�|�����;��(R�"�w�5���&��;,]�$�i��	3"�9�ɛrEn��}[Ah���m'��C��,uSL��$a�Q<7>p��IQZ*wOn���/(Ō�av�[�9��Q�kl��o�����\�����|�gq���Pm3��<�o(�sΡk?̗��cD�����2�.H;��B.ЉB���N�`3C�e�Uة=� lw�IS��O0��D�CV�
�V7��Di�p���	��"�ئ}A�{��B~̱��)`��&W5ڷ��L��l2�_Jhӥ�UĿ�ϐ����[�%L��:$1���`�r!�VU�eP���=}R���D�T���9��$s,�m��Uأ�<Һ�b�;���Qfw��%k|� ��.��	/!~�I��;m��8d���k{�$;��p{�sӧ�W�E��$F�)��ֵ�;��\83�;#��q�
!b�'P
�Tw���۵�˦�`Wxb�����n�D���,d��0E>hN�[�V4�A'Z�￙t��~y�*�L]`Xef�X���؉�K�oq�,(v�d6�\D`)ژ<� =�y@w�����f�{LD��z�l��摊�$��+��.H�p����C3?�U�[��a
[�+�f�uVs�b����o��9�ʄ�N�+�-�~���%�ǻ��7-�^���)�Ι神���<�! #��"�`��J�=��A�:����p與�Ɉ�����5s��B�W���Iϭw��;,��L�C��2�e��s��[P`<6ɓ�A���'�cKQN���c͞	eAx;�s�{,��$wpJtr�q/uz���7f�i�}��0����@#I���d��n��~���G�|˖��z3+�*��o)4���`c�[ky�ȸ�F���G��s!nyu5��-�P+�2� dM���)��ڮ����G�i�����~�x�7�(�'y����2Z0�����Ob��c/t�ُ΢�et�e�ruZo�m{!��94�L��:�ᾊ��d�@�C;K�ux�t�m=�[-*������&l ���cc�o8B�9er,҅6����_�c##	o�2�Mg���zዩ�!o�a��j�ʘ@�G~�AO��bLr����a�i����N���ߞ�OBB�8�O��Z�*�S�Ux�m.�Th�-�� �A����OmT��!;߆�M^-�T��ɘ��R�Ϫ�3��B2�־�{[�-��@,hw\\�3C-Mr� �%�"��W�x�gR�32�_d�ya2?�1)����B��3�dd�B	��Hjd���TpWL+�:*�Tk\���#�&�-��7F��	�< �+�8y��b��m�A�Ζ@��y�������g&��R��� ����8 �WtC�ઊB$�$[@)�"�";�{Q��$-w.�
�w������վy�Ot-�r�S<1BK�� �1(�e�q���ⴆ�J��Y�?i������9&Z�A�k�+��KZM��Q��c��ݺ�u{����5�X �_;ܽ{��s=����hB� �uWa^�d�Q�[���w��1`�����dl)�w[�\�";��W�jQj,��2�2����灎<��ͩ���%{�x3����]&(���<ԒZ$�e�, �gz�u�L���@p_��T#�D���+ݞn�/���g^�Sl�}iDs���x魟٦m���o�k=����@�`��!�Y�:���ʋ�s�J��@|��\a�zɺ�y��	V����W�Cz��r䬰@��S�o)�y`���x��q�D8Hb F���H�.�����q�||�Ng��e�^.�ˑz�-_�J��o�ݫR�[%!������x/�w.ڡ\(�W��t��d낚b��&���d��t�b�S_�DX��Q����qJ��Y^�M`��f�����@�!�'ܷcLS�݈z�w�c�)���[b:���I�P�P�*�i�mG<��܌��B� � 8� PRt�v�h0�蘧�(M�[�t������B�ً5��2p7H�i�7�у��g3�H�{S���]|�c�S6d��9�
��W,�X�j�-N�f^SY�Z���`!��0�x�K��Ï��t�kMa���l�b, )�U��7��-Cvm����Fژ-_I �>C�/tV]:�Z�2��w�4o�g_	㌭`����� g�,M�LCn��]�UY
z*�&|Wd�J���'���}�λx�%u8	h2<��s��� E�%�\4k���Ld4Kֱh�$zϋ`��Q�>$� \"�g�O7U�����枟�ɱlpLOq�ق�X�x�9�ҡ-h�!�d�5c���;E�hC��̶�|I'�X�W�����BB-����bN�MkLY��)ge�E��e�Z]A�/�a��j���-����V�BZnV�t8�ҋ14Fѕ��wS�}`)�Ǩ��x��xx���v�͆��d���0k-��I~�9�;��C���\}zKl�
p߷��"��c�ʒ�#!�QI� ~D�	�{ݦV�d����|��c���qsy��T�j���c�K����M�]^��c���T����C>E"q*�s�{Dm�R�:ؔ����
Joxx�V��M�]���� n/.�zo��{a ��(�?�8�h�u&����k���\=�;պ��{�dNO,��@P��mu�?&cn}R��-Umo��WEiI����ң�I��Z��<�|���dƍd^0g�i��b#tʷ�zB�$�Z�0�"x��}8
'8��Iم�J��R�̘���r4������lԵm�*��CG��(:(���>zp���]��V�?J|����]?8_��y U:��N�~����2d�Qh��tP�k�8Sy�}�~������O=Q������o��؈�|�nO���:L[�[���ܽߪ�#��;3k�TBs'E������s>�����9�P�㠆��VY��[�G�<��&1��C�}�U����ͥA���%;�J"���������5A�j^���ĉ��P��3%�2t�
'�Д�ZW��%����D�/b=K"R]<V s8�|[q����&W���d�ٛ�6r�>�3���^�2ڝ�����QrUP���;����sa�S��p�ǯͷ4�F���C�(9I����L��X���v����3M4��ZR7��b�r�gG�6	����W�4���KЅ���s��qࢿx���� �� ���Nd��/��x������~Uڥ�%�Q�Ļ����:|��Z���/�݉v�^��[��u��V�m��1{�r~�fYw��X=���dm�D)nʳ6�D��H3�x����~���X��:��mW�h�< ���!�չ�Rn.&��r�jV�?��[���#3f���Lы�	~�ﵤ����DƱ���� ,���$�ِiHz@`
�6F��u�6N��e-	ͪ�,��d�3{&��J�	���\�!��[Viu�ʇ>->1Y������'�⺴��F�{Chn�Ca�����F~T��\}g�x�����}k�JRC�ח���� �;�VmUY�@�R��17R��/㍌P��D4M���ǩF�O���1�*s�ּŘZs���B�_=�у*h)�RA�i�׉k�������@T��~��RI~O�a�S���;".O��u+S�{��=w�: 'w�B>�1>�q��Y���9+�Ӥ�Q�E� B�,��UO���B<�D�D��:�G��;,&Xo�3��Q�r1޷�}PD�^��7P�D���/
�sC�l]BL�6vt�c�u��'��5jM 5�נ��@K��/YwX@�aW�� ͮ����f�XǏ����Z����Wg��!S�b�@��LprA�#<d,��,����ok����K�wX�)�]�@1d���^���;7i�.�R�X(3`{R���@+��}m=���Q�j���Ne��K�QF͌�L��V����qZ��b��8���'edؔ�P��0�\��O3�f�̖�V+|0����������j�i��d@�'�G7~Q����?�_��\�������
�R�\��yC�{���h�DN��_��v��Ĵ��W��C_���	1U�=+@[�E5�� �&U�4�s���ټb��r6�(�^�ɳN�=އk��i<��U��_����0��U��7�O��4l0'�6@b����Z���ƝUa�bE5&9IZ�8��_�![ p���X�yP�|�7�����~)�� d'�:ؘՆw�Ҷ�:�2aqO�~�n4G�Ԫ���:��1�ڐ��l:D�g!0�q��y�Fɟ�*�;�*-���>�V�>
�]�N�HW���jf{����5Q��V�9{j�$�X88����0��b�OeT3�΢��2~x�-�v����o������.l���2������<�-�������F�i�6���v�*b�q�@�}ҧ8�>��^��o��g��?�k��-�2��6��7�%5듁�&�L������+k�ǒ(�nW���5Ċ>�.�6
�Q�ݿ�8J6���(��!`S��)�����=����Y:����V��D��w��Ox���oJ��H佨)�Q�!eK]g�\��5�c�O�(�{��g�&�o��ޟ��w���~��JC��`KQ�X@��;m�9ب��
<WE�)I�P���>��;5ϻ`�b,��-�'=�ϙ��
����������V.��̌+�Up���~��y�[�5tܒ��Hg)�K0����HdK�����|z���K�8�r�$w�Hg���B� �L0��f�>�R��9F�3�2���J��<}>��Pܾ!;sZ������I�*��ٍ������;����@�~$A�S=?H�.Ƽ�4����$��|W�xT^�X�r>�a�7��U�X��b߿Q�c����L�t��mh��jI��-��X2g�c`�^B763��V��D?x�c�"6C�����^vI~�;�8\����IƗ�E�T��D)���n��`]$GC��q�W63\�*N��C��V�/̺�fuK.�QO���Nԇ���U^4���<���x�Xd��S�A�ZZ� ~S�&KbfCv���n��=z�^3#�A\Ɔ�е�{=N��A�f�?�~�����ɝ�IdV�̲�>4���T��0�O���7ɔ �ю�����H�eC�J��`"�)��f�n����ڈ\�y�O�
�a&&�9��s��玕kN�	|N&���ϛZ�|��Μ��\c�,;-��Kg
j���n,����▼�{#2P�bt#��+u<b0`�P�ZҶt����}����n�q(���������c���i:o1P�zt�]�Tփ���˪ �5����HO�d|Q�کlUO^�v�ۮ��{;�AI��#�Y�|�����bcP ��^o�R����;�b#�eyo���Ѻr��z��0!|�ܣ0�{���%���l��5J��`��q3�;���?�깓u�4{�A<e'�����5w������!����YV��U�p/�8�N���O��K����Ŏ�Y��ˇ��2e1��F	��NV�'8<1���p��e����;�B�-9i$:����pv��cp9���6h�:?BS�T��xZ� �3k���w���=m�\������9�d�Ǫ�/V�l~����̔�l�|�c�.T�=4Q�+1���e�L�@�^V�b"�s;M`�b��'�J^��֫��
e�@7[����/��'p)���m�{J���U�q[x޷.�����X�����`�d�(EHs�\<�=[��B�֑�VLL���P"E����8���=��Й%\-AK1�ϛB^�[��09�q�/5�1�4ҒK��I��{���
9n.:�qY�񌇫��e�}��Eү����(�WC(o���;���I�?�Y��w|�;(�3���g���$`�pA:��D�p���Q���Q.NB���H��:j�R����I�7��v��V�A�̹�{��j��2��c2��Y�D�6��T�
D�W4w<�2�t��|3���_Mލ��-d��ϡE�R�����3������Ƙ ��x�m�:Wc�)�e���D�I���GFJd�����DI�Q�O�j������*0&}�1-t�T4i7�9�)ϭ����&�`��odq~u^����$6�*,1��;��x?\D2Sm�H�诮��	�UPJxc��l�sB��)���������n�?]�}T��$��M���;�QS]�u4Yl��@Z����14	�V.QR9zDH0"!�5��9�L�n!�$g��>}��14Tm�8NfZ��O��d����� ���'�(�l�/�fL#���P��B�QWR�<�id���)<,n?��X&��Ox,�xv�
��L
�]�J*}�g�/���
"g�MKS���~n�NSoB�=9�`iҳ��Ӿ��+˞+��T�F=�x,:�@����m���/����hq,j�аsQ<j��4������Rlޚ�Y+E��$@��(�o3�zR�$�	���gѝW���Ӝ��ِ�(x��(����`��.��X1q)]y��
�2� $M�46�KAb��G:���L�[��d�&ʡ1���k�����c�zv	�����_�"n������ċ��b�fu�Zں�K�Bc�%��θ6tC��S��\HD������x��v: �wf�����p������5'[�-G��d/$]�P��0�� �ڊZ�\��L,I3���dU�'E��m$�&9��Y�X�a�>�ރړd~���DJD�*7u럀ܐg3�abJ������l�����{wt�)�5Y�[^ߺ-��o^�{��^�)��3�����"1�x��4��G,t�+��_c�F�hX
v��~LQ���V�Y�����.ӈ�#��=|�����[�&�/7���~>�~C�INl�4�\�xƫ$V6���E*�%Sh��3^e?���?O��
57@hO������SoG]�9�Ƨ���:�����Z��Іj#S��o�cm�>��/����}��ȶ��Qʭ&ӣ������2W%0�� q� ���x��V����f���_UNN��Ж��D_/#��c�MP���99GYV(��Q�XI5AH�A-�����L��[�QƦX�;It�V񫝒�K��#��6h�p>R`��?���������zgc���7q���@E�k�[&���K����e	�6��M|�81,u?xQ��1�����V�����jAf��Gdo���b�'�(7Et���-�q)ԭ.t.j���F�UF���wɺ37�h1ׇ���K�ܫ��$k��yf;����	G���	�����p��/���2E���즊�����E�aH����	�x��)�\?9)���+�HSZ{�ǧ�����'�o-d$�F�[�ϱ�
��������qe+=v��2�	�(�lw���ɯ5��oe�o횚��d旸ڳ��)	�����vm 5&I���:%�|�P�tS%�bJ]A9�����}WU��f|F��H�����	�_�g�q3�d�s�"R�D�9���������6P�1�B}�������\�.��g�9�0�0Ѹ�h�c�R��X[=+<*�o���x� J��[	�Yyֆe?�@�H<��l��H���&
x����������#�_ɚ�2ّ�"%�7,;j����%i:�5w����E�}+��O��KY�Z�̏Z��V>��4ݭ����Y�/�G#�{���Q�����g��9R�Qd�e�T�I��a�Q����G���1e��.tr�ǀ��p������)�l��Y���t$2>�
�m���o,��H�F�RoC�}7gn���$�����=�����^M�ˤM⧻w.m�yl@���+��"���OK5T/R�VOq~��\��+0��e�tW:y�]_]-����S�����-ǌ�X� 4n��` l�1���vA�~�)��,R���5���Y�ӪY!;�v%����1q��fr���W��uDeE���DU,��.OR^<߻n��$OyQ��H�Z��q������� ��n����0�^յ���=�FҶ�ms��a�5(�:T�U�/@���^iU�u�� ���G�0�ƭF2��Ѯr�,�WF���L�h ��-wt�����lO�ƔԾe=� *��\�+O
>���M]�9ܬ��دb��>Kh-`��
�=j<�[��]g������,�j�I�)S)��p'J��:H�ڻѫ����b�� z�plJ�ڪE&�w��u��� r�������XcB�u�����e���2�C�b�O��� ���3/L��쌃���o"��@����g?w�|�A.�\.����o�TR�WD}���f�Q�"�O�����;e�w� ���1�b�5QG	++��zy��O��ϰ ��]��(�ʭ;��ý�-�=/"w�7B0���kK��CQ��jP�����������KX��7+����f�n�䉁?��Ʒ�N|���� �-F�),�|Ѳ��.��I���t����5�_x��P=r꘽y+x)��fS��X�8a�a�ߞT��e��Q�č-Q(R�#FA� �qW+1�ö�Y��ō�it��c����[	��Gjd��ʃ����MS3�P���=@��v�ɋ���qa�iI�E�A�{vv$޴�X��B�4���-�>a^��e��<<����
���=�_��3Q+�?8�v?@��i��E���Z�,v��|9��t9\˂A�X8�%�D�Ǝ���Č�^�;�'�Ufy(�i�J�����O]��6�)#�'M+	U^�2Rß1�=MW���V�X�H�ϥ/=}ǯs�u�Y MBЩ�Y�Lے[W\_Bs�PZ]y���|�%8�e.�R��(�����n���^���b���G4n�	B/9�����8���������$�=p^>����������yͤ'�����ӳz蘘&9[�Z"���?P�)�����Ȝï�}���ߚ/O�|,:�@g�_�CUF��c�;�J�����{��Ԡ�!�_�u/7�v�k'=o��e��c�Yߩ�]����t\!ҭ���N�
���.�$�`3f����T},Ƿ�����lA��Jd�lD��`�i��0i���;f�b��D���zZ�&:;��,�����_�Zח�t_[vj��}�K�@����--���I�#���B�����F��:�^���A��d���&� ��K�_%�?��E�T?�	h�ީE{<C�._���!�c���P�K��������u������^��1=b7� (��6�%���k-����
�*��j�T''J�c���ʶ=��������/_?��]�RO]5�[<��|UUs��?�n�e���ۛ�e����9)řJ��?��7�^y��0�|M���a-j��f.ae*d~��߯�e��CgטK�x��:}��J㥣���b��\�]��7a_��/)�lꚂ2�:��H �Qg'c"�ԡ$�#��շ���U�;�N�߰#��}�|+���"��견Q�Dv�M9$�L�U��!�+�nz�;����������A�f, �u��\����M�\Y���-�~�8���Q�W;��'2�=ǣRA��mX�C���!o�jfH��op�YU�)���PK   ��X7_DW�  |�  /   images/649de870-1a94-4537-ac6f-7e62814b65a9.png�wcs%\llۘ�6N2�m���N&�Ķ��ub'�Ɖ����7ܪ���k���V��(eE)d000diqU00p���p0�����<�m���:n``(C���i(�``�2��r.z`���\h����R�8&���L =�aX@#&�\#0���Ɛ��;Bg2o�$$<L��ؾf�"�����qۇ<,�^f���j[K'y@V��g�^��j/�Q���~�EP���]�r�O�M�r%D3�����.�h0,��-���}�]�U��&�Y���^d�����uaA���#��k�/�����I ��B3����Ru|/X'y�D㉷دDe��U��ս��AX����s�������cjj���Ss�v�:�
�Jh�+�AG�ɨ�]]�Ns��	������.�����o�J���I�XjD���M:Z4��� �IX=��䄇h��R��1���8��w��I|���}�;��n��(1�M��w�Aa8��������^��JZYͯ�7��8I�ܻ���Mk݁����R��YD��rRϗ���������z.�/B����}C��#���w�QE"���fJ-��w..qw�5�󞛷����R���:��^�$���Ô%������[~�:������X(�v��9�}�|�'��=|ڦ4/Xsi���\z��b��\��|�$��M6i��l=?z=F��:����wި������r�>a����x�
�씢��/(�܊6��{ 	<@��7u�8{��6q5}�Gd�~�U"����}&龙`�E�.���~}x�o��{\��A*xss�q�����l�ܦg�oå?����q�a')��MWO)�����U�h0W�	�t�����)���q���W��q�v��+x٣OL�4)��������E}�n�qg���MD��J���[������9Uo�����׮���u8[��Եw����g����<��5�Z����h���)�h���'��"�%F�DvaX�y����s4"��E���Z���o=�-�y%>�zux+���$w�U�Z6Z���Y��)�x�N���.�^�7�8T�!�Zx������mݕj,[�:>*�켳tO�$R=W��A,���x�h�G�p8E��vz��s�l� RO��N��a�#GS��	!W&�
w�E��P�b��p=����W��M����e��ѐ�:}�7t����P��j-���r�F|��C�*�oҾۏ���.���pY��� ���/{������@��E�ɴ�Օ��O�n4�9m��ę�wr<_�1�(����{<W@�^���VW�=h�]���M�v�Aa��x���V����U�����^�2�Km��f���{����Q%?cs)
�o�E�	����~F�CL~���y�N(������o���[��@�b&!-�2���V���A@|��`��k��y��d��O�+~I�D)�����p�Ta�U ����z��\�*���pV4#glxкRz�g't]����_=T����}x�8�٣F��`1c�ܸ�o���F�c�^n�I���@��k>pPڿ�I��ᘣV&�#2���h�؆
8/L��i�mM	�L.G����<6
C¨��Ca�Z�Y�3 t1=2�2���X������a�3���rOq�>>������l�#����S����<�D��z�,Ֆ��,���V��
~���	g<��ջp6�����~�W�"�����8 ��}��@#�Μ`��|211	����!T��hk}���?��w�(</�52��<��0�s�,P���@w~<Ku� UWW�OZ�
NͰ̙�5��h� :>����U=�'~,��;�g/�/B�y�q�a�
��ph�Ϋ{�P���b�]�sCX�K��X6�@YM��k��~h��<�|A����G�5�=���E�`�������h*Shxn%l������H��*����S�V�!�) B������p���t�P�_�`��yU����ꭷR'?խ7�
8�.)R��)E�����Nm��J�+�yF�Ќ>�7Y���i0��۱��Q�;t�������s�N[]^��9: �(4F�$(�ǈ�c�|3#�i�҅��3D|��To�b���|�sp@O����M�8��v�G@9�4|�����ܲ����L�L��t`|��(�$�����ܨJD8-n��1�S����w�mC9'޺��0K~���	e���3��L��p�=Z���UY�Ξ���]W�%eC���w]k��/bz����Pm�2T�.h��0���3�ꠀh�D�/R o��6EƪD%�v~�?�G��v�������g�� ?�l@���_�1�gNsY�*҉�ȏ�\/�Ҽ���j8_J�_�|E:����B�����X\[}�i��Ȃd̈́
��qh�YX�@�N]��x�j(yx���@Ӗ��)d��D��6F.0�a���BaAp�𲨨q9��̅H2d��'Ui&�V��f�ҒՉ�(���W���/@�Ϫ?�fڶ���,i��������k+.��O���eтQD<kX����1د�* CX�W()������#��Ofo���!���q!�1�4�#�^H�ڃV��f Q������Q�`��BUD���5u.?A�w�6`W��!�ޭ׏�s^~^r"��p��̄�is�j���a��[�%�1,�P-W�)4�[wR����Z��+A�bOA��pao�z�$j^�!R�u1�E��4�>��Jk�&�G�c.��8A����\�J�N?
j�$�uƝ�DE�8D��0϶@-��n�]��-L:�����n^�H̘X�zMY��`�A4;R�3u�78';x�'/�N�_���
�UY.�o۹X�����{�^����:�?�����ŋ�ZB]��٧Ɓz��j���d1�H}D;�]�� �HT�Ϟ�:�센���`����(�Ą�ߑ�/��U]wK�d]X� 8M��P#8������ľ�U:)��6��2*�� i�Cpr���� %$����\X�O��`#������j��H���>ذ��<�Ԙ��ZJ�;ߕI�4�'E�ۨ2�J��Ӳ�������C�*���[��{'���2��W� ���`��)Q��r�h��VPnP>^��TP��1'�-ei8tp���N0��U���C�	ő[��e�h� G��Y�ZM�f=I-e?�+Sr�����0 m�X�fOD1�U+�J�E�����Z�n�T���ұ� g�>�#I^eZ�ed-j#_��y �7M��@�g�2����*'Ii��}�Z@{���?�A_ �/m�XV"�@��[A{,���X���R:��N��r)ؒ<����ڈ[�!-�&M�c�Ԣ?g��ŀu3/K�b�y�-X��T-Ƀ!	AD�.̬��Ƞi��<%jk��&]2�3Y� F�uv���'b�H���§�D�zP�1G#��Z���1���FձA� ڔAm��}@�g�9B�M�@`2���fO:|�BVQb��3����iZ��|Z�=R]���$�.��Eaz�U�*���V6s.1/�*��w���U��4�Rƙ��t���v�f�F�g0Oh�B~�|Q��Dɽ��+&���4k�۬�E�o���11�i�(�N{pf�A����:�=�5f9��z���Ũ�����@pQQ$���E�^D�ݔ27�gЭ(��绲�I%��nڗN~,k��ը2ǚ�����È[.��jH���Y�_�ED������u�A7��_����Lࠦ�x���o7.U�.�_?!XO�8I���@3�"��bM���*��g�7�Ď~�&�Ũ��DIN=��X<9���v�	�����9$�I��8eQy�Q^v0["��$"?�^�3{�3��voH59l��nLD�^t3'",:�T�ƫ���:h��	����U�i�[p"\��ɞ�]&�g����F���4�H\[~��M,:z���j3���$h�%r�����X��U�*���$y����#�E�xeD����4/V�_Q^�O������('܃��	Y>%�+WK�Yv���r��Ę��N�#�X␙��${ߐ�� �z�>��)v���gf��NJ|�� �.r:�p���mZ�a	�;+3.�d�� ؆1��U�o�*E"TyҬY!��dc/�T�p!��Qg�!"��T�p�^IZ�V]dx:\Kf���9g^A�e��P�D�Io6���|���z��2	,�x#v�暄�1������h��9|�"x�0q5v��*&O�Ѳ4w\/
��_�PjYa�9�S�
�[���훤�HKࠡ�T)�(QZ%��ZPe���@�	��Z�m���݃�U	��MU������dj������@�	��U#�fBg�ȺyV�0���v/V��1��N���F��s�2��'��YG�L��� �F�
�Q@�J/LT�e���p�;�1��%���S[������S�6G��q��i*���[3+c��8��4��"u�f1�V}���6(�M�%�&�6�fY��;��|�O�'Y#k�2ôE��P)���<��:z�(���:D�K�	�v=�`/s8����C��_���Jsœ��&�zP�Q�k�>J'c�K,<,j�:�2i�ݗ�0�»�$=HDRu�R`rE%���|E�4$�MSF��CKQ-�!���#*��U�M�j��|�����a�Y��p���$<ƹ�U�Fk)�\\�3�n��%�?�2�%���\&�:�9�o��k��*	+���d�qZ�مA���JE?ح�Uz$z}�Epq)�2�k�[���j������e�R`(��hƳ��y�+;�����N�k����G��@����у\�]'"��&��6���$�t"�f�C���~���0��B���-c����Y]�����_��ۻ�y�Gc-4��G��is�j�R�Pn����c��~�ݪ	�|�y��9Q���_
���$�s��5+�z#�WI�L}�k�!􉏸خ]jh����w	��߆L�ɒ:%ixTC�d��$��K�G�xo��l���`�UoRBS�[!�Ê�?�Z0�R��Ӵ1ܑ#��-S^�+��y@�i�������\��Hl6Wa�zǺT�-���F���F��8�lk�L��CwS�� V���1�G�����^dy�fȒ�ӋK������YOz��{�������/�$����s�J5�$f�%�F3X�3@:��b냿���ҕmѨ�V!�\�i�Y��/9��)3��W�-ؤ�qn!~Ğ�0~��*�q���Ҭ{���{���M1���QL�h!��N���Wu0!��م�@hHvӠ�9��Y�f�f��1���A��G�>G�AG��0|_����#C�@�$��۰�XޅL/^y��� ��g�s�Z�Ч�\��C��,k�;���V5R�4B_���0f���zGMʻ�@	�Ȋ� i����ƛ�T��ig�,��2�w��ĭ������W� ��j!\�t.���^[Ĕ�C�1>jZ��:�K��w�	!gz�%މ�݄;I澩��Z��X6��Y���|�6�|�Z_��^�	���&y�D%�yw��CM;I��n�XC�����E2��,�B�pH{2�H}1�
ƹ�R��_Q�$o(�co�ciK+9��.êp���Ѓ<iUb�:V&C=��,��z77�sbLs
}��(y]����d��3���ċ�Ĳ4��ػ��6c���N�j�d#� � �%k�O�bFe<��ζ��)��I)ѽg�sx?�0���^�Ʈ{2����S����;� ��P��d�u��s����G\@�Vm���2 a�o��Ď�ٛ=�� '\�>�O�}�i�/�3g3fJ/ӊ�ou!�cE\�͛5��th��E��3�R��!"���1��aM�8���G�z���p�no]����i �d�Y洌�:u~+�$���� 3�"irs=ǯ�Zz�� �CA�Ck�+�XN2$�/SU��@�`��.=-�'��1̴ 5Eg�Z��mC�>�@S�+�M�kL�H��4��#$ڋ�����%*wb�zJ[��4�K6{�zY(��G�7Uo�`@�=l�QD����l�\	�S5k�L
��*�v��].���)�e��?���"�}X9S��s4'��c�I~=��1��x8�5���rVJ�5��>n)�Cc�Y���5̲�.��س����Ik��� �S�ğv�C1l�j}ot��4��I���мD����N��,���Q��_����&������Ѩ��3L�a��Y��td냣���ᮼJ��LjVh7Wo�Mm'woD��Ǥ���f)��͗خ��H�����yY>�o��`�bL�{�Yqb�2�B��H����Eݰa��>$�$x*�>��8�os�:�u�a�U]@�'��4>�(۔FsC����K�jf�Z������Q�%���c5!�P��J�͡W�ϼt^��.̓ Dz�5�cr�>�Fu�X���#�C]�Kw�tFC��^���վ秗���L5��G�d�:{3$Դ�У�3ȓ�2��T��/���o���@y�y��ȳ]�)6a���r��a�tyC���%6n���\��C.�̥Ywa�ٝ3��f;-Dˉô��f�O'��s	o�.Nl�Nq:p.Y'w��62Ū��_��)�����o�ߡo�n���(U�;%�ht�[�2��G�s��N��.sҪ�����ө����tOn��eC��s`��c�.�o(Թ��&�8���0�ƷdO8�
I���&�
�t����1᤭�&�F,98�CNV=G�c�%�!���2y��,�Ե��Kek�]��e���Fy3m3�� �N�lG�Y��+��5<��v�m�§���}쾇D���]	52��	Qz�ϦC�fh���h�V�֕J��H:W��Ͷ�7�Q��%�����=T~gw&�Y��>�"%L�%�9^q �.������6ʣ���[��)-F���}|�6Z���z
,z�m�?+S��c9慍~�v���& >�#Y�NQ�X�����W�,y��79*բ�Co^���#��=Z���<��+�W�&Ť���r~��q�	�h%�w���c�\�[9�\�a��[=����(1Ќ�N
����:��ˋ O*5�@>>u�V����W�	�"��̨�.g����������ɶ�b�#^{�VQ�#H>��6����N�Kb�B�wٟ,n�d�_2�9ZA!�S�~g2.~'Y���	懱h�ܣ{PEn�CѦ�O���/]3�X�{�x�0�ܖR.�up��}fk@���lE�)�"
��|���HJQ�4��&��dU䇶���V�5`���R � L��˾n��8�����dX=Fc�{l
��4�j�f�s�h叡 =MÜmM����(�U�f8���d�l���^�֙㋭�qG�ߖ��P�B�k��]~�f�%��T��պ��{��������^��V�����y��ꑻf�_^�F�N�<�~��7�Ԉ�)ׁ,)*R�*S+0���y�c�R�bNc��_d;V]U���V��s�+}�Hh��v��$ �_��M�����cK��B������U���M��S��� �Hn���T>�)vf1FHQ0RK��0�cg�?��W�?`��8}����N9�����v��~ei��>.s��z�mUt��)3���C���ױ���o�L�'�gEnjg�X����k;�g��Ȼ����9�)mTAO'�F�dS@�y��蠲!���ln�[��0ƴ�0)[n��Gj��:Y,}�Nu�����oKb0%J Պf֭s�� ^E]BOK���zI�ݜA�����o�,΄�i̹4Tl�,�'E�Q+m���R)��q��"='��F�Yk�w�RIa���s���e�Q����h\��ϩ/�Y6=��g���̴��nR���XLL\v\�Q�%3�����ܠ��)�F��!ײ�_���E&�
%����^.E���ؘOe>z�����x�|"8`�.�M۱���Ae�6��>���=�3t�2|����XCC��(��β��Ɇ;7d5�ا��ל␗]
�MdcC�����oݛ�tE�2��U`�X#�ѻ_&,��x�$
c4��+����g�TD�@/~�ST
^WS�����7[�cX�,EԄ��(�1�]���D�[�8���	�9/O0k//" _�����������ƔX����[߽��k���f��x��$����R%�mL$�6������l(�ﬁ���� ��Z��;�*�#FU>��e�6�#�wK��*�XʊT��buXF0''�b4]��S7���dkҬGvf���O�%���2�R����?��$�!D܏U_�ن�g�d�y�_�?>e�>���)F�.�sG�5g��W.��d;�+�(���ض���9�½?�6"Q�4��>\2�2B�Ұ��1gC�M�*�4�ʢ�@Uu)7}*ڎR�O��|�z�6�n��Y��0��jY]�����&��A	\�S�ţ����g�\��˫R7�cOO߭�4�5,�w����.����̍�N�Q�0t�	8�S�(��ƄH�p��t_�������GO9��b�4���E�I�x�[P6�i�}�L���i��W���H*�~��{|��?���<*���7�󱫇8W1���ge��^:���u�ORn͜J.��/�.�44ϖ�²U��|刕��������	��<S�U�J՗i��V���y�KĆ�������؛,v����.������ۆ��2���+�%�N☏�R�7d��m�J����+!Y�EL�%���~�ب��u�D��䃍�ɉ�ӔUy��x](� _�쾏��qdE�[uC���}ꗭţ7ƩJ�m��~�VU�|N=]��=����ZC�v}���'�;�Z�k��R6�;R��DG�V��~P�z��Ӕ@��4b�*�%
��.8"y*�[~�{�u �0Ugp�x�����K�L�s�ڳ�z���YX�pX��{��	�w��˓�!�֝���r�hݺ}�y�t�L0<��v|��o�����v��l��kE�b1| (�ï�Xn_�UL}��KK����]V�}�"{����Uy�j��@��|�EB�5�fn��I@��ŊN�Ҟ�����p��ߠ��Qu�ܽy��u�U�ɿы�g`���͵���p�����v��ҭ�F������}\n�j9.��²(��|��?�[E:3�S�ET��'x�)�/8��[So�,���xO{Ҏ�Γ�]��w���+�������J�a�w�5�G���c��u����a�a���-��-I�,�U�T��sw������i�F�ٱ�,u,�(�p����G���=�� �/城���)��:a]WoO1	D|wY���9�L���k����X���俄�����F��T�*� �ඵ
:��
E�$���PF&Zv�aVe}�c3�Jp7��\m(yߚ�5�ԭW(sO[���A�uٿ��}�˅�I��պ��e<=���7!�7��V��(�/,N���g�dɥ�sX�}2�
����h>e���>.�!��$}��;-�șmgyzd�[��j�Rr���7j��h��F���h�ęL�V1�>n����Oۦ��B�M��j��}���Wj����$��V�Q}X��a���Y��� �K�w����>�����8�ϏO12�^�*�y�l�z���.��x-��?�ٔ� ����ֵ�k�I��;s��������VB��y���Bg��B�߸T��)C#�Jb��,l�����G��}%�������?OcK۬�r�(��v�! ~�e���u$B�9�.ݥO��F��J�[�e"S�Q�ߵ5�4�Ur^���]�*(�o�������g<!����i�e�Y�|�QD�Nd|�7o�b���HB�uX��w�[�1�`���=<�b��r����$�~R�S��S;1s(F�w��
������S�����mE����̳��p+!г� ��s�?�tK�2�vVz����t�r)�	�P��'�G��r]t;F��w.���7�NTp�f�j��,��V;P�c��F�,_{������ޠ�C��A�a�3�Y�������h}�W�h<ѿ 8�Pp���(XT1}�vO�����Qά��k�~��~=��Tŕ�-y��w�E0��[�����PTy��Y�H��bRu�[J���~�����j ��jt�5��S�?�`&%}0���Pa��;�!n)���Oo\Ҷ]��
F�\mNa�i�x�q$��Cp��LůcиN�A�mJzp5D������Wv�if��\]<�\�E� ��������_ ��7#{���Y=�����@Y�dU GF�\��wǹPo�[k��0�����e�\dm���"��%�d������ $�)����؃B�qDWi���h<1���"%����75��[����s+����cg�����8;������c�K����:�쩹,�t�*��V@��m�R%5ِqoA�0�r�RݣDZ^��q�T6�J�8����g*�t�|n<��j�g�F�����@���x�����Wˌ�?ҏ�g��+���^���R�/h�����.1�xE��ejX[�yJr՟jN��j�����"7U�_Q��*?] ��`�8b���,H�,�]TTy*���S�f /�� ��#_y��f6�F(���d��[ v�W1%a2���iK_����,�a(P{���'a5�:IO���R��uo!v��g��
}WӯQ�z��d~�~$1�=�q���p�������2���5Z����8�{d[_OU���KJǁ�OKwGg(��!ըBL�Ǎ�v*�ϕc��N��O�mi��[L�t+�L!�@���|Q��{�=�kt��'�e￾���Q�3���=>p�� e�W��1!�����.KE[ʯ��(���s&c�lɧ�HsL�8	[��V�0�����d��d��I^�%*^@��0����;H��Ļ�2%�7UH��#��A4|+�����_�򭤱�s�5]��W�%�fr�Z�;L���&���"<�K=��C#2���B�h�2�b4�^�K���}Y�%�SA7/v|C��K�63�y�;�=qG��� ��y�1��{��a���i�T�3���p���ֻ�?ӵ��H�{n4�S@��'~�K�2h]Q,ǥ��o��\P�h-Qs6d�͚\~
3v/S`<�:D�ZQ �0�W��h��ρ��A2ƶ�Y�.C�\7va��fT�^������5��1�\� ���M~�-Y�,5lQ���d�U������@��6�J�Y$g�P#-��q�9&�2�2���F�eN��JMk�T!.��__���>'�-s����� <b��Q�NK�>���Z����_*�ߝ�6�%�f����e>w�y HfgU!C����hN���A]�k�D��j2��)�����(]������{�Q����>�ݾ�.��ud�(������ڶM�������A華!忋vL',���fT���Gv��D�h��ܯ��L���Z؝*R�]�VA	����X5�&�?��������YJlW����?m�^��?�Y>�����E�M�A���Aҷ����Ag�"�"����tb�jS�&<L���7��&� ,|�8�ǏS'[U�d����Bw`g��ir��Z��bh��O�Qc�8}�=�.����2�3C���A�� (�~�.2/��i�c4����uV���C2�C���C�G-t�r0R<R�U�aw�ӥ��h�Q�-��d�_�e����������d�6DǑs��ݦ�����2�-��s����.��m��yanDݛ��������{���NV�1��˿�ֻ�dd+�SR��u�#+�V�`x��E=׌x���q���7�,o~���i�d-�(�:nG��%�YeRʹҗ�6�%����ե�����.�"���ڵ���O`rj�O�(=z'��q>�5^=�<��x����1�z"bF
�l	�N����oN���J����1���K�՝�Љtg�9��p�����P�s4I�y��v��5�)�t��Y��{@�Y��"�#�C�V/�q��0!.=��&T�#����o97�Fg�ݭ����w�5\�k�����$��ǫ�2�U�b(Á� ������%��#.����� 0�1�|sf����|�1�%����~#{$z�8]��2y��J	�8��q.�cl'j���5*�Wj��d!l�b�ɡ�]�.C���Z��Z!~=	|����a���x��՟��Tx�����1
)���+Y��ӀE�k�#��s��pB�.�/��b�x�M�����o�e�����7� ��l�f�� RS��v�[��>z�x������8+#�{3<��@�_�_a~�:8}�Z�_��l��e�H�
�
�$����7(H�C_�4�{�W��L�Y�p����_�A0u�C>˩C��;o9e�k�_��~��;>>�y�,M�9E�5G*xr%Z�E=�Y]TAP ��3ST��=��Iۅ�i�o""IV��}m��[^=U)�����9#�n�4�0��3����߆����ޟ=��a��M���P'�ޛ��l����$��uƴ���Y��5<�"�N�M�D�)\��O[��`@�����JjT�,ĸ6��ǲг��m����氖~����ښ���K/8v��o��ABŞ�jC�2�k�;=�����֨?�u��Dc<v*-a�6#�DۆV�[Ky_����<��6�?�U�67�����}I���*	нQ��&�@�����g2���oΧ�j�v �La� O}�ks��|��<��8^o�_^+���Y�;7	N�}����9�����ꖳ�Y�X���cb%L+䑚B�y�c��DH>:G\$�X�lL�H6p4=��q��l�����?<�}��_�_W��R�_o	���+�ҹ���e4�s�Rr_˛վ� �LrV�8?�A��׌����$�����2/d{��ר�O~����(i��h�A�s��w[=��聧p�R�I�{tՓ�9e@������ar3X�Ѕp�Q3ȿ�uOء%k��iq^5^��:�-�Cˠ�M�+n&�������3�;ׁ?o$�Bʪ�qJ���:�T�T�2���[i���u��	+ea�夰�*Q,*I�9_�ͦ�u'��F�m���f��`%��_�>AZ{����qUp���#	��_�5�)@���W�*�z�7�[������V��u��y5j�NR�RL�Jﱓ�v��6푞Z
~q'=�'?I%#��6C&��*ͽ��3t��C�dpܼ}3m�
G���!C��.��7�c���V���r�w���	@d���ʇ��q��"6��Jf/g�%��^f�;��S�n+ɥ��y�k'�zR�����F����S��}��0D�ٞ,eg��Q�<}	F�J˻�?y>ٜؖ+@��䝷���=n�؁Sw#��+�t�,wy<1p
4"��rf�K���$A�`������d�˄5��T�_�?OzL�e`���	:�P�S�/����� ��_�� �5N����gӝ^��ߓP��=��3b����`���(����������^�i�;�w��>���T0�iJ��Sd�]ul(i��=~�^�F�Qb
yO0j]�p4��5����`aß&ۋ2��tH��ŅS��k�^]� ^y�o���a��:�f l^��`y�b���������d���MN�I)R0+
��M�61a;�D����D�b&f�X�6=��v;���M�Ժũ�2.UH�8��w
:V'ݓrhɴ@oٲ��I�k���)+����=)sË��p	���L�@SQ�� -��"��@x�4j�+F�z��� fс�R���Q^W!=@�Zj��Y�P����
A���j��ǋh}2��吇v��4���|Zs1�_�y�E/���`c��E�]�%�k��`$����,;�5�~�m��5���}˱�c���d�����Jl�C�
�	�1PO����w�<9�JC�7Ζy�/G���h�.�^�w�oh"N"$�9۾���n��xк�cB�U������\Fy��&f�
~���kR�t^�����ʆcץ�.�
��#Y�8|��0,���{�4p��/ �k��(�/G��Z��O�T�Tʬ\�8y�MVYi�⑈�����?y�f3۾-��W��>�c��,Nl=mh�%q�7��=� u_Di)-.����C�N �ÛR��w�s��Z��$���0�����h�t2&B��2���i7�x����Ņ�o��޴�EU0ޯ!7�������]ٮ�W�����&h��L�#�	�ofXR3#vD�:TTy�p����ƵϨ&��/�f�D\��m��\8c
c����Hc>�i�<	R�V�Np����C/W>{���3�;_��C��R�����ım�K�v6�d[���B��u+�7ɆE�ŎB6wR/���.��\��ׁ��
n��ܝ���l�{�O*�t��M�Z; �<8�$3������:[#��XvF'�Ð�z�zl�r��A�	��M:����Yv##��G�<k%��\���z�k�[��b���9�45���(x:K��$t��\�6i�Ch<���(�Z�Z`��Eʪ;8�c���ʊ�
_�	(Q��d�ՉNb����G�Û����h'�|�c<<�k�����)��r�#Hh�-QSj38���.�/�1R+���5���V�[���	Gy��Ϲ1����+� 
�q����5'�oE�T�Wd��x��d�����K\5�A��˻��NZ(t�)C�"����ikՐv�� ߟ�C�g�0i<��q�O��1:>;s�_�T(�+���=�lqQ�	���/ʖ��7��-t=�a�A���V��פYtk\�.��?1�2�wa~+�����Ոꍵ��.�x �oV�'�K�p�ι�WW�Ot��#��ۼfP�VY����u򇌩�U��3�3�M��������F��)�(զ]J��+���)�2�j�"�g�jLk�{�#KV�o2�4Mc�jIՆ�g���	.���JU#�6�*4ȟ��'e��<,��� ng�4C�cb���$�P���4�&�Z�l��2�&+񶖄���ݔ���7,W�?�����'������n#�����%Ck�Xs����NwM�M��nV3��7Y�{����B�{�b�N��$��1�g�u��<�����\����Љ��ו�t`�:`��K��:�#P�؊���,�;�5����R�#`��Xg����~���K��X#p׃<u�&<4ZC�˿��[�\R�N� �k�P�5>���|޿��VF�bjϫ[YA�
>Γ �R���h]�ό�����+��ڜ� �*a_��E "��[A�@yY�H?78���`��C�������E�/Z��\O��Ά̴�[B<�a�5� �64��_�W�Cq��F��*T\����nU�J�z��q#����D:��S�"�'N<ҹ��$m�[([��u���ީk�@QJ9���~��ԋj�0{24zGX�i�\m����;�/�0ZWW��Ӏ��da��ݫz���Lx����Ѧ%��1b�V晣��Z�?�[Ɩ!Q�����]��[��AY�</��ؚ�7����{Y��w�t�~�ޢO**���:7.;��������4�|�_��6-�m�,�~��Iy��.�:\����+e?˭TOʦ=�:Ĉt�Ln�$�Ա������h�ⲻ>�pX�T�fK ���,����b,e`�d:��It��R���� ��]�t���I�_��M;Wufi�����l�T�־��,�J��D����>�t�����{8����?����>G�� �qt=�&�1��-�{�{�?o�kWn��9��J�z?/�3rs�r�5�R<��o���<��Y.��=�Fs���V�1���=44���z��]yL31
�C�>_uh	xڜ��5��������յL�u{'�>�r���R���R}�;���e�O��[m�Y=�O�O��+VEՑ�!�17x�zr��9,3K�wB��9��o��������<�c��Dƫz�Axa�zl�j���2B0����<[�Ct��ze�Q��+ҧ޻Ǟ�DB��r �����tB�-t��\܉0�L���uZ"���;~B�bc����(�1� K�_�xϔ��!� ��q��P/�-�5T��TN���3m�|r��|�� @�޸��
|?V�6���/��Q.�����S�ȽO���\�2�}c�OY_g�̳ȊZ=F�����
=8�����UW]5�������R���Y�12��[O�僂80�eO&��`���\n�2~������uHK�M�>NQ�:��܆��[����~�댦���mo�=~�����]/G_����:N7~m\v��n��&lS�����U��~�7���९��	���*¨-Z\�h+Q��>�YX��l�9O�QX��r|�\J���8�w����ǐw�����e�)�a��`�هG��T����ଥv�'�(���
;
�A�����F�Bj$�"�l�u�����7���ۀL����33-X�i)����@�1O��qIn&�w�ϳ�B�S��-������څ믿��;z��wqC��º���B���<.]�L���b(#W����\%���9$�|76ՠ$��4|m��s�=�'� c�1�2FU�KL/��h�i�|c�4�����n�q����]Z�涷�4M('y|�܉y���5�P��N0I�-�\��]@Yߎ��5�k��r}\�d�Ǯ�O��ۓӈCh�rΏĸ#�X �k�s�J��$����eB�n'.��Y��h#��� �KK���*����j�K҃Ș�S��ĀtP�Oɕ_R�?g#d�gi����AL���A'�Q��Q���S�4fZ�&��"�_" �c����q)�i��*oV��F�<y-�K/Z�3��w`��+���}��o��"-����٠IY`�Q8��*2��M�c`W[�ewi�nmS�pHS����ć�_��8���&��I��W�d"v��#51�Q'���:���g�S�Y������[��Ay,1�>�iHc�11�P�h����K$���\�ѺȲ�,�p��#i��y,,.���8AzٮK
e�ID��;�C(��� ���.Q�g믽�o)�h�o� �r�sf^�l��iֵ��k@�~��	��̨)e�#�Mh�Ҭg���Xe!��I��0���F Ä��C`�l0����$��PLG�&'��?��%R�f�s�W�v�����2�m``�L �X7���O5U3�l��mZ�a�_�4>�/�r���l�p���/{Ж���Oض.$`{��LPk�Ak��Ԫ�W�p�ʸ9 Z�E�Ã�3Y�_D�m��+��t��tSH����Eƃ�~&&6�s���W�5��]�=��Z^�T�oN��ڼ��ڷ����I�'N��2G���O�1k�qY�ZA{:U���%�Ǣ��F���@$�Q�����Ep(k�P˶]k�L�T$���̔�1�z駉�T�8h<Ʉ��)�)g�hL�|��Q�R~��t7j]��1�C�E�5�$i��O0�&����<�4�o�w���2�v�y���2W�Xö�ϣ�����_'z�;j��� ��u<k���D�ܬ��'���q�'k�4/'[�}׿=q,���w����y��$���׼δ1'��|�Ϣ`�9L���z�*!�f����J+0'w��xN��G�����(蹴d�&j��\���8:���M܀#��_�,3d�]�n7����W��r�6�ʮ�].	N.@v��K��ˡ�������]_���<���B�ɩ�@�B�t�'~�k{��߿��p(��VZJMfd �f�М�(q<�SȞ��7�\�k3���Ic;S~dX�<r/�.>}�Ӕ螗�6�-��R�b
��(���N����(�c#��>yY�qҾę	����hlh�����,����&5�w������X�$.hF�a�mN�\}-�+5�䛍����,�q%m��"sU�G -���iJ�4{uHX=��p���J�3wZ�ՙ���W>�.��ղ5�S���K�<Ϯ �>2��3��,+��5�b��Ex�n�rv��n#��3���:�^��]^j봽��l��PhY�yLz�qã�F����JGv��md��]G��d�p<>r�!p(kP-l�-ۧ)� Z��Na�b"��Bh�?Ô���Pz�|I��7���
H��"���b6:9���ך��,9��FsО_|�S��K"�hsN]:�l��^/k�F9���G��(�
@�b�k�!�#j<���ځ���h~@n%�BkTy�p&ߴnOл�$Zf^@]�2B	Ik�&�
tJK�H̆֠�3¾�1���皘;� 9ٴ��\�����=N�:��V��W��^�Ao� М��D� 7 Љ�C�9$���<�i(�y��o�}�zGJ]��c����]{�׿�lϞ�c9�j��e�|��!��c��+�#���b�+Z ��[M#����}ߣ��S��/�Y[M�0���8��0h���q[`�t^fn��S�hHJ"M9�5@A!���h�'�#�@�c*.��ąb�L�r� 3|����l��w	�Q�7a���nWV�t�ٳ�8���j��T/_�ËHs��C��l��q|Φ2��%�]ϣ�S���Z�u$��B����ʴ��+ZeZV�^�tiA�;��$��&��t=Ћ�d�Y�K��)d� ���x�����y��D�2*�>�4̑��>o;v��IP��w��(�#p�/�1�MY����u�0e*��ɍ�#W=��䘰}7�<�n$$����_������:�:��H]�1��.��3��~*kr��~�}�]>�^6�ۮ��|�,;����?N4ὺzV�d>�7�xV�%��hnq�D�AG����NE����)M��˞�T�R){�8���''Ĥ�&����q�����KtY�|Է&�]�U�����z~�� ���md}˞�r�����ڠe�7_�eRt����<��7�_e��3\B���|�]7y^��v��SC�.r�sL�m#����e}a?�v�#��V��a��l�2~���f�
]�q�R2�U�'t���(�c��P���t�s(W�֜�\dw��q����]]6��Le�Ma��]�$�.j��2N�5Ё+]����c�3�쥱��-hd�،,�)o����v�ϕT6�V��_����lP��Ajx�����s����K�p���R���(�D�J����*W˱��r�/~��HRa�c$����{m!d[.��l;�+�u�\�/����R6���g�km�t���v���Lv{ ɴI�W\bv�^�7�����L�^YY�֢XdV�k�����r͖�R�٠Q��d��R����.���L��%��'�b�Of+����2q��N�������26�
����:J��bz{ ��v����ϑec�	�<���q֘=��zN�$y�LIp���/�c���6P����Y��P�VL��fb����l�� (�`�lsY���县w����������K�]���W�W�L\�����EY�BĜ8Α-��v{jnnnf���m8�4kU�@�r&�
�z/��n������ut�Vm���h��$�d��v��Xx��T�@ts�i��(�Z�6��6�˨%�S���Hv�>^�3mWY�P����m��V{e|Aq��.;��L3�_氶ۈ�%�_��e�H���;�J����y^�%pu����wȺ��7�dlE��N�=��[�)XIqu�������	R����r����{(&|�s��ر��G��ߎ��Q�=C��¤/��?YP���}�2�dJI�FՖ���䜬���H����UvL���C�@Z.��<��R�Ɛ���$��c��9�^]j\�y��(.p���^0]�p�oyL��ܮ���d|��Q��qΥu���jk�;�;��w=��/�o�[��qJ�n`�6Ca'�9�����m ��e�e���5����\f���a[�.~��%�~~��$l�ɶfޒu��}�H���������p���H}�_�t#mH���&_2����')�� �A�`��f[�����ڽt��<�`=�YZ�m��<�����l���,[�&�Q^#I>���O��K�s	��n���ئ�,���%�� c�m���2pu��5�̡w.���)�d�q�r�����=��e��&i%����4��l��|��c�N�g\|%�|*�m5�~.@f𶅑T�dyx�K���#�q	ֶ���~�~�u�4��;;;���9Um3�:�y��e�����z���8�;����X�f�rp0hK�Eƌ�;dǔM8I����$����G�5S�y��D���b5Y{���R}��6���e4�#w��rɺ��Х)���6�1���k�<o%s0�A!7��D^i��&ن2���\��\';��l�����g�2��,�>$K���<�5��7p�Q
 Y�"���<.��9�Cx=����$�'�=���\])'G��������̗�e�-�l!)��q	��r��bk�1�8�1գ��$K���tsp��q���gH��Vc���Y$�Q:�^'�����E>KK+��e���u�b�Z=��l.@��pQV!KC-�����>F))�>';{��yX/��4yd]9r���yٶ(oh̳�Aݩ}�3�v�P�'�Y�\Z�k@ʸr���p�;\Z���6��9���4.[�d� o^�7��>''��\&��c���G6�`3�=e�K`g�ī�;/��ö�ZF�ha��m`����++�˂��Q�T�\T�֮�����eױ\��]#ec�%\�H��{|��=6��3<ΐ2�Z��AR^h�� v籉"7ҕ�U�2M�y[���b8>��D�I(�s��ػXHmI���sl敌@׋k�W4)e���匶$y��>�=�$��]	v�X ����t.�5J� �n���׹4�By�_S�eﰟg��v�]��ϐ��5"I0=P�g�ua[7^RtO�v��S(Hv\�%��AW�H�f+rL�c��c$��%�]>�����.|�u�����?~�q���l�3�i'''WT�l�h�0�=;��4�FM�� #�w
fuu��S�Hj_z�]��m�s�$Ic�܅��f��@��en�qژ���.沟5N�ti��g�
�b�����wig�k�a���L��-��Į6�%��}�����w���������kh&3�e�q�*��ٕ�
]���e�\Y���/�������m��V��x.+�g�da��J�C�'��	�Vt\uw�Ѷ��vε�tDx��\��=k`�F�bc`B�q�產6x�~9�(+aK;I�λ��t4�m������סy� l��?]�k�����m��q��%���ڣ�zp�����ylO�1��}(��e�̩��n�����
�ePܣҥ���t�?G˟M*[��g�`d�'B�>(���5G޾��� g'j�@f�`t��,{�P7e��&U]8PFr�~���e�e�����;[q=��n��./�].s�I����[�)[��I?zq̨�@���C[�(8 g��H��'����	W�X��↯�	g"�%9
+ޜ�LK���fX��媧}��w�/Ξ�p��.�$5K9�6�]d�YY�س��}2b��c0��S�[���6n`��؞t��sYe��|���ʇ$-$$y��7�,�S����.ps]_Ԯc.쐼`�8�ř�x�mE����c*�iynX˶���}~������Y����]�"Z�'��̹~�h �=�
.��
�_����q�1���䤢k��5�{e�G�E������{m?�</;;/��^9���j���S�E&v��qu��s*�b��c�c�k� ;����?n���.��5S�0����q���.��-�=�w���XA����q$�kG��@�LI���u��e�2��K�)���������2�9
��l�������YO����@w��{�B����t��3��Qqy�uv���	y�8F��x{ٰ)"|��6A߶��+�S��ɨykG�ءF�Lۅa�Qw�(C��%Sʙp��]u(Wy�Ԯm�lٽ�����r����#bʴ��%[�����/j?���lP�m�ײ�]�*���I�>֦���f�t	��[.A���l��Kй���q���7$��\���8��T�d��ui�����ș�Jn���
� ��ٛ`�����i�$�ֻ�$�\�:Փj�kͼ�i�[��C����ƕ��Xq�?[*23�q��'&������4"̾�(LBp�0�.�/Mn$!���n�8�,�Y�[�G^Ǯ;RD�3����ߝR>m�=_Q���|/\��ܵ�'�<�7>��(���Q��r��<Ғ�v�btn�l�m��+2eg^���o�!�����q�IU'��W�1�wաH��s`����F�<������s%f�����ߥ�u�V�|���@��	>�g�<����5I1&���b�F�65���&��#����l帲-4>�y��0� �No�f�r>��,��F��J���s.����aO�2�d�|N���8�G��ӷ��ݴo�P��p a���l��C�·3�����A��Bw���m3Ɩ��L�M�2sC~�F"�)��Z��`���/��2���匝:��>&ﱥ���	�&2�I	>���4BZ7�_�y��j�RS-ӈl���dh��G.��1��� �~�4˅y.�|��NDw.jn�,��U�������W��L�e�Ze�A
�5o�9���AmTd�K�D��=�c�v!�ضI����u�T��Rü�+�����h�ec�u�t�[�/���}i��\?c�o�3�l$�Fe�*��s�(AĮ�Ԅm�C�/��T������������ '�Gb�SBy�\�+�C��廥�`��Բ�)W�>rbVR#tx7�)�֎ x��칶�;Ϲ�x.�aן�j�-�$Xg}�m久���;�a�L����G�qݞ����� ('S�|���|����6W?��$�:IG�-��l�<�[W���?9'���*.�5����4}�F�o�r�w�r��Lir��B{[J������͕P��m�� �� dz���e�m��f|Yh��e����ˀ ���Q6�-Q堦k̆�`u����\�$�خ����mA�u������6q1��6��}�k��ֶx`���㞻@���e���3�5jb] A��S{�,���;$��m�ϖ����2A���]j�rp�ӵA�9)g��~D !ٖ�KC�`��y�����v[ڻ,q*��tQ1I?s٘�ϔ�v���è����Z�=�pxv9!5[�6J,�Ys��f��B1I-GH$�,/�_+�C�l�v	��3�{D�J�WjE�<��L;�惏/���.��/�4�,�kRD~gӮLh�v�{l�(AA^#'�?�5!Y&���L���)T�y�o�o��M
.�#_�{��<�l�)}��/�,.�cJ�+���g�Bbk���ݥ���Y`t	�͛��3V�#���I�����pH��9f��}+�+CR���rF�r?����s�yGN��_���O	貿�Z��l����J�ͫJn���r�m��DNz۶m�]�ImW��x���H�Ⱦ^j"<ʘ[��J*dk!�3�䠲kQ�A�-�G���eRu�&�u��Ɓ����}uR��ϕ���f����Ej2.M��'�K@
W[I��j/W�����%5L�z�L�~�T�d@��>M�"�d�\Yg}�<�K���z*���r����V@��`�����y����۠,-n�|�p�P�W�0��@��}��
%�����;m����,��D��ڏ�ӻ��6��*>[	nn����m��$��Y��L2C��{m3���p�l
��r�ť�ٌ��<����}v��$�]���w;@֬~��wՐ��]F�cˀZ�����EM�z��*�IF��k]ϖ��:�bdY��~�'���n�Z%d_��v���s�Ų=E�;�##%�0r���Yn׏�'��v=˔!���d�\[�p����"��e���u~�-N�8~x�"��x��B�%�9y�V��s\sp����~_c�
�ڔ�(�{���"�h�lRK�	���,t��/I,`��0g����ԑ#G`yy�l�B~k]97��w|�5e��mͩ��%��`퉤�.P��Ϗ�1z��Y��&���]�Q�VRC��E�LlGi�s�q���a������M��)�3W�%I�����w�v�'��v(�#+�� P3��b� "��ix])}e{� i��N�/�r���O\Vn+.�����Y��+�!X��ɩ�(����n����rW�t�IM���r#�@�yw\�*���F٦\n�?%�����8:�
�`yq�$6�P6�k�z�.��6���TV)�l��.��͂Z�/	�{l���I��%���@4�d�n�Xa-�Rj&�q-�k�'7�S���Q9�<���\`�0c��PU&
oLY+����H�����^tI� �I`|�w����G�K�%#2�ױ�:̧�f'�07ϔ��e{pT]�(l@�s.w~�2���q�+++Y;��	��n1*l.s����;�<ڸ��îl�n��݇�����b��6�6���ؾ�!��k���MXJ��~Z���[h#i�K��s��U�;%/qTG��V�zn�����A!��5�_�|���8g8�y�<9o��_��矸M�_�~��������v���Z�S��R���1�����7�o[f8��4�f�"Oަy�7g���l<�<H}wJO�(�eοM��/.�Q���[�F�1�y�ݻ�~ci�P�
_�93dgHMI�Ԭ�n��g�!�;�u`��1n09𹑓4O�.�Ã��ı_�X�(�a#c��@ ��x�?�kH��ߎ�.*��`�=��7}���e�*<������{��\><�@#]
<(x��IJ~�]n{�.2`�^lM��-�z��r�TP��������/�;�v�٢�>����)Up���V<y���0���@ϼ������� {.��q��v����rIP�DeS�\\��� ��^��R��06��d�<�C�&�?|.Wx����7�ۙ���[4�Zn/����þ�q*%�����V��ung&2�Tn��o��b�(x9�r%��N�}Fc��=ϋ.��2���'WH*��)	��?v:W�58 9 \��c����8��9+�ľu�����l��$��$7��ls�J�&Z�F����/��۷gLp��� �O���Z4ރ�y1���4Ӳ�/4W{�3X�5AV_��c��~/7�	ˊ�ƌ��e�J���D�F7G�˾.�K�[=�/<1�5�Ѽ��W�q{���l
��y��<����VWWi�/..f���V����}q�&;~�xVv�'(�.V$X@�������m��KM�?���¾�gr�bb��R@˾c@��ѬAsyjf�)�9_�5�|��!9�$`KK'��wx|I_=�s�����R��p����|�u�>w�9�cܗ��3��_/�	}���8D�}����΀Ģ�w��}#`s��"�F�v!���̯'E�j�R�!�)$5J[�ˤy�+ٴ��k�L{ŝ��Qs����s�N���Ç��8h�Zb�X���hX��w�2e��r����$��HA�%�f"M6P�0�< 05���V�qJ����5_$9Q�� ]@-�iO I�a ���M���8[f-�[��a�`+J�!��>*!��:"O5����;�y�ۃ��ے�g��ֈ�-���B���|�.)\��#�O��U.
a0N��>O���G	������\ne��ca+�X|��s����mֈ�G���]����Ί��¼�
��Gi���7��e�$y��g�i��\�^o
΀2��03��`����u���������Nd&?2km�MK�3�����u~P�_�ɻа)��o|��(8 ������Q��nx@k�I���I�V��_|.N��6����� �V�dt,GfndZ��(��D��j�"��;W3X1�+��lA� H�(��'	�Z��A������sH�#�O��v�w���Ҭ�\M�c�Vϴno�<�- Ms.�j�̧ڊ�
<��a!�����M�$�(N !�ߗ�3�����[�|��	������m��^���#-H8XV�Ҿ^\S A��z\{�2�'�]ǂto��!~v���7��C
X�/���ؒ@��%['X���r����)��V%�I�-�e�e]���]��*��N�}v&�8]A-�
%29j"�]�9�D�<����lf0�K�J6>U��G�	Ҷ��P�nK�E&`��.��ǹ1ѢXYZ�A����*�.:�C�-<Yc�u�^ѿk����6˿KUF`;����\�G6�7n�H�>8������Qӂ�����ʜ²|4(`tM��h�v�~�W��r~�7`e���5r����y99[8hr?j�N!���J��'�q_d�eYFť�4m��K�L��� ���)�zzV��Q��l{�~q���Nj��?m������ƽ���2�1�`.�_|c�y/o�ł۞W)P�uKa��=e��	81���%ͯ�����G���Wv�PR��[�n��Az8�	�d���@L�\B:�c\�����qK���^���DcMݧA�y�5\�����x~Jg�J�f��"?-�9�ٷ[ht�H��̵=;��d6���J%�[__ܮH��r�#vG�����/�;v������r��eU���'��B媮�t��
fA��ڊ��"�1 *"�AEP�TPAuf$����AĀcb@�4tC:T|��M眽����k�}�=��Wռ�޵�W}߽��{�N+��"�j��fsA�Z�_/��rI�S��BI����=����+�I~3�>�_�Qu��$�N�ނN*�8�Q8�𚰭[x�<c�h���j��Y�FV��wDy	�Z�
���m���OȌ��续���L�]7b�r���di
"{S���~����XBԞ�p���9W{?w�M�bф�{���{�6̭��]!8Y8� M'~҄)�)#����b89!��<��a'�=Y�KwPŝ��Q�_�Z�sjfTk陓�Aҁ�:�6,V�	�u�.�w���q��	�"\�E��C��k���3�#�ǀLY\@�N���P�����P��]Hh��w�	���
�
���T�S.j`�����-��?�OpȈ�;tYy�-4%�U�rNQ�1��/����V6����l3�P)	��vv��+�Ì�y�\Pȴ�����@B�43�d�d<mfm��Ϻ-����Ґ��D73�m� [���Nܰ�}���
a|B��[o�~e��=)�#�5�]�!삳�Ve
ǯ7��9<w��$7��l<+���&W ����]9����ĕ��s�3��`j���ln�u6�~�ۄ���kY&��41�?\t�T|��5��G�H���M�3+������!�Q$��~8����sA��I\iN7�����0��� Y�xf�Gl�
�A�6S�̈́R620���+��p�����'��J���8�S�dxn0�H�k�'%Qɜ�B�&�BIx���L�P�&%L�}��5Z.8V�t[���ח�K�Qn4�����kH�`��D�*#.�'�s����
�["�9�hd�ʏ��i�+�W2d�~d�B�!���3<����)g�/��u�ΦU��~���F�ۧF1�7$Rѫ|G%{��g�U4*�����W�PƸ��7hSW>W�}7�?3 P�/eLba��b��z�^��=���x����K��N�T�Z���-����x��')�s���oq^��K���x��%	U��n�-�~.\X�{A�f��D+r���M�t���Z�0����"u0�K}��o�K����1|/��Xl
���������4f]k�!��-w}W��t��1H��K�0�"D�k��>7GF1KK2�=�AT�4��%�V\;`�$�{����2V��@��)�����ڶ�}�	tc��υ9w��ςy{2;���Y	V��/�-�+xۥ!����pBkIAs���7|?|l|68(���}"��=?a�B�|�{W������k^(��� �u	�uC����6Y�"���Z�<�V��{A�dC�l�pr��f֠����2xY��D1�C(�>��o��v��oH�'�R`�!�EMK�q����	���(q�#������{��&�԰[�)<Xa�S\V�����U�x���5���5�i�X�����C!�S�-G*àt��.���O\�������!��b���&-�Z2�y�}�����15�uSxw��vJI�2�Gd�b� ������o���s�Z��a	T���vۅ���n1y��OH�n�`��s� ���Y�s��f��&����}I����qV��7��2|���|�g����4n;k�.����(&��p`��Mn�9��������vǘmb��χ�ZX��$��n��i}o�=	SZ��.:�ʙ�!�^İ�E;�]�Q�$è{c�I�V�x��XĈ�B���(c],tz~\� e���J99RCX4���w�ߺ�'\��Z�?�%$�����m:���s2�]q�E�?�d[��Hصi;a���.?�>/��d��]os����
�}��e�$iڰ\��JR(˹9�'.:Ǽ7�^�g֨}���J�@m��Fɛ3�tUS8�$� ?-�;��`����4�e��A;8F��`/bb���]���.�6�n�Kxvm^$Y�v�{8H�y�sn�k��]��Jp��y��y7[�-b��yʴ��'c
�U(��7Z�vZ��<��u�n7{���8��d&]�,��|p��"�״������E���w�>�ڳ��w���F)��ס�
?��|{��㫕��[|�����
��?tu��Tg��5��/W�� �Ȱǣ�''U�&>�Ԓ�ׂ�%U�~�v�u�f��g�!���梍�����ׄ���7a����mstѽ�I����S�=t�Oxo�ki����clk��u�o��.,]�:to��&�)���o��_��^���h3���"a��������B����
��P�-bt�q�)\��~V���h֋�3T���s����^�&H]M�R���q����R�z�K��{p�P	�ϟ?~��;�\:y��.�<�>xpu�q�$h#�[���@C�Ȥ��l秬ym+�X�7���;yAd��w7n� ��5����n��
XtHѢ��V�Q�y?}kH�?��{'],d����K��=v��yg�p)"��ϖ�o����3&�ˆh�9��vz�'U��sO;ר}��s�v-���E��'� �� �P��3�V&L������b�~+$ۑXOjWk�w5�������W .����'2�&�k�T]���,�s�Ϲ�h��Z�
�E��m��{��ֲ���M��$̫� ,	և�kPL�z/O���cS"�wcq5*�e��o�\��J���튵�_=qm�%d�I`2Iڊ�/��#����e;j���/�=e|!&n�t��P�ݴ�5R[�5/�4���ڿ��6[��.A�'d�Fu�j}����oт��F�.~�v �KK�������U�|��"����@	S�Ғ�Rt��ׇ���*X�y�Ǿ�ao�^[�S	ʶ�%���&�},Ϲ�23k��)%ͥ������ؾ��=�v��v���w�y��yn��������RF��#V"�Ǭ�o�AH����;n��-��-�3I���G�U@�U�G���ͼX��aM�F�(`y��X� D	���_[#x5�M}�y�6;Ut���)]/NP,�$!vG��2�`2V,�m3��\*maо^^o64��hҜ/Ɋ��=K�P����a��ש��J4�w֬m"��da&�0m���J����),�N�\�����PXY�*O��KiJj&�X&�I5k��Z��f��)�G�����2���u�~�PjF]��H��\��.~�󫵤媅�P�7�{����s�c�ss�*��N�B��}Ű�J�����@��9��^W̴�M��%�AZ�|��;+3G3���e���")�Y�Sq{�#�,����L�0�%.Z�Y�A��ӱ�Z�g�F�ڎ�����������#�M��B�&��m�!�Š����_Ҙ v57�u�^�F����U���9&̓I�(f�������EZ�v�N��]�*���l!��q���b�˹�-u��b�ۍ��B&]�gS�@W����2��0��=Z@���U'�+S�v��xM��s�fi]�.<���B�*u���nZp&�C���3륥��eMY�����C�Bߗ�a�\�ݔ�dn���>�|J������Q�Ki^K�w�a���ޮ>�Z���$<����$ܛN�zŴC+�����Ҋ���	���Kv��w�л��B�}
�;4F�e���'�qe���Ģ�қ�a	��$���r�?v}��NBy���¨���g��zz�CY�]>P��m�F�����n���w�.d�8f�L�4uZ)F+�AW�v�d:�o!af��Ңi����p!�pkaܤ�-�ڛ�G��2Y��Ʊ,kAϩ
�Y=�L5o	ii�ƿ�㫑d� ���s���{�%R�4�_��"$bn4ƾ����n^���.}ı�41À���׿�/����l�E��>���i�Tn�4�i�2�fz�y$��!5����Zo���T׼t]#�.�h±��&Cm:I��R`�p��wz��b���������϶�Z7����ܥ���1,�����mf��c�Lu�q2^��ɪ�~�͘��j�9�~��ܶ�L�S軜pB8�P�������t)�"������;HV��؆<��?�v龷�jB�
�
'���l S�)B�-E�C"w�r��b�ÿ��t�,�Yj}O�0�Q/bz�>�TsS��~_�׹m'�wҔ������:ǘ%[��/u�k�&�\����'�m6C۔@��Y��=o7�E��v���7�J���z��X����sa-�������^��|7Bk�o�s�.�f6i�nLZ�p�X�ErH*�����R��,pv�񑶐�!h��[�f����KJS��>nS��3K��}-���>C>��_gE����(+X,7��/�<���������p3�nFj��.�kKe��%�7{����޴"��[�P{�Z��j1���l�f]�i�!׺�{s�@K]*�ǵ��<�B�l�1,_4_e�d,�h���w��m�IP<�yO�q07^)(� T3 ��u������Q�]"��7��aL��˚��]�}�ՙ���t͝�ǀ `�{��{��	�n�_���a7__��{8x���D�����c˰�]�ă75���0��n��&���4u��`]$�I���su�-j�K��6�e7��6�gdc��K@��"K��b�q��B�0���=��m�m���M�����6��z�#4��r�<�:`<���0?�Ļ�y.�Լ ˝�2 ��Ab��t9����FP�^&F-}��p_뺷�@�����=��g�N=�����@�k}�D��Q'ɷ-�,Z�n_v�=
��nm��nw�5fc��P[=!�
�&�q��t�� b�m���'����=��:v�4\"� P�/ٛ[�A��لN�Ka��̍4Ch�ҥ��{)#�Z�.*�$�"��g��svL8)�iI��L��	�&��d��\lzp�5�^褉"`{��,a`�z��4X�Z)ы��K��|ݷ��U���o���Q���#L�a��p�,�)�iii�p����X�%lwv/y����������)��Ub<S�uOI���EQ�-��;	������C;]�f���a��EQ���Vu�v't?`����G�S���I�o��I˯-���
S�i�����)�fK8u]�p%�� z�}�q�,V]�/�$���d���v���C��)�D
�5�9sj�"�NJ������L&,�@���W�i`��*�f���#�L���\�P�+���8l�Y��F<�ieȿT�A�5�g�+�hrQ�iu��^q�{�Q��tݲ+_�O�XGR�a
l"n�.�0k1P:��8+�гKQ)��zг��kx�X]Y]� Kx!frb���o�{�&&�e�4�]*Wa�I�2�/B�-�e�h߾}���U�wp�_c��f8�>���:o���!�禮3���7��j������e��mJ����RE'�r!T��J����4.lI�&������8�vy�32q��k:�c�����	 .@ѿ��������'�PE��JT�4���aF�@��֌r�y��ؖ���O��yv��#Z��<,ɗ��_�������1����	arWG4�vemC�֭p�b�D�|��e�=;��Yݗ��+�g��cX�Ʉ�v�iC�~X��$�(�8Ch^���=������݁̇��D�\jf2澓(�	���t6�5�_����vi'$C�M<	��F�@��YF�3`�2:t ƣM��VSVW�^��sg�k:�2r��Gc�G�(�����sj��{a�w�ukp��`��]����~��;qw�2Ԯů'h�]����V
[�p�yϗs*V��.��3��ؑ�� 7�q`���&�����4�����d�RP+�����Ȍ	���P����<��]��kMO�c+������\.�T�v���D^AJ]J��a���=���Ze�Ș�K�����Ba+�°q��5�[��TJ^�+'�������\�ٔ�~��U@Y�~a�������~Z[�-e �,O�����Ch*˼P���qi��ߙ����9U��F�'�Z��p��Y�U�t��#�w�s]D�8�R}E��c@�*��Kd�]��`逽n6�'����{�� �;�Jb�`�?�l�bٶ��D܈�G���=��v��<�>w�m���g��}�0\�ٽi�`^����#w�๷���%��$�42ζ�k@�� |(�-1�SĚG!+��҂M`��^d���8��_+Z��H���L�o�R?�{x	\��\���)[#Z��l��9���h^x�S��K�>�f:�>����,Jl�i
�2k3,m��e�;�x��m�84��,�*�Aƌ�**��e�G�ÖQ�,q{)\Pb$J���$�Cj72��ڛ�߼��E�j&�Ӫ]�gì��0Sބ�OY\I1���I��$Dr��Y/{�}ɲ���$ဠ�,��1�AF�~�Ԍ$��n �=<�R�J�/�p`%��2�=sfv��f0�`*�mW��\i�cC指Z�I�\i��$����j��_����W����oewN?
k�KvC[Mhb��*�`��\� KRҊ�9��sR�E������\V�4��;�ܢ���+ϥ���Հ��_��.�z�E�Ɯ��Da{`�
ؿb��kL���p���?%Υ���}�c{����6F\�n0;���
����%t{����E�8q]Î�� ���Uʻ��B-�6�������4�g��n��z��qz�����1F�j]��!�w<&k�}��o0�N�
��Pjc��oh�=�X~�f��B�,��~�xnI˵��=��W�-�ϝ��~v`�.�����>����b}ȡ�:�$d�[B`h�5�ƛ0�J$j������[�NB����*��q�ص��&�[�c�ֈǏ��6x�EPC���?�_�,]F�ƨLpM	�vh�S�2{�Q���/��q�p��)��3j�C3���b�`sk�b2)�MPv2��m�I�A��^��:�n����Ë����C������M��Y�S�G@��X+bp��Á���߯{;ZH54��7�l��?Y-l4N�������ٯJׇ� r���=8x_¤pWvN�K7�ߗ#�%с_���wd-����KV�X�f��|�#�}��w|�Z��XZ�믿����;�$&�ώ���G��������&%�jR���ږ��E�k���4Q�{����#3�^��V�$y;"�Z �ɇ�֗eVG�����˭���,?�?����Hc�6Z��;�\�}�����>�����E1�s腰�)���K�N�H҆M���A���=�-��e�}�C^[[;!��DXK��F�P��9O��!��~7^����X%��
�ύRwVxN��N� �c�l|����>cX���`�@p/��tk�i�	2gQ�n���x����D���)��ٻ���/]{��3R]��fn�09��5�tӍ�5_s���(Y����'w��h�
B˷�9g�����O��gx�n��k��{�
��d�V��7<K�u��������N1����	c�fw�}7~�k�8��5��(����`�$��b`��=	'����˲��	����ʲe���������U�!�1�I��v$v�d�,R�`x�Q��%W�H%�x탚 u�
1��ƬYW��*iѦ���G૾�fX�Z'j�ȈQp!��nkMƪ��������v�h"W�eP���1k�c(�o;�@�'�U4j\7��mb�0u9�,f�0mp���+��d�����/||�g|�����Q�F?��]D(N�[��:}�,�ʋ~����#�Q��5�<�)S��A�qN��pI�"Y���2H���Vx���n�]%���H�y���Z�FMҞU0R����|���!�y�rzԮz��N�m�ǥ�x������ί�ִ$W@Er��R���M]-(�-�<H���|�+�ӣ���/û����}�W~�(�b��k�T�y���n0>y�����2q���Q�V��|�o�[���a��)���Q��§XP:���p�	8}�,���x�Iρ*�cI��K͘�o�|޿@�b''��~�IOz���������?������">{$���ȝ�֧X`q���/�}RQ����k���@;;g�)ŭ��bI��*�6�� ���Ò���O%�������pg6�CIX
��e�^�7�������y���<�Tj�EY���^z'vI�F�T΄)��eᗑ$���}|�#>�9@����0)�A-9�53�P������PZ���1��} 6��K����`B�hQ�9ܡ�'J0i�^��"?o>�v�ĕR���.�o�2�pݵ��_�p{��@�߹2�r����ɘ6U��{���&�ykZ��o�S��I �SJ��Đ(0�~�7��/?$;v�#�zի��2,m��8_�z����o~���4jK8bJ��9�)Z}l2l-��?�x�C>��vO���D�{��e� A+ Y9䘃��=L~}tg ù@͘ �L�6	��e��տ�{�����"(pl�s~�g~���x�7H~�v�L�o� .���1������t�{��4�Ҫ�X�@M|3�NGּN���[Y����vO(����.u{Wia�dΆ�x�F��~���f�H�����x����;ح>M��� 6�[�s��юij�Zއ�\K��3
�g9*V#��)�`�~�1�kM5�U�d^3��+(�ȕk|C�:�$��H�[����7�籏{���Z�W��w��?�t+�^�}���eX+e�&�?h�QA��*Z�Xٵ�<���q��u:����o�Ƥ���=�+�0�L�lF���3�Ľ�o|�+������'�Y9|d�6��o�8�Κ�����GX�h'��
ʙ�)"��)TZ	�����ϵ���O�f�eV"BS\$�)�e�
��v�ZU'MASj�/Q����
]5e�P�L`h�,��4��w|�z����f<���x+��s��/���5x-jC 5Av�2Uا�R�p��2�*R��Il̢`K�d����HOHx)_)%A.��ؓ@@)���Ph C���kϿ�5����<�!�ֱƏ|�Ӟ����=Ȩ����&��fM�Z��9B0��-�|0�	�J蟧>�)�BQKƀ!2��a�PoM����,���I{�Z�;�W��~K�:f��Q)u�^����c��^�җ��_u�;��cx̏�ȏ���_�����n3��8�+����C��ĵ��r{e�ߤ�a*�P��ah�3T�5eHX�f�a5���"��X�NزJA��@*� �.�9��n�	��۾��;�㕰����'���O�����7<[,��iҔ݁î���E0AA��*1hZ]��T0�:a?���2�yE���r��ޠ�%ç���kB�5�
r�����o�����Q��7�6��_��'^X�����?y<�=kV��f��4B]{�$�+������Y8��f}JcF���-��5kRl�Y��M����H�>-1L< �8������?���iJ��k��`����oz��ث���kQ⅙mb��Y���JQ0�4i<)O�2��=��.h����Tt'��.��5k����|8DK.�jCL=��|��L ��G���W��e�=��|�k�V�}�=�� ��E.�Х"�`ڃ��d�\L���)��qYF^�IKZ�&�	
7d�xP\,
	��]+�-�V6
՗��%߼�Q������?}��W��I2.\[ʖH�ږ��k�Ԧ͎�k�ts��o)�>%����k��"�12>
0;�TZ&�)h�3%�c"r��Y���'��7^�؛o�g��z��=�~`�/��/�+����&ϵ��1��X+)�a[�En3M�2Nq̸��wO'��0/�i��\��wҫ(��*E�ܬVe�K�jN���e_�e��g~�g^;Ћ_��?��?���׽�uO���N�Zu���ρb,j����t�8�\S*(�׌�mZ{�/%�mt�q��� 	��?s爹��d)�s��×~�g}��v'���'�=�ܱ���m_��^������\�t<����T��B9�V�bH��y@k�\c@q�<�V�Zb }t\o��e�'O�|���~��������K��+�zmm�3��;��[��a�Ud����隸�j���p�-�E��J�5���e�L�4W)E3@�J�6D�'DAm��bl�K/�9�*q>`���]����y�C+��<��?��?�"���Q��<�1�˿��_��_�՟ű�fRNgC��U��LX�D�3�f.�P�h��&�����rm����a�)t�����rgہ2������Mo��ϳ���vZ����?��g<������$UU�*h�O�n�����oe5���
:Uy=+6�Y�pY��Bjh5(r��
�����lR�ߝ/ap�V��/}ɋ��+o��ow�������z�o��/x�/�{W!�6R�qc6����8�@y���Ҙ08N��{*���y�8Q��y��+�C
�Ө%��B1�����������eO�]��^��?�����ozӟ}�����ij���+oS
�nllH�0�!�}}�`�ffS��cE{��~�<�AEd���!*���ƥH���������ڽ��a�c�ޣo��w��}�������0���6�{��x-*��p��,�f�HIc~¾���D#�`2���~�l�Ɣ�<ռ��yϻ��E�]�mo���}�B��E�\�������}�o<�U�z��I1I�A�\ b ���҂sA����{�f V8�����t1�:I�,��NKj���=+4����� �2�����6d�l�5���_��?��?�{�W?�_~�9���_���E/�|.�B�F�f��Ks�
���z<��Z&y�R!�6�g���IIJb�b���!s9�m�p�m�oQ
���A����/��zы^��v���a?]�I*M��&�(��L��I�$(X5����11�&IE�{��.p�w�?��l��i�&��i���5K�-.\���]���^��G��U7��n��C?�C/|�k_{�?�~�~g*�Ux���wk�kH�-��N�]��w	�ҹ��wL���e��ۆ
�$H�V��q=�
��o��ߵ����Eҫ^��>�s>�3?��=� i{�}�u'$�4픲i���,�0e�n-��)f-
�G�\��2.�/h֬9�^������u�~��n������;t���S�<�я~�?�矾`y�'��u����(�<����5��
����ލ�".�V�����?q�y�n�R�$)���d.��z��^��!�ɢ�yMO��{�����z��~��v!W08��qaݛ�Ș�jJ�R�M��	�%̬d�C]w"q�D俕�O�D�e��m$G�M�����3��F�����$��_��_��_��_|��H�g<�??�������^�Q�l�6:Kia\��5/B9�kcNoQ�Ď�?�w��Ʉ3B�->���8�U�먃�[�ü5�\Sd�i/�����͸5��1����>��o~+\97�O����j���E^٨��J9˛2_��5@���O���	���psc�nnv��JU0E-�2g��i��x'87�߬���/}�7�|�������?�����3����P�
Z\8�8n��^��Y�-��D�\e{3��Ɠ�\lE
��f↋��������X���;-������؍_�4+���1��S��ԧXf}�C&��x�������>����\��2P�����*tV���:s�-�>���#_���-��~����[�M����z�n/k_�b%�~Bw�#����<���]2��ծ��?�{����}��/�{^)�L����r�i���~o�^'��U�R|"d�-��{�&Ďy Vh��%��E��̞�Mˤg��V��_�̯��W�f�'��H�&�>��x��ӧ��O}���z�����VV}�Qf܂+Cw��mS�hF�kJ�&��
'ziž�Յ5��]h�V0�D�����J�Ӱq^��eJ�����'?�Y?��?��K�����o?���s'�����9�1oIñIyp��l�=������a��2cA�$���i��H�V)E��֤R��'�I�st`�?���K�Q�U�o�~��;�O~�S���O��_�K��=�y?��?��e��F�D������fI�5s��2�,���LP�����K�.��A� L���I:Ŭ��k;�ڮ�v���i�)|�?����G~�W��-�|͎��E��G>�on���������7��?`�*���
Vc7i�.BwF�l�iQ�X]�f�����@��si�%��<d<��A�?\&^n�{�3ΔU��<I*��UVU�%	&��n8v|�}�?�����3���_��M.u��������m��������5��<#��6�eS����ӹ58��If�a+�3�϶�O�`��K�2+���Q�3���p ��M�����[�ޤн����lZ-��ƃi1ͧ�Y����3>��}��G��½$�G��~�����׽�ɺ,-�,�3]e1_xbr;�*��/���R��c�j;M� �c"�Z��욎ϯ�й�k&O�ާ<�ko�m�����<y�cǎm���o�>ٔ�t�ѣG�_������x��~뷝?~��(+\i��j5�Gt` ��0�:u��#�vXF`7�ֈ��>gXD�)�jB�	k��a�G��aF�M<8z����L�A�ΥN��@���5�}�c��n�Omn��ӟ��	iY����V��佔��]�:��'�ц] �NC����;��>4��3�Luaet��~���z�2�����f�Pm=�k��>��\�����<�_�җ�~�[��H��z�۵�Sr��.5��[chV��$߷o�T���%���ٔ����M�����a.�̶�������}�g~���G|囷��O����П���_��C�=�A�ۇ^�g��5{�+^�_����ufC��+�<���w�f)<�k��?�S����~��~�������zֳ�ޒ��|��|����X����Yk��X���@5��� ��k+�,���z�w����7o�{x�K^�,��M�b>��7������|�^�� aX_I֎�r��Y����o��'�� e�K����?��x��|�����hE�ǣ���wWeo`u�~����#�V(��&јS֚�ݕ�RN,Yޢ�́����ڭ��閆�����O}�ÿ����_��7�tӻ�9"�G��M���w���_��o�/4%��Ps$�����s��/��	�y�;��������@$��dt~Lu�X��!��zhA<�)O��'<�Y?VOJc��u����޵�zG�V�ۻ��qN~����>�+Xو����U\z7����VAϚ��_�������zoӗ.�.���VU�K��\,�jҨ�N7��/��v������ё#��sg(s�p��tc�N���D|)�J1�b7���B��傂��Cs5�Ч�Iƭ7�ΰpF�U�]��x�~�ԩS_t�w�h�Z������c�?~�����-�?XZ~��n�,��1�ǹ����B�a�� '���x��=������=�{��g��l����l�w�D�������p sS�z�|d�@��K7l@
����ǲ�qN�����0�G�1E��P����d�F$����w��ǘ��|�/�acժ�KX���L�+�
Wb�Ef�8�i�b���\;Q�-��xm���\z�w_�AR�y��(���Knx{���b?��3��E�֎G?�u7��x�+��t�yA\�  ig;&c$�Ħ%,/���v����B��FI�EM�01�O�ʑ�|��"��:t���á՘�\9wxf�q�m����I��~v|���)�t>J�t�a�1��%I"!�?�_�\%��6\:b�duu���I�2���n��� �<�B5f� �'�M��@��N���ln	x��b*���p��cP��qUTI�B����%%�$%P؉�(^����q��C���%���o1K�@�0��xwL���8YPW�= �B8�}܏�_7`+��Qi`I�+�%����0�"	pqJv�nP2և��$�j����DD��Q1�9�	
 S�68�PQ��qLniطW�F5|"�C���1wM �t��7�5�H�-�~_Q�i���W���Y������Ւ�6{���2�G���@a��W?J5��\�b�)�@A�+cRfn�l-e�]Cp���t_��v�C/'�TmI	��k����4)_�0^��:�5R�b\���\%�� Z����5z�fgG�L���Y�B��˯�4���{�<N|�$W��	��D��p��Jy��I���tTCJ�A�(b��LT�����tYȗ�.� �>�˧o���A�9
3%��e9DD(�j��kE%�-ɵ�s�B$̺��uef��ۂ#@8�Y�u�5Z��'#��biO��T5�5��9č��OVi��$EM�vo �������R�;l>)Y,���65?&��/�fD���}�&5�����	�2��)ʇ�k��c[׊ s�m��=�M8�sk�B$�����
��x���48w�Cd�:�u��1�mɬj����[��?6��y�]����+�M ��[����2�~#��&V$f� eDB�^2��vj���S�T���Kͣ�"�򼧉�]����uks�DB�<�bP�
���vD��zJ�����]�#�:������vT�լ��6\"��W��jǬ��̃�9�X�4���Iʣ˗wD�4FB|wF���b�܋6�ZJ�,�S�6e�j+
߼P�g�����hҮ�Ty哐wK��V�Y���b�",�ʨ������2�W�51k�P��>�>3k?��Fw>�NW�1�x<aq} 	Ҟ�@�����0'1�"��UQ�O!s	-A�P}0|�h�e`Ӱ��EVt���d�W4q�� =/U׻�"p]I9I��o�6��ì�f��x��Zu`)Vf����|�9~��#�ՠ$M}��y�dK����G���`LSrl���AaE�+F����
N�q��=Wz���P��=l �fi4�zu����1M��9rg;���u�b�(�\=n�,�M;AR�921����Y�=� ��n%�L�S>��� cL��G��ǤyЬ����J��5C�9�=�(�\k��h�f�1��H���_w]IA�Bg
[Ca���rI�x]���_�0����yU����1i�V��@����N�����|t\ؼ�}o��)���K_��Ӳ�}ة����z�����zve�>{�q��m�2��@"�NJ;��3$�
0Zm�5_o-����p�&��Du�	��wY�|`+���Y��gU����E#5�^r��B�f�H�9��n��%':�}����$��
�]�����N̺K���'WD8�	�F؈F�^+�^^�O��̋�� *ͺ���n�K7�F*NP�4��k���Q_IعP���ҏ��/K{%S=|�{#�ǐ���{�p��4+(~S�A�ig*������.���u:Ȯ��d29�XC_��1�_�K[�jd��>�fm�`��u�7�I�C=�����f�M��i
�y�rR�+u����b���M��Vv>�t�� Ɠ������Q�گ%je\�� H�z� �o�L "�{���JUM�%�5�:�`8��+/���4���7Ȭ�2`N{U�Hn��ͱ��ګ�6�Zk�1�h���W��M&7�����k�U�1`4�wZ�I���'�V�0�&�?GDV;��;ԨPD���L��R���`J�t�\�)Z�O�:? ]<�d��Q1���3e���P:f@����u���ì�I|ƀjN�l�:����䈏Ygy^i�=U�j�X��N�.��ʷ���ǒ5��2�ds'�- n����d Y3����`;�Z�����#��Ԕ�¨6�}��l�6S�����UXgyQ��4*7����E@�{��E��.ʫ��u�Y�+Н��Z�������r>h���؟r��CaJ�N��2�ϳ%�U��E����:��	eY^����HP:_��!3��T��B,
�^/�}ʐ��US�����/ j�.����a�2<SU[A졻�ï��W(��o�^=� �AM�g�矆$�u��#����E2kBr ՙĚv��4�B��m�3� "����Ϧ�r�����F�BY��*o����E*Y��s˃X)νvݵS���0�$�F�bJUOzf�C
1�0��$��Y�@���VC�L��0��p��.	,��ɽW�r�" ]{�g���e;��Sj�K&b�6��N��D(UP��%Y��ڭJ�qV��?["0��il9:�9�"�{{�)2�b�F�g��h��y�v\�VTQNU�x�5?O][�A/�����""k1Q���|�)U��&��"w.㔣���X���C�8�B4.M0p��C����$�+H s��zjN���E(�Gx&Ap���`m�N�!pŚ��-��:�bV\=E1ƞbn�AC��w��Q��e22�5�P>�J��5�Ц��A��ܐ�ҬM\@N*���N ����� �3�rSi��7�Q�?��uAfD��V�q3���b-�.�Ҽ��
�wd^\�7O�����*��	��3�7�J5㻸���@��A�d%��gmL]���ɷ���uQe���\"�e���b�������M�F�����#E�}"v�$J�nv��_�?��5�U�76��XY^^�;U�ᚻJ7!Y��l��P��[���F|���#��vTq������j��!��Ƨ��d3v{���)�#f����[�Z�����z|ťY+��*��qB:��c�I\r	���!�ng��q����h�BZ^]>/�;Uk��׶�V+	��޹]�ϷHA/B����<uvr��!�}����c�?M��+P�f=X1k&ƥ�8	f8��@�"X���Ar��D>M���\I9�3�f:2΃�����P��-�;��6y���pZf�6yU�Q�6����w���D���^S��	E4��~�%�{��!i��/ �LT9�����K�_���� w�4�H�z���l2�"J�i�5�b��Pk'�/�5k�FŬ�<���{�q�D0�!&�A\JxPiU�=�S�A��*�f�O��p]�,�ʹ9�֪j�1��6�X��2v/̒�/E��+��I�J���)ܞ�1q��TB��]g 8�����v�4��e5�z� !5 R�͎�����'�<*,�z�IR�1͓�3�)&4в�Fs���=oR:���x�k˩y==�fy���*F�����u)U<������a���U�:D&��>Z՝~�TT5n`Dfm��CW��F���Z����[ 55�Sɼ��\3�f�$�F�&s�@ˤq�c�Z|�`�j�[���ed�2^$����i��e�i�E���d<����}���b���BI�
��V(vC��׋�8���M�05i�7"��}��z¨��mM]b�Ճ��u�}T����AFG�_�iׄ,ftT��t��K\���&$/l傉)Kl,s�C�$�5�	���f��&`���}]�9I\2ej!�n
{��G���{���׆���tP�F8��ަ�w��R�SS���@	0 ��j�����)b��c�
U�|\Q����⦵���]=� Z��� *{��K(41k�mթF�4�[� �����]ÁG��T���;���mkU���g�{i>���L.սƂ:����9tq�?W/F�Fw�U��b�e?�Y3���S��;�2N��z�bV	�\�&��E���y?up(L¤M��V����td����ǅ"���!�d�M��p������,p� �R���8݋K��ć�;o�b�ϬCP#�vz���}��RQ���ϧ`R�b���T3��,r�!�d�P��S�v/�Z/((���0��!ZLd�{��=z��|ō����55��ƪR��k��(!	n-���¨��>��܌*�8��4���w�<\ￗ�C-hH�Qy�z�t�[��B�K8r<k��<�i��/o�2�:�kg=R�W�������>?Ȭw�z��;jf����MSs�:FK�u�r�:��Jg3�Y��0�k�[E"�ok4���_�϶��v���^@W:�}l�X�͛_]z?�6��f\Zf4ӧ�$�c�.���I�[����*�ڛ�s�2�;QHk����� ��|֩�N�'a�Z`B5(dt���r6r�r@��y�����Y�`���B�ZZ���{��]+E�K�J������,	�n:p�v�X8NkY�\=sߢ*�����\,Yj��լ���<�B�M\u1���	���`�,2�F�N�&�Pܭ����8���ʏ@�ˇ�
|����:�ƕS�)EU�w2�v��h��mMn]E����)k�p�����	�o����w	χ�Զ�C��2���20{ĬKc���
P�	1����L�'%&��c���\ݗ��
 �\�U�%LJ�����\��q�Z[㗭oM��Klf�3*8X<���<㴼��KM`��eK�����M��������e�J�U��NWmAI����D�����b4�Qs`1��Z�;lrR��z��c���l!�rN�Lx�7?���VL�l��߃)L!&ҹ�h��H	v����)��KR��Օ��֬��o	MT�ɘ�β^��yj�����5j%;B�t��@��Q� �DU��{��3`Ww�,XQ�������Q.ZU�BX�}<G��d�W���<Kn7.��I0��J�k:a�(�,����1�7�ƛ0+P�}�Sd� ���!�Ui�fV ��z����T����)�F�c�pqCIwR�q'ί�Ȯ��p����*�`ˎ�3߾�=�N�H\�'���YY��ˢ����·:J��r/º²�
j�ɩw��j���$Ep��|�Y��NM% \jH	5��lDi2> .�H�{��ر���1ox��r�+�JƊ5k��4k���C�n	/o��W��fV��F+���t�p��OG��u_���1n$R�|���^@��<2	$ˈ�D�?�J�[pu�����3������7B�8�II�3���uAP����2\o�+V���+WuYRy���:ޫ�c���vWpr�HK�n?�� ��o�СK\�-���j�g�$���P��K%����Ũ�q����=���,�Ĭ��z����A���Y�ԽB��
�yo*� u��?S#e�"6 �c����Jb7Ѻ:�4����A{�%����FI�bFG�mz)Tѧ��LZ;�n`yKZ�s�$��.��evXB�KN�׼�����]�qþ���UI�͕����}ii�����H�^c+���S�&#������3$�#�y7DB�,���έc���yWn ���:�fmn����'&Ē��.3@5sr�� ���4k�4J�	C�ldH�f�`�Fqƨ3N
;F���M.�$�HaΓ�ulB���V:T��^���&�u%c%�ZG��v=�[�ޮk Ƚe�����7ڧo�Hh��|����㬏p?{7��d�U*{�ԩu�����=S�1�Y�V���5?��b���g��|ȯWwO�&̓C3��Id����̊��,�W\�D���K����^�Xy6��H��	\�F�N�#��1�ض�U4����^��(Xj.�0�;�:�����Yc&u!�t�2fn��ͤ�e	�҇��-Cn���Yqƃ����a~c�zW��fme���`X��f��]������ĕ��g�,Zq������)U$� J���5'>0��r��lbaPU[��;��{.���E����Ɓ��g4���(��������"u���4��އq�6S�i���U_�Z�7�TG3c���RIP_�fR�����x%�R.#�R�61��
PQ�5�Q����P����|2�����[�=�>��p؃3gp���"�����(�X�ࡪ�:D@��Om\�񬍁�r���Č�x��:$�2%�O87+++��v>���4�;�Z��Y����RM58�@2v�㺒K.b�޹A��m�_����$)cc�H�w��m7�o3dfu�2��Qi_D��S=�\�Fmufm*�tQ10a�zq���$�l6��N�gX�c��5��*2�O�(R�_�<xw_�4La����Y'�/7Q�������CRu��R�� U3��J�FJ�����,�����lFu�M��TJ5��HV���P+**����FU͚{�[�ֵ��**���_� y���V�1�|k������p٫S�0�X����~�H:E�!.���?��A����CUn������t"�C����Ü��L�p�fCťn&I:�C���M�F:�t(*QQYM�vϕ�C��p����k]E������Z� WJ�X�˜�T���.��l3a*ۮ RU]<"Qi�N�4Ԙ��}k+�cޜ֮����B����"�Ot��.k�;�J۴�Mܫ:�u��LT� i���VK;�^��۽�A��� �^�}�ɜ�6T6yOk����zz���T��U����>�,.lG-,���0�1�q�:*��e���X&��U㸚�b�y�l�MW�[w��Q��$�t�_<�� c�P�ұ���+l��
ù��Pok�\
�V�P�����e�Ѵ�[�7�^I��H}�H>��%{���0k]G�M���n�� -Т=)m�E�KP�ЭI�� T55k��b։J�rd�Z����B%�����})u���ڢ�<���9^A1�]v��=c��^-@���r�O�74H/DF��B�KI��BDQ�$8��tZxdE18�d&�b�� �*�qKi68\��5��gm�͢K�P���n+׷�QT��n�:$m�g�~8�̮<R�#�M��@��fp� �J���.�bF��*�P���/����f�ㄲ��:j8��A�+/��2��(ah�t^̢s�$I����²4�$c��tV�����\���

bl6:\N9O��i�*(CWΚ�J�LG�ǵ;w�� �e]�	��)�6a��	ؑ�$\(���,.��ʦ�B�~
����u2iڊ8�j�Y�;{6�uER��uiװ�ۑ>�+V�6�����,�ƹ:)!�gPN��n5�D3��IWKj0#OVNN�J�s�p�����A��NG��F�n��@�Q��HV�R�L���ycB-�a����k��WYQ!���3e�B�'��"��i;�(�AU�QY�vtu
��O;��e\]C�td��N� �ޥf:�83$��a~27-\��xd�����$i�9��&��
��u�r|�lR����qu�fT~M$�=�	�?`ְh�ZAd��jcf�� ��R ��[@�ZǕ�W%�(�Q��̈�_gNSLb<�Ӱ��W.���9u��š�Go���'Ϛ�\.M�p�;����|)i,�Y�=�}����])���Pρ+Վn�Y��w�C�$�Q�,���g�sa�)�4���ο]$���e�p��^> ���F�m��z�YR߾.i�Q��bz�;��e6H)�m낮�t�(z|ɴQ�� Z`����4�여�_R�-���>����Q�M(�+Ijm��o"�<W��Pw+��p�vm�s]��MB����"jݜ �NP�8�L��U�g�,���ζf]��(g��ߕ������P�=/�i�p�r eiJ�
�4rĩ{�4Q���<;?��%s���X�mdڦ�=T�pqLi��3R��.;B2}b#��d=��8�T�F"�ΨY���g��a�yj:�m�o����WPE�ə�V#�U3nC':�d����Aϰv�9P�Ŭ�l]k	}�]���ȼ�4�jSV�`��`U]�`�����f�f�7�3���ą�hv��y{�Y�&ѷ�� ���P*��O��E\��gf�X��q���x�#���c�x-�*����I �M!�MLd���3������Yt��O��TZJ���lW��\��+ծ<k�"���ƃ/d򭁱b��7�Z�f��Zi�k@kC��W�(9��tT0�5
�J;\��� �å����M;S�g�u��`��w�o�����ky�L֬q��_���9��r�N���L�]G�޷�,�
1��e���Dd�kl�`�®�	�>���{ʽ�^�a� dC(�qK�{�r�Z�Ip�b��C���WS6��$�"���6+0sf�᠔rL�kf*��a��A4"|��ZNs��sf֩�D�Uyq(A�}Tc��m �X�������@�U�b�TC����*j���eE�գYS�K��h8�:L��cn���4*�đA�OmNUAnj�����e+_�^{�\r:�g D5^;�i;�+D�co�5�f�qP���7�.�Y#6J�[�#�7�<*�d���+��1t�/�t��H��}%�� �oZ�G��|�J"�H�wZ�㫳_i���K�*��9�z�p��U\Ht�T�����)�~�����&^���2�r��)K&E\��I�g�jE�"I䀜�6>�."kQ\=�� �T�����ȺT�E�BJ�ZUJ��@+��	j��q��ß$j�.U3�]�$�>��lz"")�	�"�A�� c��J]T=�i���y���b�)$���n��Ta3�g�T���|քR?7;�۰l��/�Ԋ��ڴ$W&j^I]
ɘf���.a��=n]ؼ�he����ٰ��F:�>]Q���eg��� "�i����6n�XX��e\�:O6A e��S��W�Vjw�3ʒh�KD�Yc_A���h!��J=�)C��(�b�\\M�d�N�D����@��F��^��5�ݷ�p�V#�R�<�s|<ړ���·��y�YT�:��{�u���[_�$�����e�-
�?��^��F#o9���P�L
~lf�0�d���}�dh$���`��5$��ԫ�:�9@����yJ�GNP�����0j6���R�����ۂ-�rA�y����,�QJc�Q���e���X�i���§�ֈ���HM���˾�{�0�d�rk˖����8֎�D �LY�6�P5I�Ҏ�
�0�ReR|�@`ٝ�ژ6�ә�b(���g���d|���,3e�����2��FS��K`c�BT ��.���N%P���Rt�ql���k�F{^4S͒z�e��wc&��3���\�f �JEW���2L��QaZ�,k�{k-^�f.PꄭV�W9�L���-��L+X�/�1�WO6&KKK�(��d���O�zCc	2� F�T��9�E�����e`牄5�э�&�4;��
��W�xeS�����bTE�E��T��댣MS��)�Aʞ����$*� �JsJ�$��.�DTT
a�e��dDg����"*���&Z���85%� 2N��?SC���y}�"f�6�ɏ��Q��%A��P;!40l��Z2�e3j�{����ևu| ���6I5��+8S���ƚ��L�_��͗��u�2��Z�BG�͞�$3+�*�р������
`���p��"Л�B�u�~IW��y8��*F�
51�L ޓ�N�O�!J5L���D�A��Cǲ� va�E_v�{K��s�����I_VS�d��{�M�F�m�2$@E���l#,��:X��BA�P�RW@���l��2�1�ħZ+��۬��O�Εnv���YGӋ1M��ǇPNʴr��$ 8�,��O�]'�͝]Ѧ֨�4O������'˒u���ϋ���X%�	�;�k���Y!�V�Y����W��S��О1E����v�z��V�9Y���=�����OmS�ˮA���	DB�0ߤ�C�}U0��$�
T%i�Wͧ*��a��<G���eozF��!m��EAa�_��z0HP���I��V�
���ϾR8�{Yn��S�(���it�J�
.2σ�o����* �8w���P29'uƗ���Ҫ��(���3PU*�6TI���2y-�e��f�E%|�(�Ҭ��������IKހ����w�UĬAM�p:
���9%����,-(��Zk��5��Qi$��E������'�)����t��:��h��$fk6����֩RE��x�$%�4�v�k���,�v�(�N�A�eS��qk��TcN�*ut�r��1�4�(�%�(��"5����sx�:ª>{߆�S�|z	H�ily�i�Ofq��X���/��)���ɘU��µՅ�o&0��0�52%�_h�30�`�Uhj�b�R0�e������,*f���GU5mח���Z��%�.=r�s���w�>w""to��=EEf(�&��r6��XE�4U�����^v���1{I��������A7f��9�rS=��N���UU��U�?���kmj����n���L�Qe0���rzWz�E�+H�r�$�:�/"�ƣ���
����B,�z��y���8�����l����u�{`�I�L3v�z��H�y�j��."��W��4k�A�=˨�%�ů�b��O�@l���rq$��!���$ޢ0�#�1뻢�ىJ�d,Z\MtE�������,��T$�|��#�`dʎ'���f��k�z�����c��^��ܼo�����kyME�f��E��h]k{�&�OAG�Y�b�T���'/�_W�:���h3:����kz���#�i*z�:��|���,�0k_�0�.�W����)�K��P�'q�L����敗��
�=�H��9�e�Ę�g�������	�������"j$=�S����ո�zQ�e��Y��:����	u�Ȣb�&S���JC좰��^�� I�8�n�@j�����>��uuY�/{���v�����"�a�Qљ�v��!�;W� ��"�YC��*��ؑB����6:���.��PC��u�0��O�A$����z>�2��7.>i�Uݹ��Ww�jW]���6	��l��׽d��D^$�ib�z����QM�+��5p�ք˳�zb���>N���m�VU��΢H#t� A	x��]�m9+��??��ɳR4�P��^ 7ֲ����6N!O��)�)�����S��U�Y��lc���=�z��L��[�{50�@�+��WS�
Y��;�������T��I;� B��N���5��\ �{Kvo���I�� �)^�/��]]�=��ь�CkFUNn�v&iq�VUdJ��q���\}�)c�b�_�T��)+�,���}Ϙu��g%��jkfSH3E1(3�����;��:��+I�&����T}_�������Y1�A}wc�p�ˊƅA�u@>�!�mPU3H�+�Ŵ��Y�Xi}�!(I,ܜ� ���[�������Tڃ<�gaF���t4��Y�=�m�Kq.¹�6���"	gMTU؆p6�A�2�T���q��f_1��@�q���t�P�v�J�����f�;���\��k��~>�xDUT�9">�$(pS�cڳ�`=Zei�i�q�,Dˣ�u={�777N\�{ݻ�=�'Y��)�P��ƞ�I!��f/.����I�/����b���㣇�H�f�>�6ס7���˼�ə.��4��N�hF��ح�2b��U3<��X`2��/S���f�pڋ��0y�ݧ,[�����:�}�f�ٖ�䓵��լp_�)?��^�u��Ԏ��jT��Ҳ�_9��b2���oX��Y�LVV�j�n�O��d�-����¦T0�k=���߷ʆ��h��4�x�����&گS�tTŌ�2��M�p�(�&ܔ ��kj��l��w�1_�"�=c֖ݹ�y��z�Q�fbXef2���-mm����(˨Ϟۀ�nx�y�����A.��W���e{��2s����o+��PC���S`�Ш�J)}�{�a����C��*�X�}k)�y�irwl\8����H�ah7���#�\K�+�����\����$j]�m3�\��Vs��`��Ԯ9��2��yW���5~����A��m����2e{��Ϝ��զUF66.��w}�W�Y�{���!2ڜL>���~ ����6X^��*�1�5��ڲ{{L���~0\s��WS{v�����%�]*��Z'������\Ék��.,n�sk�vY���Ο?�OO�v2
��~��v>��	���,;u�m���}����y[�D��vm�g�tn��Lh>ruca���*3�Ul�u��g��_���[>Ǯ9l�Ю���O��ͮ��=�þ�%�暣p����`	��&:AlW磣��g��kT����zH-�.�h4��n��C��!�"��=:=������9x�`�
�5��S�V�Z���-��2��<����O���M��V������kV����gd�@����PڴV�p��>8t��~��
Q�I~Y��1k]�O�>}��k^7�p�w�I���k�6��U�*X[[�{��'N^ǎ�
K�2��DFv�n��> ��`���Y��[3x:�z�� �t��{�X�[�kg΢"���-�+DF'N\��믿���i���'OBi�ׇ>�a�0A뢘X��Ǯ��0���NX�ճ�L�$O�w����çf7��j��~�L8k�1Cf���f���#F�a��7�&���<���c!��?����߷���'g�58|`��+�=�N��QӾ��Q��*�����K�V�eѠ
�,�� >���U����VWV�������©Sg���c��A�|��b�����e��{��g���߿�7�Z	jVh>��&F����df;��"�軥&�`��di"����~�x�?�;�̇|
�����&U��/p��=p���8�~ۇ��?����a8|��{!2O��'���>�Ϻ��O�c������cǩ7����a߾}���aH�>�it����gϟ�w��x�;�
g�:^=F�!��L��ѧ��-�b���&��x�gZ��k��#�n��&�i��w�MV�^�n8��6{�s�a�s��MG"�����DfF`o����
���OW�}7�5ް|�ܺ� �!W�;����f�Ї~�U������+��aȞ1�����j��S��p���`m*�y}�j6�H�K�p 5�'�����we�q�U��{����W{V�d;��8j�%j�Z�FE*TPx�P�ԇJP�� <�(��
B�R�B*!�DtK�$m�6i�ر�-��g���{�.��x`�bG���3Y���?�|g�#���m�ؗ핍��t[m��Z�:�c�6�#,,,0OBA�977�J�8�i[J��$���,=�c����d}��)o�]�z�,�+�Ifw�>JDi�ѭ\]�5��A�F��Do�	�x��Ul�gJ�aHٚ�c�.[�ؠ���B���Nx��Wa�\DٜFr�b�ڳc�0$�t�.K�ضcg@o/D�N����}���oH�����2��CGkC>_�R�-4�$ˁ�w[�Ԗ)k�4[�����,\�e��Q6�*4�}H�Z�@l|�(�2�.�o��Z�;fMÍ|>�511�����/@�Tܘ���y�g�����ː������ �3NJ��w�:�M��p� ]Mc�\�߇�l��"�l �v�T��sܱ/E����ڨ�3�X��DO�b��l��o�A/c���p_'�L1���]���@�X����
E� ������R]�]�FH���(x�FJ,S�D�zARֱ*d���d��Y��b1�TƬ�|B� c��M2�aI�ְϖ)kE����W��E�C ED��]__���cU��魎�.�ՅDk[���
��3��|}m��2i��[;%*(u��i�z���������/�K�)���2浼433��l�Y�m��@vf#��8.�Bi}��U����#�tN���K� ���IbY�1vMkc����p(@��Y��f�з,��&�8F�fp0���`��Z[[Ce��G���-m4�=t��6W24�*���gzav���G���݃{��=G��2�a�h�ɴ�7F�V�o?�����XZ\����̍���-��l:�ͽ����-en�#�D����5�}��\���1X]���OKm���<��0:2Ƅ`b|T�]跌m^~-��*���O$������J%��i0�5~���"Kf<(��U*/\��[�Ǔp��7᝷OC<�L.�p���&�~߃�C�U�P>�)��3h�.Q�%?TB�B(ó\e�!�,�)YN��+�����w��I�)Aĵ,-^�*��S7A1��8r�rQ���5j5i4;����3������k�]��O�L]l�#=8����Y����:p��~�d�f�O`�MUU�o˨�$�5A�d:gN���X8ǁR1�J��X]�(�{ｌ�L��V����-Ӗ*�!�P���B�RiP*ՙ'�T�&zL��#��j=�l�5O���KO�#�k���\��1)�S�V��D�(�@ ����P'Y%���˴,���,�ԩ���敹Kh�S@�^i���g�Omd������zd����pQ�x;�'U��۷Dj�D�<3üa�Ӟ��?YA�� A�a��Z��u���̝?��ֵw�!������F(�«�;�r {cnee�k�؄(HUI�<1M'N���<K�К�t���z�a�CO�]��Ϟ~�Ş��fr9��K�V�̓�9�Z��6���My%����c�!{����"P,ae�*�Pi��(-�D6�D"����;Q |Ъ6�G�Z�;�{������7�cI5	I�
$�"��Y���'��`;�E�F%lc��V�� �m�BPw&9���h�Qg)a��ս=���uK�~6����t�3]�"�6j���2c#���W�(j�������=�N�HWkk{ӃYh�V]X��T��R?
x¡�=���F�_NO$�WWZߢ�1hbb�i�ݙl<� jW?2Q��s'��#�Ė�P����2tz]�`�C���=���Ft+	�ΐJ����~�OC���v�����/{(�����F�Z���Ey���j��=�!�������N�7j�tv�f0���fBS��i���Qf= ���n��Tjh[���TY�"�Ο~���Ţ�4e��h�{�"�ϛ�	ɲٶ��ܳ�)��̯jWW�m9��:�ݞ��X5��H��A�V����378�$p�r8���܅G{�^�:���&r6n��5U	8�jbr��q��d"����<�@B&�A���8�kq)�Fg��4�-yO���lvh���ѱ�}��#���$1�zL�no�j�k�)�t��9F�i��ߌ���h\뵥�/�w��*�"*�$I�^����$�a�ꣁ�A�0�׏�����ny<mx��Z�~�Z��YgPG��C��/%iRɓ��2�M�˳�N�����c]dQ������M3��]ݮ
�Y��z���1(N?���Ϯ���)�A��"U|����Y����W	7�y��)���S�N<^Ǜ��=Ȱ6ΰ@��	�͘X(�k	^�9����l�X���:�����_kZ��2-��H�Ǫ���+�)��k��9��+��clN���-p�n���H S_�D�A�ڃ���>�k��=�\Y���s�N���S�?d�8��ʙh$��ИM�O��h��!��
���7�n5*^�PO�7��
�������J��p��`�'3���k]� �!6U�5ꆅ��n=�tlݑ^�ڑ���Џ.�<�E��n�LA�}�.�e��%�����O%+�?�"]?9��k?�p�'�KW�RT����5{d�bC`:h����I�ew|ꎯ���æ{�[*%��	��#t[-Qm4$ɣ�~ꡇ$��e���d����7*�V�ۨ���-�|�dJm�z���,�/��%p!Y?{敧�=�S�E�+ʲ%����ɖa~����>7 ";/���}Z�'m���=�i=_7S�(h���Ht5_L�8����?^�t���נ���-�����D��@j�6�2��w�0���]��c���]^��^���IJۦ��>��4m�q��܆.7�ƖJ,o�O���S���mQ����<���'ػ��������c�~n$�;N��I��!��;'_��z��@Ϡ�6��-����v��T�.���'A��_|0�}���A�1��-�dE^�$iy �~7�-��F���1�3��u��zb�P�-U=^����fX�Dɰd�4o�eA�����%����@��k_���v������O���9W�;�
�ӫ���5���]��F��|�n�>�*k.\�� ��v��*k.\�� ��v��*k.\�� ��v��*k.\�� �r�$�    IEND�B`�PK   Ŧ�X��~��K  yK  /   images/7ac84256-6e9c-40ba-9a9b-c812e48c1c94.png 8@ǿ�PNG

   IHDR   J   �   q�   	pHYs  �  ��+  K+IDATx���dוvߚk�U�V������I��9�)��5�%�!+�X�
E؊����H1�P8�3�0G�Br@ ��. �n4���k鮽r�|����w2���*k&�_ċNd�[�=����s\�6R��Fl�Ԉ�W���
P#�_j��7�'�|�E�ق���/�v\��b\.[�0��(j{��ݮ��~�'��a��'D�8���L�X,������F�X(Xnōb��@��>+��Z`Y���o�ߧ_�$CG�������;<ϋq=}�8^.��t��j��gϞ���P���7^����JG�������lGD��8AD��-
m|�:������0�H\7���4d;j��n�Vw�^/8}b�Y��6V��g>�~�Z,��ٹ����v�^w	�v�N�D6���n	�q��§O����88n{	MN�t^Xbbb*�T*�f�V���w�y��^|��W	���Qo������Ӌ�67�.	+�H���-:�]�,���+�����ZM�z=A�)�Nt	�k��K�繞399e�54��	��	�b[� ��H�c�V,ױ
���Yx_��4o��c�Fkkk�����|����C=t���2v@� ��������?|�l%O޿w��๾Ł:�F��")y���3lT`��W����q�0G~p��@���1�C��V�����-7�����s��1�[�:33[��:Ͻ��W���㍱�^�������	 �'��nz�D��s�P3`���&Q�u �9\ 2�@8ƀ���}yK�lv����!ە��ͺ�y�x�ɋ����bcsm��?x�?�ͯ`���Fc�D����O��?y��h,Z'OJ����b�d��1|� `�)�J�����ku�a 2@������̀�c��h��=���c(�*oz�hܚ��!�H��ck����Go޸񟀜677�_�]���e'W~�B�����m�s!�����@���D��6�.*���ꀑ3�R�E$'l~~V��m��a����+ݼ{u1I.�X��� ��ݻ���~�[]�����[���?�C �sӁ)ÇIPo<@�E����0�>�f �տ/�����*@��KR�,.Y/��[(��7�_?�&O]#��s����<��/^��������w:	�V���xB�Q�����|)V$C���.��d��C��k���p���q�p��
b�uR&��.\����o~�_?���,��H�4�N�\	���zl[wH'�: _jY+��x��a��%��]&f�uyM���L�����'O% ���$�c�*Ւ�h4'����!ځ����>�i�T*.�{�J�x��k�6I�';�D�������>p�ɀ��2���ߺ^�N(���y&&��C�'�J�����uq6��S@�3��۬?N/j��Hk�(�E	u$�(��>h,�pÚNF]��a�����x���xO�X�~�������X�Ei	P��եwm��������c �-��t����*�ɀ�&�ӱ��Iəb6�t,�$o�>��Fԣ=�_�Z�FcO"2/�+�juR��!�N]d�����W����˓��w���Ki�6�v�t�굯8��.�,Fl#ꩧ����O^+|�;��f��\��l*���5�9�	�+��fj�\�@��]
VM�X^�;y���/��L�E��d���0p[����o�֍ۏ�KU�%;��v����ot��C�Y�Ӌt��ӟ\��
y>���S!���v��t7����1*�FTڼ�O,]��҃H�t�֓VV��Ԅ�Z��p��:�M�Dc����[�uO�<�%��dfj�3�! ���@�RGI8��h�+���y�� �f�纮���J���3s~����^Z�$����7;��8�|-��ցi��I�y6��t=}Vڒ�m�و7������N�'!ѻ#i�����h�dJ1s�N6���_���=y-���$C귷��Q��t���#�����������<�	�.���}r�0��� ��3������&��{�o�%`?�`�>�����/<лN���{�����8q���g�ݤو,;qڝ�2܁���u��Àh2�<�1������y	 |0��ϟ�?���?x��W-����b��~�����������m[	�S*D�\Q��������wl��̦�$�Ml��3�R�jU*��a����텅ʺ8D�gn߼�q�0)M��I�
�S��<���%�os�y�K���1/Ͽ��Ǥ�0_�t�+:��a$�Fe���D5���-�t ;���n]y,�!}&�7�ә�0�ӥLr�X�X�k ��FJ�M��,,,�^'�}��v;��&�:[�̱^o�v^o��2�9�0K������~��}��*'�V프�8�R�h�N�G��X�-0�^��8}]�� ���n�q3=��[&6Je�u2�t�>��G�w���G�wH6���z��&����ba[��#���^^m)���ޕk}[.�<�[�]gz����c��ԑt��9$*����G-�aB��N-��+��͂~ml4lzy/١3�Qʕ��Ey��,S9�3viP��G�	H�c�O�(����0�K�����Q
����ٴ,;�{��R���?�@�ac����"�����!�h`�a. 433#*�
t)�/�V$#T�;ׯ�7o�|Ĳ]F�-[D9�f2���%|C"��^�0�.9�=�49���-$4�
�q�L޸q��	��+++�:u�5
F���M�O������œ'OK�y�R%�W�s�~��δ����;5b��tJa`;{�::�Cc�����~�{�����{K��;����/��=w�{��'	i����M}*O��?�� �Բ�)�U�rИ���"n.�D�fV��O�\����K�:q�d�������0h4�ӧϴ�}��Du����〇d��t���#�G�ُe�hy��t����9�@��j����I�"��Л�c��tmx�^ ���BePa9��JC|��s4�n��o���6��B������8��K�X�Z�b�������&���X�f�%&_�t||���v{Mn��ð�z�N�
S��b_'/�Xcf@���H�l�L>�sx�0��b\�>Dn�:Jq�)¦/�������I��]�G�q����fj�:)��&�nj00L�2�r��w��V�%U|��;;[���J�������U�dml�z���{K��mnn�qZ[[2��Ѩ��t^��u3�ԑXid����Z֙�T��I<���9¨f�T^�K�:�]1b	P���烵�ť�����w���[[;����p�q3�!���7 ��0f0 t���\�KI4�����l|��ZX�����^�W}���g��ݱ
}���	��Oָ;55!�5�X}�c���7�4� (vH���I��3	2��$gF���~����|T���i1��h#��l���8������R?fsX�����r���¤�:���q'�1�����f&
^� LH���t�QE���xI�ѽ�W��d�`Hש���H%>�g�J�G${�'?כaA:��w���I�{���GbS'��E�	1��Q����W�XR�b�_�v���z�b�p�(�S�s��:_��{]3�\�H�?�B���� =�Z�$ ��Ǔ�S¬�T�Ȁ�N���l��6փ��P�&̰�S������c�E�� HG�Q	1�)l=zí���d޼W=��4�����n�sy&����A�Ea,�l��Lz��|P�R��v�(JTH2�^h����b��%�0>��v�>NNNJ^H-ƥa�zk˨7�ͨ��������-8����5��sހM������k�40s�Z���O�<�������G�V��dЊ�ayQv�)�06:�J�9༖�u�fm^o*��3��ҩv��j��o����v�N�$��[@>�ŋ×_�]���{_!E���ӟ!S KK˙��1J39L(���M��%oJ�;!� �;wn�޽{���N�u����=��������t�lt2���m������&�9h���s�����Mf��z0
Rܙ���������w=���c�>zoei͚���[*N�\�Z:;�L'�N~y|Jh�)�+�y6�����}a��J�k���<3���G��$W@���f�����0�ӱ�\1�����2|5Dv�ϊ766�^�Qr�#-�*4�0�15c��b4o@��a��x����L���l��`�8s���i�v����#�{��%���>z�񥥻zihY�`�G5Z�=<d�b�y�{�b8u@�q��k��xm�w���O�گ�.ѩ�\-#����o\y�ը���ڝVk�4[A���.P13����a=&9�)�:����YBڗ�ٳ���>Z�sFl#���٪�j�������w��Ƿ6j3�JI�O`�b/��M��!���`� �6�!���=���k_��W�ţ�^|��iMmd�jmM���T�ި�c��0Rk��%O��2�:���<eJN�?��,���o`X�b�ߑ�a+����s��i�M���{�A���yX��<,�7���S��H�ǔ�KE4��Z]�����,��An��<{��$Z�y�x���y�&0,K�~I��v��!`��v�cĈmdg�P�I�����]D^��d��ޏ?�u 󞵟.���-�+����F��ɡ���#^g��M/ú^���`ny��a�<�S�.U�{�k�X� I���#�8��t4<
�>�7b
��F�$	2X���p��d�<W�������H�{8qG�zvb���^��K�r�5]lb_��an�s�߆�<&>�9�x:�;sG��v,�dwIQ>�r:�Ȯ�nt�6}���)`�}7Y~8�5q�S����wnr��I����	��A���ڪ�Ͻ�]C��n�K�.>���ȠL$C�;�A��0 ����m|-#�����Dv����㯼������u�܏���a�
_y���׮���)� �ǧI�ΡA}��E�ʐ��p���$�$ɒ���^�V�����?���g�z��x��g����Οۺ����z�8i{3������=:���1]�6�qƙN@Vc`�����z�Dt��)�T?�@2�<p�܊��[���XY�/����`�eJ�|�g؎v݃9�k�|7�������x���i��	�Ľ{+دgC����-^��;������<����6,v})��Ò'�����6i��I�۶ƹK��t{x��&&�byy)�z�b���*�T
��a�0�B���������iy< #��k�zawww�.)9�H��u�V�ڵOol�̀`aA_���2,�H��ӲM�jb���l�p4+Y]]�_~����ַ�~G�P��_�?���s����$=�tl]+�CRy$���c�;��\4y�])�H1;;+��@v�{�?����?�����sպ������]���{_�җ���?��g67�]��\��3 �y��mSL[0��Zy^35u�KPM�ﹹ��/|���<��3����zn߾NO_,��t:r� T6�bsy�$����l�<�օŠ:�*�)�l>� ��k�Q�0/��R���b_*b�κ����f��NR�}�3���Y�|�AX�� I�ޣ:�p�2�3 0��X�'���G�$n#�z�-�ZH�P��<�3d�o��QZ����kE��Xj߳�L�`�J%�x����4d#�R��a[��d�,�<�$��A��Þ�[fS��T�S,. �G�M�k�(���Vx���XG*ڄl&kss[����ɽc?F=L�&����f.���d�I
&~��
�Rq�6"�&�b���
n�]�0X;�Im?>��<er�'�#��y&�ar�����W�
��F��/�W��qWO���^�+.A�j5�ر�������=��i��ڰ]���+>�����|�u:=�&�X���H��O�w����\*M��vj�Օ����L$����(�����<��d�H�ӑ{��ML��V�:�y��sp܍P0/_����_����KW���y-i�G�^[���V���$���/hqf�Ș@�}$��}�}�����Օ����������qw�♻���nDw�.ە�T�Qux$��5ȋK��8-�)�x͐-�Ph�y��P��v�q��tEƻ~�����;,��̸�~�[.<z�G?z+���:R5H3Rn��mJ%���:���Q������ԟ���/�����#i�LOO�w�v7�s���OH�!5?I����>A���+���T�o�Y�)� �7B�Oڻ���C��	'� !-=J+1#��PD�^S��
�3�C�i�餧�1�R���[ٴ��	��-�ψ����tNH��)n:��G��������9P�4�� �󀕧3���dL1�?�PG^�o��8��3[�����	a`�ۡ����ݻ�4I�34��Eܽ��[�������w�ίO(v8!��[[���<`�Q�I��q}ˬ	p3_��/��*U�Z��$^�zv��t�����7���Ԕso�ve�̢�T�{n��.S)u��m&`�a�����Xϻ��k��QȢ�z��-�mZ)�ӳ ,ο~���3�=��c�=�����xw/���ܗ��|�v�O�._�Z͎���N/_g3�S:���<�bF�X�U?�\�OR�~��[�%}��r���fK�*��3O=����m��1qd@�B;��i��"q=b����BWZL�����z3vN��������k�^b�rj�^�c�s=O�|�6�
�vH�+�Z��-����z����Zr�89ǝl>F�$���%�e*�L��&o�%�Z4\��j�P}q��ǬH���2��I� ��y�q�8}O��"o�Q�C���B'�����+�qWԹ �ɺ,V�U(������d=���Y:3fI �$��l�������k��PqG#
H�8I���!����,��zo�ԁ��[��@q�k�pg]�b��$ȃ��D��2%����vF��r,G���~nA�S��<p֣nT�˓��3|���wvS���T/;��b�k�*�ϗ�� B���x��/}\��ml�L�����u@�yH��d�A
2�] ;!� ���Uy�\�^ej�|�%!�7�����6�5,Y�
|4J�\L��D��+���>K$��n���,W�0���J&c7U5�@[�Q�X��p�b��C�n�[��*��$!��lj1�^7����C1��s�5{��ً�۝ ��Ct�Ocj���ɜ́�'Aϰ��Y���Lu���B֗�r�GLdӈ�YH�t�zm�x4�ň�`(�ލ�W�x��+o��]<#��م�h��i J��miz�{X����K�%%^c��L��u�i�p}RO�E?�R���J�n�j���Uo�D�������f������D������.<�rz�����m��Ïɥ�N��� ��D7bY�KH��ax���̝^v�0�8��%|��ہ��!�T��T�6ӗO������Sb�3�ʥ9g�'�!���76&ӓ�}����/�eQ�
bm{W��QAH�Q�K�nf�< � kT��@�Ii�J�@���T@S F���N�5��T��w�9$�����v���&��S,���p{����f�M�Z�'s�	�D�8Ba/҈�&&E���])ѽ��9�8��n�,�T(.[�W�T ��e��)1�	AŶ��E��&bO˫woj�zy�ر��pN�o��JA�)�d��4 �-y������1�Gj��}K8�~� �q�wl��i���I�oW�x�)t}<�R��!!H�R�6+�#�Č��Q,ׯ]y(���`�XG,g�^�������������1���'��Q}!ak��
���$�ecz\��,�>���_�T��G�l�Pׯ_������/����'N��Sǉ��6k�4��`F΃g�b i��3��s�4� �ș�+�"T��0���RYj�:�m��9���aF�Ν�SO���2�������3���Ok�.z��w�SPEd)�J��!���\�c��e�\��@R�f[�\%tdɜ�@���J�����\m�����4��|���
E�i"`�,�)1�~�B}��	 _������?���/>v�'N�	�F�g?�ٰ^_mLLTw�?�=dK�m�&)d���҃��T	6��mm%�4��Q�f�P���fٕ^Wt�*A��%�bYL����A��+�Ixt�[�^暪ek��$����It؂ޕ�vW$����r�!t� �Lo����=����V�'���-2����	B��XQ��X�G�e0`�R�"V3����Mjp�D =�$��\*@wIO�s*���ltD�$k��jy?�1��2P����^�"?YN���L_�I���r�H��ɜ����h��C���,��[?L��$A�A]L�̊p�H�=D�n��e�&q�U���Vؓ *����	� J'�l�^�+��e�����@��Œ(TKҟ����J�*J�"�Q�&w��[�D�Uo�R���T@�����-��.΂���Pyd@3w���N��![�mwP��$
�jeB��u��bUZ����P#���V�M��U�̀��0�'e��ب�N�0��M\��[PYj#�%�D�,�K�@�
Q)W����\O4�Q�҄)��u�=Qo���
'�@>V��ͅ�b�&��\7�}�^J���dw�S�gٱ�RUc;aW8�X�|�ƈ( Yt V9{;4�6x\H�	M�45B��a�Qb���F[��z	ن��%�;*!�`��������D.8@�a�#	p�4Q��.������w�!�H��lm�M�솑Et�6h^��2t5[4kMi� �f���HD�^��Z�`�����30S�B )��@�'0�c��nؖ� f�#�� Q�Q)�yiv �
�Yr!"��C���O�t�.�]���F��tcb�8��fs6�'��(Dn�ْ^E�:��u�!�י �H=p��k�ds�o؍��&R�U��Va&P@Q"����9!�&�;5SbO9��b�~�Qip1!�E��2JKG�;C&LXhy�S�=��:@JU�D�M
#R�c ^�e����&�L�o(\*�mA��]�\�+��旄B�ÈX�=���}�]�q�ir�.� Ɋr&^Q����v���4 �a#�P"����߳�Np���5�֭���Ϗτ���b��?n������X��,
Df%�8���p��p���(,a��i��L�����[(�4�l� �C+@:F`�tO���(�J/�����dǸ �@w#l�+����KOt�OLb �L^I���.M^R�������Z��ɓ߻|��'�88}��n����������_+�;� q�L�����y�TIo�d���g���<N��"�'��B9�jt>��,j�r�IjC�0��M�#,��ZԊv�=M`L�(5��B6 M_bb"'ع03#��n���~�����U���Ϯ�[Xk�6Rh��]���|�ؼ��C�O�MN$�`��N�\:���h�Eʠ��B�W�J�
 &��@I�� 
��.�b,/�����8��`
 �I%��Ä 8�Q��@%jp�2Y��!=�\t�c���O>������+�F�(<p��Mϵ�������([��RC��!�sZr�&���qJE��1@��RXҒ�N$]��_�:�N:�0����˞ �T9DO��8i�t��%=/!��u�2��S��-y�M�mF�z��;�J�A����;��* J�s'��+M�+����0L�<V�8R�>
�sKŎC $��ɕ����`ҖZ<(X\�Ws\��Z�ءr$`�Q���jםN��:���h����)" R�S�\*hA��(� ���X^J��]Pb;� �K$,5p������^�cΕ[8:�~�hRn!ف\����MLT��풀� p��-W�WW�*_]��^{���÷���G��6	�X ���C���R	�cɭ.�$P�	�[Y.%���X�A>;�,%��D6�$M��(;Ib&��P+�N�h����qm	�V�K�M���jh6����=^y⹛c�����/ޚo6[�'OO�JƧεЋ�ő�n�{9�D�n�uÔ��r�����$� p�EK�cK/��NK��Ldi���}(�8�f�aSAX�'����k��b�9ލ�.\+���<s���~����^!����_�ӵ�P�
�٦�Y	M��IƖ� )�5	�M�:��Z��$�|L��^Rl�K�}�'�*$��P�X�I�y7��]����o|�k�痿��[��x#��n~J_V;����$��^&\RI�x:��_���%�Yl�5���L?�J�Ʉ�+���a���%M�mp��)l�m�������CBh�\��}��{�6z��Z�`caL-��/�pB����Q3������z$��{�x�%1�U<[�I�D�~����T�Y�B�đ���
��Z.1SK�r��җ���t�~���%��j�^ˁ���U�r2K�}�h}�cBՋS�$ͽ�!�*�J����¦Cʗ!+�ĝ�2���1��
��R�0��Q\���"�G/��C���x5���4�p����Bė\��Җ�?R+�W=�d�kkKx0�D)�"3��l�@��hB�?�\q�c� N�����h�m�Vj�`�+�]V-��h��Z}a{�x$a?��UV��9��	sC�=p����|Eg�jЃc�R��͘�?CZ)C�LT�]*�e�i`$�')�~{f�
:#���ݻ��G�0�8�B�ب�M
�e��cEE?�c߰L?\tG��;0�f��&�A!=��۽8SWn\�B�T�^����j�D0�WNw_��e0 Р'q�,m��=����|x%�I1M��?ϡ�(�UE���B�E*H/D���j<;;{���Z��p��7�������̜X��я}�cK7H4st����[F�
ց�KY���iڒ}�d�z �k���_����3��M׼n�{���|xu�z�嗽��~v�ʲ�2;t�g�u)����B�a
1��y*c 阢��c�Z�"�Բ������_���GydA�Й���'�x��v���K�reh 4fؽ^����rp���PD}W��Գ����.zcc\�����c�[)W��[�N��j�v:������D���&DQ6BW�lR�b�����e�XL�y�f"u����[�%x�U�W��=1��=Ǳ��rgzr�&�h��juf�<,%E<I&��@ژ���.�`3�&�j����AY��>��k� ZG�d�� e�c/-���C�ccG�����cT�^�XYYy�#xQЙ�E��d�U[3ԀY��σ�p3�Li냮�:!u#�ң���DV��*�A��V3&�y����M�?��#$	P?��ϼ������}�ϟ�?=D���������c�V�E7�m���}���T�$��셑�jYֵ�	���+ѵ��?�%�b�6���bw�����ƵO��W��Ul[y5�V0�hQ��r��kpX�������lK�^E҅����Tm�Wƶ�!̇˛��X�R���b!\��n����������Ϝ�m�P_��W�Vks�~���_z/mnlˁK>�/���������";h�j�����<��@���4��䔈�1�h@,H^��K��8}����}�̙�e=<�:;;�N��>�j�
�)h؎[�c��T���o��ٙ�
K1��x��DK���M���,dGL�x4�;�p$&i@��
�k4,�&{|Lz�t}�Qw�� h���	�0H]H�?V��:a5R:a��Ҁ�ey��K��H��+����U}��FQ��d��^L]��5g�&N�<�G��n��d�| �(��qm�=��� G�����&��G�
��MR�w0{:#f�N�(fU��L�+g@���67A�i�y=��7����<B��d�� �<�a��qɌx�Λ��䦓c	7]u��1��%�n���J?��m��	��n�P�ٷ���$o}�kR
%�]��w����S�0�b@��9����3��VT���Yڗ�Vv<�O���S�?
����[Q��m
~ĳ�o"ԱKw��>&����p�-���@�r�z�y��	U����>�	�����A���FY��*NQ�����%�כbr��Ǚ�Y*��F߷ǘ�$Ƣ�I̴�Z똄!����4��_dEzIRiP�-�_�j6��?��?闿�2���(:R��~6��2�2i2��Y�����<�}LJW�p]�Օi�Ӻ0N��=�������ݭ0I���e����v��ӛ���+?��O�s���RQ �lv3e6S\�c�X|=o��In��u7������ufr�
�*��WWV�-aVB�<�wy��/���B�����4o�X�=���R's!����ճ ��yM�U2��
�t�Ɠ��(�Z�Tz�O/���S�Tc{{��D>�h�Z�����ׁ�@�d:�M��tL�=r_����@Pl>�q0�{F�B��;Ns�? P�V}V1F�(7]/��c1��k2~]E�c�l����2�*`?1�'�m-�f�
������� 5��i�F�����d�ĝnKbB���P�@Z�=nI'KS�ߺ�ƿ�8*�>V[J�qHfIK���\|�8)�#���S�z�Ɠ����F
������?��^��D=����3�\!ݧeH�TuFku(�b�8t"����ڠ/�2��Vc��	"C��³SS�+�����v��^�ݷ�y�μI���Ν;8Η>�p���������g��7"Zw�/Y���(`y�τ妣��|������B1�v�� L�R;'X�	?v|���ֿ|�_�#1nfN���V�c��m��t�رc��i��N5����z�KQ"+��3r]ߒdLMT�(+M����[[[��(�m$�W�dv�e��+6�9�E�<:͵��JD~�����ޗw�N�y~u]������ʝ0��x���II���0md@��fw۽Iz���j5U�[RE>y��u�$8��*������L�M�Z$I�ib���y؝�uHl}���G�B�0��ѸYJ���nJ�37� ��6u�,��z�c�����	�<�q�5v6��G��g�,ͻi+�!?�$8������*�𣩹�q�$
ܨ��F��������S����u-u]~U#ـ])���?��z b�kY~�H|��� �����b�u��~W˒�	��7��HoL�rIS׻�0�o;�Q�;kis`�]I��Ť~�.��B{�E]
���!0
��Q�V� 9��=f�@�L�|Ӣ�LǠ��!� �l!2�v�w!�[��R�"���JVWt���ʤ4d>���^�A��zўg�@kÊ�C�`�����q��֖u��B���@ش}4�d���V�
�n��Q�W��^�^ߓ;:�5�ײ�k1�Κ<�+26��lkp�R	pX����p����ʅ��$���e���W,��n�3�������juZb��!ڤ�aP�u��ߧ_�_oӿc�cY"��rx]�%�!<��_���v������wŸ�bRܚ�O}���T���جV'�Y�O/g���t"��Ub�p����k$&i<y��
�O9.b9aY�>�НӧO�w/L�"�C�I������&���;h���T򎛀e�Ϳ�Hy��a��� S7r���G���Id�9��;���&�W���10.4�70���7���ғyG�6c��b�x}�T�,�Ն�U��ъ��tt�����nw�:�J����b�L���)}��T�Z޳���yӃ��	N� a�0����N������)Fh#�����;?{�%۵J�U������D�����/�1gT�g�$�������g�����y2�a^urB��j�Nm���{�p������xF�*��?�����w_@A�f�.c�ʕ��7{7��կc�t?�?J�C��	;���J�/�����$]*�ն��m�@�������o~�㏯����ns��L�֏�j��<3P�~��Ǐ��y������'��7���d��9 ��8�îK�A��Y3���|��y���د�gf���j�|
�ȁ���������(��&�e�٭�;kJ�< ���F�����b88 �3�EA�G�լ8LP��6� \ �8�=g`�N��!���_���Y5ga�񣈶s��Tl�=�q�o|��B˙��zGu2��~� f~��N|�)��^	1����V��xP;�+ز[�V�-�"0r}�H�Am��Ӽ�{V��� VjIԏ����|8�:����M�L"�=���|�F��L��K�r�0��8�HU��>#��m'��!b0BN��#����v�ym�"��vZ '[|��4��dj�x=�E�~p�A��Ȩ0s� �BK���T�Q��~}�j�f0j?���{?2͓��]�m\oB��㦜���|Z��x��(/�h�8���np��K^y�U���.�;�q��L��P� h��)�|.k��7&]^��ݭW��7����ݻw�}�̙���!�^��{���X�`��=���0��< �i����sk����4�ÿt�ұO��~������ų�ӋZ�Y�㒧�s��0og�uh�r>�}��|N�c�ȏ��������s��G6S�:rd�i �1�Qm��x�A�k�M��l�v'q,�4�U�|� ������rgg/��ydb��3����B�͐"nI����}1IK�0Ţ�O��[Y1����;~�]��>s�����x���e琈��igƃ��3�g����u�"_fc���{��L��u�Xղ̚H�BBJ����9��Yz�y���nr_}��G^��~��S�5@Q,b���Yw��B��:�t,ӱU��D��YI�D��FS�r�C�Kw���˯O���:y2F ف^�Q�t;�^���3�X��=غ|���Pc}o���כ�q����o]z�>�=�����x:@�ǫ����������x�e=<�JCH�Vr��g�y��Տ?���+Wd�����ă0�����<����{�=��k^T��#)�~��'��/>�C�Z궍�۽v+�Z�f(�q�����Z���a$�̃��<��sl��<k𼔌���JT����b��MZ�8v�bҵ��� �LP�n)>���w�{e��+O��'�O�V~~�:W���&''G��v�����y�}�PJ{���@�ߴ��u�)����	�*����F�����>s7h�{whfԁ�n��
����3Q�5S)�c���l�����}�<ԯ��4P�3.��^A������:2�A��ng�I4�ҷ����`�:�5��w��N:@tC���I��#�pj�-H'#�躮ϗ�G6_(�N��Q�`�U��G� i?џwL�n&`র�����|,�
kZB�v/�^B�h��EI�TiV��Z.w�S��v�)�=gπ��S�"S�0���و=�FF~�I�C�=)JĮc���0nu����jJ~In闝͑\�yL`�qݛiJP���e��Μ���`��Ǻs���C=t��}h�{tq����N��������Ͼ wV�dj�$3�� ��M���`��o�e��s��f�xi�$���7��o�������o���4�:t�E�����c�NH$����H6��I;n�+�^<�4�M��7>�}�5�m���R
t�1??$��Ђ��n�$I��b89�E�MSY4Ig��l��Ϗ�ɛıQ�`&�����Hv����R Ӎ��M�^:7G
�/��c浲(�P���g�g'����RU��1�'4�#'DPسG_���f��CY� �[�I\�Q'#U�|`��qM��;��<r�Y2���+�C�<:�w�� N:�^���@�&t��Q{=	9+c�yN&���:E���Cj䍍�u���KU۶�jh���~�c��k91Tb���)��sz]Ļ؅�%��*K6Ń4GvN�����TݥB�aQB��KKK;6s���Z�
$k������x�A���;�*���Y�����c�gb�lfi�Ѝ��:a:p��\֡,<����c%YzN��^�t��./�}faa��ٳF2FGT���p���3g�<.x凯���=�H��̓�m(��K�駟f�뻉m;�H��ʥ'�p�K��7V^����:u�{��^{��'���珡��X���LMMޱ�Z�݉�\JeB�|u@'�N1��Ů'l�}��=�u.��	�RD�y�'@��p�L?�ܫ�Q09Y�YX8�%Du������w>��Z�t�F��챯YUJ['�y}fY<�1�B�`��]�&����WJ�0fҔ�-)F
��i�
P��Y�� 4ҩ7w]�j;�51~�����e.[��T�yS�=�̳���%:���,Μ^��Tg���k��F�m�Qr1$`��|5�P��P%Sع�s�nGŞ�#�%
P��k�{��S]���x��x�J1��qP�ܲ* ����3g���6'd�c ֺ���Q����@�#�ƥL��<Hpw]��ݣq����A�7��¶�#��
��:�8�4�h�tj�fj0�s$�Q��l;N_�1�I�@�I?��-����T�n��c� a/��0�-�>��z4�Va�����j]��U
�Z���-O�����y+{���Z�\|Nb���#KGN
���vY1�1���E���Y\@��)$R%/i6[joZvq�,���^K�Y�J�oX����XR����{�7��q(��>�^¾���q���VYd������$�.
z��w'�L�r�#z��t��iD�BG�M��A�d�ߋ2��5P
��
j��֊���ё������x�'�-�]�|"]u�	����)�yהy��~d<
�E,���T�=ϛ�A%�Gݼ~���O=�t�����s��u7k�����O�n��>��EY���0�ُw��O3�{Oۻ�F/����C��v��.�q���ƯG�K�_��'O�ڽ~�:����":�� ��	2�Iz�l[v�>i�{I��8LS)ymρB��+B��%��鏺_BF�r�*+�v�0��oV
��q�5�ϻ�J�9��%+�f6W+���J与���rQ�v^���
��Eӓ��v�h�[$Q<�:M�FEk��b!J�4u�ʿ���k��@|��Me$D�S���ĠCH0W�ش/���++_;�4w®�vPz�2�N�� ���;;;{n���+3��"<�wS/���=��'�g�%?]*�Ma��md�a��(�#���w��M���G�X�Ѐf�I.�8�Q���Y+�ۻߺu�i��AE�G�'�|R�w��W^��~wii���̜'5s2�Q�_v�
g�H�
��B�D�����mGf���ڷ##��+��;������V&L,�X^�[۶�����W��׶�^���|��xw�ӑ�n4O�|����>��뻮�޴m|�Ća��=z3�V>z������(��גpY"-N�긣>2i����T�����b��*N���H���qzǏ/,=�����oݺ���S���SE%D{;+�xp�0_}�� 7��J,� VR3��,��S����~�J99�x����疗��\�x�j̨wэ7jԧ���f��nD�!̨)������MW-Ll�=m[K/)��OXS0��,2_�^v=KI٧���I�� |�C$�8P��\t~r�	���|�TZ�N½�ׂ+ V�U���ldľ�2{f] 1�JB�U����Q���V��-u-'K���������@��̱�s�����(����p}m�Hr�6sm���
��A��a��Wy2t�)/[��8�y{�ʸ/���M��;�h��~׶kK���RJ@�v�ў�E�ȍ��M�*�����z�i���y\z�c�X����+C�u����l��<ȮX�Jc�PLH2&�o��I�t�;w������/������RC*�2�p�jf�l�q��~y�헊�.J}K2٠�L-o{�����g�</Qv^j��8�v�kݼy���?;�{��r�ĉ�fҸx�b��ۛ޷���"����#��h���j�vhR:���k����j�ł/�v�A� GV��UmaY�0�%CF����	�A���Lv��㹝vϾ���3Ss_|�?u��5�/M�̶��B0֞��k��OJ���ĳ\�T�������'�a�a����:�
B,L��a}�L�nF"�J%��I&���OO�	�����'f���% ;D�4vk}]'�2H�n��ի\!��^��^�T�e	 ,.p9�4�K;�6N�B%�KE��'�����^'݊��x��8��x��#?%#|`�ȻC�:����߿w�M�巚m>)h���&{_�1J(�[��i���ͪB�E�S�t�ǁ��ky�;J���uX�����S�dss�So4�[��?��z҃������3b�_B�����M�N�#R�K=����N
��]��N��J��hؤ-�}�$r�� �pM�"ǂ�:^��u]�}�)ѡX��w&P����.��HaY�-5���Df��xxknv���<��Nݴ,�h�Љw~�Λw?]~d~~�4M��_t��;2�I�[vB��%�$ͦX*Z�v7�Vʽ��3[�f�&� �ְV�T�t�q7A��f���n}ww"��r��vw���-��-'!��-��"�j�z��H��cǽN�"L
|��|䑇�J�O���ϼ93��s����΋_~��Ǟ~��th��F����մ[-�y�L��t��6�Hќ�4�hrrRf��_��}	��X�ܰEV�Ϙ�K���8I�xg�1�Uo�T����?�vh@���~�ۯ 5b��Fl��An��ȧ�    IEND�B`�PK   %�X5�3$ �$ /   images/8251b1b7-c97c-4929-9682-a545aa133660.png<�cp%\�5|b۶&vrbL�dbs��mcb۶m�Ěض�=�~u�]]�?��w�սzG()H"���  $i)q  l�?ゅ�/���#�?g/��  ���%�#  ����"j�Y�҉6:��MO�ݑOGݩ�*Zf�pf��pb�Q/BH�Q��Ef�8�q��8�9:�̶9�����Gk;�^f*�Wx����y�=Ow'��W�������\N��������/�������rb,P}�_�O8�B�wG�#�6�����e8K�Ż2)4������] ���( S� �\�ޯ�s������?�����o*w]�z����s�Mv:񛮼�B�Xn�Fe_����B[�	f�W����f�I�����Z��2w�is���9��F;��Z>!��xS\ْ�s�ݏ�M����3����7)�U'O4˽Ħ>�Ka1��ҕ�G�"����P����QK��?_g��n5_�x���I{ڡ�﷣G=g��?)�]Kۑ��� P�����E#����f( �r{�j֯e�wjY�QȘ�:���`�]��RFԊ��&&�y�M�8��<��s�z�9R��[O�ȡ���*�	^OP�oR7�H~�Zo�ڌ�.�L��1���&c�2�4�C�8�����[9iӔ��rܝ3'
G:��~����|~�Ef�H� x����F�gs?&����Y�yhK?��Y�x����s�v�m]ߕz�Y�>i$��oX�:k���^���\__������}B�����'��_��T<�ɽ���`�u�J,���֪�Q9;�W���Pp?�v&#���t�b��)����=�����y��p�v��BSȵ���Y��|�V8'����UE�����U!�%/�X�#��*?�6X�\ͶnԴ�G"s�����Z�Oj2����g�j��Ƈ%�vmk�犹av��0'� 䘙V�
�s�|�=:�gK6�rB!�z���{�#eؘ�z��#�ǐ?"�uJA�(#�t��+���!�]��7\�W��g���_Ћ��)1�V��ʭ{����@��H���S�����Ͽ%�ǰtP�����1��w��c�w�X��i�B gvy�e���e�u?؞�宪P(�i�.wK1rK�՗G)��3�	J�	%S*3��th��C�5\��or�L:G_@��/m+�Mh�Ry[V�0|��������|<�4�ZZ�q�`��!8s��H����W"��m�Z�SD���4�Q�/?�a����t�OiVS��[� �_�걝-�� ������`<�[#���������Fe��F��6���Q��6uc��ޒc��L���ς��& ����_J��;5��8����^��5~�7�\U���+>5��O"B�k͔���[I�������q~�Q��s�����=/{��(��3���rfT�@A�W�%�Va��N�v�h�_<54l w�����kQ��.Z�h5U/5iB|�jV���b��'���y�*B$��dGf���us�R�HE��2����B*��,�����O���X��Y%�!.����b��S�kw=H�O�n��-�h�Vw�8�����_	�t��Xm`�]�!\��R�q,1���^�h���<6 s�o�E;��7�`�ٲ����0���W�ݚ����=�p7�m�CZ���BNk��~+ܢ1��TY�쀦�[u|4�W�76Ma��إ�i���Ke�bԝn��MH��	��֨���:��'��Y�о\��X]�L^�#s=���v���>�U� "�����&�K�@����G��i��C�j[[�V����}�U.M]BN+�b=�޿C ��g�t���`�y�^U�+�jG����X�e��j�2�f9�%���XJ˛��v�~����l�`*2K��t�S�]��L~-^;%����7�����v����%��}���.�U��5���ԣ�y�n\���z�=�?�ǡ��W�$����O�9���a8�^Y:ð:T�2��n�?o>���@�����v�=fϦ�'LF\|,(������G��S�}�-0�Vytk6v���W$�O��r44�|���1;����L�����j`j��_|�G�<kN9��{�{�` ȓ�����0����ua�/"�aە1Q"��U���ld�dI�Z���q�&�Ja�:�$y'l�N�DݿS��QF�XGڧF�o�si�H=�D�d��$��!��{|f���7�knWK5��%��(Z�?w��b�mq��$��t{��&9�m9f�;�]��%�BbF��V��m�6�=-t\�dk�������(�[���o�=L��h��-sb7hg�~e?�W>�h��g�_6�`U(�_�~l��(,�fo$�6юv��j��\�X���r\$����$��\U�:N����P��$��Pڕ��'f�T�dN�希;��fb������mj��4��KI�?��W�K��WB��e�(�OA��O٣��ϫ��:�p�^�՞�]�>���`���	E�&bpeb�x�1&���&aA�}�mX�E!=�J^B���?�׬��ݣ�\0/J*�c�q�?^%��{B����J�x�
�ď6+��U)���I���П�5jO��PҊY]С:���%,�ϣ���?�����V^{�GY#۷^z^>o;�P�vbw������#ο���0�`B�tFT�R�+�p�93�8�K%G��B�x�}k��Usp�l�C�\�o1�o�˃t�z0�!��H�jf�];�2�Q����B�<w���X� �
%��MI=���CAo&��PRg���*{Oҧh�	����� �ϗ:�J�ϝ5������rDE�<UT�%<f7��� )N�s���&k��s���H!���-����S��n�C*�Հk�{�8��\���:7���_S%�5z��C�D��1l:磹��KKM�w�~����tI���c�n�Ol�f���`�e�
���=?��9�+6U��Mj�z������q����xY���<� :�0$>M�i�����MO*z3{�e�W������_ϝ�]:��i'DxX�PW�%V�"}�C�^b�3\�ۗ����߶���uoWU��~[ز#H��/�ϲ�D͌�+�ëhC9($U�A�o$Q���"�ʻrr�+O#�ҩ� V����֤A]�@D쉥�9��]NN}
�~��Ax���@q�@�!Q�kc�csÀ������P���tQ��)d2_�di��mZ���cr	ljlC7�4�t�p�Ѥ��^7�����9��H�Dds��ƱC�	Q:ǿ�AS��1����Q$n�����y�|�X
��LK��w�!Q�hbmhY8��*f��H�D�d��2���I��s:z؟Y<"�y����~ͷ�Q��K`��@����_��x�S�7>N��Q��UG�ֹ_je��y'�F��l� �0X�L�p��sv�9�?�r;�ED��#�!?��E2�Ne�~������J}G�}�2�N|�;	�c������ϙjaι�[��>�X"����.89�m�z/��9}G���3�ْsf���$�@%��2]�'SZ��
D=ݨ�~NZO�2��~� �3���.�ٗ.�o\��w�=������W}l�Һt�ڜF�����U�m���0@F��	ߝ���d%k�P};�J�<-A���
�x_Mn��j�d*V�Gd�Mr���[��+�_-�/z�^�A{̔7K����fR5�UX�J�H�W�%Ջ���R��h�F�b`?�����(�8��z��J���e�'޹��;;"
8��ቢs����=7����;r-c�OЃE	�����iA.������x4 \�:����p��v]�~�I���]=������b̭>H�T^��x|�`=�1�#{m�ód�+X�	CO{�eE���
�dgR�'{!�+���!r�'<�����l ��HJ�p���6�X´z�t�!V�CD�������� ��hm��햑-�:�=�U�0Y|�t���I4�v�v���;!��+}&7�ݖ��^�.��Oc�3 �uĻ�r)���]1�,0p��I�P[`e����G���bU�/����|`w'ڳr�8�-k��5Dihe0^����9��V;Y6�����p����]�+LX��E�:�ܞ��U*�;��֘Y&��±�!=����.F�w�T�Lcc1����>�����,�[��y��(n�R�^��M�������k�UG|k�)�s��}�����C�ag���|�j���4��ۨ�ѿݭ͊�<
ѹ-g����'v��v�.�r���|9Eގ�a�����iW�7��Y\���㛞�L�_�?��$�t�mҴ��!U��P� @����Y�����o[�DO8Ԝ}����*�|�U�:r���G� Y��>E�*�&�4lxլh�_�wy�I�se��['n���Jw�:W�ޥ1-9����Ks��X8`�D=dܑ�ڋ�b�U\����9�POʍؓ�d\,��o�ʦ춸`M�7��ۉ�֟�Ce���ry��V�x��X��-�aa/� 4 0?I� ,��R�k�6��?�q�?q.���]%8e]��@�@���O��c����֝�tBjT���,�_��IN,�� >  w�ÂY�qb��=r�j_�^�vn9��:{+*�`y��=�вgc��7��@@�`���ᄘ�c��
�ƌ\t��v<�k2y����hpd�ѫ�l|�|]�M7Q@��\R�u�1;
��K��YW������;&e����֦6Z�����`N�r&�Ŭ�ǭ�|��Z�<F�ʣzV +�ܰ�D��[~��y�ə��ũ�J��׻~�M�*hnc���8�ARN����L)�~�h����һ�sD��^?c6�������8��z�Գ!E*���gv}�z��A+��D��G-��ϣR	z=:w��|q�h��ú0P<�͇-����?쓁2j(�� (��	%O�7���tX�r,V5�,��߾)����:
nU��R:�r���͍�p[T��kE5�}��'�� ��z V�A���#YJPB�Ya���n�ow��!RS�T0a�������q���?���3�b��M��b�><=w�a9;P��O�Ff�0��l�.���4+w���h�39#紶Pg�cSB��Q��я����a�v�Gܹ�g�u�]�� 2Z�/j鳓��"ݐQ.&����*?+������A���-vf�[ߞ\$��Yr�GGe"Tio�6�E�3�x�J������{�܉@j2��cj
�3�{��lu��VlіT�F��{�L�,��Y��]6�q3���Ύe�'��櫑�%�UFa��q���[�B���x���6�g�b8ϕ�y��"� �i�EJ�s�˷���q��F��q{���B�
(�;#���$���p�I��'\��W֑B4�^rV�=���+��U���tn,G9 <�TT�o�D� =JB��3v���(��������$$��B�!��\��2܌l��)`���`k&�j��H�X�Y��z4Og݁\iDe�#�d�^m�0f�PNn�!�^���[�l0���Ć��h��nFٶ������1�D��2��G*��/�e6(4�"�����?f�]�K=��=��=�� �<+�(`��Tg��B:~Oڇ��?˧�M!�e��e�۫]�_怋�ԡ�g��Zk�+�8�4�'T��8�������}}LG����U�R�/�)X%`z S?̓��$��J�v.�Z�{.����� ��j�M{��g4"��y��l_j��������"�>�v�@�������7���[]ί�Y�vT�zo09�9P��^1+�[Qf���?��+�7��|�y�o}�������>�2B,Mw�-���Ay͏n�=U��^B��wo�(_�7�� o��+!n^������'�%����#����q��*�K؁�>����k.a�1L���O��~.��F ƞ\?v�ÔF.5buí?!AN�^� n�����F�j��y��ʾ�Ͽ���=�sjT0����<Q����B��_kW��'n�o�D�8{c�b�p&��\��d9�&���pǾ��ظ6���;����9�]�ӫ�4�,����ԑ�f�p�)���(�D���-WD�եD�C];���ܵp�s�s93�-ˤ]�2�ii&��,O�����r���c�GU2���ՅD:���e�r��P@�Q����<���՛tm�� L~�@3\MU��������eW���6_.3�  
�B0Ze�ʙ�튝��о<"^F7ٱW��V���%�V��m�,����׾��=%bA���f�֪�幔��74ha_�̰�&H ���vEb��ս����chjV��z�xp�Y�w%B�ޱsuO�E��<��}����[���X(u}�����`",���Z�J��Cs��qR���q`Lt��ؚH�������+���~�B`��3f��?֎�m��x:K�_��z}K��!�����T>Wnx[q�nݩD����g<���h�j"�c��i/��h~ �8*$�Ku�b;���x���	��X-�k��g��"P���ɕFrϹ�u/L#Upn�q:���M����F1�C?�wZ�!Q�(^�g/��K �M�8

qb�.�{�5� {C��e��f���̈́M�2��zp�o�Q+�Y�5 ����<�a�P��7 W[���A���0�jn�YJl6�bԃv��4*%e8cVGVg���4�OO͎�a��*7o�	m/�}[���B53�b6p�L��\�@؈[�n�O#Zd��C�;��0J�o�����!�T�П��W�}Іuh-�,ďۋu" {���P��='f$<��}c��a�9��߉��Ym���2ϒ���ɨ�~�>wcX�/��W!v�]m�]�E)|��}N��n_�(o����2_.�	��t���5�KkO�|6�˰\~.�ǻ�/^2K�7��_�31r}�Ю�ړL,n���jhA�}���C�럟��<&�x�ŷ�2$�Adⱐ6��U(sR�<��|"�~ަ�݉
��������'(�`�*<�D����n{T��D��8u���v,6l(.lY��Q.R�xs�-�~w~���=��ǡ=���1'2�\Ҁ���]�ts�+$��T*� ���=v���Ddܽ�g/M�\Lb�Uŷ������JB&�nvIi�`�}�2�yr�/�Դq%6��%��q�v�>^r��ڹ�/fy�{R����O�Od�.�˗�+���zWbz�h�8֞�{3=��'�v�yh�|^��[�G��-�.!,4/Q���/V��ٵP�]��\��_Hܽ�P��?S���>���>��ri?���#k�N��J�j3]�t���^:�~� 4���ٶ��9�U�Bĺ���y,9�D����,��N�i�0(K�>8�"
��\�Wg\L�H�F��MD�[LK~7�%�o��3�� I���Y�r�z,f��?ڰ�/ϿQ���A��@k:�&�:�D_v����?�3��Tc�t�@��g5��62�������#�ĩBXIפF���K@4����3"�D�pg�a��P�H���<�Pd d���ª�Kf;c��P8�օ����]I&r-�e�ů�7�Q/�Ԑq�2�t��Xl'N�]� ��G�/�9�kN�����S��H|�:�/ܣ�^�����Dg���_�Y��N\cD�D����NJ�)z�|�a���d�Z��X��'0��Z��NoZ�@"έu�k�F͉�Cc���I�I��_�>$:a��mtWA`X�kވ����ʘ�L�S�f�D�=���N�"*�P
a�vt&��(HR�|���+����o��M�4m��-���m���N�r!�$`��$�t�I��-2[�{9�����S�A_�v��̠�~��1��(4G�S�v�k��t��+�fN���gObK%7'���X�{h9L�&����c@`.�T�6Y-�zP���g��r�'_%���y�c2��k�v�ҵ3
P]('���Z,͹����4��lQ���uľ���C�٬z?�Z�AM2s�1I�����dQ_��Q��(>�*f��C�J�:�$�\��JP��<���J)k�y���H���1*dE�:����,�sDmGW5b�����)��'�r��,m��&�vM���moy�%�VeI9I����$���X䤣�&����Zgm���k�������@Rw�Z'g0�R����� ���Cz�#%�*��ÿ�|�5%cl��	<n��=׷�"/���ߧ�&���$�~VB[Ew����&�u��B��k��G�Q������*;z@��.+
��A~��	����(���2P���6 ���9Y������Y�?O���9ߞ��6�X��z.�D���T�k��t �x �Is���2tf�R�Uf�wâ,$��!^�7��js��s�\j�	'S7$�n�Hj
m��Ϥ���a�H�d���n�)g�X��]���S��Bʜ�q�
Ѹ'Gq?�f+��Ʃ	f#ax6vbS?���*Z��Fm���w�xVhO����7�8v���l�E6�Pg�w���-���h+�����!73/5:�0D+�m�5��s�k#�֟��4Ģ�#eR
7�II���~�-�]�(bNffg�������!$��,�R�0�a�%�R���À��g	Hyf�,��� _|��\�!������-F�݁�@���c�-$M2��M�۹I�M����gn��f�x*��!�v��&,&0-l)ѻ�sҠ�o̊L�zL���I^|��Rv�6fҍ/Α=v+�j�	�]A���{��?Q��C��]�俴`�|p�y��7�0 !ΩYڨ6�m�f�� Å)%�s���U�"�W/�O*����LU
��{N^H���ϼ�C��L���Hx쩈@��4P�v�g�1�3!��J\όut󒅁o�����v�}&�w\�\�7<�RcʑN7�V��z����!��y�w��� M�%��5Å�Z�E q��Ἒ�rd���0;�O{ _�̙X�+<�h�N+W���)��4]�e��_��gz`�(h��6[V�Q;�/�g�+wroo�#�Z4�ύ�媺-`�a�����F�K͚Z��+��ңvl���4���: 5�A*?��x
� y�#qTN�'�����p#���k"{@��F�Lꔑ��+��ϙr`�����dϔG��zd������B7�J���,�7)r���Fl�f��^�sC\~6�h:�K��߶w�t���E���m�Ϥr�r�g�I�l1_kH�1;y&��zZ�ë�����޲˽�'����Y�������{��,���.��7�޺F2�<�7����qǧ�F�dɁ�k���1�ą�%ޒT<�M@�ҋd%�p����5�O����Oo�����w����F�JQ�=�JH?dK#�������lY�� ����Qu�"k�Fi���>P/x�l�h�1�;LG7�������Ҩ�8q��@��dU?�� >�	<���P5��1bh�5�N;Y��=���ԣ��t���`v�������4��% ��x�5n�x;���B2lٴ�x, ��z"պ�Zi=D�E����D�{�ʡ�<�a ��:�[!��Fp��	�aX.�:�|1��NB�U�,�K�)=c��Y�4�	�]�,��ß�S�L~�����t�P��z��ϻA[�GbćfO�l��2�D�(�ׇGG\���d���kv1�}^��NĦ���7��Ƌ�+�OѦ�U����7.?���!�]�]����Nn�W#Gچg�5z�7�>O:��r�$�硼����i��&��R�D6������1U�K-�N@Ln�{�6p/B�*m9!9�>ìx9
���c�� :A��C�k�08x=�r�=�����kS��>P���^A��>��B�k���޴�N�T,iP���8�ә3��8+lK�rه�,���㮨�������QA�ZO�k���dt�^r��:�}�h*b�����]��j�f�\)>D<t|�E(�z��k��80�gS]s�
��J�.�FD�&����1p�����j�v5�)������f�g%P�:@b�I����|��Ղ,��z�,%>�\1�H���NvV���iz
���A�iс�� �@�d����EF����13vE������圇=��A� �}q��B��_�����Z�m�p.�v�JS��a�Nc�\_P���E��Y�iz�	�!�\V�"�9+�~��Թ�Y���*������?p���@
Q�0�LB(]�+s�1���1��%G���Ȅ�R�(ui�X��G>��/��'�*��S
J��f"Y�P�b��O�p�x�Rjo�1���%�t-+{��8��T%�0s�I[��Ǜ�3&�ǩ~�˨��Y��>��a�7�|��q̅i]����Ғ���@�y���W��3<{[><����79��]��+zdSPp�MG֖`fl@#���-�ْ5%���I]�X'��u1"���W=f�VٜQ�k���GØi�����솶��,�cQ	aᳱ��}aBdщ����Q�����9.d~|5�p#]�����¸�%�=�}DY�:&�.�Hn��6���&�@l����x����Ǡt��c����6������0<�A��r����������B+�!	����U�o	1�oPҗ��߻/[�U�-����)�_^�8?3]���W�R�c�m��iqƓ�(KŻ�q��#Q�-�!h�f�#
���L���ʆ��գ������@��ŃnhW�܉���2�Uy�G�W[�,m��K��Ir,�8fJA�@N�ӽ`����ɤH��g�C,��X:�&P�v�<Q�=��� =B�JH���1��&��N\��'\Ҭ�5ȳ
�ñԊ����쉗7�Yix��	]�M���XC�f+D
�Q�6���	�d�r)
D��F1�޻�I{�d6�q�!���_��G���N{��l��nY8F����&��'��B�-�jxv�� ��ص�t3�`�2*���B�x���9F�߫�V>3����),z,�y�P�i�����Iq�7�5O���Ÿ��d����s�iR·��J���귪��ү�&�@h*���qa��.�c�� ���ݷ�u�5�A�	�!!����d��\�|�Ecx�W+��Ӯ�1Q��Z?���+L��i�����.J����c���G�6-�`sj2��7c�4�ʒc-V8�x>C}�pN�ߠ|�[��-֞8C-���M�e͍�c�"9��V��}t��U|�?i;H���V[ѫtu��U��]�cծ�侻i�WA�9��J���I~�3"��צ:&_r��	,jr6�)�:�(��m��� G�}�%l����0Е�nb��y݊^��5w�ڻ%	�$��DW��Oœ/��L�U�k�O;�T�s#�qZ�G���\e���*��*��A"eE�-h*#��ⴰF�e���}w��bA�h�Je���F��"v;�/<r�r1�!<������I��S��y�B��6�t�cĵ1��z�yQ��0�Ay��	V��v����n�8���?X�ʮe:[�����E�ɮ����d$ھ�Di���������[$������!n�~*�@���ˬi�n���h&�]b[cI�� �^0��hץo���T#7����ovN����k0��y�ݟ��bL�!Gx v��������7�-����1%�R�c��?6@ \����k��e�u4�wC��A`/q׉�S��dȈ�URѵ��"�A��y�ّ��ߤj�5��Yb	T^\�!KXׯ�X|RF4�9��n�{�Ɓ�V�ʁ�(W<���[/��:
�++�x��x�0oB��t\�(212�����X�_&��ղ@*�Yټ*)����^��sJ�m9�
��v��G��N���aC:آLMBY��Y j6O|�-tke����(y��60�����r����Y~saRX�׋�!�h�j���y�Z�<��lQ��.�
0�s�է���6
]Z4Edu6�MzsZ����☪H��d��7� �m������k�Pg����.�I�@Íez-a���e�h�9���k�����&���O��uz��Yt����'�@���\��u�H�r��P9Ù���=ƮҪ:��"}!�4�!�Ta�(�������1��P_�>�ˊ����h��9b�����>�WR�2!�M!��ϔd7BaőV�/���7q3�mc�L��I����)F	!p�%��s�KBx'��d�iv0>�s�"���������f��_N�A���e=�����蝬ӷ,.�?�\�h\�t
Cw ��q�hj�&|�놪׷���S����[�����_C�i���i�r�[#���"TȋR������T�Q3H����P�!V��u3H6���cD0�SBa��Cp��n�:N�2�7]W��z���R�pA���c�����\��r���x�G�Ʞ��nI>L4u�YY���ތyd����0r�x�0�R�a���S%�Na)̒W���7ȝu���+㉁7(܈z-��W�_��"���E��U��ZE���ú�mLp��j���츍Ȱ�3k:/�$2%Ư��0k� _����D����!��s`�#G2k[cl^��V�g�Gύ 8�F$�8��l���a%Y0I�4Ȱ!��!�I��nJ'�&���ķ �5=��y��x��Ӆ4#��L�<kK��9m�rީ�uK�ҮŔϣ�Ӭ�B�����-[`l�-����q\�h��`"�6�1	�Z���E]�DŎ<-�����W}ܜ�Y�[�z�4���E��5�Ph�� ��_��^YD�g ���8���y��~��n �$f���R6��UֹV���y��:t,��!{M�`>��\q��q�6�:��z���ڲӭ��s�;X.���%j�:�&�0�����BC��� 97#�.��r��0�E�cN�\~��{��	�&#G�� b�z�%�Lb�ے�v6,z�^BQ)f��HN27��H.1N:
-~l���mu��+Y��|'�/:\'"������&��V����WƸ��`)b���H��]�3���D�Ǎ�6ч�F\����˹�<�2NrVT	iB���8.�$Ƚ��nKa[�'���b�!�W<�r������hr����~��$
7�Wmi����W1vn�a]&6��3����H�d,V2k�^���&7�X������XzG/._C`V,wm-�;��i�F`�`�PEo]V�!fB�'��Y��߼	x���n
���@�h��X�Q����r~�m*�����&tr�a��)!�/j�9YTR(��(� Ơ�FEw��LK��*���֯邨�S�"cC���β&�>�U�
��MԒ�C���.d�R�٢�&���c+gc,$�g;�����H]�.�Vt-:��*V�XczFǆ�̽ʸ��]���0�&d8���֧��`(<M+�6�yx���HnH8��������R䩐��H�,%eM!�����k+����B��ޫz���;V��6��5�C��l�$��PM�gB�����'�w5<.u2��%��5������	�M�	��`Jҫ����`����j ��;fȢ0�:Nry3����)� �EȨ^�Dn&�sV�h�#�3���`�E���W$�] ��,���`XiRl��Q����s���p?}<!�)*�����}�3�G�%H�D��[�0q�?@�.��Z�Ktڜ&5D��6f�='O#4pβ��Jf����z�IKF���u 9�=��Iv+H�D'Z};�4��;�%�bL1퐷�b�,枹�M��|�9��2���Uգ��W�'�Q�%������/��0j�^k�9����?+���:��b$�\�^�썶!$/��s�_�ޯ�4�J@R��������k%��2�����RP�>VCi#+s�5UU���A���y�Eü�٨x~���t���N[�hT����_�}x:~HD_�E�᮫G Be"�� ̇�GϝNOx*����-�5`���QY��?!�歐8C��K�%����<K���I��tg�CkQU�wI���o���('����#��|@��[��qu�|U�����r�XFgS�MO��3D���JS��v7@?rؑQ}�Rz[��yY{>?��f곀��՛e`!���h�D4m��Γ?�~ы�����~��@1�{�0�r��X�_w����B���!�$�o�k��m+�Ǯ"W@�!��KU�#t��0�2,m�e�nRZN���>,�Lo�D���C>9Zv1�=0֣Izj��k$V ����S�ԃʢ�.����tX����`�i�����^�RZ=bMbD�$�L��W�7v��b�</�7W�0�kp�HDќ%m�]��e;:Y��e����uM�����v���u�U�}��k���wDH���~;�I=���WլKcEm<�s�*���P�S��hԃx��?�懋�D��5 �C�Tmc�kI���1A	4��]����^,;oު)&)�H����T�u���G�m���AEs��nd�M������-�����ɧM��e'�^���.��"7���؋,�߁9ٳtA�p�mY�[�;_�(��p��%Rb�)'�7�GF�������DĮH��κuOF2P0< �$��͠iZ�K�P��lG^�z�m�ռU<B�R.rW�����VOC����v��bI5�iW;0�p���G6fs��t�]s�$5�/�[8�h�v�!N�4���&Qh$�(�����`с�8�%=�b�!����!�ʬ��pa(��i�?<Dc�3Ex��O�M��'�ɍi�ӱt���|D��E�p�=�֠{��b��ܓ��ll7�g��ʕ$B�r5����0�M��©ߞ�Z�Υ���ΐ��MZŸ�/")ȧ��F�j�ֆ�t�\W�	����~r
��ڑ+{lx<Jh7��y�;0@S��Cc�6Lx2��@�7{5�J1���:��ݓ�ն��W>@����G|�W�d�;�{�	��	�M R���k�8����c��-~�qG�=%?�\���[J��{�Q�y踲X�G[i|����r/U��z�U~��ލ��}��@�Eg�GRĘ@G�5��ɕ�"���]���[���^�KF>�e%+�䣰��"�q�p`���9�R��ʟ�'}��`�`�G*�3�|U�;�\�P<o�$z@"x�5ͱ�|���X��z���;�Xދ7��nw�eʫ�m}���^�~����UD`S�{��Sz�E�[�.ß�%r�p:�A=�F
bp�v�+@Mj�E�F��X6�����ZTO�k	;����y5�$�h�A5`�s7j��%��]����3�}���ȡ+#�nƤ6�_t?�Ё��W�_�H:�AjaU�z}���Ϥ})�!)��C2�?b���^N��bƑ�h�c�L�����n���+���I����J̸Z�}Xx��Rݘ���OL���2Vb	�Ui��)�c�V�&��*;���΁ư/JD�e�W�?�6P�v�O2R��(��G:�z�h�7�{g�,�O������G��~Y世ʒ��a�>�;0-<��k�'��m�] �T�>�U�Ёs�w�Kd��e���-oG�E_�3�ȫ?�OCͥ�����v�(��NG}�������!��y��ٵ���X�G�:.����u=��HK�����1Kޔ�s���Tk��姁�}_�{"�Cq�@
�E
�`��'�#�&1J�����n{�n�L		�c#nYn�V��cﹱ��4����:����<p!A!(Y�O�j���L)h�nAK_H����4��r�f&�Yg�B��£xI��N%fu�k`�'��i(��V0él�V��>JL3 h�����D�U89%��T���U�a�|F�򅯲˙��1t�ƺ���$�Ά�|$��g�ܭ'�Ǽ��lo&���/�!@th�盙�a���A�s��W�d���^{pu��Yb����l�5�^
ŀ
X���~W�%�����1-�U��O$3��� �I|ozjVHBO��Y��"�0<E�g��46�	����uV��}l�+�j�cOp�һ6{ݚ�7�{z��~D�:�.2�����K��yq�@vV����p�k���@�@��taLm>u4r��xSvj�=cAbqA��P���W'cc[Uȧ�AZ(H��~n6-�(�yS3(�ձD��X��H���D"����#
����L�]��n��H趞������n>J��������4��n�Q�;�va�Ka�D`� L|�n���b!O�hdd�5������J,J�����A混�^�P��"-ʌ@��G�G"-���v��Ʋ,�u^_���_��E��@F�	��� p;U����J.�����t��������A����G�i�9�hɈ{T�6�)B���T^_��WW�4ܸ�`RY �>4�p=0�_}�<:�W�[��l0/��+�cܶ+�I���-�;��۶�`�I%6�@�/�/�\�pgUD�pÙ�9��joOSNӲ�a8���y�U�R�]8�(��>mEV�˧5��[ ��� ���:抝��OG;#j��@�@�p���:�\�A��Z�~��j@���{]ОO�5Wj3'Xg���������@�1�Pv�B��µ��i�e�:��5���$����v��>�7�����P-~`aX���;��@�:��q�a?yS�ȉ2ۓٙzϕ�r��tƨ�u���[�r�F�+e��N�Є��WЛUkF�A�5�wȉ�WֱY0���cTU�|5��U����3�\3Z�1V6����^JV����<�ab=D\L�������,�gc8)�L�s���{�j��w�˗_�Z���� �jX���M����syyq"g�؜�1� �瀒�F����� A�n[�%�g���R��,f�,g��8l���f	C�����!9P+O�{�kg�Őo|��f,�YW����>ԛ�
j3)Ǐ�0������u�4rw{#��/�\���e���p��y��c��y9;?a�!Y�2h�s̦�{�׾}�V�zۗ/�b��'�gs���A�1w�q?ڄl�-1wM��8^�����# ��w��#��g_��,kC�h���>z�u+��K��>�󾾸T�l��;gB�����!8��,�oC�ʊa��(���0'� q�BՂ���6\�"�`�ZJ���vw���b:�S�� �R�h����ŵ\_��]��9�w��ӹ���Gk+���x!?��Od�v��G�³�
�
^��rŭ���7���c��$v��iF
eS纆>{�R~���x�	���|9Pkր{�Pۅ�G�}��Ƒ��
,��X��l�PF�(���(s�>	l�Y$�MKR�R��n��g�E@�Emc���&�2(Xj;�Z�������w��֤��X-"���w���9r���j���8.y���O���G�	m�|�!b��B�]��Lc���A����tg���#Y#����hZ��K5���v��5dJ�ܺ���M/.���;2��8��<2��@�����s}��.n����D��7��g�}��)C��C)�2��u�5 T�}3u�tani���ۡ[�zK&�dz�V
�
����@p��EΪ޴w�_���[=���$0�>��£V�3X5dg��}^"2<���Cޏ=K+e>
�\���&Nu!��߯^��@~����b��/����%�u
����|؎��uD��7���n%��G�AeI�$����ޮf���7�˟�\A�b�K3L8->[�{�0���؎8�aS� ơV��E�0<y�P���Z���0T53�$�ٲT��C��0t�${!�����+z��i��!�dSJ
��c��^�m�V�C�V�lfrhA�\.���F�LJ���̬����A�0�&T�%(+�Ѕ���q:���r5ГQ)�'����zs9�,׋>��>����K�p�f��Yx�m];��a�B�&�[l�����V��:�u�l�c�����.S9���	����Y��Grrz"ejM�c�p�RrGfvD1qo(#�C�����Pk��*S<`0��S2}~�-�^k����;J#�=X���+����� |���H����b�_���m}c�Xat̐:��4���@��iԈf��\&�)#Poաe	R����ghB��Td�'�<֟sn�"�=e�9���x-�f��,�
�-�zEq[��
*�Q��z��=��40z�N�3��FJ,C���P��p?�#�{7���;u�d��9Z]����.��.x�b-p�%�M�OK��ɧ�>$��9�"S>C"ւ�����!�E����ñ��x��^��~-痧trp��d��vA����c���[*��������z��ѧd��@Gq!t��Et�*��Aj�A 0zy����E�����γ=C���L)i�'�u���r���P���X���Bk1�D�,W;٬?r�(����9��Ȅw
�s��Qf4�Q�D:�
tB�2��D��#H(e�X��v[�a�:<�M`�J>>=��~.ˇ��kn7{x��$�A��1�g����F����&̠�X��M��{�J�Ņ��IJ����-�+���,��:��f���J^( _�\ȏ��^��(�AM	4���5���cNF��ݦfȿs�H�qؗ%�ZS�u:�żv����}hb�"������&/�
A�
�J�-��Z���Ҍ0�;��5��S2eJ�]y��z&�;X  �������)�M���K��l�y�B~�/�\_�P*�S�L�跺жd1Xlӑ-�qn�E����Y�5ƣ)���b%�w�:�7tP���gz:����p`?(����=k� B�A�b���K�0���5�������#̖�5C� 52�����W�����KS����_���5�p��Q.F����s��md��NY�
n�=h0�ʀ��F#�T��p_>�+��S��L�L=��21��7��ulw�+��-��J���@�!���[��X�^�˺ޱ�ߜ!�,���:յs��� ׯ^�� 8l6�DUHG�-��2�[��BDӞWo�`c��A��0��l����Ϩ���͋�@�=hk�ґc��ةDX4	��
y�� �CGB�r���Ш�!�V�~�������g���IH�Bҁ����ղۿ���q�S���?4L:f�" ��j:��u bi(D8{SkYK]�����ěp:���/�Ky��;��Ws:ܸ������C��c�{,l�49�q=��d�,�[H(��B�֩$ϙm^b�y/u�1'Ԇ�]V"?���L�*�Vt0�n)M�����p����u�l�X'I9!�d8Ԯ�@�z�޾�(��'Y?����)|����Cn��<���p��9�4tX2�%�Vm��栤��u<W쀄��6� /��N2_�~����Jp]�5*?~�9+���!*��Ll�iq�:����P�Nf(��Dd쐕��ˊ�,$����Pg��?�����?�3�:*��e�,��̉[�56X`^%t�)ʰM"r)ȵ����i�?_�3����^W�K��� �Hj9.����zܐ���v/iC����gS�DIy`G�vI�Zq6u��,���J]g�3�W'
�������ׯ�͛W� ʁ���|�L�Q#��/_�O�5`" rp:5ȩ��;� <�}��&��@�����V��[ș���YfWr�)C���
�9Ǵ���~P@}R�s+�e D�Uj��!���`�^�:լ�Np�-��GP��9mu������G���  h]!�^7X�":��zo3������K��
!�[�H�
���L�!΄C�%>D��&{cƘ?<](���x7�Tכ}Dɓ�����:�*�M��.n��x/�����K��qM�� �X6���{KpE�![Ȑ�������LǬ�0N�v��#���F�!��T{Կ`� ��>�E����uM�������Z�@�������F��S����ø'H-���ي׹ �6)@t@�M: 0B#WV��M�^5j_|�#qo~B��_��_�J	�m��Oe�cB�����8ο&I�	�����㽅�$�f���M����F��=�xE"��F��[W�o�́mEt��Z�˿��/��/^��}��W`T� *�:pc��2{����%+V�K��޿c�sߥMP�[�ǣ�X�b�:�c�c\��]�@�+?���u��GF;�c� y��y���4:�F�z��n�"��8���>����!>�s�H�Ij���X�e��gS�v�>(����6<`�Ibpj>�I`Z�O��4�hϒJfj���B�*�AI/J��Js4�ʫןq������7�N�ʓ5��T��P��ȅ�����r�(xSc[8�o�=Y�!O��F&��m�:�%M��^�1?��}�}��E��b�Õ:��0�a(
�'�m�:�ء�6�p���$�X�*���ϡ�#� 5�%�5�uWB*7[�}ǲ��8_$D�����"�[���oC	G`�u�J�����X� Ǚ�%�f�s.���齝�seR��"5É��!
j0ȑ���?Q�$�̆N���lt��m{��F]%a����5���}n6=��L�~E�N�7?��,u0��@�:?A��!Z*����{���>����4kۺ�i���
1��ķ"-���>��T�`�gj�`����M:�<���\{밻��i�\x/c�n���ӑb?a��ͮU�K�0�.�r��3��O�탽Ŧ&�����Eqj_n���5%�0�N`=�`Ajl���[��|ʶ�'�l��:T��1V<����%��W��D�6r���� (t�vv�V,K!$�\>Do�h�:�g�
�:Ok�u���w�N��v�������ڙÉ���&�a��̕��k6 ��{kF�0�32�F�c���_����������ޟ7m �_���+�|
6���#�F�_��Sd�a����G��w^񳏙u�덟��=��yІf��?jH|��
s
���Ib�8FP��D��`}���:b�
������ l|T����/e��H'�7��3~J�!�=�f-I�|����0��ݷ�5�ɚ��L��+}�N��/)k�1������V&�5lwKy��r�����H~r�O��ҷ4j���Z���z04tz���P���\A���M���������t�C5I�h�Y��	IBR�3�zst�Ø@��il���t�.h����eO;�	C�R ���ۏ�R�7��;s�+T��e~{����D��PY�A�YZ� �%�Sc����!���g�Z�z�1�&0���K�SC����پ���?>Ƚ^��C)|����D�~w,��l�-�� �Y�0UEP�(eڱm^b�����[�n56�zɼ�X�W���6�:^�mބ�X��CKϞ�-q����;)�����<�-�X��e�[��[�:j��w�����`�7��.��B=D��F�O[���B�leZ�^��s�ٶh��?(K4ʜ��B*WQ�0���dzv)Y9����|x� WWjfgJ�mW�]�N��I^�w�A��݋���%)E���|��8U���0$�*����D��_^�ۛ��_�U��c���o����	�)��iݱc�6��Kq���s��/��8�1E�eヘ�"#��|:�Ym1v�2�齮�wO�$���T�^���I���y2Q6�5f��w��F�a�!sk�b������m�����7�H�@��_��D�B��lu�>�#�� ��ܺ���Wz�P��9DW,SbG��B(�m^�w,�v����}�qΟ]������z͊
�*��ȶ������k�m`����������������6,�ĺ�|@9!�T�����\ǆը�:ĦK�!"'Q�������j �m=�����q���P�x\��cp=�S��@�-#w�ׁ�l0��db�G�&%	�T��}!��1����V�vB6[����S���d�?����X?�#w�V�~����7߾��x��P\(��k3Y�k�+��c�~_��:�Y6lG�������C�<�����A�O���0W�3�p���(�7oe��e�&l�v<+��}-�e-�>��˫+���`w��ţz%j4�������ԡ'��EM�J���j@0�I���3�d�>��T�;���/h@�`���Ã��[q%kX����X�v�{�'/&(�����@���1|ۆ:h��Z����c�{%�&ƀ�SA�MFF''l��;�/�B��1E�0�6"�AmC?l��֥)a.9	N]��%4�Ol����6�G9��cr7����`?��
�������/T�!SdZlc�$�������S�~��ދ5q�5�7(l�j�X���
���C����{K�A���iDv(g��;�
������t<GaЙa7���&,·��\8_9(��ЇeGp�Ɉ��N��[]�\ț7o��յ,�-Î�OM��� {,�����5�en�0�P 7/�J8���c��߼�����^�Z(�v6w��L�;@!��t<G���9��611Kl�	��^Z����+3U-�jXl�Z*��s�[��F�:��T�*s{�z���`/�hT����R qG�F��Qf!b�;���b�t�w�r�`m3}�s�i�	Zd�DN�	8'κT�z#ద;da
(h��iBG�����D�w9�%W#���~��v�T���ק&|��w����?<�V�p���q@�%�韞�������ku�f��&t&p��q�e��~bTV������g��齚LӰa��+�)pJ,R��oǹ۸n�z��v�����1�m��������c�G���Ci�
��ވJ��)�\]�����;�w�&�+�٢�7�)�u�������쪸j
`�� ���s�����NN�c\���d*#�78�DyN�3J�w_�t~�y�cr��� �zS��*��oe��7 ����-�Xw�p.Z᥶~�(]�q����E��yb@t��7h`�ۭe=)�{�� �*a� \2����B���~���Y���w\8X0�d��P%�:
����'t��Vz�.��7/�SN�>�z��S��.g�RP���~���X�F�^lr��Ęx�P޼Etm:n��zGg��b��'��, 
0?���\l�^��8�ӱ�}��ono����6���
��Pl�t���e@�!'Ǟ�YP�b�����a&&�kp���i0:2���J�4�n���/��a8�-�߷��&�r�mgM٭�ZLBۆj���`��D�!�N��<bg�|eq�X$�j����1�w�[Rh�H� ��)��(���.<Y٭P����W�z�=�s����O��g>�W~��׬7������ٿ+��S#�����z�l���% 4At �i8P��:w!�C���ým����
�6�5�����ؼ"��tSSK�aE.��؃2��1�N3��l0�6r�XCȧa�ݰ-�5p4a!C���$�M(j�z>O+��QO�p~g�`�<��ש:��&��E&��:su�D���o���r�(�Co�f�3�.&�,B��6�v�����Ou(0\�H��#�~&�}14�B��a����z"��l,\�Vm���YA���_q����O���}��'��|�ϗ�p�$��L6��n��h[��R�%�~�߸��-KmͶ!�L�M�=�M�OEW>�5�|�͡s���{�6���>~fz�ݱ��uM����wAc���Hk~�y>>3G���ɔyv����d�����,Wҿ�F����/t��B?ь��$�U;	!%��F���/���BN..��ťEu��g'����9�>��L��Ax�\9e9){sK��̴VC�R�pq�Z&I���Qf
z_��3�ԉ͜M�Cc���Xą�\nh�N����I������m+w�(�f�K�5@*K����9�<[o�Q�'(Sf{�
J��H���%<U�ZV߾�T�*���vz!Ԝ���d-6����k�;��]!j0�F� �b3:g�T�2c�}�X�wQ��J������}~���|�d�������� �]��6%��x{��F��Z�#3p�r8SU�Rս}�z���/ү���?�ͤn��ΐ#��I�CD���v�Yj3�2���<$<����Z�F��f�������{˾���9| ����f���r3S�כ�����?ې�k,��NB��� �u�`��[�&	��{�=k{���@I:��{$\zSɍ8�8�j_"wM���S�aD�~٢;=!(����1^�wRyM`��Ӌ*�{�Z��10�F�)�Twx��g���J#K�F�O�TI��g�������R�e���1@S�zg!���u��9��Y��n-� o3�1-�M��ݛaO
�O8�{ws+$U# H�Iz��Q�h-� �{�����>�
N?Ju:������B��ܞ���u�z��*ߙ tUV4�Fm��?� \x3�M��i����>'�n��L#%��r�瑐A�3�$�f���	ƨ�#�U#���T(���{����P�|��u�P	�B���	��pѠ����*���mO���A�����cX�kj<{���R�OP�zF�<n�gh*�v�>��y˯�tg����v�ono��ew��.+�lW6h��$�UQ�f�`(��F� �������lV�Z��[j�N����Ktt�ٗ=�����<���Z�X�N#t��D��M;/-���?�[x��g���T�h��>ƅM$ SE��q���S���}X�||�`� �}���>�9��]��٢�W%A���ڽ���U?<��O�:��o�}�b�����X�����>�T����� EIR5��]or7\�c]%�8�z>Z�h�dzo���c*K�A
�L��$��W��w�,5�5Z���e;��R���96s:Lʉ G'�� �0��;�=�m���/l#/](ڲ墳_U����K@�h�8�sT!A�}�Dc�*T����Psb�I�XQ)*�dRв����:���xSi����J�4y�~
�|7vЯ��C	Č@r{�g�"a��>qB�E��٥S�I2�0eQ�DҔ��N��(��ë�~ @q������� ����JNb�?�y���B@0F9X�TrD���e�v���3z�<0J|&�=׈���4��~����T_>����|��ѤU�i��d+T5��J�q�QHdA|���m=��P���9��'�A:���	j��
В�i�3g��ə�:����c3P0�-]&T��"�=�I	�D���dͩ|N�+�;�;�r�dʦ;��2>M,��;�}t=\G��^��lG�44;�����\\�m�h�fj�����[�SӲ��d�cɞ� )�	�s$��[�3����$�K��;�nhjK� ��W�R�:U��(	#�{U���9W����"8)H�t�"T/���D�41�)�X1�02�ݞ�h��
����u&������{
�3#f2�P�2�b��®��������X8���Gsʣ03ak0@�
U�u-6/��ݣe QV���A�f�=p�pqo�<��U^�����۠*w���S~�N����K2�����������p���⩢X@�������/j�|"�,���u��>���\ڮ������L؄�W��^�c�m�2ݎ������5�����AB�z:fci����鮇�9�/;�掆vW�cf��Z��
�=P���!|���p�����6����	�ꉣ��S��f��<؇$2���~%�^�)���d <���,� �a�V���X��R^;���\3�z�jn��(
�V�r4����O-��~�PYc��'"�R��Γ��GRwQ�K�خD"1�=]�����o�žb-#_���,���  �h$⨐9�Y�<��0�|xt;��/,Ki;_�ЮՋ"�t�1χѧ�ѝ�
@���� �dv��M�P�58�,3�5��Z���y��@��F$���ݣę, I���I�!��E:���+8�����Xe���e8��A>8I@o2Ɩ#�AB��A8yy���N�(������~0�Ms^��V�W��\�a��̳���d�j�1��o�����T�d%���{��Ə����t$Os9�>fD���'�,5�Wqaey�q��ӣ0/��"��}��x��i�0�A��	p�BqKj��x�w��ï��>����"m"��_L���d֔~d�3��5�jY@c�7��=���$��*Vx�k���������9�ޮ�,��Y�x�}Q}�%�$��PP�`�?ص=N"4�x쎪�#OA)��R��7����^'dA��gHt�E��Ŷ�=<dX�Ah��g��[�������� ��_�. L�
�!����^�z�vŏL e�i/h�!\�߇��G{�;�AM�q7�tb:���h�v��}��{�j΂k�ظ��Ƭ�e�kmیV8�����Xʄ��'Sf�%g�v��]�~�C��Ke��H�X���~�4h�q�����	I�	�����p��M�;S]�9>���lcܧo��h��������f��)���k	�>m�}*X�
U�h��(�[��w»��u+/�e=��#�z���S����"Lw����}m�Ug%�(�8�U�p(g88F̡�+�`)�eљ�9zq�$�+�0�^���7��.	�κ�����vA���	*Ȧ��);TM _�ٙ��"����Ύ,���tS�p�����l������{���m�ٌ��W��á���Z��9�UR��J��|�FhX��AKE��x�����_}�m��=����=�fj�'m�:e'��'��4��XQ��������2�f�u��H�Ԯ�!�X�m�6kN�C�R=�x�xQ�����s��q:����'Zz�J݃�9s=���+J��ζ%k{�u�,���A�n�X=�w7�ֲ���[�w��/��"�V���>��q6 �[�*��+�G
��Հ*�e&��� �Eל�J��|mYv5���H�^�և2w��W��uZ&��KA'jID��ؓ��t�K�.	�� �!�/�!�ȅ�],������o�������GH�(�5��,�h�����Z+���Xr����\���uP������2:s���Z�7��-%�q�ӵz	��F3 �L��t���텽ݣ����2�=�|�'���Q��e�2`C��XT�҂��`G��*Z2��I�4�^d����f�?P@#]���LSr<��R�0��8aJ�cF��A0N�*7YvR_�з�{���G���ʲVJ�RV[�d���9�������peA����-�y��TN��q���z�sU6�Ւ� ��@��+�)b>��4b�G"�y��������~��};�V�s�9M=l�(��|���G�Nt��F��vBc'�j�Oo�(6iL�)Di�����5uqm�SCX�,�1+�Y�Em
�7�VCx��˥+mUT~��څm�9P��^�T�D秬꿃�u��<�&�$������l2�������o�03C��p}x^�2/�A�TC9GG�>�� �0'�g{�e!# �bib���ޓ���b���f��;XZ�׻�£�<��
5��E�͝q��^�Mxt4�P�A$/�_���S� ���K�N$CTy=�QE�@yZ$�G	��b�)���eh��D��~����� y���0����cs�{B�Hٴ�P�|s�04��Zx���76 7@l�N���ZI.t̀[���Vd�G��?��n�o��Vs���e�yܦ:��,��gI��vD�f�kEݕ�X2_E�9C�Z�V>�ۙ���{� {Q����\�����<�̱Y�a{n`�W���(��+�F�ío�- k*�ڽo��g�ܢ]^SABQ��J��J��.�eSFqa�&�e�r��Hvx!�(@�[��{vvN�4����nB�}��ޅ�Ҳ�L>CM�'��0mu�sQ�t��'ar��hiF9)@w�h�9�ؾ�}�������Č�BU��������`�;D ���(�����ɞ�Q�|����DԖu�U ��`��,�ݨ�vs���)ޗ:ɑ���X����IX���6�~T�	���pg�2ɵ�A�G��k��k���u�Q���s�.�
g[��@0��{��ٿe�c��0�I�|�3��`-H[*]KB�p�d͍A!���6{��޽�2U���qE4�pG������>����ewbp�~vaj{�ͩ>��@�rgӊ�+�6C)Q%�j3NԌ��^!�6�g���B��o;�/��I_�����_:�m��I<���	�V�8��,��ڙ6��|�GI0*Q	�����b�Ι �W&B�D�HN�
k����R V�X�o�Q�"��D[���V��>��N��������9iŚ~I#qZօÉL���-%�cƣm%=��Mv`wzmV���O�J�/���pR	���%�t�Q�Hʟ{o�B���7��e6�)�Ǌ�����[�fhj�������٫�9W�c���ڮ-�̝�dv�C�;f9�^S�����L"v3�U��@���]vaj�����T�L�Μs^e���Q���l��*J��g �j�����*Ef� f"�g�����q۱�ke�����
�P�l'9bJ���E|4G�
Nͧ������� ���@��@7V�N�H{i�Ɓ`CS^":�\ѐԫx(��#��	g-�Z��A��:��j�o+�A�"�4	��Xٸe�׌�������lF�<�,t��C��0ǘ�k3^����D8��"��u!0��=�L��&z����TaT�ʪg0孬���	Mŋz�2���R�	%��h�_�����A�>��]�!�� hn�*��q͛�e왱�`�-�[6��T�,{���W���E�m!֓i���H��Y��U`�߷��Iۡ��?�Q����U����~3������`k�5E���-'�OT������!+g�y�)�8E؀0��;;=8s��,h��}\[�����,�{C��3�E�fE)A����qo޾G{�a�3�;;a���'�&;'�Z��!^g����V��|VeöO���}���zaA/�Q�O�>�gx���/U]��u?��=�X�7���vMd[T!Ԯ�HU��l��}.�y���Ѝ�J�IMil��ɇ�vSh���a,h͖�<'2��� 
��2��9�L>1����m#M&����2��DI�F�ܰ��1�U���8(�m�c��\�N�ї���6�%4���z^������١o��U������n@�*~����	�	(�آ���A:��.b8"�o�G^��������݁|C���R���L8�BYt��=�������e������,����W��9\b�	�P�ǈ�	��>�仯�SI�r3��˪��/V,��W�ی�t:���x�M��*�$}�G �68�w�g$��1�ą���3��x�����#̓�7��_P���_��ӓ�]]���@C��Ő"�ilY�(T�)�bdCIo��������~�駰��#��	-[9A�h3WJ�PE�:#����=I��c����w�i��YɄ톢���T��d�C��ss@�rPEX�0��2C�k��Dq�0����f���f�1�:4�gj�
N۞�>.ë�_`��{��������<���]�^�ZЌ!�����bD�(��A��C�rvS�s�@��vm�������[f4��KG��F㐙C�!���d"�Z�D���XG#��t
�0�]7Ų6�.D A	�n��R�K˘f8��l�u�%����vw�����ك8�K�Oߩ�bc�xJɎY�8��mա����˰��G��.ȸFc1U&���p�ƾ�� �]/���C)�/�=������ؕ9�c�=%	�F2�%�0��!=OHl�P8K�Ϭ.�<ٙ�����|vo���ݍ�D{ʪk�������dg2�^�/O_�- 	.
���������ugd��3j�#�}���W�#�߿W�Ү��_���/¾}ֵ(	����æ�Y��n.���%#|�Hf��Q��φ1*w^u�N{gӫǦ��q�tU���L|�#�	!�$�'�]F|�x�	�vjo-�ߺ��.��oKv�Y.}�S��������A�2U/S?;F}����ʄ7Է��f�C��5�Y��ؒ���	f�(��F]k��gQծp<K#�{k�H��a�U��&դ��{����ᖲ3,I�针U�W���d��C"e׻n�_4����yXv2�8��0u�z5hִPfG������>��ڽ�������P��ե9���A��*j����5�`4�P���^9�nfH�d���e�"F[8a}_JF|�m�qb<uY9�YK�NK�@�G�LpAײ��9:4U,�X����m��Y����^��W��pa7�,s��8BGY���ʲq�UD�
Ӝ��oxe�eY��EX�܆�FG,2�ol�f�K�d@EO��.�|\��o���!I���2���g�.o�G;�fNGz-���yJ���7����|7��!�̰؃�V���=�Ge��*�g���5��uP#��f�#�ej��Z�u{B��(I3o;��z��裙s�0�� 	�8<�A���-��C˼>bh�E�\p��Eaf�����#ڳv�&��D���Է\Ę3�!�.��N3�7Ͼ�e�r�:�^Vt��.�9�4wlǾaD�Svcz�\��*3�Yp[��P���#�`��0������2P�����QԻ��͸���c�K�������j:���|�k`T� ���>��j~߲J�:�)'O9dj�Nd�c;�Sw>~�D�89x�BP;�Ӗ4hU��8�-����*x��}��	����'��{{���똙�pB��[;.�L�L�*�������Y�֮g�]a|i����A�4{���l���w�D9KB��+������)�ڱ_&r�h��U�9 ��q��|���џ�1Fq��shK�� h��.PjJ�Z��"�[��2:g�h^~�m~��Ϝ�v���i�,[�rfX6}�9�g3�_:�d��!{֚Gށu$W���x��OVh<M��g�Y�κ'1Ӧ�q-�_gA$�cP�
���ch�ۢ���k��
'T�YU��/G��yfIG��<B�b*O|#B�%� �_(��2��m.�S�&�=g/�UU�ޏ�(���Ko�c�;g�������3�y.5>S��������~{t���b�ΰ=e5И�2>B�W����؎<���um5F�Ъ"�pg�X�����:������ݻ7af��]CRvv���e1�0�8-nv10��46�	�G�lx`�3D2�Q�8Bt֎%�¥���G�R �QE F:(�qfI6��K�cFqjH�C<O�#���7jG-/�kjـ}�N��@	���Ht��8������̛T&�͐o�������T�[:;Z:�i[�9�DT=�+4��0_t�lf�ԛ������24�k�q�-� q7� �Yx��Isx�:�2�jy,�=o�҅l��Z(���9�����5^/#������Q	!�-��Ubt�
�;v i���C~u��o��R�3SX��&QQ��p���f,�һF�-	����&!���0�<��#`�K~�q������ٵFӰ�§�H���=<��E�ĐQ��=�s������z�S��po?�-hI�EB��p_V��q�݅9�Oח������w��f���Rk�,(SS+΢�s 
g�DA+����֫%���^�
���&�f��W�fR�"��a���#��ڳ&)^�Jt�ij`�oԵ(w*��0[]T�O�")�P�r��<~�y��K٪�NE��U��;];��{{[�2:���I/r��Ά�~��e�[��%F�Ϝ붓��#O�eC����~_>��%���icW���pf+��ת������%a���-�s U�@�B
�Q3���&Z��*~$m��x�R��Z�d���%�m�G������Q��>N8����b�tQ�!�<!���
`���B]z��v)}�](�Ț*�fu�P�ax��2�԰�1XO��n �B��%&�\V1j�n^싨��YTi	����u��� @�� >�_B0y�%�&n+EF/1��'9J����I�ֵÌT"%,�2 �{��e�w��J��sQ�S1� �=���s�6��$z�Ͱ��6���g*�8W�?���1׋qiwʍ@?#��k9���u0ՌMgC�����(/¿�1gm���9N�/ކi�*%2: sSy*D>�h����N�?�#�kQ���k�eN���PH��\�uR�NՏL�;i�`�-�!0�sx���8J�)[Ks5���5
p�l���^Y��j�Y��p ]<�I0�LE�Ӎ�E�+�+0z;��e�tw ����Q�پv �f�A����c��8d���M��,�-���o���Ψ��./8�U�`�N�O��;�]9�YIYӂ�o�Y\��A�ZW�Y���g������y8>��9��QF�o��3��r~�9�)�T,�v ]`���I?=���װsK�xV�(�[/#N�%x6hp�����T�F�o��4-�3d�I���]�+=qMY�y�رτ�`S)i�Q#�v��y�����A�Ƕ�{�3��<cj %�jF����}��y����M=���H�J���h��:b{�5�|��I����5�3\ǲ7�άAB]z ��h@G���y� �7E�R�V�x���7�ή��y6��=��PcUMt�1�L�+�"J��8��;QH]?WlՊ��h¦��&B�Q�(�q]��� �[N�	�̒��;�2��A�E3��<{�`?�O��T��7�3����ރ �v�~������,�����}ݽr��u�9��/|�"'\���j�g�(Z���h�X$�g&=�t3|3���Jo�)���V-��Y�@f��� �_{?$�j2��fi��e�4���8�v�_����=҆֯R/�^��E B�N��!�;}JҖ��{��A�����cv�!��O[:X��=�4�YD(۷k���`��*�PR��Y_!�BjQ?�l���cw����k~�6i��AE�Qd�%�*���9��s��W:1��ǜ �A�����J�d��A{�,'�UZG�ʼ���zD��b3����K��s�"�h 7� 8�Z |Ԉ�Q�U��:�ّ�e��r�v���N��	���,��,�wo��Օ��P>ho_�֭��4��Gfp���`��}�ғG�d�r$�;:9�G�B�Bw�gQ4R��Ž���]!��'���e����\�^�ǖ��L���z��]��-��no����F�iw?tv��	u���iq��=cg~]E��"���%�vtpN��.
�j����`�^��g3&K�՗�̹�l_�m����?��}nz���|�z�G�0����n�A]��k ��N0�5��<G�Si0W����U�6�E2����[R�����ꨣַ}n@g��[@fs����jG�b0�S����	��$���}F@�'L�ǿV�؉:�򹢳��ׄ3���I�YԻ�к�:��w"�����2�lVE2�����]F�]F~�:|�p��lSV��-�ѕ���nn��SF���&'��~[�a��#��}9S����>�J�� ��e�5�}�i4K�:�̞��w����ԊT�O`�BD/�T��b�;O�	�`:Z�}� w�f8/�dZ��T�-W�Z�h�ש����2�(m!+π�ﰮ}��Ч��>���X��T��s��P�����К(�r�WA���/͊1~�� ��y,C+M4�I���y�[�#Q�nu7�z)��>�
��E���#�A�j�n�hRsʉ��^Rό�=ϲ�tvv��O��\˞�	�/އ����oB��)���~o��YIn*%8a��4�g��$��T" ��ȑ`$�Æ$��	#B�+@�ܐSG?��z����xnx2O7���f|(�u4��P���y�?�/^)+:3%�>sR����0���HS� L���0�׊�a��밙�X�w���@�5�|#��!HQrxV��S^W�<��(1w�,���eص�udAV�E��̣x�1�����!<~��!�@��G\����kehdnD�
*�k�\��U��NSH������a8{���ʮ@d���v� �Qҳp���!���!$��Ss��l'�%��J�Q��v��r��p�o�U?֞b�5hRa9�����Y8xq��V�[ ��d�,Cl(�r#D��ϙ����������V��J��'rΡ�%3����ZE���W��l'�o V�~�~|�N篿R  ��1��g�����yؿ��`�k���7߄����C�����pfg��=v��O?� ��>*�l���B�Y���D7�>"H�x�&^��չ���;ـ6����=���������6����Q֨@��ډ9�O�(	���
�d�|�ϳT�A�v$�'xtN�Q����}�L>�(-���	�t��Me��b'��#����������6e������ʖZm�<��3�Cq�G�������u�۽���Y��45�0{�il��z�G�^G�ù*v��Q�8�{�x�PLs�k�ԭZ$1��CQ��so�dè*��۰OÚ9m�9*v������������''�vڣb�^[�2�+�T�l��^�!�'�G�1g2s*�3�wu%�J���r����E"nF�Xl�g.Q��,n���8P���(�H�1E��4���γs���Kg�0��Nx�a�9�*4,���{��W�e6�.l�d<�QZ�>�7��#�g�*1fyU����:��#q&x�J���TŲ���k�{r�(�g �N"�﫼(������)=��'���d2�r�̈����zz1'l�Lh5�F�@�R��]>@�*�?@$�>���q8D�Mx�#1F���[�v��52�"٧2L|��'+����ұ������b�g.F"J|koFK� ��i�)<�A�-�==��w8pI=h	��d�.�'�tw��_hi��Ã�p0ܕA��Md�r��<����(\3�h,K���g�k��	��R�K!����@ڧ�{� 2흝�m ��f0��'B������e�Ex�ؐ�d�3��J��l�ý&[�w��/[]�d���C��	'��8pJ ���^���8�>>�}rz"���Թ��`�'�VQ���H�&�kWt�ʮ1�h$���o�Kx�fl����+`�OBd�K2�4B��D\���"�x�Z��v���<��bVF�  �Ү�������U^���`x@��9�o�IJg"��|�,����N�0�;�<��%��	>7�������k^�Sv�`k�1ld��`^��F�Ҁ�˃���6+}��1{f+�с��zUB/���5��S�#�]Y�F�J�&a��~s���S�������� C����(<��R8�f����V�����ml8JT��m�8�a9� ���O�Q��5vڋi��q�e�IO��ES1�M6\��jC�Mq��a�Q��
?_�߄��Q��;L1*i��#���YXH�X��E ����U�Ā��H�)I�L
CO0�o�K�����XT3���6���e�u!�n�B�2Ľ\�TB��_~�_���w���C��J�4��P9��|���)#2y+a�*�p*�㨋��uT�Q�P�Po���hƍ��w�w�Zr��AK�$�8F����wO�\i�H��"FO��҅'r�e�����y�i��Z\\]jV� FT��'�]�̵y��P�B��&/�<���3ͳ�Z@�0SfK�(*�5e�rg�P)/�|@�Ӱ��[���*����FtZN;`;�P��96����Y�z�X)[���s$f�׶����B�v���J���@(gu(b�*D�SG��14�'! W�AOӭ���?q�y�T�/k�"(��+X��B(��98����99p�a�+*@��+��|!ǀ��cCL����e�)1�¾�5�� �lJ�]<�$�=���I� ���S���̿~�]����ێ����cx{�>��s�WfЖ���p�0<yT@z��ܮ������g��������ʾ��>1�S-sr��Q���	��0htÕe�3{���~߂%�뛷?�D��9n1v�e+#iG�7e�%����)d�L�&���>���1y�
`3�Zz{��mfm��0��/��b6�
F%�j�~����~��Φ�[�@���G��Z��]�Rf��猯��v�=9h����@�rh� #�$!E����P��i |e�؋��Q>b��pg�����H�+[ѡn�<��ڮ�y�<9ֈ��������@�QTU���?Dv��۶�������fo�Uu�/�q��eEu�H����#�	��o��y�U#P��N�l�$�cK�3�oA6�q�����E4��["	��١E�h������EN�i�:pG��gm٦���x&\I4���6�۟�~~�s.+�΃� �N�rL�Qd8>&���xQ�M�D&Ls��ߘ/]�9N�q��p���iwv����o^�C3��?��ǁ��y�se�V��Z� ,ﯮ�[�4�,Rz�6��=܉���������T�֫�R����K����T�&��Ne���Ml�p:�dp�g�d\�?���P٘��G���2�����:gjRVI8A�U�'0�p��N�+�c�uh1q�V�eZ{Z"������ ��/�ۑ��g��^w>�|f�C�t�����Tk9r�0W=5׊�k����Ux����� a�������Fdh
۾�ۤ:s��,}NY���ف�dl���j-cH���j�?P�� YD��m h'�G�G�ҲE�C'��,bo�Q�9E�Ct�����ks ��a�Z2���>\�*�#����վa����u[XVԨ<��$����ah�kU���zk�����!�;�?^������G��gZC��c�Tdw�d�w��!�/3g*�|sw����v��Ë��4�Էk��t��2�A/�-� Cм�}I����T����V�3����D��49㚝f�)c~��/a�8�x���p���狏����UY��XXۂ�Y�Ld4�F�q&؝��k'ʱ�p߼�ßµ}6���ٙWdZ]U�R�^A�����8�a�b⢕�Tҏ|��܂�����8����m�[�
��I;g�O��<|��^���Ǐ.=9�v���Y�I����q��3=�5�)�f�dS^��$��
x��r���X���2�8���a_"����d�$Nm�m0�&��T?�+y�﹢�S$�'���*&��ul�����M��?�6t���{��w��o�������`�~��)4iA�h�P����E�:�8u-�ױJ�p,"{AP����7����eNx-���2�$��:�vĹ�T�,]�`�,��T~��D����=m�"�p<,���}er [� $8n�`d+7��l�qRO`�r���՚�4����S;������W!�aS#�n;�ȴ��Ņ�덒�^"awZNsvy�)��x.�׫�d�fd��h6�>^BE<L��ܬ�j�S�c��uYľ/��vG(�>�����ڝ�Gp��UNK��q�Dh�橳�b㠼ǃ�f����K�8a��gu=ZG:ɤ5+I�TƊ��d		]���R�c�4�5��� �pe9���L�_��,c���������Y(ON4k���F�b�;�j����Q�d�D�iNk�1�]���|{.���,C�z�-���!*�[��߿{'��#y���z��8�����Y�qn]�S��ڋ�ً�|-��KIKvNN����ʜ0��R�Y�5�K� ZQ����r����PA��j��l�u9�?�T ����]�Y07m���i� }j`=���ޛ�F#��S��;�l�/?��_����/�� �>����P�����>��H���������%���S�1�3�۳!��aR�P|ek�o�G��[�g��	����ޞ8�����;f\u��e_�&OR%�d:��YF?����mt"Ǻ}aR��HO�Fu$�X���g��H���^�s[?o�9(�L.��K�X��s�d��c�h`����=>�`?Ae��8��M�@V#sT#�ʫ�\��#�#
#�-�2$���<L��4�J�L�����$(Sf��'�/d�V9�3'm �%,�~��*�25�pUbs�3�-��P�mBO�p�S)�����q�(�ގJ�6���T΄�M��޿�J��[@��z���鐩��Z_�ȼB��.i��f�N�pn1IU��=04e�W��
z���ĞJsD*�f(ʛ/"(k-��+����E������O���P��3�Y�n�D�11�0z|
�_�6���2���m��-꩎�H�	n�"�H�	i	ٺm�1�v�Asɢc�aHB��Y���͛��凰lfg�� e�:����PYtg]�z���KkY�7NR}����"�EwGΖ95]C��^�&~c��-����@K�A�|�7K��"߬�6 b{����o,�ˬ G���	�lR�Ɣ�I��ې���#&C�9Q�84��gA�=���T�a���� s"��F����y]?N�����ѣ^��a����޼{�����)�129�~S���_����s'���:�y�r��݃Pͧ�\���C�f�ub{�1���M���������s8�33�"\	����2��ͽOZ2�X�6��x҂�g���XZ"U�pd4e伎=[�"��|�5�[T��ĕ];,eIf�8���n�w�a�0'�(TPo��M��.z�+˴LN���������xmY�P}�`IZ�Fɜ��n�h(mm�w{C�s�	e,�r�JOB��^�9��GX�9O��{���q��t�z�ڗ
j��+]�>W�%�_�maz�6^F�6횣#Ϝ��s���^9��BYi%&1z��� �v�?�^/��c �Mҋ:k���h�)D�4{v
a�'�)�'����\���JN� ��JM��-��)s��9!���p~�������d��-�6�ѩ7���<S�����@�3B����Ly�k���w�j��+�8Δ�:m�$����NG>GX;Q�97$��"�&#�h�bhu����s�ģ�Z������yh���ٶ���"��Z�bљ!�脿��p���u�r��a�HE=�ύ��!(��De/��K�h�Ɉ���Oë�W�l_���\���{������/᫯���B�(����EĽ�����V�ф�� fh^���OvA��d6�9۝~�ن��7�{
��2��2��B��`n1Xf�7��)O>���Q8؄�� �B
��~]��f�nԞi9� y�ͩh0T��{A3_X�L�����k�S�3e򷟮�xY���0���ܨ�$�5�����2";��U���ی,2d��F;@-�Z1�~J�\F����vnV���2�C3l��������^�އ��.�ǫO�T]$rv��F��w����>�#\s_{@bR��{?����۷�?�{���P�D0yǠ݉��B�V�\���x�e���{wsn-#�����?�=_��R�4�}uo����'3�v_�oO0׉�]]���������K2��]?N���+��޶C���]���D*l4{���X�v�{a%�,�ؤr�2A�~+��h"��r�
s Z*[�4�_m���7��F��糥擵'bh����XS���0���?��C�?����"xd��to�fE�K��R����]��� ���\����αʱO�3�,FvɄpFi�FB�ƈ�J�R�@��c"��j��3z�n:W����uߏT�������L���2b֖�������q� T	��-�{���t?�x���zf�ml�$�뻯�Qٝsy��c(��� ^<��=�î���#���g;S+��.����FB����ٖjn3f��p'�}�զ{���9��q$���g{�����Ib�,����w��\��9j� �<�+�*K��>�3��`
	^x�r��݇�㻟��ƌ����;_A�l�Ek�}�@e/�6�p�cV�r���f�R�����e�8!\��}3{e�a�%�-�O�9���S���PjlE�>F3(��ܒ�.�Q��g~#N�4:�{�[�ZFE�J���u|ʷ	
�Km"n��՜��յ]�DB�D����Ww�!w@f]JӅO���#�Φ,�S�(���ӱ���xd�k#�:H&�-���~gIwmf�zj�o�	�i��SG og݄pUo��̝�D�lؔohBJ��`���G��ġhl2\����s۠z���9�^��z�x[����W_}��o~�y�"#�g�{�p~��
��-\ܵ�T(ڃ(�ĺ����T(Z���h���p�p�K� x�y<��h@�|��y`]�8(�Y�LS���Ҝ�	���~3�%<s>�%2<H`D�NƂ O�	R�F3�v�����T�U`�� ��Z�/`py�/t��)@SLG@˞�������S����)����('AKf����t"�
��W�c��f�5�r�|eG;�R!T-��s���3��M�@U���ԍ�����P�Ȉ��, >��=���}�S��0� D�..��o����򵸔E�R%����KK#K���d@���Jǿ){�G��v.
�+^�(��VU���j.%�����:E�Lŋ����R�2n�/P��� �}�="SfĈ���i쟭Z*C��Fu���Ȟ�-�8�ut��Y�Di�A�'�N!٣2����q���(�m֪�HCx�}z�m{���E���忿DYo��dY�̐�߯�vP��+��N��z��ᦂӳ3�HH��ғ)�Zr�ә�녝����{������&0���ަB������I�������`�͑�M�F+OLWE��D[٪3��iф�˽�_ƨ��63�R��e�,��,%���s������a���~7�^v��ή"{ĳ)ǰ�v��	��/�`�w�`�� �1���F2i�����A��4�Da������f �ro�ݴ+;8�0�P�;?�({6L^58#� �j� iF��Q�������F� � �4�7z�R��@�D|�MG3��e�7?`Z��s�T��*�Sy̤͠Վ ��ZQ��0}/��j�?��%����՞ظ���@��K⡞t��\Yy)�|v��ٵ�h�ʜ���v/|wt������A8�u��}��C*0Wf;��3�s�Nk��=�ʫ��ʴK���o��*Ý�����o;�)bfm���P̙k��́?h�6�����b�s$+O�3X�F���Ƙ�� �Qo�=#�څ.%G:mn�pRT��rv�(�>�Z�*@�W҅�n�{�*�),��}���S�ͣ�}��G���|,��#;#G��$6bS�R���axqz&�:�n�%eV27Fr4�����Y��X��0
]���8�^q���h����a|gN��%�`��0!ȃ�j���HR8E�r�恾{cZm��ڹ��~�JPhk�u�vOZ�؞|F�͵�궅�e� ����Vr�-F�������κُ�5���!(1�$%$��ImCը��;����'��Y�e��F�l�a ��0�}��q��?���l�өg{�0:v=��f"������
����S�
�3��U��rz��B�Z�<�#�!�H\_8�"J���A���z�\��v�:Ù���F�<zNL�eX{P���,RS:���奝	;���,gZ'��
��̶ߡv�ID
PQZcLn.~���Sg��1#p/�}v�I�vJ�}(i-a�M\#�3����X�׫q��pȋ֪h��;Ԃeޛ�܆�P�V�C��m���@�h�y���Cx�>�~������I8�?пYh�+><�lǍs������[6�w� !_|�P��h������k���xb��&r�3,�#it~��zg�ԌƽE�h���-8�]	1�qjx��o�<�}Ec�;��b� ���vb��J��骨�3�r����gI�F����i���W�:D��?�����J��2�@����8��C���m��3����p�z�g��1�]���]z���{�5��	�,�����f8l��.4���2zk�Z;��[��^ڽG�G�D2w2|��d��e�����lcY�6�'��R�j���`���u�(uM���/���B�Z	1�C���]����_�?�$����d�����B�4�L��7`*F�P��1�r0�� G�����Rf. f 5�	/Y��#E*B��*�",�b	�B�a��G Ek�.=3��D����d��D�>@N���B���������*�g��ue;Qo��f[\�+0B��o�~G���V��b��Д*h�d��ik��z�d��E�Fѷ{���w��M�'k�V|��Wv�%l ��S@5d��V�}�d�K�nn�AD��ZA\���_kl�-`4c���+���OOe����(A8�4r���u���ݯU�ӛ��{�㈥��ʾ�+�*������:7G<~xT[�}���� �̨��S��ͩ@:�%�Ja0��`_d ?�ưtMЧ��)���&��ck�ȋ�@���.�G����Y��G��*K���lS�H<63±2���✨��̅�[��V	������������71��a�*V��lM�H�j1&�h���i�W��-5nvc�So�\j�NJsPݎ���/�����}��y���	�ڽ"ೠf]������	[Ըj5�sEI�tcɅL��mրC�ʜ�29 q�ԎzQ���%k�.��	�NO3���l�a�,V:<�ww!�����)�%r���}�t���o}�)��p��j'���=YT$��-� |��8CF祈(�,JW�$f�[q�B ��r�+~X�8$;$8i�nz#�XkW�H �<f��sM�ţӥ��p�=��r�(ɛ��1��t,�5c0�t���A�[?��Xף$������?��L���\���H;�8C\�i�:b��;\�2���l3��-��̉@�ݎg��{}9��� �>��N�L�Y���2jc��ok��{�4D	�o��<�kEA�H�"�<�Md�*��[�@�,���=N�Ƚ��rr||�C�,҅�s�������?�7�7���bn������1#�(�dP��� �Y�&�{��P��x?��J��ӛ��$��	Ls3ƔѦ���QMl �f��ͫ�0��� 1�ߟ�ވ8l�Y`��u���֎�l�$ǃ�d�Gˇ����XT����1A�Y���Ἕ��{�(Q�<��>31ӥ�����1V�+%);{���G�V��Ͼd}���Co���LU#�k�蛲�OO�	-�1G�R��7`>�{����U)G�X@�p��<|��o��W��.�ۘ�NT�go_�Gadgl�muxV7�m����{��}����0��WO{e���ec��' �h��������Hs�ث��]�,*��Z�,�v�ߋ��²�Q���B�-0�uE��U�<VG�X�����*��N��ǗNvS:��9��T��7���jd�kʄ�3�Y�#� K3N�)�	�ǩ
拳|Ü�Le��&T�~���йj�����V36�
�pb_p}P���'(xkg��_�h�V�f�Àb�i���G�Y;����"��c�|�}��/����7?~YO�,�,�K-|p�g؏�b�ֹNd$�Gt��7��؛��m�2��� ��hrl�(X��XF�r�9<� ����
����Ĕf��~$��{�ȗj�8��4R�"�vˁ;��)ݸz	���L̹����J&��^���S:k���B%��_�ǔjw|	�E�7H帆)��]y�v�zS�f!��r�'��:<�?��=�MVI���H��������C�.]�>ɨi$�ֳ#U�M���aia~ya � \ǡkWIowmι���P
�2�526��}@|�Fxa�ksX��V�#^>��)rS
�w�E��)k|41����MrU M,�}|�o߽?��1���]x0#ɜ��.�46%�H�rq��`�c�Q�w�Fe<�!�3��c'����2�����D�|����>f"��B��@=�<>�������s������1�u�v�!�	��/-�IF�s��\$e��2�>$pW�w�?cTd��?�g�4
��Щ������^�m�~��B ��會����̃]Tl�0∢�cϒ�gQNe��}��|&�V�N�y�+$La4�xL}.^|�0F��[Π�d�\��,+���S�#j��9g����x�s�)&뤗;6�Ț�s	 �')T�г�z�	�7w�#�0(�
`x/�W�Ӫ���ES]�Ŝ�)�|.,8E�܉�hwd��!9 �:�e�D�����Kض��ۏ�hӾ��S�{�W��mLz�6�:ԟ��#5�2�M��4-����KU��������R}��2�>ˮ��T%��w�eNŁ�7�����n�k�'��N#Q�3���ݮa�J��L���-$�c�����4����iN&���<"��T�E���D[�����&�D���X�)���͋��9S�����N�2Yr�`�UD��w����W��)*� $�=���W�'�gv��D�Yȑ�� ̡���E�+��Pu3X���#���EV������5����E�ń���Hp$e(��a�X�I��>,7S;`׷w�i�mj�J3=);3�X0���1��2x����LpyI�`�n�|W"Q6m������C��s"���j{_�}�}�����_��e&o�h�B+��������̂�^M�xN,C�VO����:Bf)�&�a]�447Z����A�<2�-*BkGL6��A�Fe�w��>}��l]�Ңo�7�Y���yƑ;�S'3jM[bw�p@�����++���K�6F��m>Y��
/��)C���!s��a�������� ˙�������yr�jLmo�wʂCD�GGiY��L�s`K�QKT��Z�FvC�/ }=��%I5
�$�m	�m!�v��UYP 1@��޳�
�
^	$�*�倛"쏆�����#��{/)Ͻ�<իN'�b�G�H�*��yx��&$�'Y'�v��i�7�X��A���,�a�ݏ��r�T!X-&���X��+����	t�ٍ��ImnN��2VH7P��s1�ts�I�kdNw��Й>��^z����A_�M���(�
f��eN��2z�6"�w����o�.j������:r9d�Tc�U\�t��:	')~�����L�01�H�6��Qv��%\Q�7L@�,�V����ݞ/ָ_!��X�Ȉ!��W򁒳0;��Sȃ>Y�;.	yٖ�6�)��~/f�~�-�,Bڣ�[p '`�nS@Jt����U�|���	�u��,jʒ#��(�R?Q7Zs�>a��A��˶�eN��/�gYP�(d��X,=RR��
�k�OO�C~߲�}=�v�������20ܖU?<���;������$08�A7����@+��\*���末v{[=��K&�͵�W�J�����w�Q������2R����_^��z
[T�U�H��2ʷW���l"&��U	����8w���	�#�z+�H����H���mEƉ�*��8������I�ݷ߆�e�d��a��KvyzpV'UF�+��8�����{!g�n���JZ�+sX �V�q���IPHJM���ƫ����Ȏ�����~��P����Cx0�8^LT,m_���XVMs��?��i��它��p��^���S0	��
��=��1ԙ ��Ge��[�Z��Q�7k���΃e�D�d�����ؖ4��Z��ul����F�{ܛ�l�8t��\�oAeI~����Ո����%oA3�� L?~� �U�~nS����;��/@p��b4�$�<'5�C�zt^����e�$M�-{�?�S^�
X^2�-�ׂ�.�лFw�i��,���������u�ԋ0������B���۹w�؎#��i'�eS�;�m]F%o�5�>S���J�
g��v���g��V��Sצn��M��N,���BR�+-�gZ]� xu ßUmٴ
��ƱN��%1h66�x6��@�	A�ܧ�"k��SDL\[����Β�^nl���6�����:�6A�#^E�Q�H�'�,�{נ��L��@�F��O[��8O���3WD��n�n��_n�_0#�)sJ01 ��.#K��ҽ]s��Ph�\e���<~wtX6��j%�M%�Xnu۰�I��f7��J=(��|b1��l�E��%_�:�][�ٰ7-��o�mb�(1�c�M�&އ��hy����9+^�ޢQ��>%�񻼹��ͽ�~<�<�M��,ʆ)��)ў��=��]oIt=� ���%یqU.C6�y���<o��깤�S! d4��*��Ĵ��R�%B#��v�� "��*
dp�����j�}����48�z���T��._�Y�^��Jd��c�m�z�P~��e����&��peN��>� T@
�L9� ��6�1���:=ǖIA�����ûO�4��4�-V�.�zR&B��ʑ���u�S	��Sͦ[�yEVy?����o ��zꩽ�uC�T��������u�yײ/xɿ������ �#G�V�8���И��ӓ�������ɹӆ�nlYW2����ж�f��H��ݡ�Qp
�]���ƒ!�RQj��> $U����W5�RtD#�pa�J%��iB�(&��C��(x��	s[�;s2:�z�{N�(�9�.�}	#E����~ �y�3����M,H�M�*V#F��B�`�����A�S��}Q�#Y��v0�+�)��8r�p�;'�	
�E^��6�@e�,�#2����Jck9[{@�J�
����g��s�ߺR;��J�ɠ7��@�����ګ3TX$t�Od29	e���W���]*7R���DFP�R1r�67ם��y�%e�ۀ�M�x�ʷ���3[��DR��j���1�B���ͣ�~�*S��aS��kJ�!�l\D7�2\����)�mBHR���v�F\T�j�R��t��m���;�^�[>�V(��}5�O���`Z�^'�5�=_YX��f�����RI��U�'��Z�D���x'�3Bm�?��c�~��2s�A��˗����.�f?\̜S� {#���no��� �_2a���b�A	�Y}�r	|`�d�?���8�)K\^�Y�5g''�����vV���+8��F�3�=k2]l�+�CXG��g��th3�hζ��{5��ن:�ˡ��n<�"�����¹֬JB��|�Ol���R��� (�(I7=���m�JPQ�,�;��b��K<���hȉ< ���rS�K�x�������{sH�z�:\��6,�hN�*�A!�8��e�1O�_���F*���;ݝ�:.�jY��Ճ9�g̚��`��G�v�BdW���	
����}����6��W��p'�x
�֮9���=���|�A��..ã���R׈R�L�ʽ����+�n�}���0�������)���-�q�3�q�Q/���ю+75�����%����������;����p��� ��n�G���
G��unn(e�\�|�4��_Z�9�8z5�u�Ɍ���^�o*�cbB����{��|y'rU�$C�������/�'���U�G���;����G����9��f����	�֢��Ϋ�����3-H��9 �A���l�N+I�y[�%�T<Su���y{�rd+�A��^4��ð7�52���Q�a<Kc��U5ڎ�������K��^O	D�.���R+!��#��� ���l����,]LA���2���
�X���핁���ܵ~ɐ��N����ec��3aMhl%_��$����V9O}�d���\������3۶�zcP��k�3�y�AGl���(����BV�U�S���@u��b� ���n3���c�|���*-�.T����J�"�
I�U�:���i��ʆgE��[,���������a�H���m^���8� ��lVo���D�40��'˂�`ᄶ(pg���0�9�hDs��+�?X��T6�������f�;��*��
[�%s�+P��гC���{:
W�WbM2��9>J�;s����~+�=�e͉f. "@ݿeG!n�*)�M��*�W٦�Q�nKrn<��=Ē�X�I��*� "Yh
I�{p��n�?�S9�ü C����jD*�z��Le��Q=c�b����ؿ�6�'	��G3�����]Ϸ/_�����d� ���E��(��� �f�U�Bs�d5)0�-;j��4ON�E���G!�ga %���%i�`�_.u���_�|^��2gy0I��K} [�U�>o>������Q���N���%D����,�(#*'H���B�r�:=����@80�N�\ʊ��ܵ��s�(��� �8�oB�_��8fÖE=����M���+����1(y#���[aسH�2���}/�]�γ�Vt�!�Mp��ƛ��z��L�����j������{������7cf�3�Й��'(w`�"�����_"ۇ�u�� K��en ��@ �i���_#ή훏o>��ŵF�i����F$��|�/�Gh?��|f�n����_m�]�����c��=:��r))��L���r��k�%b)�5\���,�A:cfyrN�&'
�[6�s���>J��5s\iܲ ϥڠ��K��Ƴ�L��w��[��&!����*y���������3Χ�,kN�w�L#���.��L��_K�2j����;�䀫�ޥa>|f��+}R��#�5�vB>	��{\V1��9�V�9��ng�Q�$�t5;x����q/8��T8��kk3;t�YGe�> �����F��R-.�J�48::����;�oQ9s�s"�ŕ�� �Z�؁C�Cw؜�
Ҁ�X��拷��էOr1��tP)�P��P;�6��{14����:b05����|�!g���2�ŵ�`*��ic�x=SX�8W��Kt�6˯'xT��l8	����&���G����&kĤ�f�{���������ɩ�{����{���RF�I�����R�_��/��𑾋�*��6�[�utΠ�Wq�G9�ed���CE:Z�S�Ǜ+e�ޡ�:��۵�U�4Ԧ��2��U���YG��mƤi��?I��9`��^R�&H�b����1�����㴦���<J�I�Ȯkh{�����<���%Ty+��h�Įe����Q�)�����O��cCօ �@����@9����p��7�2��N�$&눌�Ϻ�7�?��ѽd�\J�񐅤�G{a��$ώC{��kᖔF�b�R����z5'��|�
=/� �����=�N��ݖ��y�d�WWW�ݻw�~��޿��>|��xG3a!�<�l��7|���G�'6�	wt�|��֎-�p��~Cקk��S��O�8=�;R��}��r�gN��y�@s;g�B�đ�P��?�z�&�wfԝ���no�3k^
��[,l��`�#���.�Y�8�Μ�o�.l5Vl�Z
Y[��3ٖȼ�4�^�O��γ8~�z���Jh�M�t�	�ϙ�h�/���0�[���f��#����3 ��*?''�D?�xΥ� Na�qǂ�~�EkS�˲�x��4�
,��&��L �,�\k'Q�]��W��]�=0`��*�{�?&цX��^�B���kU7�\���^mU������/#�4^��Z�I�M���_0�T >̱��R�4;|gF���N��G'���\s���}(;�q����?���,�L����<d1�^���5���f�R�>[�Q��
����H��	����E�Wz����$���e,�83 m{�6�a0�HX��]����z2d��
�G��s֧4��H��V��&���3q������e�w2��Ly��O4^���q��<���_�Ɠ0@��m�_9`HJe~�6�[(!J�V!@W)F��2;������F\�6 }0_G��&��/FSe�߿z�����2��Ry�b�
�9Y��&"�B��W��x��w���Q��ޮ���4t./B{�U�Qb�N��4+ae�ײi�:[+0&b٢��t�͝� ��Fۅ��A}e�²8)���1ː���C�2��M�ȵR=�j������H��˂;��S9�����Cx�u���cW��UGs���x��8��о}FvR��N��3�,�Q���L��,闊�۵^�kz���^LS ��R�]*�*$f�d����γ�V�/��q��W{�����J����qy$h��s��~mg'���!���Ƣަ߷��]���CI��af�y޾���K�x��v�{���\*[|*�&��Ⱦ�W��=��a����7��u8�����0k�n�ٛ�$���>��щe�����<�I�Ƃ�ڂ������t������
K��&1NӪ+ ��Z��4�-�]��l%��F��vv�����L��8X29fRlb������]WY����Tʠ�r�^pMY��r �38*��$G�'�3Ͻ�1 �yK-�R7덣L�������#ɲ+����Rg��.���3�;C3�ښ���1�p�-�U]*5�v��w�{��-4��J"ܟ�w��D��Ν	Z��'�4�C�N���c�ߏ�c�K~U�t[�̂ ��s,�e
���YP���N͎P-�Z.�5F$�	*]��eǖT��fcS�~��[gً�q�ʖ��ӻ[�����퇍�/쿋�?���ݲ5.Ƭ^���{�vޒf&_�"��i�_��A��yG΀����A�����u#���ڻ�h�B'��:�C+
�E��2� ���k��=q���ҝ�4�>�m���<e���=���.f��9G�#{��7k��d�o*drx[!eF�"�2�}�r��5WB�����!����c�a<"�[:��F&r!�ɒ��D�1��۶i����f� H������pl�/m�,�Ew�і�|D�I���a�~�.Ա̚g=��Db_�'җ��H��E�s�Y,
t$���=�<�,ۄNo�7�+i㚳�XWν9:����Pd>�ô �ʲ��=7V����Ee,�XP�l�=�z�LAE���_T>u���W��@urs-��0?ϯ�(`��y���;T�0���l�*���;׿���*v-��l`B��d4?��	dXf\qXK�f:�Bo����p�ټF��,bi�0��
/��7aX��t��5�3c�6���
�5v��><<ۇ�a`�oNٍ����-��Q��,��SQo��c��3`eY�/<�����[,(�:��-��r|�!�ɥ�K�k�����'���F%m��%yI�aF���*m���?�liG� S�zFo�v����n�y������Q��}�%&��*NK���m������n��ޱLx�c����~	n�-fO�ӳ�3��'Ol/��K�ް�F5��jTך�R���Z�=�$3���5��Y%�h$0��Uo�$�l�hWN�3��U@[s�i�f?�+��&&!�d���!�9���2�(u���{��ٌ��$Sּz��K���'Qi����g�E�׋-?o
Ft��_�U-*T�4G�m�B�8�
I��vصgu�s GI�&: r"�
9���l;U,Ͻ��Z'j�̃��'W�.on-� �<~O}����9�n�7��vFx\���L}���n�j��Cep
 ��7�
{�j��4P��c������Z$ۃ���Qs[�[�F��[E���ZyQF���r �r
�����B�6>'G����
�l1�9]��RUߓRd^҂��c!��L��z�-��Ĉ��o��}�4pB�㼛�i�b���[��R3E�%!|Ŗ	PVő}��?�Ȝ&�ʓ�$t��BN��.�D����gDE�W��A3�m��;@�TP�*�*J-����P @  蘻R�4N�X�3xrt=R�DlYf�jS`��iC��J!fD�q���_xl��|z�������kEI�uO��ت��o{��o���%`^�{Q=#�b�"��>�it]�U���d�����^Y�nU�j�CjGb�:9/��F�+�F�Ԝ#Җ3˒�_;ا��r���]����a�#�j:�#%#�mw�P���^�Vs��o�%j^}aٜ���FLIbs��]qvom	,"|����v�!u�j�LF&̆�J���<�������Sźo'�Qe:����`]���Rl�E߷}3|8��eW#h��\Mb�ՒA'�MJ\�(R9��� gg��eY��!�n�;b���U� Ԍ틧�Z�L�>,sd��.� �Z�HQ��KUg`v������M4����B�pڔ�A��3B�b�����8�?{n��C��s��y�'��zk��e�]�&Wu+f����VJ^6�#����!4J,���@���*0ɴ��G��ѵ��i	 B��'-?R��L��U<�'J��v�DO%h��"%�^	����eW���O�2[�|4�Ը�G��w��_��J�O�Y'����K��Ad.񚅍��{x��$�Mbڭ�y&�٩����6%_q|��R� .	�CjC�{���1`��8��X�Y��� �LK",o�'\d�E�SeO<o{ S�� S�(fD+U�l5Drn�S�s���/?�"S�/��>�/�l}�\ڔ{q	}����!��o�-j���}�2���_��}ѥU��s���1�"���YF��y�� ���ō��K�tz.���2�!�ly �U�*�M[��E���ce��?�!/p[@�:�71`��l\�<�}d\\���^�,��2ܱ�?���8��w66B57a�I�V�I�� �4�ɂ�h�C��R��_rX�����l��p�����hcS����gmk{su��p��Q���~�Q!����E����0Ǯ���|r�2&�����l=?)����L}�n�Z�8D�F�9`������P��r�2#J�#�X6���措ǹ����g�����iͰ <:y�6�l�t۟�/>{��a�~� �����-8y��}xl��}��:����5�X����T��m�;�:?���^�y7�A�v,�ꘑ������M���Ie�L�%T':�?��cgǢ�Py����GX	�ⲓ�r��pr�*���3s��R/���^rm"����-�[У1�θ�7���-e"��\�#��+1a:�=r?�M@i���r��[T<>V`�z|�~���0�Ϟ�g�B���e?-s��~z�?�jTs�fp�K�){G�٫Wvv�a����F��d6�R�?��<�{~�8<�g����_�,����U�����gD�.*w�n_�˻[6�b�=����9�����v��p�k�3���LG����vO��\�rj���M���Y������ӢX�a�ww���ߏ�6}>�A ��^�A'>l]�����K����y
�X�kd6v� 69�[P$'���z�	��t��>پ���Ʉ���s*��*g�i������[}�`��Ix|�(���� Iߖ����)4�/i����G� g.��R0FT%��g�H��/f���S�n����nՔ�HZ@���jp��GdN:S�@c$�Qۤ�{�aی3�	=�*�=VN܁�e ���b���\Q?����f�W�dx�Y(/.*�l�s+�sf)v��v��0?�m�M�^s� �"
�Y~re��n�X"�a0ʤͣW���yrq�Y�Ү�ekWXBƯn������X�*�-0f!Z63�g��Y��O���~�J��(��݅8����Jq��ٽ���	�5+��e�DPǽ\�:rV��E$=nD��x��s����C��Y��y��G�-0nV�4�4M���s�2�vu��Q��?��t�m1a9á�Lc5Q�}��	������ E騿7O?G{�>Z�o[��g�l���gI�^T�]��FZ�4+��(�4-��	�b������ot�B	[G�GfEo���F� �Z��^ח���ݑ;�V&2�溜O���?�l{��蒠sل���e`@硜.�Q`Ш\Y�ʜ	=`*��P�P�V�\��d3Xgd�L�O���j=��a/
��Ȍ���~;���ƙ�s!U�LL���ef|s|�u߽��限����[Y#�ݲ�YI���q,����F-�����uڿOf�f��Tfe�bhv�7ꇻ��'��s.�n��`�û{�������-U������f�tlg�O�F�������8p�.�P�8(���£�Ga��U�Zc~�ք�N�1˸�f�3'o�DF�XN�5��;���L���,��DU%?+�,ff��m)�J#B�걊�m�p����?4�\�0�,��>�z�=�W�L`T��:=��q��`�?mm�PP!�+Є{�g�Ng�ɪ�Nc���/>�<�����#�&��������mo��\�e:O�sә�t��}��T3�^'qlyaC�@�-�/ ����a��Y�`�Z��7�j���6��Ff��S�.�80Fc�g����f��V�q�C˘����j��/F<0�<���Z���6:Ɯ��2Z.����� D8��K�f�{1jw�me��.O���~H:�;8p'*U%�@Ap�n[�v`���ᑐrU���e$�>K'�|�O����pD��v�J�����At>~r�rݧ��U�A�P �a���0f��ZO��=q �P=.c&���q�=$!my@2��?�'3�������z�Q�����q�2���POunF��T�"� ��[cs7�Ѓ�e�%Yʂ�^q��^w��!�.&3֭�t���b�d b�����1cI?Q�ϟ�y{���޲���E�p����#�ڴ}���IJ��f�5�Fӓ&��7���%Ƚ��вlil6�����ɫ�9�.�9�ϴN?��>��JX���`02��y�ʶq�.l�3;Cx�m�������gfh��ڇr`z�RZi|�KS��C�]��9��#� 4>BEk=��t�r������tV)��[��	��3s�p���	N�Vc�f+�3��)�����8B�� 	�';[˻i���m�G�gV.��]z����F��,yik}gϕ�������Ȍw_wA%�������^�S�86	£�ii�26�7"�Az��eA��g`?{||�ZչOP@)�C����a�s���W�_�/^~f���j��pɪtQB���ڂB�]/,h��-#�*	�9l�܌I!��������׿|���I��%��
�����n��O���~�+q|2���@wU�'B������v�	%�m$�C�H^�x!���n�V�̼��h��a��\Y)�#���o+��?~/�46������}MelmnH~��?{�=[�s��/��)�HI"���p5Q�L��j5�,�������ww��~��/,G�I̭D���>:��KЋD��~�<��/�����f*y�$��[���4z��a`8��9�m���`��<�"f��9��`�	�J\�+�}�7��M�Big!��eby��}�;�����i�8���)mon�/^���,P��������k�,||�d��@3NYˁM�3̼�����m3�G�N��h��Ӈ �^�5��2$tm���H44�nG��G(��xNd���xt�"�Y�:�TXKU=`2g>�@BP��� ��J���C͞��w�,nG����\삞���..�6��ʫ1�MLK��t����VI��c:T�U���y��O�[cG�R@=���%1��3�?�m���o7���[�{����o����L�I��h���i�7?�� d>qJB���*�ީ\�a���k	?�>bU��}&�M�'0�-���k3�=o Y �ږIQ[�h��q�u�2���=y"�]{.�مR���ef0�*�y���N�p$���8�3)Q���(w@�hT	 �o1�����F�6���8f��G��k���T7�8���c]Iǁ/ʾ��u�YC���+�<�7׷꣒�n�:Q2�T��7��f�����3��vË�G�pw�Y������w�W�X���<�nn	D��5��	���H;,�adN䳗��S[���1�In�RP*�l>}�<�����O���|1�����]/|��!\|��o.�|�B� �}�����ٛ�\�q���&%>�����O̹U�̢��P}4J#Hƛ�X�|H��ճ�>��6�jT��*��v��UN�6D�Ud����gZw���oD�;�ZgMY)�C��q���0"�C�\���Mя�����c�_���o�t*R����-�X�S���E$��5�ٱ ��}�˫{9MyS%��+V!rD�|�N�~��~�2'�Ȃn����b���o���m;0e�m��;�!HY��0�E�%�N�J[e�6�ٚmȞ2Q��7�dV�	k�b؅T����|+(�Ւ��+΂#�xndIk���[�6��˕�M����?��G�@�甎*��@�hD��r�R����/��ac�>W�2�i��,DfDp�߿�)���~|�&\M��)4rHl2_o�C��Ç���d�YIy
�L�[U�U*���!"�8D��9�� �#�P�@�D(=�FY/����L��9F��@����mIB��0G�P�-E�l�m��`���?~"�ʲ8+��|��5=[�]�v�&��]_��O�'h3��*�ޓ�-8���ǟk~�Pf���{����[�qr��ՀI�y�Ҵ��2�Q�����B�L-#s����u�]_��M��5�F��~��{�����[77�2�
T, �<#ϴ��̘ �	Ҙ`���.Aj>d��v_s�:Gf�_�QC2����f+�$��R~a_�!p~�m�Za�>w�H�i^N�j�am�������ֳ���0��?�:�c���eB�1��ږz�qse�-� C6o��H~M;@;�B!ci����q�o���N.���������P
�@pQ�Q[��?���d�d��;{a����:v���X}��}�uX �AV݅p�V�$����o����Ҝ�W³0O_����&�ƪ�q�M��v����pEp�\�µ��/w8?��}��"C���O�7�`tGǫ�!`Dz�0������7>��U���^�����ϪG)k��s�?Sk��4[�Z�3�XQ��G�	���� �~��lkG&*�wp��p&��D��ʉ��� 9k	�P�`V.����t���T�j�++��ؤ���������TN��rn�<}"g�=LH�B S*~����s�Āԃ�u2a��̴n�lwv7-�<���~�,c̀����C`1�z̬I�W���}QJr��j�YbDq���٩�"�p(�$��à,���,%�.B"��\Ƕ�T*������/xR/$o�h-� �l�6k�U�L��%a����P(�?;<�}������sJ���NTq^�#��9;�~�I�/Gy����3�ia�b�cyZ���0� ��9٦��;�y�.��Ԑ����	m��s`���9O��l-��Q>F%`��$d�E��!�XZF�q%���5l�Z�kAV��5oݎ��c��?ن~���4�!��=77(�SN>99���I����FJ'5���1�s�g�Y�z!a�Vâ$�f+
�C+Dj�r�0�M$��Q��6|6�Nx�Hk����3�x�)�%��T��|�u��GhO���<)��}^�t�}p$�����lؚ��_`��TzT���N��K����v������W5�k �O)��5������9/��ʬQ�b�%�d����Ap ʙ}ތ��I�ǜz���=�Ȑ;��m=/���������Wt��2l�؏@��@��U͂OV����[Q���M`;ן-^�~0�'9�L�gk�� �g�=Иd�lVДb;z�n⨋Or�1�������0�ӄ;�$��<��H��@�!M���h����c��q~6����,>� ��dr���N�D�j������c��߼{k��:�;y�+�����g��w���ek���}J���<3�l�)�l�h��Q���6�R�ZpC�$pV�Ԏ\��IP�ȷ��k	��EE��g�\�L��v�@ >�`����!%b��YM�
.��|[�-$9��?�j*����HR�f�U����a����*�~�V��w�>��x����pf�58z�H��f��{��eXڳ�M��v�;���/s�u٫�-�e�kC����f+�Wu�\+�R�-�9��.M�c�P�G�bT���s����-t�a'j���`��z��n�^W�w!�ԥ���(�H��?��ۃ/�g!��y*�9�O�Rd��u_�Ј�O]��R&�b�-']B��,Lm���T�ڴ��Z׵�;$ٹ�
 m�Y��]FD� �`i���YF�LwP� ���a�=��(�!sF��x�-ZN�8$��:RH�ZA�c����8w����m���6�mP�:��1s���У���p8��GT����m߂�c�7@]���a hA����w4�/TA@9�l6	w7.GX!�E-���4��Eӎ`�{����=�fɰ0�	e�w�k��-�O���p�8L�]��@��g�b2����ƥ�����4cO��^���E�[��w��I{��y��_��:����{t��H���mK/k{����ր�PS����@�<9p��]ŽG�I�������q�OJ��Nг�3�2-<ݒ�Ђ��R��=ǅ��܂�!�����w��BT�!+<VG�h���Z{66��:��|ӱ�]N�SK��Q���0��3���&X��tV����<�����၂̀�
�a����&x���( g�\�i�R/8P4�n��J�ќٿQ������w�k� AUR�L��\t�t;����B�*Gт� B"��ʧ	��g�^]�Û�{Q�(�{�!�ތ%���9�%�#�)g_c��-u\�K��9 ��
_��Ԃ���`���9[q%�n�R��u�I��Gz�}��T�كru�-&Tt)��*[.��;�5U��G�
�AU�pO㫹���G�l*;����>o�"�h�,���ӭOˀ� -�F�A���Ŏ�Z0�m�Y����&�T��pr{��ϼ�m�v�� R�{t�v�93Ϡ�-
l%j����9�(��jS&;�4'�w�� vq��garw��tJp��d(�,jGD����u^�z]�����!3tn�d�H��:�XQRT���	P��DX_����|n��*];V����*	x!��Ȥ�,��5V8RŤU�{$�~�7�T�0$�C�azK�X��:1?�C`�Lx@��/=�"�[z	�^�|fN��PP����f5�`[;�1[�:J�%t��!"�������u�3C�p���C圾S'�Eߊ^��G^GP��������R��Vw('��d�)3S'%+�>�-}.U���݂F���hUI@��4����2G>J���E��h	`�sx��+����O��a��16%a�v�I��e=FPa��m@B��1����_���?���7_�}8�t���A%��³���~(�"b�2<�{��������5<�0J��&oF���e$�'B?0���P�è��:?�ÿY�~�(+� e�>H�М�6Z���e�����8c%��*��1�����X4��h~�
����;�P �D�#k���4�.�a���h�I���5���������T�) �l98x���M��h-浐�To@�/�W���3w��'e�,sU��J9����L
?�^�y��M�1ڞL��|�+g�"�P��L]�����" A��������&�F�(+��!L3�K����}���$8%XA���*���
�����,*�H�v��^���)Aa- ܩ�<1���2 d(�L߿�y��sa{��9�=��*����\�4io�3Kr����U�l��&�K֡��'�V��U��MIC>9a�����'�7��J8��l\
��idqq/�C�oHn�h��j� wv���:� �P'�Xro�7�ˁ�+1���)[O�Y�-�������߆���p���M�u_4a<7��q�b�
o�݊�ns{W�u�gWr�,�ٯ䄕}����"#�((�n��￱������r��v�VՊCC�����[��9ڒX�Nu֚Y$�ZDf�M�MA��ͨ��m{d�9ec�	4��,sXΖQ�a����LR�ԅ"
0��ԛ�s�W�a��H�5�jܠؠD �N���MG�%{�������F��e��k�z��lor|x�i��H�ҢcJЖe�!�`- '���Yt��p3e����)t@�̐?9:�U[e�U�{��1�oCW�������w����f������d��� �7kwy7�ى��}��{��*ϧ�ۀ�+A�^\c�d&=a+p�s�V�b�|=�*0H��^�1�J���;d-��9;ֆ���%��E�8��˱��f��E5���V�V+�]���Q� v􍘁�:�`4��@��3=��3��	������NT&
BVK�׾ߢ f��V��j��:]�V�$��n�~:<86'��,(l��	s/�|iM�h�*K�XC�����Ջ�� Ns���hEJ�ё�/�N� ����e/�ᾃ��V'"����N�P�{�����\ k쳷F�7_|)gμ+��
{��o
{��N�h�μ��hT�H�}e$r.�gܪ��Gș�Tޯ}�"g�ȶ��MyB�r!h]��5�z3���w������Y *�2��{�nz�Lڱ��!�et����l$�ì�P���ً�@�znb&�zo�\|�y��;s U*}�`#�Q
��}>X ��tZ�{����
qj T��V��d҈QZ�ĸ<�p*O�٬n֙��,8}n���bt�
�:�cQ8K���ňp�8�*��S~&!)ʎ��Oo^���lS�j@&��(!@Bb������E蟼�����w��6J��*�� g�1�A�]w7�#S-w3KΜЈg����]��_iD)�PڜQM��|%�_��뫫��7߄��ONpO�FHG�4�(0�0���=��pWH?2����2���Dk4�D��Đ���^�;J�<JT�k�N,�:��)q,��5g4�yXu\��Q�JY�/�RFP"j�6Y��s��d؝|�q%'��e�&�m1����"<9~d��Fxn�mU�X#�X[:N�1p����<�3e�j��C�Cm��F{�Ik��b�ك����A�h�U4y8yd��;��h(�"��� 4C�o�Վ����m�sv�I)�\�mQ$�y�_�I��6��:�W����=��"��0��iY`���<C���ϙ�µ����pv�|��&@)mW��Q�P���ЩD�z �����c{�4�xwu���k��Ζf@�.u8��V�L*H��PQI�=W�X��,�Y"f�W�9@��Ϩ���+3ʗ��/��
�6�g[��߅7?���`�&'R	B4OkO|8h��|t�X�*����9�A�~�q����\�^�Ha���\��vm�U��{AC�؇�,XT����c5Qƒ��|Pʸ3�F5�o��h�ݸ2SUy ܊%`!Y���9H�����o��bf��8�gEi���uc��2�C��B���Dכҁ9+�����J�� W��S5�2ۗF�(��E*Y�(��΄2�p'��y��{ﶄg��� k���w��b�м��� �Oi����%�lZ7Ty.��7�P����pP�^Z���}��؟�N�l�%e�l,�;�8$/؏����}L�{�t���7x����D~"'Z��;�IO99aٹ,��&I��g��4��j�Kة͗J�1+N���).�7_�X�J��髬S����q�Q��󮩎�3%h�G�j�i�Ǿ��S-���
��]GR/-�����٣��]u,#����n��ys�=�k;���@Hxc��Zs��<r�6^��~��.@�oz7Q�W ��|�΢���gO��?|����W��Ɍ�J�|P�K�W�M�Ulc^_���Ƅ�r=`������J˝q�w	V;�p�Y�}p�0_AG�R1FjE��O,�8E�/�Ω/��ݗ"�Br��5��*��W�od�N`
1�ֆ�ٸr66���v���ak{W�f����\�x��jW�a�kw �|dMەm
��u���MuM]�Qz�E'�$�f�>�?|��q�*��v1BdB�#����ml����4�@�Y�Җ�1ݝ_��3�0��a�.)�]K��l��/�f��X�
�x*6�|�{���BP��`�"(���vM^Nk�E,�E��g���+	���?{&cĳ��2Ck��Y���=��k�	����JR��'*@��V!�k72��~:��á=˾�iy�s�@?���9(9�8�̣Ofw"���CBo �������0fw��c�� �۠�a���tl�ON70"����1
R|bܬ���:'R���N��dU(|NY%��eL���4d�Ih�^с�������̃�%��ʃ;pF Xt�o��hQ߼~N�N�M��xq��*�޴�8�������p\M�h�Js��]�mjq~Ȃ��i���_��p��7ډv��uJ8�1��~�v�ˢk���Z^�i�>oK[袶@�Z(�&����>�k�����oOO��ݲ{��;~��K��'��*��˱.�'�&H�2���!��[�G�t�)^�W�,���_����zzʷ��}?'1;e���R~��^;aNr��~غDơ�`�o)�-�����#��
���&�l&�K]m���_�Ĺ�Ut��x&�j.[�(^I��	��aZ�=����Bt��:��e�j n*�hY>���N���8����ӕ�3{���X~E��vؔVϲn���U�WQ�I Ⱥq�e`�2aP�����"�����l��:� �0�;vÿ��U���Ke"#�� "XP.*�����(�H��p�\o[��g���2Rao:5��	�y����X�1d��M�#���%�W���R��qʔ�Ч��7^���
N��l�r1c��FUk���/ʃ8g@�%�IBd��ix���E�R�_iOrg-�h*%�"ғ�Ws��X�e��6�h�&:]w��(՗��
�x�)B����-�lEŦ�yb"��z�>��!���2���.��7/�V�Xâwz�.��\+����HsJ����f嵕Cln�(��S��@��e7x��qx{y���u�^���؉/����n4��N8ʻ;�5�Ƞ�Q�y)���_�s3��m
���	��H|��gN�����qas�������@ws�8[�L��Vш��6څ�5���
Ǟo��.(.�1G���`g[�6�H$A�ۀ�L�"}e���F��bEk��������4��ԋ�J�x�q����d����z����;�̸��V�����d�N�f0��kGߑ�E-9��m*?ϟG��:܌�"��q�Z�zO�y����m'�~���K-�����s�	!��J�7�����4-a��w\*8�}�:�ť�N�1be�<k{�O�OP������$�����V�Wbf�[x/������n����#cvt�3 /1�Q{m��G�D
\�e�I8�`���_pL��p�����Y�ź�&�B�I��{�Nc���?PFzȈ�v�@��	Х�eQ�5���Y*���k�5�ߎz�I"I���4�$#X�,�NU�Z�s\a��W#p����ni'Q�A�-%C�v�G���Boo+d�o���KXP�-ll���G}��l�
�w��7abY���,�-������p��>y�;>��34�T�M�а<�Z_~�Exn�ik�)�+F(�=z���Ȝ.� ��Yj�F)��VS��g�/ڳǏդ �1�:�6\Ӄ������ח�=��MD�lTлW]��%qo�H�qЩ�7�C��R���e���p�5Yd���N����_��F�+�<U�B���簽|�E��o�.|��KGc��h	⮎;RO:>�L	O��+��;��x�3
A�P�"D(��I�X���c�8�&DRMGҋax���r9�U��T���b��h�{e����$#�� ��|�3��-Zo��ڃnµ9��}��0�3�@6��ށ��
��E($+zƛ�{��<�o  ��IDAT�(v#`�ӧ�f������CY����Ks�R�M��Ђ�����l�m��U��S���婮���s�6��Ȝ"�S��߼7��� @����������'�~��=�x�/T4u�ц�F=�<64�a�#`�v��ɽ�����FɈ,�)�<��{��H� 8dl���2�s���`;1�o������ܿ�0���i��eg��`k(v���J�<�9eƆ��-U��@Z[�OT]�M5��R#e���Щ/�K�-_�@�����ǪUǞ}%���ǌt���E�=�Ri�Fn
WJ��p�+Q���j
�Ӱ�	DS;jZㆪ�^�b�rE2�� _!�2Z7�N?	��T��r�,܎�Q.�P]��5�1K�� �ru��$5���Iʪ�*?��}��^�W��v��!��#��g��������}8����b��a�f-y�L7����^t�a�,�v��F�E�mX�`H(s��e�8���s	@��U��]AM��s���a����N-�gcw��Q��h���̸��m��z�tE��e�������+������ך�f�2��҈J��^jU4�B��"��S;4���|�g�{�-�]ޘ�=��W�!�[��b]���" 77�q�X���5���1Gy`��\�Y?J��W/^�ϗ�{q�>��|�,��a�)|��1{�ӏa����=˾�'�.!@ m��w��z��P�����`M�]��=8�<�p�T�<3����[�|g�q�5��v���:ux�m���Sӏkҡ+�T�q�n�@(�g����cը�[��o�(�(�!3��}/��bP��6,�Y:S*&�M���X$>U��`5荆�^�|�?�-���@I��^Hh�Y��2h`W�y�Ne�H�'�-[?`i�m[�AK}��Ζ=�+E����Q���کo8/][��M)��@�ೊ�YXdS�$�t�<{�@��ZV���o���[�֒uxb����WrT3��E�J�B�������ߩ_ة�DfB�B���4����q�7 �,j'�`_V������d��aW}�C��F;a�����e��/G�� U�}VM�����%;g⹚s���0_�����
�p	�8_���n����Sg��Y�c��s_�YA0��7c��0��Cm��^�4u��k�DI<7NP�.о;���?��)|��f�K�GgEG����N���7��ܱl�e�+X�86	p��I��x��k��`J|�gR}k�I�r����C 4�l�s姖�+�K�	8�Rkm�I9�%����Z��l��#�B�;]�	%�PP��ߑ�c@8��2�{*��NUv�S�
�b�n���?}:���5�mϒ]�C\�,�j&���=�۪4ҙ���,��׌Y��]��>I���6�[�r�Vo�=Uq��6ռ<�CG'�f�����%�_�����x	V�N�2:o�����ɀ�UݸvF)wF����;j!��5���;���(� �x�F������/���m3������F����*3�������1�����2_*�&k�gQ�8s�-��M�5)�Lٌ���`5!�K�D���OO��>�o���2I�aw��B���Ň����[r��f����۷za�P}�Ϟ���N��\�q'����F��ϔE����o�����5�*~�#�4�CL��y��A�5�L*�z�=�|�D� �o�D���� ��.3x�c�lrg]�c��ch�^o-���E�D�P���N6�9.,Ym6��ү�8�kd�l�(�D�(�7@&�wmc���D���û01g@agW-�k�.fk�A���sAo�c��8>�];%B�j��Ԙ\���^]]�Z@�`@""��n�-�Vk��Zyd�rcw�.�@í���-�[!Թ�
"�F��d���W����6{[}��G�j˒0� x�`$����ţ'�l�=q�w�}/o�$DrԦ]'�'׶ޢC�<��͉`�g��ak�7�9�=�5@�#��r-^����\kL�9h�W�������:�l��)����]��a����%c�`O��Z� �#�7��B�ӻJ���]߾��]\�[Jh�)�hĳćg]gWҨ
���D9ҽ���ٵ��Gf?7���
UI�|�,Ļ.�����K���i��TfΣcDJd~�XC��Ț�!Of���8���m1/_�k�e��8C�]ab@��Z�rx�o깦��,w�]G�S~����T������PW�ZF (��i�g~F�r�9���\텏���X��ɒFN�--����pY���Vp��i���,��@�d\�3^%Nк��q��V���#~�S�~����N��ƥ��[_�"9���ƞ�g6���4ʊq��s�yU� ��χ���ܰ�����J$-�ZZ�� �o9@�%\	���d*���~�����i��0�Y3�DE�������g����efn�Pg���a���f�CӦ̚�����<���䏽ai�����Xv��B{���� �<��ž%�E3C������	�=Ԃh�]\<����2�?�����R+y�,��?)#����}{������+�i�Ҧ�}��I
*8zM�36N&�e)2?��8O�������o������9	����d�,���1.���� �,���U�N���,j�E�z�ZC֝L/���(�Q��{V�����i	d� �w������+!��=W6��eޔ*{Q.��u�{��jp��k����#Rvmo��q}}kF?
�gIZ�A)��M�/� ����W"z����������"��Y���d���1�8�3��k�ﮮ���NƓ�$%��R$Hz���R�{V� ��8=ۇ�.����|��q}�����?���@���}쨺��ڞ���-{o�ڷ�"Z�C_T>w�����{ug�`?��I������.�;�.�(�ۿ�s4���J��>��d�H�wI�]D��}���b�<܀����3+u,��{l����Z���Y���y��斪�HP�	�؂@���.d/�D�S���ʇ��d�����"������b1�H���ek���s:_��ܥ�V+x������!�`�k�ݖ+�)���6���y�Mp�{Ԛ����˯�9�3�B�[q��}ć=\�S]%�Ѧ^W�Tyućh�{F�_8j��L�ĽL �R�拳Xr���> `i3��\F	安?�]ơ.�np�W�g!�pe��0��'�LrҺϪZ�~r�8�N#��+��,]���m09z���S��Jrİ�Q��$�s�~o��~vley���x�H�}WD�Mˢ���D�����Xݤ�hM�U4\$!��D������'�\��*2Y�}vyN�iA����'5��^;1���2�T��![F�]fao�c�1��ŕ�נ��R���"׹#�7\������y��C�>�[����c�J�]�k@y6$+3H3���=T5�Xl���"n�1���>�^K��>3G5�������W)��|�#w�f�w��������,*�M�l��6�<�������=��s�*��xV�U�>+M�L)�qȘ��-��v�s��(/��\ň��cc�9~�@-3�gr�zh����GSpP��ڣim�{�J�	��/T��hٖ�v�r��%�XҞN��P�0e��hE�|����2R�J�PF�����s���+��d�2]k8u�K� ՠ��tu!'�9����2����ެ�����eؤ$
�a �D��\������	���}���;ͅ����27gy�l����G�a߲TD
z�2{��A�Df{6���a�Jں����E��� h�Ar���;{>�����l��;�)��;g}��������G�]��Ϛ"����p�D�9d*-es;;�=�鵽��LB��hm/q�=r6�.͉�B/��X�g��}8���~]�������7�!�c/3�YD�&�����3������4"����ѡ�H!p�8)���I��2������S	Jb`�r�r�f�(	�OY\��"�ɬ�����+�U(FU�dm�� �Mgpn�%�A�"$/�1ֆgAK����e���o �w	�{L%�&f��ݤvV��*�'����l[r�����Չ��i�W��j= ��u�:9�����=H��2��>�^<3�Q�,���Fwij��E���Zڋy�WubQ|0�@��d�Ί,~u�\RU%�5����_�-R�ʲ��'<���iv�ʇ�A�Kt��[���jS�!�\NE@~c�NO�%��+Fð��\�|ah�f��X�p�v{r����mZĽM�����!j����[��<hi��u\�1��7:t���h������(;I>��i��aN�"�)\��15�`>ܸ�ÞS�\QT���o*��
0i�O,�8⻛�:��E��J�A�+���.}����/2�[Gz���8@:��lpy�0��s��^��hP9rX�nx(j����;�œ��o�p�]w<|���^ht��GS���ۄv��=��D�+ߕ���}91wv�&�0	A�[��Ï�������d0!Lɛ���2z��(.�~���Xn	E�^B!�2k9�ח"I�f���v�G�lJ��;�1�Dd���I��_-�����j=RG@PZ�U�۳x}�Q�=�'L���0��?m��n�?�-f�]'����3�$�8��~����W��2��m/�,�c�*@yc��=שj��@$)R�"[%#n��gYW�ۄ�hC�2{f[�Q���f�W7���q/m��@�k�۾8:ۨ�l,����
l��_EL�g�zۮ�Ft w5����x�m&/Ȋ�+�O�E��0�2C��Ι�?D�Fs��m��do�����W���'^��b��d;[y�S�^?N��#&5zq6�c�g�\��0*�[L�_��QO��pߗ>>����,`	�5� ��{��Ը�	��˿���O0O%,���j#Vj��+�둡��'"�`R#�1;���ԉM�N��y_~o���W� (?%��	I�����H}�(?�4��h�|����<VS���@��r����P.]K�g�#�*R�ӒZ���	�{�B���W>���v���l5��:�,�+�C��v��T*n�·�T����؁�N��c�p��
���|6��^F��1��aq����WB9X��e'z��p�{=��Q�2��T4�Id�7��q�|ߎ'�?)�s$}���?���f�{�WJ���p*��|Du%j��Ћ��;c9g��pbƭ���O+F�lT��HB�6b\;�A�hӲ[�(Ďtx���m'�z��gt���µe܊��ZՑ>.�C���\�f�&
���§�'�M~�� Hw&���E�@<ϥk��8v2nT��>zr_z�Mzqs.m��捸��oc����y	���wd��gq�87KKd�P^�' �����FI�Q�R��T����u�
����C��˿(S��G�o�kسg�G�dk��CT{n����d>�P������`{���k�\^2$߹���!{��>6'
��� 1Fn�m����5Ϙ��c{��6�����d�)3�#V�e̡�IS�L�d@B���c��^�2�L�f���pz.�9ա��=v]s�p��FE	2�ʜ+m����������csTm�/-���΅N�1�Ǚ�Ʃ%o�+af7�a>*آw��S}�o�F�RE`d{�xg�iL����w~bk6[�r��'"�zΜk���~�b�QAb�=��X�7����w�Yg���>�ci<U�(��b��B�x7q�@=^7�����+��ÿ������S�h��rX$縡U��<h�"��%�G9a�N,���qw:	I3"�yU���n�$[J)���@�!�U�����6�.���Ri��'�����V�GAw1I�,%T��J��JY�c%�K���˭ց��5>!V:��<�5
4���x/	Vx�S/|l�%���BK���a��V*K��-,*��7���2'�~y�`��>\I�5��-b�����g����e��ή�����'�
�K_dFU`o:z�D��<"�Xt�sfN�l��/���Y���j ^D��/q,�Y���J=(�L��vS�A�/�˗����]��GGf��Yr���)_ W6�O9|���ui��}v�������u4.�����2R�qH��u�	6�ٶ�#����P���(9��,E�I�(����ۚ�ؚ��|6��,]c'3H�l���AH��v�d�ȁ��{R���������|R0����ǆ��|��w���e�P�����&�����!`�"��*�j)!�TQ�U��c�h�_�^Je�ׯ߆���{�G�D�pO���_��gn����]���T�� %���)h��)�*�!�)-΀O!@���ii�]gt"2�	
N(��Uz?��q:UovgAX�.�-\��H�MƗ,jo/��o#e�ʁXS:Z����c�5�a)1η9a�c��$��L�%\��۔�ww$ Y����UTr���	#j=��oޅ����Gǚo��}���v|&Nxn�E���jO2M=\���� �8�������|�%�1��H���� ���=�3�-����z�E,������0��ɆHy�y��3�]kGT�G���/��G[�a@�B��#�s+�U����8&�D:1s��X�4�*����>@��ףp��0]������6�$�dG:IA�а���Ŷ��Ź��~��Aꗦ>,U9��V�׮{�1�m's�l��X�̦o��=k�8Q:o��	�l]"�{G�u~&���cŖ+��|-�?����1 HR���4ݐy���O�TD[ ���uӛ�g�>8wgӱD� �(tR^�Ҕ��s.H]�=�ħ��+��f���z�v��ob�� ��z���|%��]�0G�؀��yx6���V*�,�z}�����a4'W���	���܅זq�f���O�E�������w���BC�0�W0VI1�l��[d�0*�O§<���W�^*�x�|���G22����o0\Q��O� ��)�3͖ڐ����|���p�d�E�I��+�����^��P��x�J���mS&���,��̽?���	8x�="¯ȟ^R�,��`����}���%�ƷB,S"��f�®���L<��)�u2r� ]�(����#�����kE���m���اi|d��� @�!���p�d#\�0�u���C��Y��֒�QfP-e�0Z�v_7Z��YA�� p(Ia@)��3v��Z��m�thA%D��dm��aRc���-����N��NeW�@�ܞ��"��ߴk�2#haƁ1x�۬�T� �)1J��	4�F�0�+���9����s�XP�Ѿ���/>�<"�T�$�����c�Z@�т����V�-͹V��-�����p||�j���5�4�o�{�ioAk��JU����)e�U��	Fn�%�z ��C�,�C��L��!�R�H�0�!���4J8�:P9v�av#N9s#�� 1��lA�L}�I���D%�T�b?`�^WA�Z��y0�VM�c�.�w쁖U�D.�aW�@D	P
��{,b�r���4�G?�N2_����^
�@�lbEV��lz�q�{M�`�a�q��;8I�(u_�-	����u����2�_���ys��o��*2�i|��ɒ8{|-9�hk�)	p ��S�g��&���3�4�Zڽ������K͚�e��t�^���������mV���h��4������9�&d"��EbBvƟ�Q�.F8�户�����w�z==H�>WeWd
�OCnNU|�D{���@��20��r�wʩ'N���o��h��1��k�vɩ��|]3���L�V� 9e$�0N�|�o�1�/�l�7"�6�!	�7�^�sg�b|)2�ןޅ�(��[��lmi��*g֓ٺ�A�	����<�4)�7����O-p�_aM��,����O��O���b���k��z�s�*pN�q�,c��5x��Y8<z���^J��gO�
�va����T��ܣn=㾓�t �hwEG�zNlsCF�(=T�B�hM��v�du���F��\1eQ٥v�k��ӈ��������X�y��Č�`M�G�6�-#M��{��9A����������-�ߌU7i#��9�J�JzKw�U�[��PQ7}�[x�7������X��������:4��Js��H�}����S�0-xB7�[2,�j1�z��H�;s��JD���f��I^bq���2d(���uDE��gbh{��i8~���F��7��}89��������u�n�5�K;���BT��}��2\$���ե��Ee�!Է�}̬kњ������}���T�鳳�v��F�#G#\�ev,����K	+�pz&�oH
����MT@�+e��$�L���{�Y`Gb)s��ﻊ3Lh�����tmW��5N'�yc����v�������.4�a� v�}��~��䄖���S�UҔMKA͜63̙g��d�-�V�] A �XE1����C��O�h�9[�5�N��N����	(VĲ8�;v���զ����_�ѻ�eӧq�#�Z���X��^�z�FB�@!.�I�-��QA!X��iU%'L���hpR^�}�ڱ�y-��4��
��M�A�C@���;y���	W���x�^\kT��#�R}_�N���'S���m�_���z2�塓v�RE"�vd�L=�q>#�1��\n0��|�c�lBnn��d��X��QcO3B�!>1ci�D��ƳjT{(�}�����D"?ڰ<��g�����L��h���9��2��|6����>�"'�>��������Q%+I����Y�<"43�<%8a~a󎲶eg7��һ�gf���Q@�|��`�u�ahYwF��v8�I%Z"���Q��+��gq�ϕ}{oӳJ�W_}����޳L��؁9��Z�=��L?H��؂/��*sԥ4�#�/i1������I�E� �kVx����س�D���[�z����P��������Of���eF��"
����`����e��_~��0,�/�h�55}��cV��h~�t�R�H�ٛWEZFy5�wƌ�3F��p��{/3BEO��]>�6��(m'�߷��I#���|aʂeiᆞLd9�(0�Y�E�:����WfA�j�=�z����ty��6���p� P"��Ui̽��	n��U��	a�������	������Jͫ3G̗(`�s�;���7uC�c��y��@u/����BGv�ע�pe����6U�!ڳu� 2���qbO6Ӟ�r�!Y��g���R�E�
M�\W���X��>e�71��������l�<�1UM@1�3�(Gx%�����(b�N��y, ���c� �U����	X]��f��]}W;�8�'/�[�i�����@$m�4�(�	�b�_��B�!μ�ىҧаOFQ�[v,�`��\��;�3|>�����W0q|<7�;���u$A��>8V��({%`n�/�b���l�c���l�;T�����TD�I���%'���C3�߱}�;�, ��hB�'N��uG$b��oM����Ty+����K��/SQ��z�b�(D7N�}��aA/��txa_����)���N61���qH�At�)"�O�]z�6��� ��3���?>V�}�t��2�`�,��q�)ѳ�&Y89;-�}��T�e�T�I��=�#���e�C˔(����)/]��nA�����$�f����e������k�>YH�M�8c\lA��&DpV�F5���r�S"g���e����R��%�N;t8d֗�R�m;H���� В�KKu���0W�T�[k�c�7�b�]��dA�^ڣ62�ڎ���^����8�=��p��$�u�s�?�v��<�(�Hi*�l�f�	dw���.�Sn��^�zA�C,�����'��B D�9��՚h����.�����g�g�E��ǛI��q���:W�Js��p�"��tڵ;�5q�q� ���T�aӲC��-��N�hW<��H�EjPq�R}�����d�I�����#�[����ۧ{��xe�_Z��k�P_�����O��\���Cx#j�I��D�kYi�{'�-"�H���e�m��.�L���=U�^>{!^wph�~��p��c�j.�z� �S��N6���ke� ��],5�v����l�f��kZL8�i�|��^붉e�7X	�T�9�az��%�g��7�u
ԕ�8�߆�Yʀ��$��7��0�ߧ=CŌ��B��>_]d�1�|ȯ�����E$�q��ή]Ȁ�J/֖��M�XCZ �"������3'����a3՞!(Ej��a-	e�#U0=pF�6̆i#�)�'��H �3�ݐ=��0Δw��U���D5��C���Py  �,ͣ=�k��-k��;�ɩD����`{�k!�`Y�9�#�u�T&	@���TᔵSζD��n1�?�y��X5He�4-FB�������o��EN�6�틼�JI\��"�H;	���E!@4t��7��k����;�PyP�prS6�ť� �ې��D5oߪG�� ��=�"Hx��Ge��j}��[fz�L����6#�A�^�h؝�
�<s��oz�֌�R%�3J'v�..,�U����J8�� u������Q���
'���6-C +<�@�Bߚ��%�VQ#pnS��-{%~��I�%l?���=��޳���~.0����8�B=8�ڗ���v��"F?X�,�"0�L_WN���>��A y���e���<����2�b�S��r��D�4f�3/�(-)�BP_���u;��ּ�Yt̅��V��<��̪W�	#�����Ǫ�F�(�Y屽nv}���޶"x�T�gsd�u�@ᘐl�Чϋ�|��ɢMY����:{����t�*�1�����@m)�ˀ��U�D�- V��3Ҋ���,�[���zGu:�sJg��^j�d��G����#��Q�܂�gǇR;B���& ~|�����p�R���	�z{>��NFf�a�+Š�)�nC�`k܁���L�.�����=<��l���X�0�r�B��������Sę�B����#H]�b�v�1��7��2��G��y��E��W2��wc����y�f��8�|٨�R����Ftd`Sۥ�҄�(�+������|�8����O�䛰����H�Y�Ey�>�
cP�*b�R$ۭ�Ȅ������s�9Ӆ3��v�7��QME��S��)?�~-��|�J�q^����Y��S����#ܥ��5�f�]�-�`N΂eL�W��Ӊ&q�|,��c��m��%���=�PVk6�"�%��G�ԥ�d�hONX����$]>��h�4qaP�5�gS�N @�Nx�������s�i:E|A�,kx�A����H_?g=Tp�jw;��/rnV����5�Ԙ�&���՘z��6�n�������G�'D�d�|r��II��f�ᮜ$��!��G�*3��0�p�8D+�\������U8=9xB�;��'Ї���uZ2�.{�墅e�C��_���&����4��8�d�ݖʳ���f(Q���
�4����0(��.J�W�=�fDp�t1����,܊�v�(����I+ �3z�[�m��'�ݏ�K�L���BA��n8��g~l��p d48�2���d9`�N/n����X��\ƞ?	�v�7���E�
κ��g����]�(w,����J�^�mW������=���3����L�9? ���5D��(���f}��� �$h'm�z2˫��PZ����G��Dv���������B��v/S��+�gNl�ߚ�����O͘��jdIP��;�j!鷳q��2�jC݊Z���5R[�ke�EY�l�>�dDY�1��!2u�aL���5CslQ��Ã���Ga����٩9{�g����Yt�r~�64&4�Ϸs".b�*Ę���|�@����]�f߲�.���(�]�s��gM&��."! �
 `���!��O�{P��O��I@h�Hx#�H���?��]kK���[�f�@k�[ 8��1����u1i��t|����w�2�Q��vrr�*JV]f��ʚ�_��=U��\�åo���ھ�攣��KVD=�L�z>Q�8	Q�{�k/mZ�l6�����|��1�����٩kض��@Sۃ��ۻ��ע��*�������-�B@BɃ��3��@4$��Nt�4�Q�k��`w ��Of�?�K,~1;UI�{��":R��o֣�Ǉ���P���D䈘Ded��%3ǎ �j�Y�H9I鹎�W`+[�+UrN|�+�u�th���̾�ٳ����s9O��h�^3]�2ظN���U>.j�p(8X��.�G���g�����?9a&��g&od�q��A)y���@��c��G��D4�����3y� ��޾'��R��< Y5{��N�)-����'2�VX�0-{�����*�
ܘ�_�3�x	/��o��r^�K�YZ�>S�z��ќ5v�&D����T:q8�E�K��7��~g��2!�*h�B�R�W��GG�*�K>M �J�ȇ�>u��ٸx5� ��-:�/
Y�V����V)�k��^���,x`f��T%@�͜������o�a��e�zۮ��ّ9s��g���q����9��֞�9k��h���>��H��-��Vk���E����p2�L�O�I� 6/�Q�4~��cwe�l,}v@��L����0�X������\){��$Ș�ؠ�af�*�*R��n���C�ߞ+AϹ_g'����.t����7ڋhmH`��h{�`b�����;\��3��Ým>�0c<�hI�T%��|�B�h�2#)���&\TN��(E.��F}0�3�oS�m�ed{���vxn��сD��E8��^cFg�eZp�,�,F�1�M���l��ǘt���}�v�E-�������qdY��	�	�Ul3=v�ht��,���HWwz��,@�����a��w�H�Z�R�����,�@fd�9g��@�F�swЕ�9��ڂ��򳸫�k�Iik��0`��l� }>��i)��󫧚��`��pձ5���x�C9}��1�d:��|5�k%����G�K_ctB����f�[�I��nHڰe=h�V�\�>ھ�&)��i����3K�!�������*�~W�6.A��3����.���F2�{�+���鹒u,a5��W�s���hʘy�<J�j�]��r��]G;�pS�*�?{�J�^� D<R�R	�tܐ�^��g<�g����j�b$&�:J_�����T�MUܴ�Y+t��J2����ak��X���R	SH��Y.7��Tܜݬ0w���#�$y��\�v�q� ���:p�m��1�OϲD(�ݭ~�J8+�&��+l<I6C��$�t��O_jf�')�M%Bł�-�yb̥-^���;ٱ�sѐ���շ����UyW�K�h��n�>�hf'S��G尬��pLqίZ�p;2�E|$�c����UH�Q5<9��Y2�i����-�g�re9�7/^iij�3j3�Lc6,��R�>�d�S����Ra?�=�v~�)�z�"l�m[�x�-e��;��N-�No.]h�)��_J���&����v�<89�����(�����L�`Ѷ=C@1����v��:<y*Tǂ���"�C���&��B�giS�Z%��)
��g�N�j�C���њ/�0~�M�vm.,� @��#1��7����Z�Y�ԙ}�:-�i��qߵ�Kd!頚�$�҂��a�t�R�e����!�]��:��Tge>�\E�v�x�,h�	lcmi�1-DC�b��N�>��jl;�:)���_m�� �����,D��`x�{�o����IxytN��Z)zs}>:��>��KkKDF'����	s`���#�ޒ���`�=���2��\�u�鐩"���aT: �8�쾦K��,pn\��{�p3���R��QR�"�X�Z7zMKXd�A�vx>�=isX�^�e�u� �����P�bS�&�|]��Do�B{$������/~�!��=��)�d%�|�$���nvu'g8��f��n�1�-Kۋ������"0�d��w�S��	�<g{��gΌ�$O�)Y��9ziυ.�2�~����Q8�8S�.��i�.(�[�F3�Et�����|���f�3���.�5[��o~�����K�mI��~��pCw�BQ���߄��咊��o��޽�H��t�L���ϵ̢R�/p��z̴�Y��v��|��7��Yu���u�A�5����J��|.iL���C_ų5Im�{];%Ɂ�u#a����"(M���Wd�Rx������L�-+�#�jEU��%���y�R��U3�T���&(�U��b�E�`A�KJ{7�B��S����?�cx5y�Jl���r�(���BH�bz�V�ܙа�t����?I�U{�+�cשG���*Y5mT����ښ����c��*c��Zdv��ޱ�"��V�z��v O���j�M6��/͐�їΔ�����t*|V�s�<�"�J��=[P�i��������ݍ��PGp�!3f���4�W;@f��z*��vx��O߄޿s=�N.>�t�tOU|S�Z�n�́,��o�O+դZ��4���lA��5��R���c*Na�3�ڻ�j�Z�Q2���+�u(7�9�@�
��[� QѤ�B������7�nײt8�HK|�'�{=dKi��V��$�B�g���+%�!�M�jQ��y�ud0�'��m�+�kQș�
�#K@�,`�ߑ��GD�g���|����V����(����8�E{M eOv����3` Cp�m� ~:�jhh�ꎭGa�{�����*i�f�=+�qŒ���܈�K�9�b���e��H$W��|4]�Ʀ2��d��δe� \(�=����Pω�Ln5-���@n�j�D����P��Z�G.�9D.�\O+{o��j��՝֘�Fd`��%���a�Tk�'ڸ�¡�ȹ )�%�YXs;�.-х�ݷ��J�ΡUr<�н��$��E�P"\!�[��(F��pt�v*A��:
�����$R�<�,�� ��G���9��1YzN��/�L��*�\yi{2t��0�-DCpv[C$F�'y"ϦJX	�N�`Y�x@��z�uZ`��3�����%J^h�S!��N����.`� Rȉ�JPYh���B�}~�9a7���׃'n��b�� ������g�㌘�C�D�,��3���up�D�u���޳T�l����/��U�Y�P'���m~�B�.6�"Ze��!�g��������o��g7t�C�l��I�QvԴa߼|-2=B+�����վ^� �_��1nKRAZ�4��#y{9[ʖ��d0�&`�ԏ��D�1�+�4J0И��<u1ˬ@a��$'(�j��sߞ� ����v�fRe�1ACb���@6A������.?_� ;��\Th�Q��I���e��a&��\� \oV�Sj�iT�qA�mz�������A�W��T�vK�j�A��A�A��	5`;h���`�yx���N�F(qX��PpZ�Nsӎϔ���4L|���
�f��	����B�
-�Un�qc��;:;�	��k����v���EogkWq���Q��;Zpľr>+ë���۷*�{�l�g#y$@��|�w�<}f��k�ja�P��,Y� M8�H�  ���S��u�G�j5]�k�=&�y6�@Y�2�c�~��:{���|d�o`�e�Өcf�����Zv��%��'ak��(��P�+`f�#�k�����|;$�Yf	`�(ZrWb����_)hj[��-+'���3��琟������UHW���������u�'�fF���	gA��>Cgw�GHp>˶Z� ��{�	s�J��ԑ˛��qb�x�&
E��Pр��Sw3c�W�!2*�:F"#K�n�������^��ucg4l���6L� 	@���l���O�v��J� t�HR���t��Q<	I�ۇ��;{��C̕s�v6�:��*`O���*��N�u��:�֠+� ��>vsKN���.3{�璑�z�����M+ըp`kV�9�Y�)(�g�pq�i#LW	:%,��ܻ}K��-Pc'�\�r2=;��G�����p����4{j���H���c=�(����Nض=8���j�� �+�}^�|�={�}�k���oép.󈼖 �,ko(��=��;�q_��ES�/�ކ�$%u��:'u����_?��b��3���p<��=W��3�R-��^�ϭ�dI��?��_Y�m�
�Ge�� I��l����ɓprr$> �~�B�+r)�W�錚�L<�\�*"���MWR�rK��sH�SQ�-k�;v=���ҌvZm[�`�-Z�<%HY��1C
nV�K���d���/��Y�[�TX������k�r&R�TbR�mA�ὼ�"���`g�)ITF<�p������O4�H��A�y�:=
��^�#����Gt�\��p���<<����%�e�0�M�2�����<357��D
D�
n��-B�|A��uo����_+��`U;G��r��.Њ,J�������������	�� �<"0$@$w�"{&h
�t��,¡�
_�x�u�������q�m.���pH�bv8��R�@�`ږaԙ��*
�̍�d>-J��tY�Z(�~ߪ��*&8��~[�^8�Ϸ'�H*xP�Q��vpr�wl�m�ڀ�B�*L)-Z�.�s��Xձ��Y���*��~��65ݪ�M[�[o���0�X3׵˝��w���D޵����]�g�&aN�ˮ�vl�"���vm��U�HRI�r��2��CO����g3�\ �@����c����R*��]������,���O�P#�؋��i��4(X�<O�>���N8y�TU৳S�ک�F/J;/B� Ep��ٰ ��to]33fWFq\�9/��`|�4�JR�}��²�V.�	.k��EjZ9�,�e{a!��2
�=	�B��73]�+�21��5��`��	>�db[��v�mu� �Rus.��k�ٳ�e��/.d�އ5�cgסT�v6����I����������뿩��,C�}J`p�~���
�K��oW�K[W���z���0�k��^w�g��6�ON�y�^֒:��6�l'�M'Dݐ4*��^������jҽj�e�����H���U�Z±�� �*[�9ٔ^_�|e7�f#������������`�I�\־i؜d��
jU�~���Uq8�핫ah�am��wqۮ��©=X�}�9x0�e��i�m>�0������J��%�_Z�����o��v0���*�hep1�*���Y˃���&.|N;|i���߉z���,|����y�hJ�&;?;��C�k�M��r� ��������)�.�D�Q�)"jQ�B�\n8��f��]�k<��=�B%f��^Ӟ�I�\+-WZB\�{-���l'�d�^!y9�;U�?(:����2͡ܖ.Q��,���9�y�Tk#$��"U�Qs�P�A-�'Ǉ�7�^)4kR�%����6jA �Ё�������.�beۨ���͵��5��.W t&�}L3� �}�_�5 ؞eE��t.d.�0ޛ�d\���E.)�xI=�
�қ�`ڪ��o��s��w�$�@-Î�é���LHcR�#
��%m^$j�2&aN��b�E"l����9M�*ղ�׳�s`��J�E�/�x��F��֧�m��eAjU��>\Ye9^;n�	�,>��&�:F%G�#���Wm��t��gZ`�쫐�|T3��G�Tr��nB^ՠ��V�} ��F����["�F>��c���wVY����N1�:[�]��V�6�,D7����Ȥ��n� ���Q�F���\'����k���|fφjN]8���4���V�0K_���������L�+�����ވ\h��J�EK�q�$�(�7����N����#�c���?�	� ֤O�4!�l�Y��ٍ
[��T�B\�Տ�����V��`'`��3����|�]���p۝�Ot^�1��=��>�^��~�s��I,O���g@ߔ�3��zM��~Q0lh��#�����}ˮ�R̲�o�?�)����ZM{����͍T�lʹ@_��������H�n�u���o���s���>˴JK��t� )IB�š�Ni`�B%<Y�E�`�qUS[8�%����e���m��2����-��=ǱeB��%��!0��wgCz�R���bBk�9��NB	���a;�p˿�{e��	:����â���	�g��e���V�BmYf��8WD�/m+@4����ZY�E݀
�Vl�|�W��a��#߇2E�DB��պ��X�Z�D�[1Z&��+�2I�%��Z����2�Ϥ�q�ϒ	��&��6�$�3}>���Uv|�|�cױT�[ʠ]n5j�%�������2�t�Kˠ���6�M=��X��)��f�r_�T*I�l@����:4�0^;M^���z�KlPc�:.�m��x�t'[2:��f1�X��ծdL1I�yG�����9W�Lr�Z��BK�'
Av0oZB�0�RgZI	��'H{�,��ꬎ��e��=�c���}O-c�ݬ�����M(l����]���]�S��"�Ҷ8��0kW�
ہXfbU�*�%�����A���GH"R=ʾ�]�s;�l����0���Xj���-J�^�� H�d�@�'�I��`(��y��fV5�Tc�A3v����/���
E�����0�ɇϏ�,�~O�Q:Si�H'z`a�2���{J�~h{p��M4����Z-f)��xj�N���X�1��vVT{}��4!uŵ���v�G��v�]!����Ϙ_��ѐ�HJ�HU�d�6�źV� �[�3�=L�>���	��{�w�z��T3�/s�{���t4��u�k)�\H-x�эS@\7�ItV��:$>SU�
��Sv¶ �-[���g{N`..?+Ѧ# �e��A�I��w}�e�B��2MbG3D�/<��R�9Ͳ�:���O�D~Ư�]	7��'-�M�J����.�nڵU|5�04�kGV"�O����e>�L�Ü�!ܸ''G�hz�ٯ�z����)IfC�(���/ʥ�HY�9+	��z�U]�����V�B���\(�l�Û��¿����ɳ�.I'�w�����Y�p�)�����7m�2fRh��__�{���o�t��v����A��F�
 �
����D �R����X(�R�E�.TY1C�WtP����m�݉�p�Ro1�~IJ��
��.�,r)�P�=T �j�no�Vr��-¿2��b�X�|v�"�4���;:���{��2U�z�	�b�p��%���i�h��U���ԩa��'0D)Jb�:R֒�Or�&��Q]� �w\���kw�UK�X�0�)�pT�&����
}����+��sn&�K���q-��]Ჩ���g����в$e��5�\L(QK�@9K�����C0��D4\��D!fS���7D�O �,�ܝ�*F��[j���X�ހ;�ɪ��{��[��:\�A��{���Ī���%\v�aׂ-3��3$�T�HF�J'G�2��嶺a�pg�/�R�e� Bb���Y4:���@t�K�"��+I`0ؙу�	����Hc�>q $��@L�/)����y׸k�}$���6�c�i-6�I��Ʊ(��|�ϸ�|����GJUvn�v����w5ݪ�5܊Z��C$��Ԥ*�\��G�O��Cw�X��T|��w�I�!�e4��=��r��'m���:�tq ˲J�$&�ݮ�r�$���Aa��O�4q[C�ڍ$8O���W_Y���d���!tÙP�SL�������l�{�-�N?]���g�c@_��|x�V�Bk;�^�h�ʖ�ל}3B+я�8|��>}<M��?n��x�G#���l�Εբ5�g`���a[ϩw��,�+�9�_/��s�Ҳ��Û�+W�ܹ�<���{TB��������'G{a���M/���i�4�+�A��B�{
0"���eIT���͟��\���E�P⒝�^�%�s�R���*������uOL\k�*�í�x�@ �(d�����\����/�B-t��b���n�9-��ӕ&���K�pD'�R�)�&:�@���i'�d�g�o~�k�<�j͊�"�@��"9hY�+5ӈ�ڟ���Z�qa��sv�Ҍ�D�Z�DN��,���,FZ��O�t@�w�ނK�`�77W���:,�<wr��9/>�Pܖ2P-`Dd����ծ���������KP	���W%y�4+�@�-T����2��l�T�M��h��3J�6���FN�C����L*1�9�>���+Y�*�_3y��)3����m��Y5���\��D�h��7R�JK�Y7	f��Ү�+mM��h�-Y�ߊ��^��Z�tX���dR~�z�}�����;{ngP>�A7��uiIO:	�5(���k���X���ڲ�y��ŠM;�
��Q���V�"���gn��s,���:��Z��D`I�Z�
>�!�|  �N��̡�;���_������?C�Q2L�&�.1�slTIz�����b-�6,
��U.���FҪ�%*c���V�@�p;�&���/:JT�7w#u�&h�[0�6߻�M;� PC�iT�d�h��>�`�svt@��ψ�1
�om�;�X{G��*<{mL��qC�὘�f�FP���Z�k��@�A��,�g��J�_���P(�*��y��߷s��2}���U@�ىz�ͬ���<�+�F�p��s���3]�or:pT��_2�!�Z�~f�Z��fI�Q�T����V��ʎ�	�g���F��T�4��q\����zP̈́Y��EɂW�F�Is!:��#���n=�dZP+��������Ӆ~����pa#��\ }��Ү*M�2N rF�ޗ�/��~�
��qS�*d�J��۩�d��fɴ~o��͋��ѓ0�)e[>�<0h��S/�Ga�U�{�;NXeݱ�����2�c�9����̖����eJA�	��2� �R�j)���U��~@�xY؝V���Ơ�|I|�hZ/^	#�Њϣ� �Y�p�oF��� ��OE7x?�u�.?[0����v/�PD��ZA�q�ʥH��3JrOl���4؁�؄��oe��Xղ�ӡR��Q�ǌ�%<��q���CEϪ�7h9j��1P�~M\�����(� ����T� U(Jkt_ �(�Ϻ��3�B���L�(�+����`���v��IH���P��4z���
�&s�xݨ�U�f�q碌��E��+&�H R]r���k���ځ] Y)��4\���ե�ѳ5�ϩ��Nͯ�����`Uh���8���Ԫ�"&"��ŵ�OՂ�6���X(*����|��z)f#�N��m����{r��Cow[.Jl�uE��Ee�똤��;�����m_��J4���sYD����!��$5h�#��rz�\���3;���D���:����7v�#{���$�����,�s��U�5mp�%��ۚ��~_b�H�5^wt�$
kW�#��-�@vO��f�w*����e��o�c�9Z�e^;�@V�Y^�q˞���X�$��k�c"��r6S����ý�ؒ8����ؤq8���e�$]i��&)�=b	l���	�x�a�d�S�]fq�Hf�Ɗ��������;(���3�ռh��v���dÌ�#O��~T!��	֍?���ˣ&yZe�_H��=-�b���P�m�.���Ȇlok�~�ۿQ%�	�������͑t���%&	�����n��o0�([X��J���	���|fE���#�Ptd������]��pG@��	�s�`�{��F%-eg�fa�r1
34��-��E��5Tf^d�H���^X�v���[Y�t[.�A�E������b`�U'� �Q�S����a�8X�i��ZVЉ��M�&�/�_��Q��)W�%u����}��/j��j�����Yx�x.��7wd�5����Wz�.8���V�h5(혊N��ع�Ӊx�M^E�t0���,*�r�)����y2�r(�Y����M�?���&�q�
?s��r�1��4Q�WT��[�� �k�j'�i�M><�U�k\'z� 	1��-�l5���k/�NB�=����K�Jm�9(���8��g�뇳խ 6����
v A�B��n�4��p �l_Z�v�<�P`��v��--�k�[p�[�9�.Z�h�T��,q�Y��ͽr�G�v�����.t��f.L�+���Ba�~�m��( ��ݳD]x�6��8�!�����Ց�z���������(���ݝ����<�����g�l3U�E�N��*kq�[ҭ�m�o�%��h,]�/��R�QZ ��`��p�S=�m��.���w�S��m��#ǝ��\��Y���I�dw���fwg7�X ��.�~t��p=��� �x`�!�m�.*�&��"˾�����4��s)�V���JgF�!�G#98�D��?�d��l[�$&�����m�N������l��8F-�;�"����� �M{ V먡Ѝ�H�F����
�T8`9KF:Y���5�~��4�����s$ɼ;�s�|!䒆����"� -<G��{�����\ER֏.����c��)3]Y����VORm��Ƃ�|���zM(�|6H��V{�Q����ě�������=q��r���p����8�	Uxz�l�����"���;�l�� ����8�f�ɑC6�?��.|�(�G8@����^wv�nض�{�u�����'Yձ���J�tt?��x��;Ӊ��2ix��yc{.hǽ<�Z�Z '!��aLe��w�Hc�T_̿�S���63���\#$e%��!��שF��QHms//�, �v �<�d9s�<y:W�vz@c���v�2�Z�lPF�B�	�i8^�7� ��K���#� fg�Ӊx��E����=���mL6�R׶r��nOA�d�k��t� /��ݍ�&�v\�U;�P�<mh��Yn� ���Ul �d��X����o��W~��3���~*2�6�%��>"`�T��+�$p��Ė�_�{N �]|�։� :.HK:��$�=���H�䑴��l�$�0 0�O*���~�8[���yD�O�| Z�0[�D��5����h����?�c:��=� �U��U���W����Q�1*�d�.� T�e<3�q�jvW�t�$�<����ݽ�b�bt�&��E��P��Yy+�� ^��$�=	-[t��1�[�ugk���s�?�5:�}6I��kd��QV�_n:T:��/$���3&�+�u��E��Q��#1G ��m�Ҧf}��.�=ܩz����h��?R����0�}P�vtOd"A۸\�z^&-G�3걯{�7_}��Ei��e��0kE�F"�eߛƾ!{� ���:�ڽ�O�%ؖ nn%Jұ}O�EiK�=]�2���2x��%�{n�9���<��>�J ɱw - [�%0\�d�($s�nAi�?�5�7Y�$1H��ȭ���]Z�h������72솿����	�y�={���q���w��- �@ ��Bd���HJ0d�F����)E���{OᚲX�-< Ӧ& �(��(��H��l��V���_O)i�QJY�W����3̭����_��͛p����ٺ��
��X$��iю���Wj׬w��k���a8����%�:�ZF�/5��C0_�B~���ւ�fvR�F����>if��)/c�Ʉ���^"ص�Dϼ��KI��Փ����������
�H���;���E>���m��q�a�
?���(вۘ� ��ɛw1U�H.#�S���t�+}��bk���g��3U���%^�H7:��BtW� �/T\k[sX9�u!��o��o¯��a�n�pS+K�j�IëՁ"I�m�`
��T�y�I��taz�j�A)��9e���	/��e�[o,:��HoH3��"��
���8��QjQ'{��w<��k��K�s�2Q���C��BO�QQ�h��������Sun����  ���H��ɡ��S�-��P�p�˕���3�[�����:�=��
nc��.$R�k�g][�p�z�{��O����Q��>D����$I#:=�z+�k�1� �.��C��L�V�O.�V;��a�3P��L���7��$ni�_-Ƿ� �����Z{ z�̆9(6dC7 �?�Z�$���̤u3��޴�zҕ�>&Y?�8��1v�[��:�w��{)�U��-�B.S�R��,����DzI�+u]��^z'�5��lB��+�݀�tD�./��M��]��oFu���2��
<�P���F��>�D��$�6��y������p��'V�$�hX7nl|n�XWH��.��/H+/��	�}�%��7�F�C������j�ˍ&t�n䎿DE�k3/&������XR�?^L���"�9������7\Mڐ���jv�*���������$*���<3���T���r P흜H��iV(g�I-U*�?��&Ӆ`�۱��id�}m������즚��_# Ӂ'�Tcpn�=�������b)���}�'��������$<�9�����ܓ��?^ڡ���"���>ugs�j��������Vao-cA���d�l�`V�gcv� B�r�O�eI�R�݁�ʫdC�w�����B!�LCmLة:��q���iGц����F-�+�= M7zr~��VS�U��E�|,��4qj�Z��#�jЬ�6�x�"���֏\�F�5��R&���\m8i��Zvx�����wk�'Y>���Й���}���5c��c��2lF�w�i��vv�?���K�����ۈ�	$����
ĦUqp�q�:�<��%o�7�]��to{���GZG�� G�hfν.�'���ԓ�v��n��:޶ 2mw�cg��x՚9ZU�N5�f�[���R&����m�0����A�σ��"�.�|�M�t���S@p���[CKF�����H�X�P�"@2���  @e�E��}^��c�N��q�}�<������i�͜.������g���XF�S�)X'v��R����е��-۷�8�~v��v�*r0'�:1�z����m\�V�Y���g�a�ˍ&��1{���@Փ󁳸�9~��ݐ�Q%M��S��Vf���o�lr�X;w�[K轛UiĆ�B�;�vt�b�u&ҧ�G�G��4Di���:�N�v�v{�з�-�0Ѻ�Ol?]�H�R<f�o0��w���c>�����8���C8��vk禨RY�erOi���k4�Q[�(�x�#C�~�ٙp7���}��<b�� z*.�-��\wm-��&'¨x2sG{��9p�?�OK��N�_~��J�V����p�guc��\��@�����L���Y���_i�thA	� ��ZB�k��CHΙ��xza7�n�rV}m���,�8-�_}������]�T��h�����AS�\\^�?����_���pwu�Co��5�& 5�8��Ç���7����n(�����M(Kͱ{�*��ZB2���Q���߄��'��w-�TvP��� - �ɤ���#K"�'y�����������������o��+A�*h�� � N�� ����u��ҭ��r**���&�����j��,���t[��Z�� 'Jk��8�2b�PON��7�E�pc�� u���: Xs܄��w�5;S�jj�
A�%������*4z�Y�i�D�}�R��X ]�J��#thI���\B@=�}�����ݭ=;�ÛɁ(�=!)��GG����\�Q��s�+ſ���L�=�,ZoC�*���+�|��\��/�F/�K�?3_H��p�1OU��'��4�*�&��Ƈv@�(f͑m����?8�[�s$�TK������XI)3�F���j]yDy��7�^�g#K |~^F�f��ݠ�ݩL�-ͬ����]5�Ċ���9�|k��D����栴���7�'�a��Ӱ��$�,a�`D�	g[T�O+W�kp!�;�Y+��EN��|&����Ju8�t>���c˘��N��?��bh�R�r���ħ��\��K)߭�61m�)}�� ף��k�o�3T���"@���7�W��1#v��kfommӖ�
%i\LJ����?�^�[�F�J�� ��� �#�8�`�w�62�>#��R�����V�3���D�DnF��	�}�����4|����yd���5������fT,��R���J�{v7����7��sh�PRa�{;��]��Ϟ*U1H6�x��L��>�I}��F����:�k�E�)ی�����Z�>[k�r���tߟGQ�W󥂈���H�j�lc����W��=۽���ѹ6�Z���|��h�0���B"�����.pu+��g/����oÿ���ݨ��Q7�p(Y�w���Ls�O��=�m�S�D�%��g'����E���L>�'O�Ë�t��r4�<�Gޢ��Yf�1[5}��m��p���4���Ѻ�_�H��������'����m�c%�J߮���}��w�M6�jڬd�d�t��1oYq��Ix~�4���]Q^��m|9�� LR���n<��o����Lq������ح����w��ZG������gw��d�������	���F�D�S��<!�F�%��t�Sr<��E���j�S+��;���F:=�/W�;��'��֒���1)4�H��IKZ�;���˵z�eej���a(���QEI��[���b����hE g�25�pt܃������p�G�Β����ٳJ���!��}r��WE=�k�����|Zj^�C5!H$��¤$��I��R|'KS�J�
UK�2����ZPI�Ö
8�f8���R.�V�X�'Q��]-ML(;��][Ç{�w�Ϟ( �-�U@���޺'�r�5G�
4m8㾞X#���)M�3�������{�M�U��Fr�����_i�S�Rz��k�Q���nFk�a���9Tڳ���皟�n@�����|�$u�6�SzaC�O�̺��+��J�O�hO�uGG�s�X�0 ����eQ%���c��M�FY~^0��3�"��|G�b��Ii�X�㜓W�YX��S��m��TN_�]�3?P��s0�t�X�̈:�A�>p��@��S�2��;�Ԩ݁'���JgUd���|�"�?"���u}����������֏�y�[���:��$��\2�?�,s��-+a�0ȿ�|��jv>��۶�	a{ڞ�$Y�\]��t��n��kjײ�ON4���	"�h?[d�:�|L��,U�Wu�B7F� 15GD�*����V%_k�7��U�x(j�܊vBe�Hڛ�ji�p*�m7�V-�.~}7�v�?L��=`�FU�h��!��B�s'ٶ���{�֚[���=��~��߄�����e	K��+*M����婪Ƿ�3v� d�����o���C5#�_�K{�,��YВ.���9����Xﭲ�]XE�<��\K�����\d�9v�ȯ+�9����И���jS��ti�A��>O�6Yn5	>[S/��}��]Ue�ϮUѳ�X7�G��`-(��������h!�� ��e�܆�K��(��0��-��=o�)r�t;��r�����Bԋ�s.Ւf��Z���\���m@�d��|j|�bz^V�
���U/sgw7��Y@��˻�|�*|�mU=��>V{>^��A���D!�{ۃ�i�t�����+U����*ߥ�T��W����s;�Z�;!�å�
���>���eߞ��>ײ��M(����L��Ē���V����A�[%�o�p��7{"�����j����Ҁ5,=Y !s��J[-�,�Z��^���_�������<J�֏szZ��G��|/�Zt��[�ݯ4}�l	��� ��6��y����Y@1C��\M���_��fe����LZ�X !24��I���e:��|!S N��N۴�z����f�$�lYm���:D�N��SW����"CYFi̲~��7:̲�����tB�V�=�U��VU�Do_�>�yE���7��4�ȢkEL��F?Of���c[���_Rm�i\��%���([�(~7J�`�DQQ�Y�Z�2�p�Elm�����!e�!9�P��!��N���ت_w��])��o[�I��v��<P���r�*��M�^���e��+Ѫ����U]+�.Ve�{���"q?RK�V�h�۹X{���+k|�����$�u�dIx���Y��j����܂�]w��C���aw+�8\�[��F��P���q%&Z��[[��T�U��c���5[�̃��D����+����}8{�ђ�;u��2<����|3K���k(KMK�<]���v�$(qFS2����F�����>˷������Nv���K���ʒ�����e,��~��&܀�S!�� ��	{6NEYWխ'���<*.�5M+�.Q���giv=�l%e5Z��0Y����و�Q�P����^F�@�r��.���u����A@�����X��V�%G��%�����fO|F�՚x�k���i���hm�Q_<Υբ&���R���p���G_9�[_X�ٮ�i��Pӟl���o�
�R{�2_��mک���u�qkI�U�=�l&0�q�]Mҷ�QŊ�t��Qj���z�g������k[K��'���Z�>� �}|��lo��-U���/8�����-�-v �Z�>��ܪ��A��q�@&%-O��^����,��+)N�����{x�8��V�z�lk�(	4T~�	���(&l�� K��<��ε��D��C�K�(]��[�Y�lf���U�.��{	�a�����^S���l��"U��[U��@j����πv���\�&;CKbe8Q9�E����Ԏ'<vR}?���To��S�Y�޳ts�K-L�L�E�y��2�����!G�!����C���X�ؕx��״ޅ�o�:+I��u����K]�ʿ$�ׂ%�Y��LΒV����m���G%�Pi��)�x��,����C(�5��J��U�̼������!|<��jT� \f��Љ.7�Ў`�Y)H�*-m�
�	%Ȕ�@�r|/t��ý6���tzV��-����}�#9=�8�B5i9�PC��n+\M�ʮ������ý}���!�l�.NHv��wmQ�xa��U�ĥ^��I;�f�U,���G;a���i_~�:�g'��
��`��Ֆ�τ�;��H��>�*
���A��K���a����u�R8*d#�Q5�]���*K��`����'�O�ʞ,Z�KqGqUW2�s���-�VO�B�.l�l��5����x���Or���(��AG�S?"בD`V�fm[�Qƨ�BhV�V�	���A�jcQ���m^+9 ,��`*�r�b����F`Nc�&�I�C<]��}�s�:�v�&���R�⁸�槢�b�O׆ �|):I��P����'	�	����
iSƓ<Cl+$f��a(�fJ�4VYH�b��,��w-�� ���C���e;�^gaj�;�%�@����÷;�|:s���ي& }w�����V�v��C�-*�"�i'{2נ�^��&Q�4Z�!˃�vEO�묿!����+o����%[�$���Z֏�Q<��K(�Dj�h�ps6�'	=m�>ɭf��S�b{�`�(�1[���ʞ�Q�R>ʼ������n�u�k�<���
� ���� Q���YVў�}F D=�fF9�բ� ��Љ���ֶ����C�xw�MW֢`P!~��t$�Vӹ�	Ŗ�śynQǪw]D%�J�q@��F�3{/�% +��N�FYͦ{AqՊIUy���?��;���u�Ȟ� ����(QϞ,��|�"-��|��J��ȱ�괨�_���6M*nFc�L�Gi1U>j]�U��� �m�G�U���ݏo���Z���vφJ����K�.�)�̒�����f%r@�(�*|���~�1|�|��s�3�|�1<X�t��t3���HEzs��0�\�t������]=X�9�1"�W�@&�C�f:<�؝٫��q��Z���3­0���g�������o4���DHy���j����\��Pm���B>h)ؼ~�Jg-��I�,:���g�%�\��z�箕U"d�N����QG.�LK�@i��J.���C�k�RJu,t�he➳��7���Ҍ/��e�[�ݗ�"ӲC��T�R��#�${�QZ*=��b�nt^l��>��KZJR�՗,%c�|a�,	Ӊ��;[
|�.�~�����Y����`��.�Z��	�����YqV���j��6I�8\$������>]���c�XߋAߞ�4̸�Á��q��A�ծ%�:�@w���{��6�'B���$�^��(A��뿾��|��<���#��=%�t�=I��x��յ����+K��,�r7��"�N��Ҟ��1�>���N�^"�D�]�hY���-D9,Pp�g[ �i�N�� lw�m�o�ilb�)�/x̥`�i�~V�
��3�%j�>6Z�����2��Qǣ�ƍڼȄ�1�홆�}?���N���{����lHK7ᬛΧ
r�R	L���^�����r��G �s�)KhAtuV�L�ّXt&�~��\ ���]���;4�sB����{9/���ndL�.B+]�D�\j��u��#�"bN-�Tj�=�Y�����J\�u���$���^���9-Ü����7�j�̔�áaF0�v�J&!T�2�� ��tU*b@����ZG�,27�|����Y�	�y�M�F���q�1�괤;�yص�gɽ�K5-O��+E��z�A�0a�H����qB�d1(ɒ�/���?Ἢ�����I��2���d�j�k֐�0�rQ��~��f2�J�|��,hm7��"7-�>�k�+�7� ���-��>���ޝ��|\O4v��P+ui@M#��S!u,T�:��8L�mI�1oy�vT�èt���A�k���C��:�%������X���F&���rD%�;	H����X
8�F0��H	����	��[<�-�$6�m��KkoԪ$���J�d	�$(	}��OWN�hf3+���m]S��3��f�2�r����{��g���2�]}�rR���Ԁ��xD������`�z�����Ru� \����OIMN�Lݔ����G5l6�<�����|��k�������{Q8A ��|�k�/-k^��6�4*�,�vi#���륨u��O���Ŗs���4P7�t��ء�@܂�9
���JWL�4���R��"'�)A�k�ǖ|����б�Gi�ii����~��6��`!�A����N�͉-c:�o^�����vs����(�5�;�n��6v���@(3���=`Fo�Յ�	�����$30�بJ[R�c<���n
� ��"��cq�c	6��QH��(m�7
̂��TK���u"�5����-R��5b�C��8LI՚�e�z WW��z�����k�IQ�h��m2\� M�XP�B��	��,�?�J�쑆c����y���ߘm�Jų���V9֎��@M���e{�뱡�?A!��3�E�~�
�R[<sF .[P��l�ڭ4�Ё�3�3�6�Z�[;����(p7[�?\5��#_;�T/���y���+s�>��?Z�&��.�Z���A���T���E�H�Ҩv��#�e�V�	�P��u�1$�Z���؀.�d����Xi3K�Tz�%��vt��ȉ��YvsKe�.
�0$���ʕ�ߪZ��d�r5��N�G[��w�R�`b��Ր�M۴3K�&����$P�r�_���Z-��y��:�Y����#>�V)�T�}eY��6J_Rf��̻�Rv_�ʂ3!{0h�0�Θ��N~�Âp��ŕn��MI���B#��P�t�U	EX� @�H23�yS��������Ud��\T�c�Yg'�=�>[F���m$`��VAfe�O3x~��cg���! ��
8��A&N}lP��k���1;��D�m���h"ǹU�]��Z����U��j�(��PC�S��jCO'���������=�w�VUu��o|v��(b�"~��g��U1�3�5���ϼd��^s�`�@m�������!ɵ.�@�?�����ۡ�E�����击"RxȲ1B��JQ�Q�0q*�t�����ߌ,�]U7�^?l�wMm�^Z%L�|�j��DG�N(��h�ڳ<x�4�|�wl-!�Rwyҁm���`??o��ص����⾷�s?Oõ}�k�k��V(��p��	���PG�<��Pe�۞u����B�\c�L���uL�u�	�$/�Β"�-Yd�*��P�k��(H�y���H�w�_���>~�"�_rD3?|i����
���*h�.�{�O�	�
U0����-��'�O��o^���H{�3�@3��j�'�����d�e�ӏ��}���];�%4���1�@�%V����ϟ?w^;�ί/���a�Y���=�ܲ3��i�����(�%��Q�̙��;��J�3�ɯ�,�?	���֙��"ޠ����jL��
W-�/�L��7�<� �62�?�b���F���A�>c���5��5�-{dlx1�׫��o����4bI�z�݃p�=�6n�ygQ��4bn��_?��[^	���ɍ�Z��x�A+p�̥U�T�dl�>��o��^L�^�U����߳O�a�
�e[�������@�x�*]枫�C�$S7x\op��T�djH��ձ��<%�JYT�cܸ�8�^�~!��$�|V�V�=��C��@�v-�~��qqpo ��G�n�Q����c�|���*����m�XKDdB�g�wt7
�H��[�d�I�?}��D�CZa���p�<R ��V+�>t�<�Es�ҫ�E X�$>�H)g
z��JHh+ƕ=~��TPgn�8�B�B�Ƭ���"Z�e�)���B�Y+��k �e�M"��"=d�P���k[/i��ء��ׯ�o�|ƣ�pwy��$� AZ���;��ߘ�_^\���;�R�O+�JK�ɫY��d3jQ��J%�,�\M�/�z��,�u����Á���7SeVfs��T!��}Ι�I�+X��ǃ(s�����Q�l.m���]���B�d�}n,�����9z�c�J�����.��a�#�f������$���BY+HA�*��4\��=Y���1v�v��0�vaͨe׭Be!*����_n=���Dr�]]�J��Z�i��]'��3��7����;�y� ?�R�P������[վ��"�l�����������Ƿo��ŹӺ�$[Ec���^����L�f�ؽ���|��ˮU��(�߶��b-��3t;�(,�ptx��Y"���������E�2��x����X�	��ϟ�g/���?q��\��,H���
��LP����F���4j=�gK�- ��h:߅��=%5�4Ղ��up̂Č�:T��(�p�5��Fg&��oۃ���k�Ŧ���K]n�?>J웳D���S�8���FS~��,E�w%�E� �����;�t�0cɣ5aH\}/
��&9��u0��}9�jOJ=�B<�,��P���R��4K����N�!6�h|��l^�ߪ5��ٓ�w�;}���PK���[]e�+;��P�"ia�>+w��+l�,���}r*bZ>��D�;���qcьmY�'����i��Le�� ��M����@�yG�AB�:Ȧo� �
��5��"�b���%T#��KI��D&�*t�����6/���Z���&������ai�`/��0�zYE#ri
��FK�u�"^�
(#�6UYD�.���2��W�6� ~y}�C�������:����Z:��=��� G���;���	�PI��}IY��TG�j/�*��RU���%m�Y�J@�`�l)���K>�m�<����������)V����r��u�tCW�������F�>�	��\�,x�!X�R�v/���~�'Y�]^�
�z���^��i�����]�|�I
C �� ��%@�\�����S&4�l��dA��/e+�:�4fj���$?Y�=��=[�w�v�?����@-SU���G�U�m�q'��epr:��2�X���J:R�Ҟ_�C>��Y��HŧŶ��a�-�O�5��=ה���̒�Ҿ��M�T��n���Iˑ�6\�R��UȰ��]H�CSIU�x�V���>���)VU�թk��4O\�U!V�p�m�Ҋ�����þ]�WO����S��� ��7��t�Aا�����»%`���f�Ŝ�9L�<	j�}�m����Hջ�uu�8�ɫ�\�>��={�O�+�#��:ؗ��Lj���V��'���_��_�T�
�C�YU��%DU������O��r�
�A��]�N3/�ku������z�V���HO,~�fM6I��w��r/�2*�=���4f��C����$���7A��o�>T%��]7��&� \GFH3�8�@|�iR��ݫiQ��KY�N�(��]�����Z�M'%]�R���{��i��FߓlK6u������{�f����󒝝�p��E�����^����~�] ��[y�vUQ%(�H�0�G��jj��ř{R&�.��{�¯�0?�%�Z�ˈ �#|NhF�� ���0�L���F������(F+���,`�
�Ӫ�6��<���9��y��b����M�<|ba��aߪyt֥�B<�&�<�3�1SD�������(��E�f�M�:�^=}��n�Gq���W��f�J�a��cB�D�- �b��B�����p-æB�d�V����hgف���3*,Z����9`kK��W��kq$�?=������R���Ύ֟�㑱��h�!�e����Ax��e���_Kp�.h�F��k�t;� ��L"��3Sk��:^}�}D�p���*�;[��}�hl����ɤ�Q8RYs2S[���<�ϼ=����h��V?��b*[��z6�J��Z��&����S���%K����H������QD�a�(�XBw����+�[�gV��u\2��JL���RK@B�﵀CP�ʉU2v��/�&���l~�J��h.��M����B�JD[���:J��k�3u\��J4s(�v�P��k;�T�|�-YC��`��}�'Z�������JƵ�]��=~���%�N[������������n�]�h>�$��%a��! Ȍq����ӧ���_���}�oh�$:��Τ'�+�!�*`��ϟ?��?|'Q�@�> �D��"r���"���G��w�Yb� �������[r�.2B"�+v-����_�3V��COy�}�i8P��D��_{���]y�f�yb ؛]��������-�C+�aBӊ�r�ETDk�d~�M�F��[?����
?����vY=&Hގ��zD��Ts�5�8���	�ZNi.�Bkzf�w�P-jT����W(k�.�k-�������k�ח��ga��K�嗕��g��A�c��J��1��v���p�Ï?(��û�0�*�2h�j��*��A�ǌ�I<��z�������NO/$��!�.|���ܥV#�fz��� F��;���'���t��ζ"變�l�Y7�o��C���0��CE'��X�d�9
7�� �d�U����o$�`0�@.l��j��e���ԥ��#Y�1^Zu|{/z
Vi�GG����pp�/�13$�1�Ev�.#p,�y���3��W�D{�{�&tum�!c�Ks������ˆG����1F�2�Cw�t��G��[����v5�:�xx0�;!�"Z�d��k.O��**UӅ�^��㳟ݵ
�����T�s t�D��b�E%�X o��F��OG7�>K$�0�
F���A��A'�T�A7b���D��ڛ%cT��^_���K��@�6U�x�($v��\� zhWnϧ�x��h��4�B&޲�0��5��a!�a�Ug��Vi���v����'���]���'��]����~O���,
Kۀ`↧�-�}�[�s0	X�K:�v�� ��Be�;����a��pϱ��:G��@�����ӧI�*>��T����$�UҔ��=����}�|wc	�HV��U�� �$:1Ӌ��NY�;�@?}�.ܾ;յ%��Ǜ��Q����l��]���E�������������_�:/�/¥%�nz�R���F�
��`g�量
ƬK��+�͢��Z�ȼڽ����o��J�t�Q����΁�"?=f��]x��4���*,���s���Dv�[�@{>v^�z��Z��.�Jw %��h5	7�u�*]�����~��U��5�"�Ơ�(���$c[?Γ�o���Z�X8�U�Bu���3�8��'-im����c.܏<Q�0�B�G0�񖺅�p�,�Ì	�eC�jb�ƿ���­ZZ1U���i��թ�ĮJo�+� �(�}�+��[��{���2=�_��w2 �eV'8�"T�)E�B�����B�E���
	�����>3R�c�.��#�ڑ���zT{i���	�DU�������y����doW6hg�w}g{�UT�x��J��.2�I�Hɑ�v]��C(,�8� 5�bq��.�@�߀�A�{O� �N��|���I8><����v�P�l�q�cj���A��#K��(>���3�q�����3K��Rm\�a��u�. '�*A���ж��V]ׂ��{4��q����i���a���W�r��MD�j�?[�-H9PO��NO<R�3eLD��N��������p���ݶg�Zb 1p��V���y߾O`�(��ª�{[��v��C�%r�%p3O"hˉ�.��Z"��Z�q)�m<o�����XC����@��V�M^�]�s�<��8�I� ���� �T��4��Ձ����6G�ߏ�@?�`�~�p�W�piA����y+<�zr`�Ӫ���в ��y��e�I��%Ѫ`�1��=���<������lW���ّ��n�tw/����Y�+E-h:ܛ~�6��3^�n� [��B�^Jn�tE'&*eL2P��������9!0(�)\G
��3},��o�ُ?���$���G�Q�1m��#�����8:��г����c����#��z#%?�0��uh7����E�1�:�3K�y/��.�"wv��g�4�+�����|����	�$�--]����25`��??���>>����A�ŧ��D�L���`1h�>�ĭ���z��zu��L]�F��y����"F�we�x���w��;3:ծAW�r���o����V��EU]\7�GQ'M�1��@2��9��r�iL*��"��N����;r�"����6 �����s
�v�Ө��
I���N���W��y~������j-��d����Zw�!�n���fM(9;,|[|{=TF��Εy��﫽���\*�-�T��-�X�"��x)�P��XQiv���r��ǌQ��<���di�Dhc�EQb?7���H�Ti�H;7q}�R�)�8�.�J�O3tm��1���*]�9U�}6�����me=����YY�q��ٳ�\XKһ
;{{���H	�d�~x�}x��dSfM���mc�Q�!��)|MHPTe�����,�p�j&t�U�y��ӧ:im>�ymf�fa�#�1�%��h�w�N,젴����Ϭ�������N�l�����6/����	�"�
�F�i���&��6�4�bVЭla�>�{��a]:��9���u��89���w�n�Z���Ѻ�ܳ�1����J
�Wͳ4���Y�һ���'Yl��0�Aaj��f,D[qm����������D,���K�� ��l�$+��j�Q� d���c����ϥU�s�J(Bm˥���:�ۺ<��7W7����*[��%'t���K�NÐ`��n��ګR6��^:�Z�+�����c�M��Z��К��=��nHW�ʂ0^�IZ� �Ś���G-k�T���K,�����!\��������z[�2y��v���6R�	�O����> Tunm� �hYF1��n�u���7t�琧��إ}l����U��bl�9$�v�����p}�������������b�m�um/�^~V�3�=�["�A��4|������i8����ü�ϾՓ�P�������d.��"Õ��o��$�xo�^�/uFE��JR��^&?�@j�v�U��Ei��p�ߗ�����rb���y�%�)I�p�`�ަ���cE.�Ő���� ���u�]HΓ� w��]
)�|�V�nFJv$@��<Q�un�v�TG~� \�դ�S��3	P���N;� ��g����²��Pse��!xx�vʯV�g.��؆e��"EzΛ6.\��S�x��BPe�j�C�Е��R�A!I~��I��:j����@���=���h8f�����(s�o�tH>��ʝDԧ3>�j����c�z�Z��}tJacw�!�Z ��J\����u����~?W��=nmuT!ɣ��E-���Q��*���N�V��K��r7@�ARW�`~73�2uII��<��|�����G/^��ݝЅ/i���e�U#̞��O�]�	��*FIJ���W� �ܑ���*W!jÅdё�cމ:��?�Ujbj��_�0�)�$��l~_�Tx�R��!c���$MbL�@�B/�D4:B0��J�|N�T@f�P+��+����y��_a����:�����0Bu�H�TEXr��n�������*�d_H���p*��JkV�U�?�_S��x��M����9�I\��<��{*���PX��K^��U.l¡ɾ���m�9�
������U;:�-��h�^��B��Cb�@Y:71Qe_�3]�TIWQ�ΰ�u+�GPyJ�,RS���C��pkh2�wlC��B�x(K�A#�R�5=�3t�^nՎ���hq��{�%�0�C&���~i�:�[��z��@"�~Gi�}l�2�y�uX̑�q���m�H~�Q��~��ʖ$��E)�sn	:tK���/�(/��?�>ZR!�j.���[����CK���E�~}{���ӟ�~|�>�s;���a��cNړ�1����`t� [(�(dUѯ�A�r���oΙ:�-em�H�=�7������S+i�P�C�d%u�c����M��ԡj��$Y٨7f���q���]�
��hH"?�����-������U�M�:y�w�[���F\���2�9��W����Y+9gf�X�"�#�a�o�˫�����qU����?��ْٙ���=�)��P��&y�O����z=�E�<��L�9fj��n����yΘ�����G��NѬ�� P����{����jp�������´�*,
AJ�;�H�E������k3RÈ*�95R�������j_V�Q�Ӌ>��^ p����Z�D΋>dTL"�I*	�3�*RӹȀQ�!�$�d�'�_�vU�Bd�yԒ-�aL3���![h͝�hp� @rR���]����Y*�d�P\��x��0zE���H�u=��q�@��C�FU�j��+�}��L@�n�tA��O�D�������N�3
usw�-J�`0+yd/!�?�	�d�$h�up�J�v:�xxK�e泊:zT�f�(+I:��!��������@�>�����"���X�RsNT��-�l�)��s拷�4&2-p:�.d���Z��2�2�g�P���Z��c3Ҽ�4"�S�w����5`��;ڴ=T	]�g"b�G�}���2$k�bi�7Q�V��x(�C`A�Dw�� ��}����
@�]<�{.��U�����f�N'�pck��!�ّnr�7���̥2I[^�85r}'�N�}�1����	����v���
��j 8�6g�v
����po��}Z���ҍj�����'���3iZ�y�,�ph��\�����t���Px���c��-��Թ�,  �I���"�x���,�V����7F
�ɢ��v��LH�z�jϦ#�#�T&(��"X���'�_,s9׾٧����.��Y�rgvͻ�wtv�de��^���m����
�����U��Q����%�ro�On�&PR�?�E/��uE(����2��{v�U��IG����LY�]u_Y�#�=�2�	�5{��ԞI��e���jTƱ7��f,��Y�)�6lt�%�ԏ�pk�ny*�)Y�]�q<1D�CU��ڮ�;���!�����焛fEtt)��Z�G������7a2�8�:Gvg�"�mC.3ȣ�&N���zgs��*���ĉ�_|��VW���CT����H)8H��� Z��ֈs���"���Y�`�\��T���c��!`O��K�q���蘬XΣ�hP\<��Eą#&B��G6���J��,{*��K�M�n��c7�5q	�"��Z����hI�Q*R�f��N��ƈ�k����QXf8��A����#��fS=rL%i�jN|&��e=�Hv�2*cS�����'���?ܔ�����"9F�����!��蝉O�D�Γ���}�6E��"�{���[G�A�|��%�7�^��.���/����2d&}n (�Ygh��`qf�{) ��ȼ�b�X�
�'T������Qz�K\�1�X�Έ�D�ckS��*���:A�����V���1N5^"�bq{��`�V��ݪX�Ǽ/�A���0!Yc��-�4�i�v-3{N������7�ښ%a�ӗjSi ����>�\?�G�o W�n�^p�챽�D�(�͗��^.|L�����e�8��;�L�I�2�2�J�v� �5��{xtwy.�?����d�D��M�R5d��E�^���eO[���[ˢ[�����e���Rޅ#]YUZ��{jB�:8�	pp��S���p�l��L?ڹ���C�>��%*�l5�F����)���"�2U9:�o�aTcj��������~�S���G�!��K��r&����O�jj�4�>t�g[�����������[��=�]�	PE�F��\W��j��J>s�e�s�hĚ4*��/V�_���;80TϠ.c�~rZ=g�e�`k�~*-�ռe�f�[;��sjVHG9���.d��e���e����cx2L[;�h5�9�W�J3���R�Y�*:���oćy��_?�j�%ʊֳ\��ۡY��~�Fs{@��2�}f-eX�Ј� ��*}�:j��jBO�Q���;NE��HʱZ�����ʵv�����������ə�B��c�D����4Z9 PV�٦��R�\V�M��rX��R/��
e��k�2i��$�w��'g~{k�^[:ܔ�U�	A�(��Κ��q@�K���+��U�����*�#��ĭ��NG��9�~:���Y��g�3�Z����h�`V2#�xh���6��,֣�na�V��cd߹��5(1��-]G�R����>,|��J�����^�GC����x�[#1�tk��o�����ǰ�w�> �y(���ɡRP�rc�4g+ĵ���}��"l��#������"��9q�n�*P�	�'r𑰀��gG�p`izH*H����B.�~ �DJ� ��Ssg���h��J�N�M|꩞�K_k���s�dm�n���-���҈�y$s��z`ی:#Z�Ϟ?�W�q��e���������}lk��R�4����e�渚T��$wΑl%D��$�5��o|�>�|:���*V��\��!@%ȅ��D`=Y���mX=M�<k��0_m�]�/��'�����*V�8k۠yoh E�P��׶ F�q�����Ѩ}hDTF���-�O����v�p.c�!U�����d�?�ۻ;�p�������nh��6���am]������m�IOә=��0̝uO���l�t�7h�ý�ph���ˆ�]��G2ޭ���a)��l�+Dy9���g���qƻ���z�y�%:�8.��m�.?��g��A5��"f��Q�k����j��#�խ��7�,���|�����("�z쪓����t�vA��]\����lS;�+�x�v	DG ���.3i��&���CGwV�������SlLZ��<�Xt�A�W��(=-� ��_/��xrE�Y�T54>��Fh����D�R�ꗫ���W�s,#�@�pD��&e�
Ǩ�x\g�4�"�XE�'�XӬE�o��*�.�U�ቦ�6l��s�̧�3��ABWw��/��/�7����-h�*�{Tm��jR�3c9�F�Y��ة$1�e��V�	�ں�/���
,�vc�K`��K�-Ts�|6c1�2���g��!����=$fsq��*������+mdq���;-��%���P�hX�k{�^�k�ӝ��*���RС�%9�b(�Ѓ7CE俷{�d�A)3^�,��Ob	y���}��͝Ʃv�	�lvn�cwQ��, 8֠�y�"�ϑ]㈅�s@�����]�^����}��0j=���ê� J�0�-��� Qކn�ג�-�)�����1�2����خ����~�oB�s �'�<�=�S����wS�s�v_MF�sL+l�vm�3�/�V��/zk�k���'\��� ̶l��4'��4!��G*?�D�C��J���~m���@/O>���SD�i��QvO�}KB�_�4�9��+��́�ˮ[��tq��L�5Q0K�*�]�4i�ɨL�L��g������5�*��p��"(�gZ�Xf�=���L�4�'�i��y�Ã��}�ph�@������a��ǻ�?
�L�r�� ���8h��|�	����LA����U>c{/���~�,(�l��ߧ��&�EYYE�a��3J�c)'�WZx�۟�#��	;�g#E��|� :]�-'z	`H��h�$K��8�,�m6<����v~������4b^�(�y�)�y����j�c�7�����B%h�w-"�5͈IT�{�UI͗AXv����˄;���h��"
��Te�0���4�Xy9PE�V!��(j��W�)fy�f��*�E6!�y�ڦ�T�b�7�Ϣ���Iֽ?5����4��Aeom2[x�v!>�5� E2S��x�Sh��,S�hP%���B��*j�اH&�������*p 2�E�wy�N��|>����׿��sKe��f�3�#D� QQ����A�O��pg�β9��<��^hE�gK���xB�/�g�DY�?��Pw,b7ð	ےH*X�BC��P�悹����=��`�2l4h� q�J4CB)M�J�i�#���E��"��E6-��bo�{��,tp�������q��9J�k�J�+20��m�9;���FXX �����H���a"�/߯�8�^z�Y<�����.��;�1%@[��]��M�B��¢�s��	���?M�($�.BIY0͝�#f�A�}�2��X���7�������/d�	@�)`OZF��Đ,$pz���y\�0���1���0���X0��j{�v��2f���3���a{���a80���; ���bb�R)�4��me2�S���
�N4~�
�&�ex)5"Ҷ�]	K1{���sc�14�b���'L�<\T�9*W��:0�X۵�[ӏ�� �K��&<�ii8��D �!D���3�s��\�O-��}X���e֋�+!p�QP� ����'SU�(y�'�Z�|��������cנ�	>�6"(��*h��_{;�"יY�r�x
f��n帜���899q�x�\b�r��	������^��>'��J`D���;ܢ&Y" O#n���_��Q�<_WS�	�f�h��kL��$���H���Z��ՅȆ&j^�j�vwf?�0��h{�@/u��RS9���&i��L��Ns�UYo�&֬��w�ݢ�j�-+-=�c_��.̘Me0 �OʘJ�;[1�e��������yN�`�-sG��zq��6���8)���,q���2�F��/��k �`��|���T��a�!K�������H=�`����-�'%�*��?@�-�a"�/]��:Q��gHA�6A�ڽ3o��<*
�����=����~c��]"�4���Y����"�J=wƯ'3F�?<i'�8T�m�Z���;6�
����Y[0�)m3�d]�~:B#�E��K�v]]{%T+��]> �J��g�rǘ�R-���/c�@Q���\!G���vGcY��Z�fB9l���9���(� �Pr�:z���Q <�Yp�Zl�Ä? � �m�:E���$�kWѨR�^���mM�B�q?[��Ȱ���4'�Z)0@+�U{92��`D�����k�%���x���HA;
��ӧ*�,�l��T��h�9c�@�T��� āx�@�ư�%%y�ˌ*�ջ�;�}�;[0?�°3���ۗ���gtk��N����� ���O�vl����T��2�j�W���q|��|�vOm�|��
�j �l�ޜ���߿�漘�
���ԕ��$[[�>�4�{'����ߘ��sг���Pd�kf�]"�tJS2vQ���W�x��t	BXKz��.To?G0�c붽��`���of�9��W���@t�fK���Ӊ�x~Tͤ�]Ub;9?��/���ȡ8�ϊ��b34(AK�����EhMQC_
P4%��naY{�E����+zQb���O��"3���mP� F4sUX:���u�K>>+k�Sᙱ�F�i����8�y��0-��J���V _���G[�tđ%�Wa�"b\g88�@?��٦l"��a��ѳ�Y������]�~����=��WAk�ԩ�8�6���Ls-[O٤���4�����n�o"��Y��0�v��N�]6�VƳ�c�S�>������FG�k�Z4����ߋ�R�|]ZvV�B���uxx���=��ˮ&I�;����u�9��@�H�jA{�ۖE��ڞ��P�4�1�(��?��]٦Aƍ^Y�
4o�-�����6:�'=M��@�1f����z�Q��\W���U���ξ�:��O���e89�6�ԫU�g��pn�$Q�9g3�Q}wN�1l�vD���t���#�o��
�Lw����+&r�5w{>#��(��Ԗ�Q�BC���ENR��e�M��k�ɤ��jߟ�#�1ë9��񆔗$�$k����3�$�ڻ�dڌd%�q��d[E�**�Tr�m�}�}[%���1'1^��p�(�T�
#��e��8&6�K��dQ1�yN63�2b �	n�Z�*+�B��b�G�����ҳ��.ʥ,�3�eDf�	�x����ί���� �Z��u0��TC�C�礱=��6��k& �:;HgcG�o�q%3�v�(�n�GR����We���k�&Wg�bb������!�=�zas���)���L���	3{�����dLd<��?W@rwz��}
�gW��|���]�	�5�H	��&���1Oae�ײ�6�ad�i#s��v7�R,h́�d�5(��5=h�"%�4�[>(к}�����b�yyl��Wط�~P_�=���+?��4\S:��O�L��^��
�a��lM;ɶ�����8����p��{0&[=���p�1���;�BT�ٞ�b;!��Y�&�f陃DyB������hd[b8�}H�J-��k�S݅J��`�q|p޼<{���dR��l��H�2�K�����xd��x_e��Ӫ�m3�#���ZY��8.J�RE@-UŚcZ��HU�
oP���H�\�E ����x۶�djk��i����H`���fAa
�挥���F�I���6�#���rU��&�,K�F�71pc�����ݏo5�Z.ܐ�Z����.z�"9Ə��c|��Lc/���%��g&z��I&�D�:5��po��_����$cM�3�h��I�;ْ�+W�J�<�2ѳ;��Yq0�d�d9
7@��x��ut��XF��YY7���C�����ʚ�u�~���2�Z�N)����"���9�g##u.�R}�Q�BG�A���T�^��# +�5�����ZDA�(�F��h��!=(�Ke ���/��=uD�H�^2<��i��5=�{^��ep�e�kkc�^S��NsQ���R��=�O����Ϭ�j�3�eI%g*�M�J�)���s��0��~�����?��E��ر���C�m�vvv°�u����˩�$F���O���ť��e��Kg�j5;r$����xd���y�Y�F��c�\��o���x�{s� {n�/Uڄ�ϥ؞uEʈߎ}J��^PV���]�[�"|���3�D���YЃ��i9�b�y0�z'28�����<<A��C�"8`gZt��x����k߂ ���a��Z���B�A?�.���?���R���"�i9L��9~���c�;��\ƈhYd�<1��?獩5��Q�tf/p�#{��x�0��y�A�\X�nd�Ӽ�(nKo�$�8Ώ�HNnn�c��X����.����>L���<X�S@�[�.�c��SK6f�^��L*x0�!�B��A/[��fا�70LO�/VKi���C�"m�+(�'ס���Xm*D"���%J�mm[�r,��F����]Ά����G�W_��v����qN�*]=C_W��e�AL
#�\}��)GS�Rm�\��3	g�g�+9,D�f�Is��MB������-3ޗ�-\���Qh�����"��e� ���4�t@Y�rz�-6�Z�<�s�U�T���N�����B�:�P�5�׽"6)e��%=p���+��wEWY���H`)��r7��D
!���G=p`-s�6��Z>��	3pXt�0V�Z���U9\��	�!妅�A����� �j2���g�`{�8�V�ψF�\Eۑ@�C^|&=������"^5:xj���d�璋�<��Z�#M쀏��G��xD3��'	I6�5��!�G��󀩈��=K�O�֦��D,�����K[�,� +�D0��Ec�	
2m[�'���1�|�&v/�׿�&~y�ÞZH���^!܈k凨R�֫V>�PD'����DQ=@(��m������Pҧ�빹:o�K�:��"�vҶ��/{C�}��ٓV+hH�3��r�<#̻w�¹e���Jn��������9�˿����p)��T�#�:	v�P��Eb�:�]7�ω��4i��<D"�  �N�����ێ�y�D�C��C.4��D�˖dЊ2�k���m�``�)(��]`�*E�RHz:78Ƃ�gm��*���f�g�ƨ~��H��^�u���<��nP=J Z ��)�2J�s&��]ߜ��ӏ��y�R`�cv��L�c/o���w��ɀ��Mv�e����cG:��I��W]D�,Wa��##$�:��2�S�aX�����T~�$k��!�psy�>��ҏ�}�����k%/���k�s��6J4�v��S;����R��H��a���ӕð��3i�T��i�
F��Ո$7I�/�������x���*Uk Z��v�}Wz��`s~����?}�_«��N�i��������U�$���j�1��(���H.\,xk��,���������i�\��̌؍���J�n؉tx�������'m �� ���Y�]^p���Ch݀_��E��g>� �k�D�9K�J�N*J�g˅����~nD0;r7�SC"H��z����l"��u��
9^�2`�_�g�[�7^-�ؔ@�Ρ�,�<���2���4}DMM�Q`��,�xFR���,A1��
�ک�F��x�����r��
� �G�-��5{��t�]�>Gq+zn5�nq?��3�= �6�.E�@����߇�˟�����PX�E��4s�8Q2,"*��y��0D|�f�l�׆X�-�>_Y3RA�R� �Pj��ْ3>�@���GeP;{��`�E8x��F]K����9s�����a�q�bC*D�WJ�pb�j��z	� >{L�#�1J=E3�J�x�����,�S&#�>�n�̌w @�qJ�2wސ���*�5���/D"��"�(���dq8I�zϕ�^����ӳ6=K���o�2���-Vk ΄@~�/����J����#�"s勬l�h
}T{���˼ pa�����v�Z���t�B�lWJ���f�"�h��<�X����w$�C�|�tq�����Evn �-�:�p_�,%U��;7�l��\3�ː�s_��d�30"ֵu������>\߅�|/,;����C��7�o[�-�x�3a��- ��9z(F	�X�A��`��E�Z��IC�!-2�>*�0�h�V�lp���|f�Y.�4�)k'���'���kQQPM��K�TWro1���4�g���3)p�(%J6��k�'����]���,����9�)�r���U_A��YX�pq]�� ���_Gk���D}v�g���T�̄M�헿�8<{۟8@�D_V�wJt�Z������f7�����3ǥ���3ЕNk�*�8�W�d���Y�O����:5����aQF�g�Þ3�����=��:�'���v��3O0���H����<��K�7	)�g����3p�hj$a�n���se�h�z*W�,"fޯ}])Џ���.��zoƑ�"������t�m����sl�B�I�t['z,��(ۂ�+
G�3�1�~�V9
2�E�f�aP6�Q���/����ChX6c�Y�9��ǒJ�0�RB^:2��C�|2'0qr����F�2���e���w�ӧO곡B��W��4�,�j%Ks0�Q,��@�k��#H��4�ϡ��� ���b�_�2|��������@�*�;�#3�@�1�4#R��9ꅍ~'�ۍ0�b|왷��}~S� x�Wr>QD��������'�*܉P�����*�J��CtBI��OX2x�����-��J�U����^_X`���8 }���h�lBt��~�`xpÓ=a䫺g�3h:�D��S�7�O�O�_�9Ֆ��"��|>�g�[����T!������>�5�C�Α=3�ˎ�s�m_��� ��3��X:;������T�e���ՅO3];�N޻��2��(P�{���i�x)��(4]���e�N����{A��ٜjF?�!v����V�o�����9�9�j�q0���$;eVW�|��'�s�����eoX�O5~�ĽM(�=��ʯG\DҘ�� �>cH���wF�4fH"ј�Q����x_���b�JL��YD�c'7�m'~�4��	���g�xXΈ�\#9�L@�c+*Id	����askG���i��1c�udNX���0��%��R�P��٨d��82Z9#\���R!�z��v���^o6A�O���,\[����������}y,�'Q��Y�b$l�52��++���b�����g�U5����JX�n��z��@�[����T �r�&���k4:�C"sB��R�c��+U!�
��J��u)�R\��Ahv����?'��/L�V��1��?�F�f�a#K��-�������a�^���Ww�"	����O��
.T�^��R�R�֮-Z���^%����4�K��r���T_AJ=s��#6��Kb�3�O�%�:2�1
D�4�e޿K�j�Py�&�A��0��C�r�Z����<�>��G�^JkuT���r`�����z��8|��7aW������p��D�O)�ޤ���a˂|�,p?lY&|h�igW�i>����Z����'}��Y蒍�kl��̲,�!<�#iB��DJ.�:ʌS����> �9X)�o�=nkB6��q���&AT͈zJ��L\������I�fU��mѻKP�_��&����$p#%_Z����˰�1
��������������>��iT`|� y��ۍ(6T�=Ҍ#M/�u�'Oj��z����:`��Y��6\�b1�S ʽ�h��g��-�ɖ-�2u�e&�:��" �@��U��Z U�z~_�y�b[mW9���J�]��MHj�ѵ����83co��"�����^2�VtU��8�=:�?���;9����ޔ��>
X�>�NB�r�96H8��L�dv��	�A�����]��R��i��G��o�� ��X"�8���=]?�}_��������I���XP[�T��Z��k�>�3�!Pn9-(�c�/u�V��kUz��Ȉ	�CUTA"��F.Үg`�6���Hס3j������W�]zy5��2uX\qo볼�|�^�������P~���L���k����fn���Q����!ցXmK?_���kg9���p�{�*Խx��w�qM���!E�k]�N���P����$˕���4�/�%ؤ���J؅�=�S-i ��s��MM����v`�l�M:;�W�l�Ҳ���7}�,'<X�Y�inQ��2��*�0Uk�"X|p�=44yHd�D�d[��um!�ٯ,b����KI�	�M����&2����P�A�zZ���{'~b�N*t5��E�b/͖+���Z�j��,��kh�4�I����c=������xu���+k�W}��ō���)���65�N�u`׿��ڦ�Â�IHbs�fh��_���/��0�2z��)�-Ol�r��u~��6����ɇpws�1���=]{?
��#\,\� '��_��:�I^��Ӟ>���=۞9�'t����Y�/8�����"q=�̧�$#��gM%BH�<���CP��MUV�sWo��>�K�˞����U�\���j����D��x޷�Z�:
��0�ۚ���i&N��_]˨4Ĥ��vzy��(SS�\h�p�AEE��>�䒕��a2Ot$˘qy��~������7��kl�o����آA����zŌ=4\l^s�R�I-���N���� ��N�Oy2��g�}2<��h~őn�J��lF��Zw�rA�l��H�H�2
�Q����'kP��]����2'�Et�+U�R�VsۗWW���������ك�9��ZAg�BX3���Ps�K��i;����*d$�T���P�O�5�׶;?T��n�eP\-��Y�ph;[E�_�4���K��?��?i?��q�~��:Ro�I|p�³_0*W���֬�5U�J���y�W΁�F�]�����_' ͬ�Ԫ�6�^T�#*U�	~�BV��^{����	L���(�$&0��֠�:���iW1�M���F�Q�f�W?��*��{�v}&�W+�������?\K��?��J�y�
��Y��	V겳־��R���+�����໌Lrd��:G������ �Ͱ��n82��r�������b]�Z{6���8��&�����tZ�/��#����amG�%��!���p3���{uu!������T~��qj��F��E����Y��\�O��R�V�l�Y�!\-ܸ��2�a�ʣ��b,U��{1;��2F��g��ș>B�x��b�$�sr��aѷ�^�馈:i+l"8�iJ&����ێ��h#X�{`Yߛ/���^��;��Ks�7���'Zoл��{�8��6��@Y�ut�����QT�/_�"���&���_�@��Ȯ&v@w�i7Tz9��-ϰ��lK���#ef��I �<�^��JGWe���o�����u�JS��v����A�9�U�:J�cs'?�N%#Y�0�z��m=�N�!m�F�*�l/���Qx��u����J�Q�s2#�:�q�������(I�����z^zFzH����V3�%q[�ttv�x�M�J��_�{ ��٨g �J��S�Ԝ�t�������p�8A�����,�jv�XA�1� C$���DO&a
��q:H�NH]�����e�8&���ΞEy��zΊ�uyp ��{~��!��*U��)Μ����R��'�C�����L�EŲ8�F�'/�tا�s'Q�;��g�ߍ3��:���(O��?��?�f�ɚ$��E+�1� Ҍ���ʹ���ޤK�ܴO@DT	(ٷ�v��Y��FE�ŽՎ��1_�$��\�p��i�f'��y��M���5�ă�G#4?��d
 R�g�Ҍ�,{D����|�r��2s�c��ũD����no�@���m[;�N����SH�R�\s�L	��������������n�XLqd��	Hٯ����3U��Ib�@����c�;�^j-��|a,[פ)\�9���V�w��s�g���`�P߂4�
�㔼�_�,p���C�%,IA��O��or����r�^�����v�%Ѝ�,E�:��Y!�g�i5͕�b��������d��m�<��Ϟ����$�>|�(R���yÉ!\�;U-~fbzJl�njb3<��)Rk�⑭�S x(������Hr,£O�r]�<�U�D��3F��u,�FT5YiSs��xdx���$#���[�B�U��(;/�"��,��ʉl����-���3�2��Xd΋zp���*	�$S
y�=ܐa��\�М��Ʀ��D������~��������?�	c�^(� ��û�|#Y���s{{Kkh�)z��g�@| �6�=O��t�*�e;D/Y�ud���īqXA'����DN5��D�d0Mt��1^j���pO���`E������=�X�E)�|��W�섫����ݮ�ї�٤����������m[&�H$.��P6^��.�|�H���
P����/����k%�8�
��w�w�ʯE����[*�	��9�v� �Y���i�4�&D�\�� r�mS��r�K���$I������ΔP���1�����z�3W9ѝ���H>~6f�D��"d�*ն�2�:#8{J�������í��Z@!y�*�#)����X�\�A0�--slGo�k�S��g�d9��cFY�#�� �겱�k�|>�B[B�C���~��z��k�4�����@�9#e�h��mͿ��h!
���y��hbD?S8���v���T֕j쫧�Xy��+T�x�p�p$SU���6 �_PƉ=z�hŞGfAu�9��N3r?��i[=������m6����vU�A�|nv� `��0��C��#�([s�ɹ~�m�x�-�������0��+���O
v����۔طFJ��,��^��������i���x��;��9�����w�(��bw�����q��mP��͛�����T3��Ml��}rqs���;t�N˜My�-YIZ���U��-����)}u��v����I4�r�psuI��H�߷H-�MoF�Y9JM�`���c;���b�)筄:��[�2��Yİ������~l���9��őʄI+nRP�sWu
��g��$ν�qIW1��"��¼�+ku�~y��u��PIS��!�-�?�F�qh�S�M���z�[)C��ޘ��[t~�p�,x�;��]|<�߿�l�A�{��0�-R���:����9��)����=/���,�����tB�l��AƄQ�N�+����!�/�YPb�X[[��H�}��`��8}����ж��2R(���Yќ�/��Xz��x����X�Si��?�`ri��Pℚ望�h,����
7S�lN͈�,�j*�i��s/'�I< �N�<�P��H��$(;���>�^%�W�v�|-dl�Մ&����C��y��)7��]+���ɅӮ6��!_��b"f0N�P	�C���z�֘��5ok��j�B�| �L����.��0�̸H��M��mt�׳��7����,�pR'��L��7�(=��=Yʀq�tX�*��jJ��Z��X��:��iC$�3;N08<���bI[I�@����c[����gbn+=z��~��g��,�J����r��p����h�Z�AAE���g^��E@TN�u�r9ha)	�����9� �W$��`��"��-����PvK�6��\��P܎�H��\Z Op���,�\�w�� ���A�AשX#�lH_Z��T�l���NU�T���_H'��%����N3��HPiYz))�,�z-��:=7G��y�	���R���T����U�:��:(%�����`�6� ]�s��-$�%	Z9<�Э��������m��w6� �: ��p�zt̞���ݡJyd�������kؘ�&��J�U��f��N�I�������e]���uzR1/�l��u��o�zo�v6v��!Yب�L�ҫ�c��fRY�K�����b�*��Bk�h��L���-C�W�ʈ{��[=�[����y|B�M��pA�2��j���`e��x4���g�O��D��|T�I�@D�s�!�`��z[��m�nf��*��L�!�d:��������p`���`#��?��������ʨ�㩮�22s�d��A�l�����Bxs�>��Q� PF�b�A񧳉�Kkݛ��'ο��1��'PY�nt�3[�v� id�c����ޛ���\oZ��Ybױ2#1�y/8 A}de�p��9?�.�5���Y���d mf� K-�O��^���=8�'avo�Č��,L�'E�{���p���Jj(h��$��pr�)+s�����:��-�jV������n��|n�nm����Z��8@��!�b2�Q2M���w���Z h�(��;!�Q�"+h�1��C�41#<��>-�Hӹ�\�Y$��=ht 4eu����y�"�DQ�m���.6����R�ك�!��lf��`<�w�׆�����Ƶ�R�l)�	�Q�%4@@S:�K����=3���z4<#wX���Oo0�dk�X��w��sT��#p�3n��Dc-�e�`���/Te
�kd0sٟ����W��ʂ[�� �tQư�|��t�/+G�#H=��	�}�4�=G~��XP����۹��m����Yx�ڑ	��9��6��B�2�jK�豾}U�4A`���ɇ���^�a��e��d'����:#{�����j:sF��g�$���}���5VF���]�#-�D�tw+� �1W�~����_UW�0M;r�� �1C>�>j~�
��=���-��=�:*�SUH+��M��^:Rh?��%��%�V"�^5[��n6ZSۨy��Tۇ9(�>��L���F����q�XdL���9�f˙�0�z���J�_+fd�XnW��f:���@L�������a���<|~���p��{Epp w{Ͱ	U�8�y��1�f0��ߒ��w4rR;ID"Ǎ�T�T��EcD�axaQ%���ˣC��@�T%����E���ܣ9�;;܋ʉ�)[���H7ʝQ�gSp�&�T��p��k���>ybß}�R�,�Yq�5X�?/�΅�ꫯ��|��mx�L�@�׿��p���CG�^�x:֡����i'��?�2T��mQ6�{�����{��3��/���J�l<�M���?�g=H�� � �2�`H�x����r�W)�U��R��s�k�*E'�>�}8�.s�S[��b5�{>�����pj��c����|c�؅2��R�Y�>���^;���TW�>�A�zVeG��#�֌3۬/�BPD�$?D�s��"	y�x�����,��f��ϨW7��cPUK�B��䚉�].��S�ǽ���|����&c��X��O��LÜ9k�k07ʙZi$p������@3cF���,E��PK��q������B�|�5{���wtp^ �g��Ǹ �Џ�H�������ٔ9k=��p����6}ܦ)
�U���
g�碡�jgZk���:�f]y?��L����� TI��1H6诣����ρ3��3�����p����PU���O�*ӹ�Z�L*)��i1��Q��O������k�ᛳ�hVh�5mg"���G�JC�$'K�2�\�}Q�R-�}C+��fe��l({�q.�7d ���W��!x"sN�gnn*86i��sz����.��Ȕ�53�y$��ͯ~�j�\�uo�g�`� 1�]p�c�a/�q:��s��U�__�59�1A4��	I{� �1��B��%zPvJ�������س�͆�2�4mZF��?'̗�����xAY.azdf�p���
!�x��U���a�6�؁Tn��䳢!�೭��ճ3_���J��7��5ʯf�aa޼x:K[����� _�a��;�?Y�x��鈮�bc���F`0��S�%T�-T?u��1���{_��-���C�Ć�P�,r}�(D1���b��{o;�-2�)��S�S�Qa+e��P��R/K�Ll`4�zmSO��@	��o��z�7�Q�t%�Nֻ��+p�;��	��~�Oç�s��8��bP�9#�������砪E���&ڦ��1t)�[;�g�o1��襡 q	�,8Pm���zY��N��R%r�	�g�x�2Ld.>�T��AT��Se�K��W�E��вg�7cз5Û�s��[�c��$��Y�T��s��7�'��C*
Rx�ɠ@���F�)K@�ON�td��U�<�@��Јt�b��}� �����}BP��a��Lld�y���%�,��h�DJ>�p[y����5Ƃta�ֈ�c#
j �U��,f���У����5:�G<"
�ҿeG���)4��\h:��"�ɏ2KI�����z�Ke��<AQ��T��ަ�#yO���JU>��;��9�Ab��f�����l�uC�5#��� �O���dnY4��
[���MPەzt��zr���o߽��Z��T��zW>M�F��$��38x���F0h�z��Y�?�Q�Ԟ��O°���m�zq�^H�z��Eț�E�sN��5eӨ��0K��$���3RJ�$x_����s�L�[A��k�r�T�'y�۵���a��sM��&<�|a{}lA���M��);Ki��X�"<�܊۝�;�!_u���$Ī&���} ����eܶ5��\��N;iE���t5��x6V������l����_�MAz�aN�QEv:f/�m\U�*$�x��!m��ې-ř�'�HAbsv��2��Q�k�:�2���>Nx�X��8�H#}f�R�Z9B�7�'A��R�M�H�R,W:�_h�v�+��Y5U�b.PĒ_N��C�l���qx��R��O��)é�R���Ce��D��i2�m�tT��}19#�<�i��<n����{$�D���a�i	�E"h�)��p�?��}�c�Ȝ����.=(�E�c[��J�w#��^8��Kg�b� ��{����0���MX�;�{"��ڌm��ʁF��5٘�n�}���բ?���;Gw���޼�^=���1i�#�2��e�����X��g��҆LJe�M[	�@j�?�LB����#o��@�8�� t��L�;�ga��������G�3�ޱ=�����~C@�xF�P ���
Q W%?~�ޥ/�r_���g��>�����qJ���Z�p��D�h��O�����i�\�����<.��kx������7�Y�g"/�rX J��!Y�
1rg%�7#�}|ݍa�����k��Qq�7�C�Bũ̵jY�e�2�Щ�T�!�W�*8��l��C��!ґ�eA�Q�����q�Hf���-��':d�TU�LR%̈�pF��ȃk���3fCk���[�*!_G)��b�*<�(ml��v*�8�5Ug��RZBX��f�;�7Wᇷo������"�tk�:�`�@׈u��%�,�`�`�1�;�5�7k9]�����H�׶Q;��4����Was�ᝈ^V�������+�K�0����y��#A��pp6c(h<iSz�g�p�C�}p����l�����e`��J�����p
�݂�4�$T/h�\�&�m�	x綷!U��$���UC9'c͡?�һ�i\�./5��*�NU(q����z���(I2�d�xf��h�J�`$8K���ͭ����5���
d��[�Ȇ0S0�v ��ػs?��n�}ֈm4�L��E3�7|�l'l"�C�Գn^2{��)BEF�C$�o�¼;h#S9��N��Ă\�EM�bf7q����������9h)������jn�Ms������[e��[���o~l���`N��N�!����ц]�^(WЄ���͙ ��q��m�h�A��4�m7Т�n���F��3ޑYv������[i��?�����>�O(Ȧ�PU$&(c�C�3�B^*��YֵR���<4ˆf�PSs���kgC2�se%Y���A3��oa�bӐ�,}a�A��2z��7�on�`΢f2����F��:���c�(7����P�[/�Cw{ԂR"'+�h����H9%f<��L[�h��vp%>�=��}%L�@I,/u�(u���ͨ��-����B�]ˌ̰\߅���L����a��jL��^���B��<2��WB�yFI�8U� %�D��$�ўZ>��%�A���1(���,JW��'�g&��穌Yl]�Nb_��u7V�?����p&p_wBd�@|1ˏcR�_���a��v�D��D�2g�XW�R�R��s��@�7�{�Ou�0(���ѹz� �����:���0��ޚ�H,](�	���?�_��$h�H����룰��4�E�G~8�ic�L)����1PJ#��h)O��0����zr�V�A����e�_���F�w
0p��1i'��?54�z��z�̎�6Z�/���R���1�`Ks�C�*2��aOgˉ�c�\<����O���j[۹F"16�9ћmwa9�윘=������p���K��!��,$s;��Mi5�~���w�lk���!��������"�ˈ&E\��z&IKs�"�1[�$��k���R=��W�)�˄�=�.���I`L��A��hؾ�����~���?�P&fÀdi�p,>2G��6���=�ۑ\��6��u4�b�'�\��TF��jm B}����.@)�� ���� ��r��t{l��I�\];�Z3�A�}ЂU9�� dAB<�d��U��0�y7g���\%>�u[�CQ�����t�2��O�T+��S���2�Zv���K3��rmk��p���PyDZ�/.����X�"�� ��e�����r� �\�qi-d�5�C����Si��
������W�	��_��p�k�}���?�������z2����~��*��������Q�����Z�b��F�Ʈkck�����>�9�)�����c��d���� �rUK�u�{k)�$F���(��d4�J��vOdsP�!.A�4��)X�szM!ʠ�K���(G���=A����Ĩ��E�q�l��s|�$J�\$ݰ=42o���HN4�Y�B�Q�LHk唚� �<��U��\�T�"I���~(�5#=j%�7�p�Rsrg+����^�lz��ֆN&�
`�1:�d���G*}.#��(��U�"�2�����V��'3д@�s^�/�G��`A�g�<E}D�l��:�YiQ3�L�z�|�jBP/:�Q�R�!� �; ��^4�,s]e�b)[�~.���Iy��pĠ���w%���j1'����o���`����n����Ok�����������N�9=ֶ��=+��]��%���1�a��$ T<>�M`hl2���VN���Wֿ��pP��X(�no�÷-�
�M` 4��d'	�V�
F=�pi�:�)=*3&�Ng"�����+@�)̿����2s�~x���9
������7_j�_�\�?���j��-p�|V��S�ڟ�fG`)���n?�Z�P��Ǡ���O"�ȧ�N����}����4�k�m������\=g��Ԝ>�i��=A�
YY��s���G8��$��"���h��+�c}����:�\H>�ҕ��J�5�d#ɋ�O&�U)2�UgS��4ET��`���	Q��<���/��|̝9]n�H'��et�:���e7��P�m��/5Ξ��0����f�Ȫ�OOaǲ��08c+7��Ӊ�}.'f*gsg�*�z��!A��}g6
��V@KҔ�0�>LA��8r�1T�p3}��%���oZ�{>Ov��f��._yV糘�z��=g���cK�VtG�Ɨ�ᴏ��Gm��r.Vv�l�7���/�٩
��-�)����v!���a�^ ZmT�X:�,{?�� �������xvi�0S�
89��G�𿀏�tP�:L"ηW����a�KR~I/�iQZ����\(O�J�ՅD�}죊Ƥ}�̳��j���L��8Xz(g�Gۚ\�_�������2`J���lS�t��ͭ[\N�7P`$'[��Uπ,G�tmd��R9�P�$���N���\�ąLp�dp$>���@y��Hc?�/E����PZ�U7�6(yv8;�F�k����8��g�dN��)�,Yr4v�<ǎ�b�Ԗh��ۮ4��g�l�pe��D����6��H#Jr}ϞgvE(D;w�O)�A����u:�a*�v�E	��� �M�P��	82�V�폏�zO�����@G�!'ȱ@�}�(܋/_���~h��hH�[IßE� ,z����Z�9���7zo��ݝ�@���iv��qyqf�B��Ζe��03�v���U>�v�T������Bbcvjǲ޾=�wv��s8nD$h%���{8c�-h�փ��%.���mߟ=܆;��ω3�@8�Q���%Z[U�����c��*�o�}��u¯����ůG������s8�����e{޵��[U���Y|5�M	���I���!p�]�c(w�?�h�)H�g3Q-$�PϞ�F��jן��Ɡ]����J�ߥ�.��Z#�C�lX�z$L*́��]�����0M��CyH��R��<��]μj�v.op%p�<~�.��S9ڲ۟i�#�|pSc;F9Z���j�\��45t��7*^�2̉=���?YT��)Ά��Q8���@��l�t����1�33jw�-K��8���;s̖%__)m턮E�`J�n������7J"����_�����s���� ���;���hz�k�8=.Ɗ��9����ŊQ�A�,J4���%b<��TڰM,В�=a����n���`$w5���4��sy�G黕]��uC%��c,�\�۟��7]��'�僞J2�T�!�L���� !t�|��<6�3U����LYF�"��% [
,��IU�t��$t��I�2�2�8�R�_B	G:T�r�&A ѿS)�@�lʰ�P�@��Sb�GL�&.�O�gW��ә�)w�,�rz�Vϐ犳�Hy
G�����[��zΰ����Z۴&����-۟��l`x�;�ZV;��p0T=��*�{^�G9�����m3 X	F�	�k`�rl�9T_�8v�S/RgH�xJٹ��7�Le*'�_#f�e���a�"�)�%N\!��L�m&�UpK��F�هf�S�w�z��BV����B�d���Gn �y��W��:ե�*rٳ_
d��~�çS�\f�m]'�"�{{�5;?x! e��	�a����_�	��J*ԫd����?�:�j�YwQ\F�+�L�[/_�L��-��׿V����O���K��L}n�JƠ������
��b��YX�B�aB�Ӟ[oϜ��
�TA�Xq���#���ˁ6Q3Ui���vo3���?������a�?�Ϡ��m�_jrЙ����3gM�EUi��o�f�go,�z0����_^h�2`���$����^y��w�j�aOA�/�,~E���,P�f�T�^KZ0O�g�AM{�5��4mD܏O�h�@{,���VJ�6IS��aʚ܉� *ƿW&�&ٚ��6H�NV��a{�w���R�ʐ%Ν^���fH�!E�0�� x:U�S)��^����P���<

�H�ճ �E����o�N吼�{��6Ş�\Ur0�ʝ��5Z���ݻ��
���#�;���{/�"���WԈ�Bt����>G����������߆wWgB�,�M:��`�^9X(�T|͎S�q=�?Tr��@��ܘq8[Nm��m7�p�B9[4N����Qh�¹}٤���gd���kS6�X𓸪NM�N�"RƬ>����24F֮�ٴ�3�,���V����xaP��A(S~�?��*��Yаj.up{vp��qo��tЍm�}f��c{��Gs���abw�(\�ztR��"�4�TD��n)���e�N��z�r_�EH�ʞ��.x?S�O�+#��E|����*<�5��]#�O�ړ=_�� *T|��d�mҺ�V��[��H'�XK�Uѐe��zc��LGγ�d(�_��,AJuY�.O����{8Y�,c�
����g��-���S����F�k�8fS�/������/`g�7����S!��[�ȓ!Hj��F�Cp؞�xȫpg���oA��~<gS��v�+�O�����G�\�0"�E\ce[�8]�aj�-�EFh`o#��u|t���K��� ��'�g����^�}���Zu'�>�z9������]\����8V�8��X���(��ݖӇ�NZ��Ys���f��L[ݰh0ni��ר�06�G�,q��=Yt���)8�8>D�5�TrՈm*�/��W�� Q�P/f���=���T`�����U�ʟڪ�B�d���1�i��\$wX9��pgK	�`G(󳛫pg�ڃ�Ih���2m�3��Tf�����l��Q^E�Q.	�D��\��I$��̒Oӵ+�9_CO8�v�LW<D"=��x�E�0�eQt�rtw(	)YZ6�$�p�ƪT3"B�-S2��g,Nq����c@��Hc&�^���!��s���}JJd�g��"����h'��D+�ԛ���Y�|��ԜaS�$t�����L2GG�2�S�F���^okv����5�p�1�Ӊe떩��B��i�%�t�1��d"V�NJGxq��zð�M9ƥD�g*�(����wo�[cn��;�e�IS�JY��ʑ�2E��m���x`�k3�s��f�)�ƹ�r��[s �`��غv�MI��N�td�kk��:�V�3�A�h`M�%�Ele���m��Z��Z�\�,dZ���ߔeѕ�Yt����bl��<�N�}��C��K��X�����+�(�R"ʯ�<k��xn��c_���g=�HZ;gU��/n;�~�4��v3 ��@��*�A������]��`�ќ3��3屗G�P��i0Y��4k�q�#��2�_ZB���'Smii7��.Gא�o�����!$RhN8��:d����Oa����D��s�D���Fj�wK*>9.���&��g/�x��LXN���J-n }�߳h
a����pI!����MC٥O7@�`g����0�0�R�T�����2��hs�cMR �Z�$Ƣ 	ڷ3O������9�}A������>'��Թ�8"�dI;(d=f��x�9*���'�C�)t!
�n�P��,%����@�G�K��V���PU�n��>j���T�m�̆�N��M�	��!��s��ּ�*A�� �1s;� �I�
:�K����i�^76���}l����s�	�E��&b��t������e{������Hh�Fx��k���Κ�dE�ā���+@BX��F��W�8P��:��]�d5�T�qoQ��V''�H�F�Y�#�5o� �A�ڻ~>xt,=�ԣ`GS�ak�v�8߭��%��ҙr c�)�͈�3���p�����K�IƖ)�UV`�@����(w��=J#��� �^���B��#;4�ab�c"df.����Tܷ̙6�ME:��L��L���������&�}�.���,�e!7���e���ۓ��_��Q�20�n����x��jWOk�]p��C2/ႚ�Ԍ?f{5-�?�}�1L��̇v�����>C���^��B���{��D�K��;�$��8`
��\S�"�w:�-3�2������_3(���i�Uj/�1��e��F;�O֟�K|����T	p&V�  ��IDAT�rZ����}'�B�zow�z���^��Jg��<S��A�eX��ݪ�S�_>��Us���i����U���V�v K]�ƝY�zEa^���f��e���H�
3��Ҽ6_�;� 	@��`sG��w�N�-Z�� F��s8/�A';C��+�D�i!1�B9'.�����m�f��3h���^w��̰W��-E�O�i+�1�<�O�,;��aD�|�2�m'Q)�=*y�U�?1B�zw�ŝD�0@geO\��W^^M��hK=�`�l��=�@��P
@�9aH[��p�"�HD�I�� o<�zDAH�>:k���|�O �n�&Nv��{�9��4W���ed�,R�ӳ���\�`�\"x>��Mk��D��~��q�MQ�O\���,##W��<J��྄���k'k�ёF�4�-]fT`V {�L�P�9l�m�X����"L^>�*)\��y��}���VB����݉]<��Gl�]+\۔��<�<�;5[%�v�u���sgs?qTHY߮��-eM���}��X�
�݅��+a��N`}3����	�A"�eIц]+�yM����$<;_�^la�d2��2���dDx� ժb�-t.*;3��x���|`V��Z�V�� ��E�hȶ>�0Nn��H;F���0�UC����RGRr�ȏ+�V���T�7�B�f�!j7Ԑ��A�g��(�6��yS�r�;��mh�ᇓe?�����PNK� ,�Z��*�H2^�w���,tT��3���ۢ��]�6���0�-R�΢����Ζx�+�t�_��n�/�J�!x����BKV8(�R<�dڸb�aF.�,#�]��:�W(��*@n&'����;��Fǲ��*�|u�%�e[���l�n۵IC�s�R�A��p~^�(6b�= �@�t��J։|��T��
4d�鶖��ӣ��5��Z��H3s��U,a����=���$R�+Q�[����c���	�4�D�D���XS�)Js՞�܅�2����r�B3��9sUM�!
�2Y� U���_pN_��J�;ۡ�1��g�)=A|O�܌��|�
9�*l���=��n�u}��]YSIF����s��  ��
���m�q��F�h&D+A�'0��K��z�%p[Yp&r�T��%�.L���Z���ܳ
���P$p%q���Q ^"�C@���&@ߒ�a��J
xR�b���u��:N;Q;�L-�2��1�PkK����h�I��+�ԡ��U_Ɉ��>���j.��<+1Q!x �Z:r�U�`1f�c��2�Ǘ�q��Y7�.c�ƛ{e_������;"���*{^}{���XFp s��.�/�;4��Q<�
�hs+��|��!g�@��_́��桙�-l���R�|�]&�����hk�Q���_|<O����z�L��6���|��|�?έ�b-qh����i-���0 ���譩����}�����i�� ��x�	�mh{�Ck�ϕ��7�U��6�<Y��
zD$�bAu+)��wIX�|ΈWJ�V6�oʂ�&'�@y�>_��Ξ��E��yY�.�x�\I��KˍX�p>[!Ъ��[�5Ek�z(���q�a�yR*A��5 ��^��9�0�2��s�\A�\\����F��9Q$�[^���%�D�MW��H�!�GT����ot5��P����aN"�Ռka�Xc��s�C��5���>�G�#�v��aa�0�o��ʔ��>��j����rf!T/,".�����e������2e������=�,ɮ4���O�V�JWA��l��W�����
�k�q�F94�h��h�P(�:CG<������s�GVS��CGged���ޣ>����@��|w~�m72���������W�!�bP��Ϧvh;W����>�� c��,�����F@
�Y��\� ��=�+3���IҞ�uxC��l�nv���?W!\�d�穴�	d��E�W9������*��Ρ�ỵ@�S-A����ZլՅO��R���d�g��ݛ瀚'��#r-������|ik��UW꜔7.3H��x/.�ώg3_jg����F��.(@e<}d)Q�P� ���4�$~��i8�%(�\��^,��@�T-�H�s.�IW��(3��yDr*�s���<*�G����DA��o�v.�k���V�<���8+�y���~_��Z�u���j���7�Iˢ^*	e}�-�"h/cV�i?��G�T����jn�_��t�@Yk6lg�����huI4z��%x�R�+�ڴ�^-���:��?�Lƀ�l���>��4��������?����
�a��F���w��7ߧ��>�V%��� �0���V��P��g/S(5�LJxn�υp^7����U+�2����me�%g�֦^w�p��Z�.�^����KR�K��z��#�PZ�t08_wO����-	֠��~Ғt��v:��*�F!�{��M��E�+^�64�,��]���j�\�x�)���=~rV(�ra�ɲ�OUA�d˴%��y�+7�s��P�l������DuJ�L��ᙝM8d���9�ø��:�^�5�½��5\�q�j�<�C�I7�r�?�Of���I�����@�����N�$���8��Ȥ�L�A35�LNR\DX�PA�k���OON���+�O��;���S蔔	+�f&���-rjQ��M��7w�*��M�Jώ}����NZ�]*W!�� ���B�NU<�8.DN��>�@�#�0��woӥ}	]	
W�+Y�q�$Ȳ���$�h�Bh�����z.Cm�w�q�g:$�	N-�����
]���M���}��K*T��´�Ce��_������|��w����W_}�`��\�����-h�t�w�D���w.8@�A�Z<{�$�W����O����E���[�N��V�x��+��8�,0-aి|w��-�����{�r�`ӎ
�e�) ��VC�"��>�ˍ�1v �$�����X8/ea
� ԡY���n ���J{:W\mt 8�B�Q�֑Ǽ.�ex�-Q��Xu�I@�(��J�$r�i��$��k���L�O�j��:Hh��<���_�lI!��J9'T|�UW�E<d�^d$w�dk���U!�Z�˰�c|r��d�ѯ8O�Q�Ě��l��S�s:�$�T����$�Q�hw[�����3�׵p�i��gcݧ�Fb|nY��Z��<�'��3ivy��,�]�)Rk�
Q$�d \Ž��}�$T�B�w�~�wФ�S�pr���)f\k�N�hsO����~��ME��U��uR"��2��Y��`-P�J�$�v��<}�=�>��SKv�����W���;�p�"��v�����=�{J ��]\�[b��ma�A�˴ļ���G'*���W���j&l%��2�f�W�c�d��&@�I2��<4�;���V�'(���j)�4��)A���r�z��BҖ�����r����@oE���@���z:�J�n�}W��A3taC%�
+�6�.y�g�&,2u �a�y���5�`�!�#6@�!]Z�4�f�5ʢA���;@��,��p�t�=P��e^#o��	�e�r/�w�"^��O��A-f;(x�Q�3go����DS�����CT��@~{���X�r�=��:2{/s��2
p��ޖmr���F�~S��Q�ZXlf����	O����N��Q��J )���4s�jDY�~��F[�d{����x�z?:>M�}�yz������{�E���|s�����{ �&ȲO#A��vn~��,���b�±�	�5F�XȩR�����BF��9��w{Ko�Nή�m1JϏ�����v����3�����`�%(��%wQ�ֲ`���lXv�=} ֶ&����J��@�/G��1�h{�y��h����M�s�-D5]�jJ[�^����D{��+�+���H/�J{vH�^I����5�N�
ʟ˧fQ�����l���h�Xpw'f��t�)���s@)�ss?�i��2fռG*>h7+��|���c�Z	4�k�Ύ���?7vͥ4T�[L������S�3��Ź(7x��hC��ַ�,��~��e��uw�������|ѿ�*���c{_C�z�̲��4����3���	��:�u�KAΪj�|�墲�[�>��ҺQ��A��t������i�ۡ��_�����u W�6��lqr�<��Y�Z��Wě��Yg�;��[��dk�>#B���
�"D:H@��~��ϟ��O�>O;��p�r��BQO�:<=� �IQ����G=����kۓ�E���O�ȷ�sCkb�Ck�8�[06�B��o�]��Q~(ϗr%�|��|��ﵮ����nN�֡`�dr�&;��BӔ��r1�@ ��H���{����X��hO���A�=H�VA��N�5�V�e�}f=ᯂ������]�qKv/+�$�:<�r�b�M�G�I�N<��[���M����'�RNXhC���V� �ME�/ɹ�)���ɢaE���zc_�:ʄ�� �<�n*e�)M�I�aV7����[h���tR��u|��;>[�J�߿�z{�ꅃI<Њe�H+u&k?���V��������rU�Y��m,���W�[��.]O������Zd�PȖ�������hf�$�����g魃e�N�
��[��7�L۳�b�����X�D�IR���#mj��!s�!Y�ݛ���y �,k�'*o�u��T��[��Lp����ގf�t�b��y�<g��A���k���JZs1oŻ�B%� �t��N�'�1W8���]˶*��^��l�k��,�JKq�Z��%�3�K� 4�V��s�٥�(l��!A�׷ ���#�Z�/q����w�T�KѻQq�mqz�z��`���G�p�+@Hj��¯�AjۂF��t�-��ڂVΒ��!���Jg:�_��/��u���kU��xIl��U�_k��w��0]$,!AÓe-s_��H>�� �a�ʾ(x�_�J�,㻕�vR"E/�S��t$�\�R���~ e�Ƙj���}e�ٮS���������bѱ���Y3��E�����Ӂ��;s�D�_8��[�w��$�8�����Q�,��X�n����j��Y��,�'ѧ ��'�t0�&u�Ty�w��]�����'�S�˟����h�џ_��7�8�l��g)�X�0> RoT�&oy��L�}B%r���\5A�*�);\|Z��[;���E���o�o����;ڬT�^�������켍CG�Z$��Z��P7U��	�ҏZ���+aeDMX�X�f
���4�siF�y���t���qnAf]�!TP9�
$���%��^"e���֍�bK�<�$.�7�P�Hݩ���-���D�ڪkwP�\a�b?����	d�Uۢ����!4]/��D���6L�Ꮶ6�Z	�P�%d΀� �5��񇋢d&�us�Q�Y��x:�Ѐ��,�}�7������VG�;�	���CU\g	��u^8�Ta��l�Fz���y��"�5�
�r6
�"��ަ�w]x-����[�e���ew=�J���@|�εU�tw��N����+a^p������{Eb���Ѯ^(pֺ>��Qj�����h�q�%�.o����k x`D0�M��{)JR���Z��ʁ�;2�A1,i5��$թ�Ł��pk�Z��f;��](�R!�b�Y�>�:� �t]Fl��8)Ώ>�$����歨A�7����ltfl���dׅY���sK>fjQj�4@��Y{w��Z2Yr� no�,O�\���r���wqs+����:x58ьU#�p�b�@R�z��K�;��!�^_\����ݳS;OO����]a�U�(���0� �	t&|��]��Xf�)�QUvz|m�F
x���XK`��EG{tl���F|����R(��Ψhz)��2�	w�S7���}�>��|�TP߂��𽞺��\��u�,A��zg��%;W��,�k�Ҙ�]�$NI�Gs$�{����(	5��3?��W�l�-"+pT\�Y�	X���깪�,5����\Br�mh!��K&q�L_%�w�5�! (�B�-��_�F�3�����;�!� 6�n�/�--��"# �Y�FWv�������vT!��W���[0U]�}�H��K�y��Ӽb}Yܷ������"ra��j5K_�}�^ܜ�������IN�k�d[��%�-��T��h��o&��w�jUm�BP�1����*�4�6\I�'��.���{Oָ5�M����O[�yH�(@CY��ˑ��'E��_�,+<�C��#1?8bY�j��	�[�]��p��(�Ц� #5�ܘ�g�)�M���AnfR�6���.8�ö���N^a)a�L����I����g��9�g1�B;N��w�^J� �#k��<x;����Z� �����la�5��hߑ�O�<I~�Izz�&]`�������	-�\��]����#x���pM�{�57�6��T�K�N���+�5�����H��j�U�����:X7�k�ި�Zۚ�ɓ������v�~ש	$v1p��Z�\~&� �N��f���g�W���ע�P=yt*@��v�v��C"�)������6��qP�A߳�[v�������c�	���_�g�;^c�Tx0�PEok�ݥ[W�>H/��� q�Z�����R����m)/��vj^� P���D�	�b��KԦp��K4Rv�����6*���0�u\K�-���ɭ�j	k��C����o�������j�Ud���vI�h�W��#>�!i���\3�+t��lm�,���ߋ^�̱ƪ��a��]�%�4B@i������W��oiK��J��������I>�n�*�>T��oԎޔ2��}X�^F���ѝ�]�v 	0�Fi]�N�+dZמ~�K�Pƌ"�K
���k�qs``vtt�v�沠@��.0� +��M\0I�9��9z���l�R�p玆� С��>�x��p,<N�im ˔�b˷�1��Z��x��=��MG�@@N�z9���/�H_]�IgW��B���J.R�?���5�Ƣ-����}>����g���Y�����m�qr*��=;xWs߬�P˳�|y� �+�ؠ�=�[� k��̓0%c#?l�~L�����W�����L]s��Ѥ�)�IZ?G)x�9��?T��#���{S�^wVQ���xC��.ިtO8�n�/eb�z�j��o8/Dt�+�qb���G��ޮ�ൡ�1�~��pvy�6_��-
>Ĩ����7?�U#��BRR������L�������Cw��v��!�܅T�>�����ç���M�?�1�7-t%G��JU���z��e:�;H��'$Ϋ�8�7HZ�xm�cj�������z���:� ��-�퀞"8�W"��w�V儇���b�CE�p+L06�>Hl���#��~Vkt�	2z�Ⱦ�ş������Y�fmn|<F l�Ô���(����ѳ��-"8,r�h����z�\�����?�W��ֲ'���;�r�6��Z�B�=�����-3pʕ����&���O.ܻ�U�`5�Ŭ:<1��3��|/���n��'��R��K?~o����c�zv���Z�Et�6Eʑ���=8y�k�jZ]�l�҄�p�v����9ْQ��F��l�tQ+Z]�2�t�TE�;�t�۰<�+f�됖�|��縴sA$� ����wq&�&UD�/�{&Or�BQ4��H;��ɬ%_��h�C���ڜd���g~j�m,;+���7�w��V��������Bҏ;��T�����6H޾j̞�r�b֪��o߼J�W����Xl���0%���E��0�p ���,�gj
t �ɛt������� \�Y���G��Of{'C��-`|�⻵�?O��a��d���6��r����l�J���`�,�+o߷��&�2Y�����t���{㴾�*�o�*���lt�1�Ϲ@Q� ���9�Z���RhN�Zw�x�U�}�ϷMơ@���t��Q�i���j��7��C5j�z��q���x�k)����P�:6m�x�|�b�p�Q����T����1!��p����'}��xy�^��G��k򬷎CU�|9`�gܲ&���X7��Yr�"k����������5�~5w��﹭C��8@�d�f[�k�ʻ�ttԁ	D��`U�U�<�ONR���j_��+��U��Vii܍���EZ����Ī�k�ewW��F=i#��J^��^�Ģq��	�2��_m�`��RU7���O���Z�CF �Qd��*K �?~,`�-ISpQ����]�޹�b������I��.
v����;�ן}���=�?��~Mֲ.�n< s��zpf�f�q&�d�Q�6)���.|��O�}f�3�����<�J]ӻ{���Y��wu a�
ipT㍝{}����,9��	[���hфmӍ�<�i�7l�����￴ lI룣c��H�7��鲻vut3�A���{:R��x	I�8w23������>�l��e~�X���o~)Q���=�\8!ΛyU�V�
 k2�W�E|�L�C���0և���8?Rt�W^#�+Mvl�y��&��'�^�Yٛ�<l3x���C�����;��l@Ax֛�~�G��	���eZ�D A�Ȃ�Ֆ��6����Hawۨ�]&n2A���ŋ�����L����(Љ��=3��E�z�psiC�×-���UfT��meC
G��+W����ů?s>�}�N�ߥ���=ܖ�We�ד��td�M8�@��\����5<c�G�pG��,����4��v�tX-ڶ��h���g	2[�z.;׋,�-3�����T��� � ����=�p�Q˥t��'\jG�G�����x�Bb�T�u)�.H�N�!�ބͥ/\��0SqW���SAm�VH[���l�VU����8�cZϥ]��Q�E��a�%r;,��P�~��ߥ�w�شCkC�Ш4�^�G"���5�D�j�I·J^��7�m���ѡ����FR��pX�=�:J;�'��z�(�:x��q(q�2E��?WVh[t����"�;ܔJ7�Y�������/;N1�`P����y�.�7����×j�n���_�z1������%��2ڢI�a�Bఔ�u�z�3�tc*��	D��lt� &�)�]5��2z�[��;9<R�{xx�>��4��ق��)�����7����C2�,�}O��;�˴o{�h�@U0�pL�n���ξf�@��Tk΅l��LV��u��FhK��,�E�� n�����P��'�b@������@�O5cS����pAܫ�DAc�$�nɣ�4/ڵf��Y��Nm~��z]�F{� �y&���܍F�EW�x$n5F���Q�B.���u�BFW���:q4B-�����oI?�m
���qCm��{�ׅ�����vZJ�%�f$8�v���܅F�u̢����E�E�J��q����|���ڑ����>�o��䟹켏�.�܈��1�'�F[�,n��|۠��ƚ���P�$0��Y�B�IѶm 4H��P�:���-z;#�qH�;~/�P����d�,]^����s��W�V���ʹ��3
!iK�v��������~�Ĥ�G^����yP-� � ���U������N5�����w�v���3ٗe�AZ�S;�ok׎��-����A!9�]��D?J����婞��:^�vh&�!4/Ckۘ�j��Ո̿tKF��|�Y�4�Y��}kq#���_@=d�E�h/�q}5[m�ZI`��-�G%Q����6c)u���@�����K�@�����M�ȣ�>	A��Հ���k��|���:-ə�Qp��*Y'9��h�'�[
�z>4��F8xe��D,}����<���rJo�	!�p��6��ɡ�T���.��l��խa*:Dσ�x����Q*,8�7�YN_[��q�ͬ�,��T��^��gO5k�b^�{G�Jr��#>I�6�4]�~��YPb!�����z�4�!�@���;�����*��U�w�~��T0�lR'��+��4A+�߶��;�b���&��p�r(��a�'���JrG�D:Itȇ�- a���

{H���&�(�w5��H���C�t (��?�����*�u���H
�*��ˋk%$i����y}9�
�]Z؁����GR�R�ŉ���Y�?#�G7�5A�#��j(}l��ٞ�]L�sb���֨�,�H:
g`���d��R9R!G�<�N8q��5���ٚQ���м�!����_����W����~͞�)��$Y�����C���� �ʻ2+�%6
�`_t��nY�Fm(i�1	-��Q'TB ��ݿbk䒬�:���mic��H�R���I?��3�u��<�=Z��om�]�1�M;����|�m��y;��Ѹ�$�zr�^��O緷	;�%�{��J˖�����3��s䚻j���Ɇ�:�
�ǅ��n{�+R��{\�BN�n�L�W�~*W���~�&�]ԝ����~g��~u�bj���=��٠@��s�s��Z�{7��p$���ήԼ�	-[ݶ  kn�����T���&�k9�L{aY�v?mnW�dŎi9�0cAj����T���TN��+���H�B�YC��Md�1����3��{���r�$�hnՏ����+t���sr\c�����'<�e�&j|����+%�<SWOr�=��]��ɥ2���.L��ȍ��bc?g3ݤ���D����u0f��'�@ #�tBHָ\RH�
��Hx�sA��u�ڎ�Q��
<R�xu$w#<w�1
�����L~�4<z�>�7�J�x {�vP���i�Y�$�[��؈�����m���J���[���v�JW���.�H:p��k��i8�sD���6oS������Uz��u�Z��hf�$Q�{���JQ��Y��ӕ�/���뙤d{����+TM?[D˖ĎQ
i���q��m��{
u��� mzZ��;#������c��eYb/��X�*K(ґ��]�Z�7�kT����٨�Ჴm	9����?JǏN��In���=�@O�U�G�;�UK�����m�t��&s�P-3�CZ̸Y�6�&@��	#':���Щ��q�����.ܗC���.>�T���;�a��yTЭ��$̓�j2����Z7� K����K��#V	5�X�s�;��t90��粸WXLq���eXS��t���r�*I����{�r N��Z��r�tϮ�w���|ظ�&3i��H>7nJ�EܢcKQX�Xh�o�y�������i�=I'U�Ξ���T���.o�hI˦i�3?]��^�^��EH3�po!� 0�h�����{�ju�����s�p5	O�\�pұ�
S��"���� ����<�-������Awt��>9uA�9��,ח��/�����׿U~������E��ܺjL̃�&�������v0���VQ0<���M�{WW>��{m���7��Qq:�����,�^4�.��jǅ뒮˨������h��4��� ��E��`�c��7��E#��RW�7aYwc�9�OHd���|0ϸ��:��7�w��@ ������رѩ�c1�ƣj�Q&+�,�FZ�(���u���J�-T���N��ޫ[.&UĴU��o�ab�@�מ��0]�M�%�&�����n�ԝbv��q�G}�jmj��E��mwm��x_��&�'Mے�>h�E�	\���A:�J�|�#u�X�j���n��ͅD򡖠�utr��..u���O��T��u�X޼|����w�9�vDy³��	���r.kL�G�	�?nv'~p��]:!e-1���ܥ�k�������M��tĶp�?�ĭOroz���w���;;K����̗��r���V� AB��7NsD��v�2��H7|I��Щ���	�7VpM-���Q�B�m����u�A���Oh@-㤡U��E�T�^q��!�G�B�ܫd�gA�c�,��z��������9�.J�|t��旍�Z��o��6�~�J�[���$�Z{N���c��ѝ�Ɨ.=K�WX��^Q�K��%����ep��h:ܽwCY1���7�GU�8�\�ljԝ�F:��I'��id��
A��NaT��q�8z�f���a��1�N�"�b,
��#,�D?}��Q�髯���a�@�xG�JRJ9��YU�ζ��X�l��:@�Q���ĕ52��Dpj�rГ�2�6+���K{�;,ά��P(
��f��*����~:��6# ��U�h���
���?KG�>��7r�x��]�>���2c̈́�0�@FA�f8��&U�O 6���?+7Uz�T��x���(������6�<]\��?�������ÃG���� ��},�zm�ۢ߂G@P��3w�p$CĽp@��t�@��j�H�#kU��t�	�`Tv�2�3_Z�\آ�<���yH_�r�-V� <U�:	�לD@�c���+���a�X2[��8��@bg����v�ֱ�PFk{>�B��΂� �ЌM	��8�5��`S��������v4S��B�L2@��{0�,|�J�]|n]���K�:؏�ܰ�rP�%������`L�j̒�]���ܱxb�c��ª)I�h�Nӣ�C�1Z�h�v�h*a�د��^����[��dH���@�/��ʼE�q�d(����p��wgkW:�]�I����#�\Ҿ[�^��ڍ
�I�j�xe;��o�i�lK��*�=�d߼ycAr�잭[�b&��u��^큝�X��t$��B�6pc����-(�~�˽��� �
��g�ӓ�G�'g�<	�G�c�x�oAuI��#|7ugs'lA��9�3��;Bf�)$W�1Pʫw�Ô!3P��H�ei�����Q��3k���~Ï��W/�yF�c0x�5�M����2�\�^��2Nh��Z�;C9:��ɾ�r��hM�j!��*�Tz��U�{>?���2�{^#�Ë�/�D;c�wҳO>J��-�k�i�s���u:�ݦ���\q*ˁ߯��#_���=�Gn�c��k���>K����M�#���#� u`�zQ�h���N?���$Wj�u�ѡ�AVr�Q��X��\��h�of+ׄ�kF��X>��S�����(Zі�N�r,��N�� ؽ�H����A��y�a(�^K�N,E�ǖ�Vk������g��>�N�MR��KT� ��E����2x��tA���^�z�'�@��7������W_�Wo�t��G���)��P��V��Rm�V�Oᄱ��m>�L8/�����7�PuPUw��3�ף����M)�nb�|���X{�	jPx5��+�������&��R�hI�KoWo ����1�jD����M&M�hf���%7J��'<hM笙"���T`��C�Ͻ�>mlt:�<>=},���}��?{��������=U@�'�������!�F<�	)�ƻ7�J���	�H�{mJz�S)�*�|F��BSa�:T�21�5���d�k�+p�d��:=����}U�pCgv��g� �N�q��k���!d*��r^10jm�˹Ь��c�jìw�V7�4�l�R5�-
]�/�d���8�$(\j3�� gm��"�j��$�nDM���.�m��K�e�8���-�>:�\f��*,�P�S��]\I|��H"-��T�������?umt��wV��+Bҟ��4~��0�Z� k4{Ugr���쪭O릣�I' �P#�KЭӌH|d>Pރ���5*�j�ty-\�`�P�/Cm������\�y:�;��[1�v܇��W�H�s �ɸ�r)漲��ǱJ8�P�(%�Q]�5c��aydH�aCɄ�]�,�:/!.0��Ŋ��Ȳ�йܙ��/�����_�
��ZR�UH+F%_�m�����,�����xG�<�'�<A�(k�_zHM���fl��o������d�m�le\:x�#څztt��?��ftW�/�"LY:q}a\�È��J��JtؓU]�
t��U)H[2 �<`�$��S�<����4�J���{��k��8���9�r�*�?t�*ti����B*�l������ԍM����~aA�����EpfQ/�X�*����u��k;|ik��.���p����N�����+�w6P},����A��ls�[�u�P�9J=�
Y�t��
�b����V��=�
(~�\��RI������+�d��LP�	ʼ�ĵ��L���W���������7"UxUwT)U�V��!e�C��d��#��/q)�`�H����"�?{'ay�H/6g�!n��M:hl���4M��^\�p�x�V
F��K��q Q�5E���r@�T�옓����l�z�ܘĀu��:��֗���J�;��_%<BbbU4s^����E�ʿݹ�� V�{V*s�%��<�L;=��ǅ�y������D�%�v%�>w�ɾ��?����}�:�e�l�m'�� ����RvE+�Y�ފ,3��?蒱\U
 )H���|��+Q<�V-KU�vIȦ��
�9����ʒ�M�m�;��O*F�R6л��ӗa�?����ܣ��������7��)���ӂ$nFg���4�E�dtSDP� ��Gn�k}E�ݏj��F� K�����\��<R
ի�ݎ61ߕ����N�(w������v�x6�ɘoGW]7И�o���.��ga���z��TN�sW���X�I�q������N+d3��N����I��F��k�wڢ���ף'��s���G����=]׷V@A9ݵe���(nVR��$��x�ֽv����?���y��I鲔�I�	ylAc梱���҆�}<N�[�v ^�]�B�I�ށ)'�ӑU+��(ޯ����N��p�R.�)���U����2� k~��Uz�򕐲l,��]ۄ��9ܳ�o_l��tr��v	�}�[� �ℂ�mF,�_�
l���AS�S�u���(d�}d�E�v�����ttx,t#����
���m�E��о���6��~�n.C{�U�C{�C;��m\�fi�P�5ai�siٌ�RZG۰�D&6�x�T����d�� �r��;���EՑ�^̪�³{���8�Cg��y_	�P��������{ U5
�B�P���ֳ�C�p*a�Ch���9�P���;{�6��"d�0wA
0�=v}�:���y��t���H��pH:��bpX�6����p�U���	���W��<�ZT�u��D�(!��S�,�@5YW=w��~v�cW�7�}�wm ����reڄ{�n�Iڽ8}y�����.��x�W�]��%�fi�<�^M�m��}�*�
�Q�s�"������ByD��`�ֵ�N��ϼe��>ढ़�oHn�2p0�m�S�]�e��,�����@<��t���u7���p��2��TX�mT�hp�񾳾~v��U4{�s��$^tu���'�GN���Y9L~օ����C8�k_��L�C�~-�؍��YE*������"f���l��<��-��F��էR�ٺ����d�Pw�fqm9;�H�,2���@e�əNJ k�!�"���~ĺaV�*��v`��z`�Q�*Π:�qu���x �tU��ė��t=�U�G�u"B]0+#>�ړ����u����Ʀsݺu��ӧ�����6F�Py�q����'r�y��i*���:Ӎ��`�ù��@Ipf7�=)qfi�� t"־�n�1��L���裏���m�j�L[TrV�2W�(?�?��b�m�2�2?�Z'�KvW�>�(I��U�e�9�̮�����6�N���z���U6��8Ǎ�W�f���rI>Z��ᵓ����LW�̯���u$��X� 
��Ar F�k4'�\��-��V*�t�9E)����&�s��(c�i�e�"]ܹ��:���mY�n�yk6�浖��zE�ilI���+���N�J%�"Y���^j�+���;�c�	��[�_Z�L�����(�c{�^.F���h���Y�mВ:N|�ߜ}�v�����P��%�k�w�x��b#�b���ٳ��g��rh�y��9O���'��\1�l|.F��gvG����PDnX�_|��ڍ�^��́��:*�wgR @�ý��T|6�)�ݷיWP�r��J���� �Y,�
�h &� T�4�C���U����<�<���.j`�׻��U�Nsh��#w+cD�^9�Ǎw�h�R�P� T!�vhl�H8���ˑ%�G�sT�����e4���<ir���0��+�h%�h-^-3g�>?�-w�Ꮅ_m�����ῧ*4�\�"��(��
#�`]eQ3�F�/u��n�\���>=Oˬ��h<�dg��D9���)t~��+���̨��5�S�,���@G���Vׁ��b��I�EF��=+*a���k	��'O�3�'�K�K?Flet'�?3�b6���8���"X�6�����Шv�c��QNek�	~����]�Q_�-{9��Y�>���l�B�UQ>�z������Ya��/�p��Ͳ�7����E�����zd�v�s�z���)=:y�UJ�Z��ˬ���sd8�JD7�����T�rȶ	y�ą��޳�!�~���j��n�+�ޓ9��yᰡ�[��1b�j�7ns�jnY���Z�ld@',:�-�����{���5h��n҉������:�/ߦŰN��wiv�&,Ze�
��,�
n�xV���UrW�^�,m?{�V[��Ȭ��C�&s�_��g�KJ?��wk_�����iH�X�s��nX��kU�?�����Ȭc��3�\��,*�Q��m9̱�G7��jn�;�5*]��Z���4� o�V@�T�p�5h�=}t�� ��@��٥b�h㉂�' m�T����K�>�͊T�Q>��(ɿ�g��SʐA�n�x��Xpy�����_�:�X�6��җT��^�ח�����q�t0ZVt��<�q�ɥ�-F�y�'�w�'�^Њ��F�Z�p�z(��G�V�IE�~���T<�S[2 ��
VAv�`���S�oF�l�F����E�� ��<���;22���H�9�]:j[3�� 3� Hl*������Tctx�z ��:�KgFh�ݸ4g��N�����=9�8[LW��j(�+1�=�g�l.`��x��x>N5Qb�~�a��g��_��ݝ���uj���DuVu��Ȳ�r/Z��F6��Y����{ۊ@_m�,ԡyj������W�#�u��~�ZR��z���l�V���Ư�+�g"��W�\cփ�lm�]�!
]����:g;�=X��ڸ�<#���c� ٞ�ʘR7N*.����T�J�ƽm�������h��ίε���6x��}�"��@�s"��ߨm7�X[I�i*\<�m�ㄾ��lo���7��~H��D�밈ku�b,�<��Lo޼K#;HD��w��n���g�	i1x�Es���ʕF捖#�3d[l��i����f��8]��I�M̕��82=) y."����2�mU�jq�[hQ�8YlU��F��vlcL��٦���a��`�>}v�Jl0�J��K��ަ��U��j���P_���ե+*�,V�#xB�[Oi��R7�z_Z%U����4:��p�l!��ñ��p7̊�f:Ql�k��T/	��j\����?�o��	��snK�N�޶ÇyX�<R�mi������ ��J�kB��|4?����Y�)z��2f�w�~����s���8�>w�pmQ����2ߥU���\�����6�*@~h��5	��U�Ԥ2Ț�p�N�Ӯ��ބ;�%����O�Z2ٷ��h�0��?{_;vF��7��+��oIIH��@4���w3�R����I7v��ߝi�Hg-h�#�k���ѵс�H[�����1�z{���	��e�)�t��D�J��ҫ߭P�ۦ�����{�9���쒐nwH@!9��Rr?c8�����t�p�oR>�=�o)�_Z�B��ɷ��'i~;��oȖ�O� |���rյ��ҳ߸�R"y*�mߩ,ٟ�㑘+�IT�=W/����ۏ�������RV��/�./=�e�o���9'���c �t�����X�L��5x���-I=�������~v�v��d�::]x�_����o�Q�s3���B�W�@ɢ{�y�⅕�!��PI[!F	(�]�g���Tc;J0��s.�
v��Ҧ�ꥁ6@}ϒOT�@,�2:T�*E'$���R��9.�Fr4����Lg��iS{�����Pe�n6�u������Mm���U���|��@B�]�X�rE@ ��0���2������u��-�
O�h�$)�b7�O�F�3*~����Z�x���v��1ֶ�[-�f�6�+�D���&�H	����I�iC,Bv�����ךּ�M�yO�y3�8�B��g��`wh��L�\ڂ���(���A��G���0]]L����4�xus���`��j�(��`A��S���Zu�;��(���b<>HO��>����6�Z�V��V��Y���Y��0�6��a��a=FU��9�@���%�	��`�Z�O�Gل��xܴ�Q�j��[^U��/�YXHm�2u�Х̄������$ �9��������qk����6�Qd%�ql����B��5Z�|�y�����dA~#�����A�XA��/;��Q#�~�
�������ߴ!��ć~�<������=o^�L���&�lB�� 2x{�ZӼ7Xr�
d'�S@��Y��#�u2܎������&ڃ��5��?H[�;�d���c�4�Y0f��	���6�_�x	0P�a�I�c��m�wЙ����*�J�"�|m���Y]� ���f�4<�{��(K�<����w��W�3�!M�Z^���	X;�C���R��0<���R=:I���o���b�D����~d���������?}�^�=}���߈hW�<|�0�b��?ɨ�R�^�6�NV�u��<?�� �D\|�ׯ_*�?��Y��o~�>��s=/�<g�?����W_}���se�r��wZ�EI��*�����|��>�sN��:��A:�Ƌ��*�����	I �	�w�sz9(�jg��-�@�r�,�!��z�8�Z�Evdj�!wY�X�C��)���M�[�6��g<~rnBGOrF�j����z�0���l�9�ww��G�3�=ae�uW���|�}ڝM����Գ*M�,K����>O���*,�A�KU���(o	��� ���*��C;�M:��b7�J��1���R����	#���% �,l$ �k��,�K3����2{[�y�wM��`�}~���M�ޮ�>��W�f~����F�tk��Rϝ]K�l���Ȃqdgkc��&.�W��Ҋ�5�s*,�lq����>r�N��'K0�����4��F ��p�*z]�?���`,񥅌�8�T�K�x2�D����]��-g��cq���h�
Kq�3�6���L��-������-HUorZ����$3D�^����v0�� �!����E/����0�����vt�Ic���õH?�L;,T�J\�  �z�=�}�c��z�Z0���
�g�.� ���H��#0j6X�;F]+��pC�c-	����>�����Q��Y�Ⱦ@���<�L��X��uf����,�aK �EH�q>sn,���U����l��C�����ko:�]3"�����U^� |��4�����#���>��P]��H@@�M,S�{��ʥ��������G�����p��LR��΄ar��w�g�Q���/Ŭ�2�����P�^��x7WWbx0>���LP{r� -iG�3���:����Z<1K�=��8��+Z���#�ԹoETuШ���{��>��3��\o~���������?�o��֋� ���a]��x�L���E{6�'�~��ϵ�4(�;�sY���������G{���
��r]�����xv&���--!bT�`>*�䬗w=����>Em��/������܁���3�j�vhڥ������O�~m��^���[�34? 5y��m����/f�����!B�Iq�A�6���2�Z�vm6I�!Q���ɔ�C�`dA���\9z���K��w�4��K;��ڵ{�b�ǌ���7��a#p�*.c�����4\U6�X.&�!���M�E�Lw�*��il�}x��w�V[6zw�8��\��'2P���?���,C\��]����͕Ͳ�J��B�b��+k�aN�p������ۖɼ�N�b�l!WG��ɩ2�w��Q���L��)�KQ]��	0
����ݜ��C�rT4<W�9s8?p�)?0ĳݸ�C�����ބ�q�9�l�*G��f���9�c�*HE�o�VR�r�1khkw�*�Qw����Di�@���v��[|^�zPu���9��w=�
rKR���2������sV�=�����-C,�6�1>�v�v�r`�a� ���ۧ�Z����z��h�|]V��h�0����?l�-��A
�)zrK;��E��~(~�ؑ�n%��*��~��*r��q �KQ����N��<�q0n#'`��EtA��y���	N��U�����$PU�͵*KZ��)g�"Mh��!4�q���,�
�w5��wijׇ�A_��Nt���U}5.������RO+���#)<�M}�. +TlP�J�P�F����ܸ޼���c��3�<'�m�EA)NH���̬�{~q�}�̏�}���xg?���k�c�t�ϟ>U%��������˗/uN|y�$���Ɋ��������������$5���|�$�9�,��IF����G���B�{��(m Ȃx�rT������(�AnS��k>{'��4�u��c��Š&`O�4<���*ܳĖPY�͜��������������E�MU
�v1�L�.�U#s�@���:ZՀD���|H��`��Y�8�ݖ��=�b#3�UE����k�ւ�K7�tP�`'��R�Z�Ұց֦�|�K;�fw���t~u�>{�<�o����2D�Y��%_����|�-2;	(�UK�v�(�DF}�ô?X������t����҉U�[����Z{a����� �4��k/0o����E!4mch���D�K(2N-�]YU7F�sk��V}�Gv���vtc��z6�I�U�L���`9�V]���8\7a����k���:/��*���SP>�����5�nP8|Q�"�J�0��G�d�ڙ+�b���xR�چS�h��E�u���[��m� Zcɑ��-�����Ȯ�2��������:SM�b��gj�Dm�C����?࣑�������Լ������֮%J#U�[�ؒ����J[Tèɥ@��=��UO���hT%)v�JzҾ�D(h�e^�?�TP�޾z�F�b��?A8+�=�Go:�����Q��������`�t�Ł
���R-��bH�2|��s�k��]�<��]9e��\&��\�k�:[��6���8�FO~hA��)IS�(+�<@���T��(|�ѭ��k��B��RB?�"$Y��i�g���� ,d'�}zٗ�A�b���6+�#�n���oi���8[$���}I���v��uo�^BM�� �se�	��~�.D�r���y����/��|x_{���	���NR���ߦ����?�)�����?��_�2݈n
�S>�+�P4�l�աI�b�*����=�W�DaL�{Q!gIk��oH��B�����u?>����`7!�K��_���,4�+F�,lK�����\�d��J!�򑚨`��6Kn�?C���[���������Ę������]���?�7��H&�3	��l3 3�J��NB������sD���=�f:;�-RQ{���I���0��u���SW�L��I*9�?:N��8h�����-���h&��ki;��_���*[D��/���N���:�M�:Bw�n(U��h�2�^����>>�NOO�ӓ�=��ýt�sS��f�b'��{�^-�W�d��/�ծC+!��A�|[2i���K�6�J�:>{��|�Iz��'��䇠4�앀p���+>f>g�t��;����؄+}�� ��lB\���-���GlW�&Wȁ�Y�AN�#' wR,�)�C�>#�f��r[Eu}q�I.���꨾��2��	��=�/U���}>��U"���q����nnId`3���:���˷���7���s�8fO_9�l%e���8��� �u�{�B�l������8yr�v��.sg���(=;},o]�}���-c�%tk��x98�����ϩb�=5#h�}��5��Mw�{(�
�D�I�E�}��B)�����աԆ�Grh{�Z�}�j�5�]� \?PT��0��l���4��L��'۽<b(~̇u̇��4Ѯ�1ya�s�$�䮷5R�}L[4�Y��du]�u}�d�7I�L#�RJ\�G����E|�rO�Q�_v
X�%����[B�p_�>�s��iź#�F�O�g�	��?�r^R�c�z�D�P�V�Wu�@�g��?��*P�J)�a(:wK�ym�(��뻫4���h�[�@_�xi��Ý� �$�Ǒ��k	�8�3�@�C���U?j�7�E����^��L�D{��(IGE�C�I��a7WJ4O~��t��bǛ;��wv_-���4��\��`�ݖ�:Te�g����sM�'	�'2M B=�mm��M*��iӫ^/��:��o�*���~��n��5;�,�Ck1_kS:	�[*��dh��g��`Ó�GV�X�\ �<�E|F�j�P5[�ƅh`�4��$;↡�L$�,S;��Oӕ��v���������j�n���L��i�7����\����l�8s�p����N:��Ǐ����N:��q@��� c�k{�ۛt�����n���%(k|[jW=�p)PVۮ���)���1�I0�;�'O��g���Ps\��i�{ ���vA?���$%+�s��/ׁv�G�:����o���W��u�V�����#�u��T���^ג7��c<ApbC�	���w��*hD v�Ӂeړ|�}�,�:��\y_����В*av�dA*[�Pr ��CZ�*��D��������s3z��-��I ���.sA�g0���"��T����<7��GOғ�Z��Ez��T�ڽ` H�G���Z�Q�r	@eb�U����Շ*Or����:�kϕT%loZ��(n�1�9v=�hp�K���&�=�(Ў�����.�_�B"���^ �T�����KByk	�t����	��,}Q�lW���y�\� �G�,/π]��g�U����>���٠u�����s�N�.�V������}νa�Z�<6�{���PcI|�{�gIp�1��@�~0��m�G��pV) ֮�EВ.	siڲ*S%]��e�  ���6t���X�!�
�����\Yu	��p��[�\{0(p�E�a�O�u̮�A+�Mg�X�N�+bKB-�Z��x%1� ��u���l�:d�sU�M���l��)b��Y���G�U?	z�u{�/�ޛ���i���b�7vN�������N�nbӔ.�J����R�zsM�&�[��n����@)z��ł�b����2|��}�XZW�;!T{�[��������7H9{��C�oU�R.�F%�y�����?t�h�Pˢ�̿�ʐfl|����ȃ�����Ӝs`���W>�Y��,�b>�s̴�J3n��������V�޺έ�7�5��nʴ;�]˸?�J��'O���g�����trb�ww���Y��Ƨ˔nI|��7��o��ާ��m ��ve�W��~0��?ÿta�lm��X9��^w�v+6����!-%��z�p*\��B.BϞ?Oϟ�k��LhS�?F	q��� $ ��bm��d��)2H��Yɫ�LQ6��A�E�Cm\ܕ�|��勶)UWOM��
����*�'���K�{�]�~i�KjQJV���}�'U1��Xo�æ�J��~��4�,Ɩ�e_d����ڒ�8T�8�qjZ/�
����nE�V./�ߨ��]��V%�)��GO��_|�I:==��L��S�nو�D����V�"F��>��j�N�z���B��;�X% ��)�ñ���[F���Mݼ���GV1"�����tu}&�D�a*��A����)��Y�ME�:Q��g� �'�E a�)��b�������wlc ��L�h#�d�mT��on��V4ma�%K�Ğ�u�K��̘CiD@JKHI���g�X򩃨��2�qR���B����
�0��K�4k6gȉJ,�DE��Ų�JI�*���%�:p��ܘF�J�*7�3Way~��+��{�����k��
���ƍ��ʲ�k��-uJKɫr�YвtV�s�x���(zT�	��.q�dJ���N3'>Flt,j��w�i��N���g��$m��̂�)�l+f�^���
݇-�;;�vGv��5���F�&��X@�F����L�=�$B�y%�69�i�����2�2�ʹ����˿I;���������~i��A�zѷEdpPl%�I�h{O���G���O�Ԥx�U١p�X�E �F�ߠ�����B�Ꝧ�u������,�*�o��Vsi?k�b�`�0�>z��]^�0�^�`Ti�'�*�U��cʓ�sZ�G����p"�vc��e�����1Xϵ(S� Hc��ާ�����Hc����8}��qz�ᓴ�o7}g�vwhu�!�������6]��H/�y����Ez��,]_ݥ��*ݭ <VCz��J��~lTD�a�,���=N{V��X�-4"�����o�w��"�	�aZ�;�⏂�Z��M�P���h�G��Q�<H�Y(ì@��-�ni�'W�s�t��N� ��@Σ.vz|��?R��T6�#
:h�P����P-<��@�ݿ=�'���,�f6�8Q2���
8�BX���ǳ���! h4V�n�#H'))� U3R�ן�E����s�:�#Xռ�Ls�Y�x��R���3�eqOmQ�l�v۲����v<U�ϕʉ�;߻��쀾�I���{�s��>ɲ��7Լ�n�:������)�󃎠X����߽t	YP���qO�� &��^��+����"ߏ�V%�4G {;e6.7�#iqn�Pcֆ�t�+��5�Me{�n���)f�'@�RuUd�X�i�]9-M�8���C�V�w�nOr|�J����wI쀖H-%���L�:�Jn?Q�y��*NeH���'�����T9?\3���'�'\Ԛ�w��`�Y�9-�JLpk
�6��6�� n�֚K)�5g%P-�ܪC\H]�Bҟ�FB������{��S��Q�f�+OX]RB'�6<�֪7v�V�R�j}��/Ա�-�؁?p]�(�,纂�`ܳ��wPET -�0�4�KO�D�n܇{��Q��|�n�lO��vV`0�o�e�-ڪ�z�(���I]�6:0�ҫo����L9m���b�:�E[����m�0��ߤ������f��חgi��e��hV%g���J�eɳ�. ����ٞ�}�X���Tvw��l�#)������\�I*M=  o��8�
�C��NyH.����9�m�!l����q�_�4��
%	���G���.o5��]˖ТIb�?� �m��!�gt3�;�O�;A��R�Y۵�[Bp��<���Mz�������[Kn�`�(T�2D�����q9�T(iac�ǅ�m�׷w�u�n��R4Slҫ��t}~�n���ZO��Z������9��3�������_V�ILe!����½sMy8��8���f��&Fm*)4e]�AF���;>:N?�P3P�͗�W⌓���>�̺'�L#�}�k������������Gif����&}��;mzYY������U��
�O/�}9(4�/�����R�nk������L�����j��Uֿ�"ñt�����JN�LT6`!-����[�a.��,����+o��V��3s=��m�nN�6>Y=�'��ڽ~H ��F(i�;+q�/N��(Wj�r �
�q�� A��w�	E4�ǥ��� n�����Us�Z�3-�W�Mx�+N����eWiI;���{W�xru6��!�0�D�U��1ʮ�[��tjgM@CO�ˠʥ�[��k��r���6����D�N[Y��i��P�x��{��_��?E�%�=�wh���HL���j�#/�c�;O���u!{ۨe��s��~�9��.� �E穊R8�V�	�<��N���_T��.#y�<P�5^�Q-�(�b�k��޽��[�=R������+ݖ�^�fL�#�]�V�DYE�Y�wO��W���[��Ϟ�>�����Ox�� ��Q����"�/�R��ǇGB�Z����s�� T���b���]��& ��{���+�;�.&�7E��C�C���2�^ڱ�x~�,���Q�L��흃<�'kӐ	z��΂�D���+���v�Owd�.�%|O�N��vP^۟7	ۄ�q�*�])͜<�
k{�z㾂o�j���wo�������cz��K�~�Ց^A��;�vq��� �:�Cvu|=}��*�qٵ���*P������̪��t��>��=����t���ٵ}��)����U�Ӆ��v0��ּ� L]��g5Ңn�/��'�0T<P%u47� � �Ȃ0V�|!5	{�z�B�*{r�v��
�$`O���?���G�}�6����7�_��i~�M���!�OCO������%�� �B k&g���f���/�j�z��8�;�:��[G�r�<� dV_�N���~`�����B��v���f݁bR�r�:f�{|t�����A�"[h����Ks��f�Ve�mˋ�!ߛ,���w�����R��p4�*�v�Y���P�Ď�ġ�<@��9�*~+w����$��ȓB�܀���"悅������HJd�!9TG����+G_OEXe�o��J�U�;�Uц���"�;��E˝u��0#�v��`Y�_^*P�	A�NG���4!��d��Hb2Xͥ|��:4�$d�;~B�V~]S�/A�}Ѯ>0�h"�1w�"��,ٛ�i���ѯh2�?f�J��_/ј�[IIYv�;V�-R��֓G�4Vʞkĸq˪�a��d{���<�+��P�eu�^��v�2�.��q�2�3傁����=�-T6{��9��'Y�)Λ���b�w�_?ZWM�S�0�1KfӴ��Պ���)��g��>�Ԫ�;�N[��	�X8/�Ѹn$�ѵ��ܫ'�G�RES��t���ic�מoa��qa��mZ,dT�B�G��}�Ɯl�s3w��ݾ���-�
9�Xv��hs�{;��Z�aZ���-��H�����% �A��������x7=~r�,Ck)�JN�!-�߽}�ξ�!���������j��.��o��&agW�r�؇W�� �V�7�����s ٷ�\®��H�%z o��Y�������*o*�T�v��.n���~����>88I�<Q[��7J���;���y�*]Mo�B�P��z$���U��Ъ�:d�b�EX|i�遮�^�Z���S���m�h�,-8IN18߹E%n1�J�n'�G���>d�|p��B�d'��H�
)2���Fy�o�?<8���`{W�
�5��Nn�_::U+JS(�}��ג�$�l�F�6�����!���j�g�Yv�u8���&�W�g�SNT�<ߩ�����x���Ik�c�G�� �j��C�a��u�ܶv��B���#��������~��4��YwJ] S�g�^����~/��$'%J��(C)�籬)��s͏���sDɸ��r��z��!�~큫߳R�?t�6�#��:yW�����&�qG���� m� ���=��W�z����`�͸wK�����?���)����Q����^��u��R��q�B�~kԵ{ݏ����tM:>�F<�46)(���޸D�TH�%]��{*�Q��et5K�����:��I��q)at�Zd�cB�d�?w�J{m�24?������Ǔ�%�=;����Kk[w���Xܮ+�L��;*��~�?�G]B�k ��:�9� ���B��b�3���W��Rf���?+/Z;�����$��U��2�Y�ju���!AK�9+��#����� |���A��V&%ZKO�ע���V�">�Y� �Z����$�]�8�u
�'�L�Rƿ^I��v�݇ZJ\�,�P��*lՂ&�Z�ʅ�ygϽ����ݭ�U*�n��0��K�Тc��i�݋�������^�����;{}��F{�9��`+ 	��m��h��]܄j����0�K4v?�:�Mg�Zoդ�RϦ+{�UsJ+p����j�>?}����_�FA(����G���Gi��ߥo�����oP�cJ[(x�~f���d�3`.D���iA���ޤG�,��{2�h����1efUe�Y�fsC������pC�pA�h W�^pI�$��:�YY�{�ln���"�߹��ZdsQ@�&,���LU��{w<��lx6UPֱ�)��v,�ەӕ�h�6����9��c���j��*�V��zED�K�Q#^8�;���������G�/���38w8��wG�*��2�@lvZH;�2�O�?I�N��T��4�����N-�3��.�%{����T!ݷ��,F���%�"�C�b{��@���u���ۃ#��{G����^/_�F�It�;v�f�6t��:1�o�h�YZ5���w6���3q~�B "�9����=Pթ�H�b\�����=�J}�u8c���֜dC)#ܫ#sK��	=�����x+wu�,�:��{�y	9�v�b�h��W��Y4~"JЍs��r;: >),E�W�J�s�����}��=ʙ��ߺR�N�n88��ө�:���OH�O�YV0#�c&;�S�ϕ���Y*9�&�u-!�^ �n�a[2p��;�P��C���b��|�׮�im$z�/��W�e��n���.�)����-~EJ�_xe
GhpI�Z@����tbw9ǩ�����Au�i�#�Җ+a�XƑ�7r���`o(��z���hTi�w�n�u,��� �����
w��+�j����(�UZi\na���H���4��������YN�,zӪ�_1�d�rP�!l՟�$%��W*�8��Q, ��d�8̑��(A4�+�E�l��rn?kN�|��R[s��+�������Ekc(01h"(��1��\^�H��T����Pg���.}�IK�llӖ���\�ڜ�NZ�{��x͡Y6�%��@@�t3QY���<���������}�:]�]�f�C����l���2H���U+!�5��ި'��^��7�@`v1׈}��f P�do��'���č�r�vۥ��`�l?����7_�E��Ͼ��n_�2�у#��k�YJ�� �ױ]�t�7��_�Ȓ�����Q.�]s��wD<��}�3Ƒ���`$)U��ɂ���Q<��R�؞=s�̐;�pٕ����\b�kC��֥��\آ��/�2���̡��9�Е�pXu�Qd0��uA$c�5��y���H=i��[�
u���`��Tzb��YPJ��pj���+�*��6[�M�^�XuBtw�<�|k�u߲�	��yܘE��e�ʘq�� �!��x0��Z�A��!=�ss}s�F���)I�#�������f^���#�-�ѢI�=���mV,i��
���:�C�ȓ���G����ޭ���pN�R�S��!:O�*@���g0Ҵ*��Pu�:�65�.ef7�Ugx3/7Z�p[k\Ezȕ�|��J���s!,~�R0k�4Hv�����FN�3��c�R外���^�
�{�x�=z�>y�Dr��O���:�i�5�^k�b+�.���db�0�����(�K�,z�Y}�(�$]n+��t=r����c�˘�Ȝ�1��d�:�~nk��#5+�fT#69��=WB?��2�ҁ��%y&� ���`v�fa�"�J[�"6l�"����:�Yt@�"�`Ϊ�͂�g�{��j�ivS{��q�;������ݼ_\��eIK���&F��ʀ[��B�gY`�n�Eg,}>"F��Y~�`wY81A)�q���91��v�Y\�wu�^Yƹ���eh�K���:]L�͹oҞE�=�}�<c��aPyz�@�f�w9XC��{i#'�_�&��������3�Ŭ�!��,h�*�4���&���1���+��('������Ʌe�ש�n����?	tun�py������a:����݃��*9a���|�N>�j�^\�(���6�玕%Å�j�v��6���	��~�o��_|�E������
z8�B!�QB��/-c��ߘS�_�����7�G��ѫ���+饁���zAK�B�Ly�`gOz�d�88 W ߠ��A�����1��#'�`�$#9�{c�6��20Sz�E�$ ��a ��Q��g�#o0[Y��	�ʌ�(QR�n��L)����je���F��F���5pg&]jx���=��se����2�"��M��#C"JE=t���}��V., �{T���۞%���j)��� �"���]��Bp��d}s���_�_��W��.;�D��9@�q5�l|F�B���Sy��F�zN:��٩4^΅��n^���-�C0Ȑ[��[�@�h���6�\����\�y�=;U@4/*ȏ��r#3�TP��?N�8Ȃ�w��G�̎dR��ŉ���N`���#�gW�H,���W�]�Y�]�q�C�e�í`��:��az �����j5��̮���6�P�2�c�p2w�鹂P�ш��X�W�=k�F�*},d�e���:����ή�C����-�{�ZI�ĥ�(T���un��?��@w�9�u��d{�%0���&�6����V��Tu��;c���?h=<иӮ����Ƕs�x?��ck���'��,'��sps���������(�(���J�ήn�2�3�c W󵢡Z���ڸ�U+�vᚥ=���-��ۢ�-������=P_�>\s���A�ަd��60�@��6õo&��G���=��k�A��z�3�T�����{���O-s@ǗL��+�f�&�o�� IZ�K�\]Y�l_�ʠ@\�:w�{�G������!�`T�C����J$�m�`lRO�6�M�?����K1wM��ZIͩ��cF bq���o�A:^zI0�Dṵ�3����_�_��eV��/�Od�eїS�@F�ϟ<S����Ԝ��H�kXpڶ-�(d"Z�Vr�1������JV��|@9��2���`����\�Dׁ��u����L��� 0B��L�h"�1h:K�'������ZUz���1'ȿS2�y6@��鸝
Pد��0Ӡ�cx�o�罼ް�/g��$Ve����P�q#.�<�M��`)T=�L��]�&!r��u�م\Uv���:�Rpm�;Zʙh>���
�E�\
fv]dՏ?y"L��_wFi���pz�����P��}[�t2"g����}��9��:��n旑�]f}r͒���*V�p$�T]> @bTs��"$S��n2 +�7�4�Y���g�j���������~���{y�z����V&�����؞6ݙh�M��#�ء�۾�>���Q�>�ǟY�G��:�n ����y������(1:'��=�=e�Ͷ'��/U�Ы��M���ߖ?<uY��)*�� �Q�N�	G;�o�|V�3�f�6�L5�uoV�#y=�3�;�%ߙϢ#���h[<����%.S����`+��I[�+��o7����~�4���gN��M��Ʉ-�]�WgkJo@. �y��m�2�#��f�tܒiNS=Y$�S�f�ƃqj7�D��8\'8���G�r�D��O������ˆO�D@�<�Qې��Pj��?����?6���Q�5ú�zWo�s�J��8���-��&'��ۓt{r���4
%���9�f�E��$��3�}�s��w 7􃴇&�9c@N���X��6��Ӟ�O��"=}�Lt�cʓ�4��:_N՟�4����3�f����w`�P�+R
:�BzUNi�X{�@v�|�<z����/��O�I��/��;�qݤ���HЇ�:����&}�٧�����U�?�����\� i9����� �@RP_�Ҟ����s��sk��GeS�����J�d����M��p�=�� ܨj����Q���U�ә�tc�1�v@�� w+����,]|<M_��b'[�3A @迠�C{xx G24�F������=9���ҋ��0;��R�E���x�}��R�ɢ�~�T�B����/͙}�씹o�=%g�$���=�p}��s��~������[��1z��R�
��x��22�A'v�g�������/��n1M��h[�������1h��t�߽�^U�O?�,�v�Ƈtg<��=�0	CI�Y���ن .��nׅ3��<V�u�*~d,	���;tF���δv�R!�E*nϾV@[�U�@T�8�&H,�,���0�A�с��]���{�|߲8exH�I!h�}L��8a��[{���*�����y��o�ԋi�Θ�k�	PT&�\�snA��zV�^6`O���͔��]=��3N�,9B��./��}�M��g��lӶ��_[E�qG��(�����tG��x�ۘ:�X~V�L/��H���
����ގ�,f
�q�s���߱h1��
�P8�6��w�J9^���%���*x{�S9�̽�>���Ev�W�� �-F�J�M�0�-`��bҝQ��S�����(f�Q�^��U5�Lز/����P;ˀ���ض���C�Y�^��P��͏r3��%�ҙL�����(���\-�)\O������?L��7����9��s#F�a=4�����B�W�Frp�y�J�\x��0}��ߧw/_�����{�C������f����`�}*�lc�j\�39���(���V��d�1�/�?M�|�<� �;L}?"�l��σG��N�w߽M�~�6��BQ���Ŏ��_B���`Ha�Y	�j�(��s���������e�8h� �ߗ�tJ�ܬ�eM�ѯ�RF�~x�V�7�	u�n�09�ѡ�8բ�ꊌ�t�z2w�^d�d\�F1vq��QpZ��8�e��Hy�G��}�wЙ��B�qm��v�a���FY�b���23} ci�����8�7��H��Yn��������>��g��知g�?p�}
�3�� �NP�8fڼћ�,J˂*��3S���7_�����w/_�j��w�����B˕���˟=��㥴9G`9���/m��������޾9����Ϟ���Ŝ����c��O�=M��_��n'm�� �,a߲@( a!��C��5��>v�\͎Wv�(k�Dx�H\@2dbA���:eИD��w�`�Q &�WϳDZT�A�T�6!�P�xI�E��o��>�Nﲽ3Ǜ%T3�1���~UT;�$� +��S�K�4/��t��/^�y\Ɂd���_oS���@�:�	y=��P~ݭdgݍ5�M׵;�����$"ɒ���&;hi7�K魢�vX�V����>�']f{�A��u�����9r��2@W)E�7eA�����#Ӎ����]��*?.?gg|7K��^�~6��ν�u��.���Ẏ�4��}��@��� �ٹ�&ŝ璱U ���^��&�	���W�۞E~#�o���|`/1':�k������ߛ��)�j�}Jon�RO&��eN����(G�y'$
9 ��@��̵&}N��fuo����>X�y+Y@z��dlv3�k�R�,���辄O*Csb��ߧ��^��o�.����t��+�Ɣ9g�"t�v/xE!�چ_�x7Ʀmz��K۰��)w��ݵ�~��Qڻ�>���ز���C���]\���o���,�}''���*��#`?�sCq�z��Ԑ\�	.����Q ����<�໎�n,��x�6��w}��P��	ӿ�숳E�͹��"��/�p�sdk�Oo�W4!�%��s h��䥡6��E�:��	�|Y��*��*��ld ��什�]����Z�r����������Azo����e����p�v �s8�6#"U�� �o��ݍp(̦3e�#�p(ہ:�������!��ߎv�bWs��@�j�q�ފ��1�dǰ`���:ؗ����Ǵ0G����SϜ���G�,7Ǩl%�Ѯ�@>������ڲ�����=%��ʊ���X��A�y	nj�׭>�r��A�I[3�GHl3��
y�ɬvn��Ց��k��e\���E&�	܌���y�VKw��#�SdbYW�
�2N� ,Ix})2������I��d3}�����d�,a�~<��j�e�f+3��R�?+'���u��|�L8o�Y�u��b
k�߳U8ɞ�UE{E�FD����&2a�j"�,���v�����vn==g�?e�)���(��k���<=����������Gi`�c���3)�/<}���)%�Z�����x�l�~��6��,����|>�u�]��JHTeo�_�\����|v�iL�E�}L�,�pIU���"`��9z�Zpg����F��ʹ����Y��L,SǇ�_��������QZ,no';��� զ�;ܵhg�2���1�lf�m�j�S�uEGS�b�*����;3�1�N�����d�2e[��q��pm̠�xc�fc�g�6Fo���y�0��X�8y�!��?H�ތ̻�o��������1?�{/ɿA[k�6�}K�ϭ��5��ڌs΄��p@4�轶�6t<�'�?KO��4�{|����-C�Ӧ�}y���}H_���O�����?|��/�0�#{���`�@QWޮ�!�Lrf���c���G�=w��aA�A�������͑�$����޷l�7�7��g�,����Mzp�a���ӕ��Uy��,` ���ʓ�3h�1�M��E��V�+n�/�2�ABw�� �>%��]�Ke�q2�#ڱ=Bf��w����B�N>x�������a���,�Ҝ+��0�H%)9�@�O�\�@
#�~e��7��,��N���;rm�j��fD	�_P�R*�C�.;��|���h��Uz�.y�F�kƟjG��]_	�Μ�ۗ����yz����Am��u!HR�I�T>�5��W )��B����s�`�]^��oΜ3{B� w���K���S��H�����S{&'u�j�\u�"ƋJO�6?����-�T.G�=�����Z&eE��,-og
��JW�����(q�s�(S��X퐯w@Q)uWAu���r���5�ke��w�F���]V���g��.�R&��&3��e6�����yvZ[��*�6��y_֑�>�U�l�ȩYC,���n<X�F{#�,2P�������T�o�����c����jS�����ҥ ��=��{��&���	ב���V����+�N!I%!m�n-�w���$�c��\�|L���D�����_w�#�|Ǹ�Ֆ���{��r��*��❞}G&��Joi����r�9�ۘm~��z�&�{E�Yi�*��$ݮ
�ؑ��JQ-�5?(~|���!��^C$`���t)�Z�(e��ŹJ�{v�����4[ߤj5�e��V\�-ЕeM�������ٰ��������ͫ�ތ����e�� <�To�,��8��D��$S�����Q�����/����>J�����^�`5B���im������|�Cz��1u��4��-��o̱��=�ü�hkǲ���x=I@e4wv���ޡ2��7L7�O�!���h_i�	��JB0NQRCp���؜ N�ܥ�g�����������ܞ3�bGi<Ļ+�-�WuN��2����tߜ&���i�{�ae����/,AB�"�<J�Q�����^��S��������R�̮3}Q,�>2'[y��ޣE�q���H�5Hz��k{��=��]{^0�h��L��Ҳ���D9�A79J�ߩ��$k�w^z6E�E;d�X�p��(�����*2��ߦwoމ�_�=c�i2+@gD�c2yw���p�\W���?y�>y��2�t��D"��L��2�~ y,S4}�`�W��gz�ひb�E�S�� O��nA
��֌~��J�0�������xw?=~�XY{K�Μ0*g�{�	�n�l��}�ֶ^��s�ṂSZ�k8#�˨)T�Yh��3�fˊE��j��Yz/K�4�_�S�ց�`�5P_�>=�O��I���3�3���N�������lb�H�H�=t֭ �i<��ћ�H��g��'VB {T:�L��M�fF��A�*,Q�i}�ׯ����3�*��"i{C��m0L�0J��u<HR(#��]�X5I�X� '{��� ����8��Ɓa������c_*�r?�^�'gm7[6A�g��G@$9�z�T� ������u��Ѩ���0�m2�Z|wZ~��۱y��O��?�	_��y�&�]%�s�;�v;�gp?z� q �, !A1� J(M�5���62���0;fF���=�i�D�ٹTfv��=�,f�>���Ň�Ԙ1����7� ��E���޲�w����$]]���	J�M��@[��v�/���qh�`�1���j���/��/�����Gi|o��I8_���w���"]�=M�^���ٛS��EfBy�Nxa_��q��C��i�df���!�����>�3'���f��R���<8�N�#jI���d��Q��z����g�ʈ98ȽQ���u��_�Helk�lSdP�C�YC��Q%��4�d����?=hթ��_�O���>cT}���=|�����W��,�##��6ٜ�|���\*O2����3�����%{��kʾ/%-i{���������� kȖm��	�%m��Rv�{_{Y��Ih
1p�.wIɻ��G\[�yn�:ҷ��]4�5����5eT����J���]Y��r��!��@��f����ˆ�1#N���+9�j�&6��)���T>ND0�`:JL �v��m��y�՛���`�jNT�(�3����\m�c�k��?zdϫ�X�k�g�{d.�o�ԂG���@���FT E�؊�-l�r��<��Ѿj����F2�nP32���lcT"@I�,h�YP�`](�C���֕kW+���i�r�9�s��؜�v�)���رu���-"�
��H��G èGۉ��@?����z�����܄`B�U���y�L������5΁h%T c]��ށ�s�n;����K`��ޡ�0 	}��.E����.�({�`HkM��<�xi��!i�B��z�>�Ys��&�7�?��a��wC֟<+�Řʨ˪��y`{y�~����V.��|1/A�B,?�\�Ҟer���,��1/�ke���C��B=�u��gXDLj����Ԩ�D�?q�>HJfȉHS�:�������w���O��0�ڳ<c���<���2�����\�^��7��,�e]ƨ� �w+�
������'��˿�E��/>O����TZ����#�-㞟���7'�������ߧ�녜o���j�~nO�G�L&���޸/�0���K��vB;�TF�Ӥ쿼��L��ft��0�m���S�c."�p0ZƔ,?|<Q�����F}�woߊ|��+jQh"�1�3{��B��2FU4oG:J���@��� nG{�*%b����g��w���Rs����2��A��^?R9GM���p�W*Je`���?:<�SB�=�\"F�4�,���ýc�B(���������C�XɱҧjD�����S�R,��Sgn\f����^�E�UY[-{��`�(]�5ã͜��Ѯ>���[����U�����d"�����W�o��G�X�y��F�P�{��@��E��3�d!XOw8=�*i��g�e�c�q���7|�M[�ȱt +�`KMI���ɳ���C[ӕ��6�q�	_�~�����|(�-�����b��K�O�����yn��1���W�)5��*Xk�{�U4��) n���O�.��`��
 *�#���3O��G��lJ��D���\9%c�yc���5")i�� i[�|9�Z�{��|�]Y�x^&��{�&�5��TT�v�@I[���e��.Dq��7\T!�w�	�GY��{����ܗ���%~+4� �Ψ��̾߬T-�K	�_wG�2S������1��f��ߗ����3n�y�q|Y*_�,؇���Er�A�r�� �?�wOHֻi��<N���M��I���D��N��p��-���"�
��G?�008!vw��rN�B�!?� �(#�*#U�͔��̘����^LJg�ަڌ��2O�`�Z��g����2*�_ͮ]�X��}ў��]�06�`P�5��ož��7�LF��{���{��O��_<�L}��4��_yY����,��y�����Y��1�ϧ��]X�b�6�lوx�`��Pn[/E�0��()l����H{o(4/���?�"��T!���gfP8��¨�ތI����~��B�.So�T����ZH^;�Hg��,'�9���}�7�x\yn�G��ɵ��nb�BQ�ʥzÈo|��H��uH��/�*������gi�������i��,ҫ�o���˗/�?��.-C����R�27�X�g4�u!F$������@ٚJsW��9�ɍ�@�7d�YW�ݛ�K��)�4������@c��Ӷ�~�P�(I
��(��r�C���1Y�d�N�9�z�e��}0[\z����(�g"V�r��*�[�K��)�q�L�,����A�`��`f�B �/p�=�^�g��p��fJ��d��0��c����B�۩�Sš��^����o�Np�G� ��y`�5l�\25X�����,@AT���L��z��m �ե$�xǑ�џ�]f5*�뺺#n���<g}Ĉ߃GilAc��/0���x/�AY@���B��J%��v���l۔�zD��
vr�ڻ��k���W����_9I���;�
��ĳ	��7�2n=����4�6����=PzI<�U�i�sR�F�:s»#�}im
e�U���n��6ۏ�K�	�}o�H���X�&S{z�
}W����rzݱ�I�������[�y+�� �9�{h����i�\?ϝ�-R��L��Fޜ �-=4(6}�C���O��x�v����-ǌ�1�i� v,����-�ihv�vE��Έ�S3֫t���As1s4������զ���X6�Z���p�˛˫4�����Ej�.�ʾ��ޘac���ReE@c��Xfu�N,>��Q�SU
���ϐq`9��'=$������	R��kS�3`�,����`3G69o��e�˙6,h؋w'iI���is3O�t�vʑʑ"ఏ���(�R���'BG1�
1܋��\m�F��Zu=�wf;�����aDA=E3gvoQ(],"G�d�d��[�?X��9��b��/�����E��쉭�N {VB�沨k62,�Ԇ���2����]�}��"����W��5|pd���в�&���7��7�4:��/<ϽC]?�ۼ���Ȭ�*��Md�^�?� ��������̐b
�h��LԦ��rcY(��
A	�fl�a8i��L�o2�y^�f !D�@J�h�����֣򠃒i�ڌM�c�ږ��:�i5����R� ��e�R)� ��R{n��N&�����^����F>�e_ � ^QQ�u��i�^�w��*h�ch�|�>� R�h
�+=w~ґRlQe�F��֜�R��[��m}A��1Me�`����Rlq�L��|nA��#7�5� 8ۏ������]1Epz�f�E�	=�s�����:�Z�{��]ẽk�ft��c�qIo)��i>�5�ʤ���8���ޞb"u�o��ƙ�؋Ȭ���uJ.�[٧�H�rK���W�B���Ȯh��:�P쇭���%e���;	�vo����c\��~�2�=#��[���W���(�J*�o\������1L+�l�s��6�Қ����@K ��U���3j��J\mZ;	tl���5U��|�*��K{F�0G�ts�(���q7�������)7�Ғ�s��^����$�=�#K�S��N.�zT�\��q'�6�A>��o{1u�R�l��yz�kt���#� c�:��"��f�ʅ����hpc�B��D�j�W�h��Q�����?�w�S�p�Y� S/�G��ۃ��/	�Y������ߧ3s�g���q�v��F��?8�x�� �%CS(+j{�����^����~��_#k���Jeę9Cp9[�G;H#����1�8�a�m.8]/o@���E�v�0�8�#s���ӓ��c����i:?��4��sp%4�0 2es�Hy��f���7f07�o�eK���Js������^!��7�k�b1fQ���v8+����B�P���ze��c�o���}���WZ����Wi��q��Н�\�o�	�!`M���$���[}�� �'�HI탵��&V1��|��CFx%�z�irq%�-�a5��k�N,0������ ����I ���kϨUwtmG�FV��&D;c�Si���3KE�#C����E	���hRj$���{�8i���̛�;�@�{y�T�����A��g<*P��5�C�akެ�:m�z+������Z����;ʆ]z/&b�H3�u#�[�eY�߻2�R,z��^_�	�����E�;JQlp`$9X�v{{��~��Zi*  J���%��ҏ2a��lT���2�(-�E&�*��V��C
�}�z�},�W�cTT12w����u��w=#�q�r�һ8�c,'g�9P�Ylv�~}���/�Y�+���̝��28������\/�M�$KZ��H�@�y�S��;1�5]0�~h��������l�+Wi��S;a�
�`�����5ќx�(�����jiY�w`�L�gA)����v�.H�Ђ�~^z֨]�h�%�&M��^���!�5TB�
���q�<2��b�2C�i�?O&l�@���|G� �-FA��X�3����P����kQu�n��5E��,�?*��)p���S����)OU�3|5m\3@��\]\j��/�M�ӌ$�B�V�έ]�'M^���7X:�g��"&ߌ3��������]��5w�wl\���,�E�Cѥy��L뚬#O	�2�'�~�������r��A�oN�($g��tbY�(O�������_�4D��o���DiӜ[9<�-&�"q\��:��Fpy�f�qfp�#Q }��� d�N*sJ��m��>L���U�r�f������'m���2����ؽ�ꅞ�ei�?h���9��@g�T-�Y�x�J�{n����R���cS9��:�`8��Y�a�.�\ Dq�������3��cϓ'Od`nfv��t��W�e�T�j|6W=��L;�0h�֝�TU�L�e� ���3�&�]�M���ɝV٣g;����#{�YQ�ӵ�8LՍ}qH[�H���Rg�φ�#\�NU�Z�f�(Ȭ�]JF��"H��z�	P�@in�9��;9kRѺ!%�)����}@VQ�	�c��]8ӏz���2z���ص�_��~�e��!;��m��w�ɯ�iSV ���'�j��"o��1˞�1����u ��CA.QYU���:�h/D.\a�����O:�q-=��W���*f��]���[ם]l���,<��FW���G�	�Jr�+'SaT�{���J��P��hX{�q��j��7���k-�BZ��X�-P �Vߣ���G�2��M[ �Nn�;��
���4�7҈�d�Y��3z�c�OO�ʜ�e�δ�����fKҭ�'�l�u�Ӯ�w��*�>$A�~�M�j׃��6�?�%���';���m�������զbјIÙR��7��0���m��S�rdX�攭��}.��#��E�f�0���ƃ�RP�k(�Z<��d��j�/'>��׭eXҿ�6(]�p���o�u�)SW��{P������+�]g+�`[40'SQ`���v�!��4��g��P�-(�0eYu�`GD�{�����ã���ͫ�Z��\ڈ8 �y��Mz����e���jz$�&� �wx�q\d�d�+	�\G�:�^FP^����,O�D�{'��,�q�4���V�@^�stg�v�)�;�0�]��g�K�g���2�����0S�@2�����r�����u(��ɬ�d,7�d�`�����zJ1�K(Bb �&�A��Ԛ�'ѻ� �&���W�]��=��{G�zD�����U���p��s̍_]��?��Ho�H��:,\��@ H����2�|s���sm2t?��2������\_=���<��q��@�A��>�1�l^OՄ��J=O���,�Ly,$2���9������;�^��=��юO#���̄=�x	7����P��a�1�Z�~�[g�����U��S#��c{y];0���Ν�]����kd]���펆�ݞ���ы�r�v��w7�7�9��6C�R}���	��n�
gr�E:�^!Ѽ�]��-�@=��y��1n�ݺI�0?���@>lK-�1o_�����@(��y�{*7��f�c\GZ��>�.�X*J��⬦�I���\��\2�.?�ai)�I��3f61�m_�>J?r4����������l�4��s�l��2k�7N�hWm�VcmI�ە��x&�E��E�,_ܸ�K-�ɦ2��lv13s��*\�Y�������	k1�%,O'Z�e0��϶N{0D�a�ƍxXUV+f閞�4�E�,6�GDt�E��i41ԾR�k��l#�E3�϶υ_��O0��Bt�(�ƙVF�>�[S>�(��Ԛ,��ӏM�A�`WѦ�:!:}�
z86���-�UKQq2��=0c~`��
"f�J9�i�\��$���~�i��?����>O���a��M.��lj*]^��������ߦ߿J/~x�&�˾9[Ѕi|pd���J��;)�3�������ԉD,R�Ӻ�/@��'�)�{����0���i�#��T�x������i< Xcrd��n>�}L��\��+��\�4*��s���P��U9ej�ڜ��z�^��N�Ҕ�#b��V��՗
���2�/��o�j�.�-�����"~�����2$���g�8g�)KЅ�N��-��Ǵb� ԙ���������O�9Л#�؀����Sm�!#0*��4��2I��Lԙ� �!��v���rN�Y+0#��!����웲��Ⱦe�%��P�3T�̋�v	ə���	��ҾZU*�J�t�P8[��m��CƧv>���W�8]�:>��t��K(���t����l��n��z���W���<�*5�<W^&�Ve�6� ��Tw_[�:)��r�� ���y��(���q4�M�;"J��*��Y�щ7no&�,)B�%�M�x6���6��pK]b���|�`� �2;~t�/t�g�E[���B{*��/��b��oo޹�X �`@�=�q舲=�V;���D����Yd��P��.�3_|�yz��~�rr�ޟ}P��Dan��tA�}ފ��@נ=',���rv�����ղ�)�ބwa��ۮW�5U�N�J�2�]�?���3�h���?,{�~�"Rʤ�v�*�|��(���/�CBi����O�ԽN��G�J�CE)E�JR�5y ��R�P�1��63���2��2�92��q~h���C�ܦ�Zmӑ��&�$��M�?��N^����r����7d��q9��/j�q����� d��+�NO��nz������O���O�ѳ���O���{�.� Jfrq�.ߝ��/ߦ�~�>�>I��f$'" ����Q���{idka'K��)�j�*	v��C���1��bp���g��Xמ�;����]�\`�"���n7�H>���J�����L0��[yu�j��Am�e-��;#M_y�a�.ҥE�(���Y�ZwlE�?�ܦ�16�yiT�����P:��JB��y� ������3���������/5���ǻ�'� �-�f�BOXd�mP
nBUH{�ea� 7k��1����h��R�7�6[*�彆�]��LOGB�����X�8��:�/���)_(���l,=���@�ʌ�ƒz"����y�/��'�gE9W:[��P~�7��]���}[�A� Z��ь����y�WQ�X��!�i;��=�<�l5�+JP ZAa%t9��3/].W�4��L��He$s;�y;Z�˺|1j����^����)�挅���[�gF|��Ld���x|�?�iݕ��p.���k\kl��?��V$9�7�� f��_]�l'm(����LA���A�/f��T4Zz�>g�y�Y�C��%�dբ��pCSt�U�������X��uv�&y>��JH�����!p��b��

Q��FqR��fNՖ��	P�j��F�-Q����K4f��D%��TǋW?(8���o�s6�F{�������\v��T	��Z�T5�"QJ��E I���N82��U(1�p�=ZE ��+O` ,��'ё�H����Y�0�O�S��Um_=J��К"��[u�oEõ���{d͐{� �(Ɂ�%� [��TO�@<��Yb0�� l&����!���U:���-#7*SØD_@���5��{���J�7@ۗ��	���AnX�(��#F>�2zEDd��Ҳ��Qڻw��?��~�4�8>y��O�Eu���ί&���<����޼x�^}�*�{s�&��2��I옑�3ݷM�s�Jˆ���-r��;��yZ� D��@�ͮԂ� �ء��#�-�J�u���j�Ԫ,�A����Z��6�Y]�0=}-��
;]����:m���2ɞYS���%��ɲR����刻�3�*�&��8��hD��]�,����̻�|��aG�W�}��z潭{�8K3rj��y�Re��g�`2�П8ae��8���9!�Z���
�lo|:��-; ��7�h�u�"�$�;�\����R�S�q�d25C��Z�S�5\��qv�[i�2&_e�L0��ٲ=�k�5m�<��u ���8���� � ���)��ѱ�n�����e }s�3�0����}7	Po?y�r:�TJ@��۫�P�z���D�S`���V8�NN�{d�v9�3 �x>Ig�jY�`��:(z=w���O��Q5c<�`�	2z.a����9���~P}��y��3#y���)�b����t��m�����W���� ]���S%�"�]do�nj=��\���\7�3;�<7�U�B�4W�:���V���Ν�{�s6��\��^�X���L���n�����'��t#nX��a�c-��,᪖3Mb��������9-����u�ݠǯɘ,��=�'S�:	�X���XUW��t�����^��2$��,�dS�agT��[�����pz�oɳyrĕ�r�B_B�ƀm��ڴR�
�I����͵�J%d���灢#R��� �o�n��Cx�Ʋ�����wv5bA`/2� ��N�������L�R9�""یY���ޠ��~w��$}��_�g�x�|�IJ�f���e#lZ��S�t���e����?�I�/-�`�n��fwv0���G�y�U�X�e�X\[�O�������'�o��
�>�"���HFKtG���NAV����J�@=xi� l{��z����|�|/c��qg�C ���|a9Z�b��:8d�"Qq>,:��
�Ta
�B�U���1�V�Z�c�%,���gs��Z����}`P~x�.�띦K��!�>%��3�,~����xGG{槔� �u!s��������#��fv�՛E������ջ�ރ���<�Yõ�ѩA�Ч{���e���;N�řZe�1Ⱦ6^&�wpNs6 �L�t�%�I�L�'	}�� }��iKy=���h��R��\��z�D�N�9_�! �\��u65N왰��c2��*0]�	�&�RY����N��a���v�=K.�q��7�{]����x%��1\����;<����].s�~ �� A�Kh�qd�:����ϒ��!�(CC��{B��0[q y]*k�����t�Kh�������΃��K�U4"x�kyw}� �������Tkw¼����۳^Jp�g���i֡�S.���X����y.���"�H�+G���u\˕%�=�[a�s2Џߗg�8Z��a;"sY��[�5�z������m��� ^�A �x���V�虉Of��Z	[�@=��?)�yR������p�<�w/�,�Zϝϗ��xB����0��<���#����1�ѦUͽr�-�*]�z�[E��:�d�{x;Ĕ�F��%�d�p��j]�m�ׯ���H9�/���d��Q1R���!�+2���z	u���q��Ɉ��ね7"�}�$'|���˯>M�}�,=��Y�{l�lZ��,���F,F8ߓ�ߤ�w����v(-5�Z�;i���"�4��2t߲���wvO�[]����j$qp�2�B�7�����.��T�]���]D�9@D5 H1"Wu�؛'�r61g51��j�Q�9�b;�N���3�IK���(˰� +\�4�G�ל!>�֕|���h�,��B�uO#P�L!�t�{� 1��M�L3�g���}"��]�����2$�[g��!��F���M��ץsJI�p��^[u4���񅲉�g��G�_�Wo^w�ګ}�kFL3� a�v�s1��۳ ��O�+��@�*�t��" K |r9�
@�J �0,0��<p��<�м�M��>(s����L	x0D����ܩG����R	�����«KK�L'3m��$�����k������g����$���d�z����/7���,w�������![yӁi�3aGO�I�rds.�V�Q�C�bM�ˮ�犋0��NU���K����֕�f��'?�zVA9*�}Qv�+_�iس��X;_����2}�'ټ��o����q�>���u �̫IPH���=a>G6�>wr����=�_Pf����y��yr^�����uhv���گ��RU�k~U$]M`5��e=`Y�5t:��1>h�si��ū��g�#~ZzUc7z�����ˊ��������;��ή�Z���yw�%�(���8�[7��r<�0��=��*l$�~tC��"���JdV8d�}����cgi��� ̨/��似7|W/cӋY.	) !rp����!�M9���[I������L�|Ak�`���/��U�Ui�B�gl|�u��
V/���x� ;w�ۆ���-6i�V2��c��6|�0}e��g��Ѿ��L)8�R�������ߤ������@�gN�^-���#����M߀�5'|k����k��kttgi�j�p�x	�j�R�Y�<���Ă!X�2 ���l{��R�4P+��H��L)�*�b����^~�e&���!�Pc�<ku2K�O��z��h��N���|d�l�����@�U�	��+Rr���s<�w?�{�(���O��o��C�5`� �U��܎�L��Շf�HQ��R��� �Q��	j>��:�K�	PUF�R�3�K�0�Iլ
Y�RA�h�5�30�1j��6���w����>u>pШ)���Z��������Q�k�H�a̦��h$�t�޻�Ի|�y���(_s�����~�h�N�c�L�e.�{�����A���C����C�`T�v���hI�����ha?e�`�b���Q	�^} �x?��U��
΁����S>�q��;�r�{"J�t����F�QM[h�;X��p����^��]8k�9IaI9�ه��(��x���X���@�U~oG�IAV��Vq��(g��������W�jC6������<��g00���@��f)H��Q�\FQ��j���n�B�h�Mt}�5�:''�Im��������0>����탡�-U ����C�ە��4�X@����g�$X�4�����ɥhpm�){��Ʊ���̯*��˲�ty�O����y�hfvx��,�E�H�\~�F��C���%	9��q��ʔ(�p8镥�����!4�>�x+*��LLTp��4�ۦޚdޒ�M��U:�x��u:}�F%h/����#e_�6����-�o�-ՋbQv�"�v. �;D����!ޞi��BO�=I�}�L>�����N.g:�8�^�H���k�f�ROZǻG�Ҟ9�j� -!��%���<�.��/.��ĳ6��ٚ���i��4h��h��SXj��iˑ�� ��t�G���v5��A��aF.P��=��k��p�UL|έd�2�럒�w�vm������m�a��ؒ���� @ￃ�&��㰐9p�z��R��Q0ƃ8��dxvo]�y+��A�eF+�08PȍB�v����@{3��;#��(S��MLZ�����!���T� ���;�Q(n2efU� 9i�n�c<����O~������S!_SP��4׎���*;a�93�.��-X]��h?Fx��B���n���v+�Wn�Ǉ�.�`�n�L
���#(�@�g�Rld1S.f'��֩;���@D��e�۪ߕ��&u�~$gb�{�2�<�|������U=L�}/Se�S�e6q$�o<�,k���b٬��5���i�W�}�.2`ߴr�ō6�yz��2�rt<�^�x��ظj�� �ϳ�#^�����U�ApL���y>��b.��޹��Gz�j̥���ĝ�>�����Yy�m#u��%��0p�`�������t�UP�EF-��;y�H��*������:�҅0��I��Lv6�
!�yd6������z�_k���V�#�97M���:a��**�uu�]Sf��l�D!B�I@z�������'v�d'l���o���(�G,�f�H��G{�K6%>X�,�^^(�B<���=S'��4�Yo�d좘��c�X_�`�7��"m��|��5/5��D+i��6ҍ��nl#�  �Bgu�P��t�N/.���uIy�������N732�n 5���} 6&M�ADv׮}w�W�cB����̎"�0��A�~��+�9���X&��z̛�ע7�Lw��͐\�}�	�V��%t('{}ט]���
2���DP��Y�I�=S�h�twd�o\�������n����k�E�����,�J8�u�*���3N��	p���4n\�P��r��?fDw�U���O�sL>>��,!��<zO�t�Y*���<|�0��?�O!|��Yb�������e��}@���;"6����v��w�bTnѹ�ep���-wr�Yޓ�a��c���g����i��VxcY±���ɧO;���`�`4Dah��qµv���I�ý�Yi�(�T�2�W����@�^��-�Z%�M̀p�E|>�A�?@>�f2wF=�r\ �/!W�)C��MV%	8�Ֆ�R�7$1�˾���J�� �No4#�,���ѝ%��<�����[�k��)�rL+��.�~��3x��g�0��
�����ێ�t@:{���\f��3~�s^��s����m(ze��~82��2�(@0��)��:�r��Z��\�ЇnCब���c���f�7HE� ����8�h��hd����tC���P��Ɯ�՞�h�s[�e#@���_xk��4l"��@���A��j'n"x�_��E�*�m;�y��RcM����k�ef+b��(���	�Y
��B4M+$���P��cT{ �A��+	W�����$���2��2��>���<�E�X��>���C8���e%��G�Fh���\Ra�����O�d�\�VT�����Zgi�t]�y�I{�9-���Y�x�>M/�EWx��Q:��O�<��2���2�k�.�:  �0|U�?���W沄����<4-w�^D�of���:a2Գ��A֮g��l:�dg� �ӹ6�ph���q�H���6�Ԃ�+s���uz;���0�A	��Y�~(��K�����Y�>['��$UZws���F��e�9��R��ZF�7�Xf�"RTi����#uQչwXJ��ޯS���pu�B��)�=�Q.]�2kP�񴂧��s
��,����ZQs�%ߢ�P2��֨)?~�$����>��3�G4�% q�����F�GU�T��۾��������Hu'{Ɇc13�8F���'�{.�������sp�����`�X ���;R]���qL���q@���cl��O�A=E���l�r�P��8�޾Q�HAX��1^�"H�,9
Z��Hhv[�jWw�B;Gg1�5�T� �f��҈�w��z�Uٕl�O_�8�ܣ��lЕ�y6[!`�p�,*��b*LK|�f�$�^�5�����rr>�*8�W�g��	�A��c�3�
�nɮRY{�t6�w��GjҀ��v��"?O6n[�NF
�Z�pO���l���u���	�M?�]�������L�2e��g�H�I��P�WuZ'�*��Rxߜr8�`����c|�1�=�����3am�iM����xy?��i�.�1c  /����'����/M� E����C<#�Գ������u�O�q�`�;*�����V�A#��a�ߗ���p�:�'7V�Z�a{�?,0�S��<_5��.�Q\�CD���Z����!����ǏB�7v��@��A���8�|�T`=����y~~iQ�sH�阡,8�k�-\]���F�[z����ϐ��Jejܜ#`����˾#W1{鈾T
�|�F|!>�R$0_��wAvi��3�����2���D��̗j$��J��POk`�����txx��X$ψ���m:��x����%"�RbV[����8�	�X2���C�(/��ZǘH�������y�q�MR;u%�Fi���V_�p�Q�N����:j7�����(φ�P�rG�)Tى�є���^j��a�(�����xS���PJ*E>P���T*��i�/���쓧)S
�SW�2Y@7ZEyu�z����d$j��~8a���Ȁ�l�t3�@<�G#/����;̜b�G�b*?)�|5�t0I�����/�� �:~��Ș�>CYC[�tlD�,o��^}A�R�Ʌ�m"k�8�Z���H��W�3W���F\�K�M�_�
!U���>�[Z11�%S$ 4D�R`���9ud�ͦjM
�4�2����n�^o&W�rD{��i�ZU�J .�l8$�ـ	��Oa�W�Z��dv&R��BPi��9�_~�<rU<�[���A�F>~�vec�`��I�Q�}R$�+r0G��2�og��X(l9��:��x��_�QA�^�8�q��.���^���.��j�֓�����?svc]9k�����絁��ŝ\y;嵑���%���t�>�-�I^��V1�B�Ku��g|JB��7W&<w����W���j�52m��Ğ?v����]�J��*�x-��}l\��,��r�Vǝ��{�#��V���p M2p����z�7�?�������R��m*��.^}�#޻�Jd�`��l��4��lrJ�G�e�vvFi�;J���~�r��ܒ��5S� ��!�`n�'7�6PbV#1����#��=������k�W>�t~�rH{d}����Xգ���н��ފ�S���X�(Go,���{�#d�@+6�8��eTf�����o�Y�(���@�xzj�{���;����y�<[��<�]���R�*h�����;\�rhN�^�c��~vNP�V�l� �y�R�W)s�آ�E����+�Yu#4��^�,��B4�=i9��9��,�t���.E��"���KvϣRnh�vY=e���Բ�K�*��)K��l3�h'd򈎰a2Qf���Ud��)��n��6��W.�i�������G�J�1ّ�z���D�v����e3j'9�ǫ�t��Z�6��<�2li�6M���Ĩ �x��2�S�W�pE�f+^½�a�Ħ��!R���wo#�o��2p��՚�n�K��D�� �m=���#/:�f1�c��#6��+�l�ό^�@kG)~�e��;:8@Hyi�B��>:׋{R���k�ɫ���r�,�,���]-�E�쐰"� klr6��Q@�cj"��g.����>�$c`,\d��V����F/����ҵ���I=B��G�dA���s?҆^0�,���ޗ��2���(=g�x޳��xY�V�$\P����u7�-�G��={!���_�2Y��j֖��rKaنC��6�+ <�K_�t4t~f��x�l?lyGfg��"���&겛X��X�'	Һ�{NA4RfF���Q{�tv3����f��A����գ����oz�����ԟ��Ԗ��G�����f�ΑEk�^��2���BFjH2Df,Q�!�{)�,?��tog7�ȏ�z��l���qp��(G�@���
�|xp��-�E�'�YcT���z��*�eQJ�� �z�{	_/90ԭ���� 6*UZ�V�l�nў�2T�@#�#^�C�%�E���
�cv�����o-��[	34B��U�F^nf-Kw���mZ'&mc��rٸ�HU�]�2פ�(�S��F���B7�+s�#'�"�D�ʄ��J��QxD�)E7^�7j/�fi�쾉�p��H@U	B
��c�����G��)�Z�}�z�a���A>H޿�@B=������1�� m�Jd�J]d�p�6Q��r����	����3���� ��x��lN?s[��Ξ:��K�:�������D9��+��s�6v�7(;�fg;�����G#����\�"��(�z��%h�þ������ڱH��<��"#n�Z1�7ٰ�����f�8@\Rx��b� 1�����T>��0��x���mctD=�;�f<��͖$F��2/t��{ 7e�w�Ÿ́<WJȦ3�Z=��P�{�^u{_��t쁏[��_��%���N�w��" I�������[ttqn��[�d�8Z2S�$>1 ̇���c+n,����MG��j���({�+�`��3��]GU��	!Eh��~��g.�:�A�z��y���c�^��U��{��B�BF�ti|�����;ͺ�WGak#��Im���R�s;-�J�K8�W����\��˦��%*{eh	t#�Ag|�.��뱵gs��g{��w�u��/�����ӟ��.�vi�1�;�Ŷb�� ���M-e�6��(Q�X�#<������w�P�UGI`�����C���ig��&��鶲M<�Ų���4&sC0a�0��˴��(�v���T�M;����qk�yc�Ԝ�z�v��0Fep��񆈑�ٺ~�z�����9���7�W�<�م���2��RgW*Gs;���?�J�Nӹ�[s��~�<�=w?�ے�Ty�����%ן�(P�-�&��)P����x��|����,�m*���dw�"�24sW*�:n����!�2�k� ��FV�@��V8ϰ�h
W�!���?ġo�(?��lX�������8ۖ�j'����7	8Ѝ��x�J��K�aL�0J�ާ��"�f�]�x��?;��g��J�nJB�o��+�	�gcΫ�'GyN���ֱx	2��"�n�'�� �6�M,�����j���BC��̟���<^Aٶp$.��z^!�ː��[����~�z� 1%��h���}lA.�{5�����lz-�aF���d��\�+Q�G��I
&�/0I�ie�j���3�fnt�e��y޴}�ʵ#�W��@4����N�N�����4�:Zg�s�;1���B	��V�k�Guyѳ�����97pk�j��|.le>�s�Ǣ
��2��Yk�a���<�/���,z�k�
N�)�D���-^<��a�}6����z�<����r�&�^���z��_w�#��v���H�9V��n���X
r�]�!s��_��_|�E�m�ϗ���Q	LE�8s��ɂ���e�Z��ǻb���"X�K}��ߥ����r�V!����Znu�	����,V�d0�ۯ���4s˄/,���9������S��Ov¿O���Ŀh��M]�S�(�J���o�7K�4��nӎ�+�(Q|�^�| �2g�!h[�����=�]
��J��EZ�{���i�����q/�������Ã�C�0r����h�Mcƶ0�:[vQ��L�P�a]G�|q�V>�!V���]f��%� +���{;��A�C�'�f���۳�tv}��' ���7e� J���^�m��T�I��Nb�)��D��kT�	}�b��t��;	3��g/lzG�{�VEiX�՘�TϪ͚��4��{�!��3b�U�iØdV-�����a(�+0״y�i��P���2�o.��?/�r��:YY�w�1��������%C�󬐠i#w�q���ro2Ӧj����L� wؕ�(��w<��'^����J/8���s���G�R�jU���TI
�y�����׻Q	!F�l���8�ֶٲ.��� ��11��6;u"���N̑��A��W��B�SLzrb����,j윏ځP�^h���" @�Ĝ�es��F����y��u<�< ����K�Aڼ*�S{�8�,vm�%������&�WULX�(M§�����@��6<8-"ku�V�΢�QL'����=�x�!*θ���	p�>��Yf=���y�F>�����s��ΫWoӕUױ�d�v/f���n^�2��ZP.��[�9
�zgvs�&3$VT%�K�Jh�����c#k3AI�m�^e��VF���e�k�71���\si�����&z/�}�Qmbn�(疽���ZVV.�3��5�u��/���o99�vM�V���>���w�s��q��������?��#�~�����/֖�4d�Uꉅh�|&�s0���`�I��a�v�V����a@��h�ym�Tn�i�8�W�\��tb9|p�z��{i=�.�����.)���ў�8
���و�R$}s뜣gW.� �m�.�T���x$r�|S��B橧�	�t�[�9f'j�3�n���2`"����<���;;K��^�ȑaH ��NT���Q�1���B�%R� �P�{H�|6ZM�%�Ȇ�T�������TWڋr�z=u�o镶�J�T�RuN)Y#�3ҹ���w�X_(�%�T�Y�xS�<qxWʎ3�L6�?�Ӄl��O�uB@d�!d ��J��z5s#P��)���fhI����P����{�N�������K��� ���{�e�}��q�޹3CEZ�-�T2;h��n�6E5r Ԝ�� I�Eп�?<F_i���� ��GQWpK��-�Vb�Ҙ���	��R(ˢ(����ܹ���g��}���>whɑhy������{�>��g�������$�ny�(>a6�G!�$dT#��f~ܴ��[<t���d��9��&�E�	�`8�����h;|^�w�H�uI�R�t���|���0窹䀈��O�����'Η�h�J&A斯!��>]o����{JO�^�'w�s��dol�� ��D,�ᇤw��e�H΅�B�Q�L�*Fǈ�ҨPU������5�P�/���ϣ��mS�,�ɽE,��t�5�i�I����C瞏D�ȇ��p%J`����܉wC:=�{a�1�wS��)�MQ�9wߧ}�|���i����E7�k���wm�C^�ͷ � @���Qr�BD�Gwܩ����v����,��{�����Z°���H��SL��WK��~�n���('�س�uSpy�zqL���SG�.X|SȲ�o)L3a?,\]���V���,n<��oo+M��hCu:�l:t�A�)hw��c=H�
ׯ<G�ܩ�'?��[�Z�&zenbw��t�C���kDċ�{�^0�se�Nh�{� ��r����N�QѺ:��(���#��k_ǧ�x �<��U"ｐ����M"O�����ˠ�t>�"�����Q�E
dѬٮ說�*�-��iN�~z��b� ���I9&��j1H/c )� ��>����¶�A�O��n��*�nD�)���'_Nk��PS�yOn�R�KW�_��Zgw86�T"�䞋��P������W1��"uY��(&�[r'���z\�D�`8�ijκ�]t<��p���'b��"GӐ�Tr���8�Ni0K�߃�'��;^E��ls(�W�������%g���k7�x�lٱ���j��t��Y�D���p�����(l�#��D6P��4jO j��|Șa��I?w6��ߑ<��ufk��ҍ{�ɇݥ���9+eq���: m��V��Փ��7e!Z�Q��m���~��o谥��V@0��@���dG"a̩6��ݺ�kq&9`}�|�=��*�soE����<6�v�>O2����l\�j��G�]jCt�T{JM��~l��W���,�\��XV2�0H���}7��L������1P�nk�cc�5(Ņ�[7�gR��5<v�Bv��]߿Z����]��>�Qh�^iK�sj���������@yʅ�p���NZ��������jA��1�*���Y�bA�I[�O�*G6ۊJz��U3�ۍYM���~��^ʷl��x[$L&�y�G� "9��̡Nًn"�����Q�^N�b��!&D�����CD�h
gV4`�]v�Z���j!�(RFg$�ק+13GE��x�jŪ4�塸�����#�7�o��8�s�m��4��� 7�Z��l1��D6F�6-�,A�w�!m�3�7�I#���:���������1�O����p5�
�>��u�#B}p��["�.�(��bc�-x1�!��i��gUe|�(��dWJnVB�j�C!��1qr�T(~_Hw:20Y�LgT�a�k�(����{{"Bz�~&A�"E��E�:����$��v�he�����(���ύN��v��T<5��7�]ٽ�[v/:�`��}�vH��bN��9�G*� ��G>F}�����\�S~[�N�wy����	�.�/\.l�<]_}nO5`&�K)>Ά���_��DVaZ!��m��lJ립���"iNUr'^��5/&� �sx��3( �L���ӡ$ú�W�5�/[�at����07:��l�c9Aǿ�eE߄��FzT���o�^ǿ
�H���ӡn]��rV��t���Q��D��C�͍�i�"����@|����14����h<HmEA4;��}�3��ʛ�P�/�_���pMzYӽG��1�B��1�s�<*91CTO�5=������(~t��H�*dJp��uއ�W{	��oQ��213G��}���Z�.�w|r��ޘ_���j��;�.|��!��)�>��_���v�M�uS9�0��
t�~5[��+|StvCOԜ�?;<4wNO��.�7n���#�b\��HX�S,R;�z�"ʄ��aԽh�8��c�~͡/���"z��|���4�oD/-w�Ņ�uD����+�qb�F�74��F����X�)m3����~8�����D�~玸}tħJ�ͧ�2�06�)E�8�!=�Z����{ts��Ɔ�3j�!�[o;��^��o1~��84]���ke�==��3��Zo��(�Vn�PaT 6��U0fg�XO��Z�*F;EL�%�'�;}MRɱ^(bt�hva˼(���Qh�g?a46�Z�ϨB��0dxq'A�P���mA�.50�t�<wbN�c�}L�Aae���Ĥ�A�H&5шDԩz�
�N��@j)beq�Cl���Rި%�����6��nX�<m��|��;޷Ή�P���E8D�Ʌ�oA�@oYy���Q��RF��)���BNb�`�(�u�eh2I�O��rEb{Qz������CtSء~/�=g|�����e~.�(��m�XN34:mk�X|D��Y	��h��z��(U�j�u��u�#$IE�Y|P3� E�#5E�9���QD%H���i�!f�Y�%@
��fH�n�.���!�|��U"�W:�]�hҿ⬾J����<H�$�[k�ނ��N�8{[���鹤���0��"�|�ѯ�N&���PTK�{7�5g(�^q%-�C��y���M��&ȍ^��z����X�>ۛ�_���to�@��:t��|����6�l&�Ch����"(:�TJ*��4�tߝuZ�b�����Si������GM��f�ҕ��w̪��W�'_x�#����>���:�R��6����#�oi�&�����E´5��i�L��4��V�s�q@rE/��Ն�Q�{Hc��i�}���*���9�Qv�>Hq��f���F�-��":�/�f�2}M+fHMC"��'�+���v���z��x��e���Lƍ�<;e�5��	cd)��K�������G��+Wy�*Y{5���+�����	��@�k�������)��R1�Vr�$XD�+�o�f����7}�l	pU��1^|C�#+�;QC$4�D"1��9�8�BZM&�Z�b ��M���,cm9j�o��X�Io���������=)�1
��-	�t����CLz�!'��pJ�
1||H�����8�^Vq9Dܚ��9~�L��1"��e�7d�ˠ�-�9EHuƚ�1%*8m��^��"V8.v��p���c��H����P6����mD�ΕJ -����zч�Q��`O`��ްʺ�V:ۇ�Ql�8���UaA�)��Ί�2�E�L�b������{�L(�Ъ-�����-~=�
�A��Z#��8Ս⨙wAX���6C8$�kp>Ӂ���!(D�\pa���#��r�n���a�O2�*�w^�e}�b���>�!�D�C��KD�Aڶ3�̚�"�c��[�0�tJ�^���rRx?�Eq�������9Ş���ډ7��ޢ��=��G���y=��C�E�rʚ����r�����4�}���Szɩ���P��ͥ=-
?CW��n������vՍ\�����t��E߫UUQ�,��dR��U���e�����/��x=*�s6[)Xt�#;�{���e�������}�[>�x��E��"aڂ�4�+>z1�|��zS2�B�( �!���ێ��lt�*m�nH���~�ĄjDˁqZ�Y����^�s�A\��b�o�����B~���k���\\���`Vs��u�v~� @J�@=�c5�Wf�+���ࠞ��q/N֜��2�����ڄ�\	[<nZ� B6��0��zKr�s�qHu���������|B�*Jq��R�"�r�b��C��v��1	�p�Ӌ�G�Ǹ�D�:�M
�% �;�f�iȉ�J�q��w��0��̈BU��K�A!�e71h�o���"_74�p#N<�n-Hy�[�t����u��M��n�mB-6>O,���HRTzߨ��vS��f���ﱐH��XpDE�x/�z����2=�9�R��O's����d����
�����*�IY8o�_�=e��gS�.{Z��@
mo��6�?sK�l!��A/m�+m`�I�qG_�q�p2�J�ɘ����"��fu�l�3���ֻR���3�?^8��������ɂػ�3�g��P���G��O�@��w�S�������y����~�u�"�S��''G'2� {"������7{3n�d��8�;z��Pj��8]��.�����q<��ӈA�s�=оI���`��c���1ESת.K�Z�%ݯu�ԡ�?5���h��Vl��֗^SU���rM���M&�~�����+&�ݻ�,�������۴�5��8�v�\j���QML�L�lo�o��窼sy6?-M��}��0/	u.�cuN7,��x�!���L߇S���Pb������E����4�ឈ#B�&G����ҍ�4�����3N[|�r�w��%�N�b��郛���ꇛ#uP��M/X����)��3ނ���\��,-�+�ר��Aa���6�/t�,9�wQU�Eq��T�G ΋)���4~�U?ՉBgo�%�)��a�pR�u�[��ЌU�>� �tf��"�Y�9�P�
c)��:����i��$e��#FQ6R�"�CA����mrº�M�L�?X EEq>]��[�.�1�s)��{�1��<��*�|9Ԡ+���8#����n"Ig���h����G�\ߵ�"�v�X��mmk:��=�od�,
r��L����O?�"�G��c�úveU�B+[U5$Zеb%x��5��c�tT��W�v{�t	y�Bc��K'�Մ�'��o�`:cL��o�X�&�S�nWM�6gD�m]k�-�ɦ<�J:Ѫ��k���^��:+7R;S9�u}okJ�t�v��xL��>�~��o�J"�l6v)eמ�uto��f��.���J��A��ӗfs���̊aD�H�x��ᑻ��n�l}�]���j=���f���V�-v���z1]�(B�cE��K�埣`�E��-z��=�>')rܛ������
Ob$�d'��GDf�|�~��^���EnD�ߒla�/����>���#?r���t;�E:�q4�m^���&�����Y�����o�W��t^�U�+�) �mb/t�yt�,d]O����[�Y�N��"�=��];���Cg��r:+�Q��"A]"ކQ�7T�s��n�9w҆)��A�*<�Ȳ��v��&� B�a�	�0#�� ?m��_���GP �K
ft7�VAH�)T*N����3	#\�\���%�Hpi��D�g�U���Ë�T�pכ�;+머.�t��7�����aJp�f6��A$���Pq��ڜ9GС1)��LN�Z'm^�(!�P��@��B�4 �5�Lp�4Wj��)��Jn�)�^3ꋸ�,(9�(���d��RǦ��>[N�f �����?���P�Ed4 �~�x��+@7�������8G��{�{-}L�v���H��'����i�S(�j�e�jM�۾����7����p��SZ:�w����t�:��>]~me6gm��X�.аT!���J~X�zZ���RGσ�C���Dj��shS�Vw~�i�qS���1�Nz�P���<�_��ž+�S_��ݹ�'��b!���w��6	`$�~�~h�Y.�o��?X7˲��ǚn�:�De��-��׋3q|t¯Ϡ��
n����=�c.vq�ɵ
�]NC��-����W��>�6�smݞݼy�Iꆸ���s�?J��;��������ihY;g��c��T�y��"˷����x��_���]ۭ���^�`�Ilց��h*�CC��{l���,��9���t�5�c&��D���=d����	_z�=��������ͦ{=�U�$-l���b�qv��5kDr�I�\��b��iJ���І�m�`�r|�Q�.~1KN�h������8 f͞�>������_Q�=ԣP�`M�.y���;w�/����$�
���k��zC7�z����2�lW"8��f
!����j:�Q���a`�)�s]ͣ�F_�!q˧K�/S���[���:���Ns����]�:3����	�����v~C|�ژ��ўk�ߢ�\�Z�t6�����G/��+�9UP7dB�{�,��z:q!2��SD�"4ZK��`1�5�u�'%Nݕ���v�^���~m�혅�n����t�Ƙ~��x �uXӹM�����Җ�ѷ���龀c3��Im�(�3�u����XWYZ�˶���"�j2�˥{eo�_���b�7
|�����'�3�k;� �E�/��(�����O�x�{��Vz=\�������fM��p����7,�+{�[��l�W� ��� ��W������+�ݛDT��5�f[�߸���ܜ_��{�~�k�R{���7� �� ��u �����}�����H�ƍ�g�Y���B���-��.M�!�a�C�.�{���k��!d��&(R � ��u.����M;2+��m���'�w��g?Aw�"����nz���B��u��� �f�cD%��bghJS��p(���lp�I��(��@�0|�Ά#A:a��ŻBj�7�^E��(v6��=1C�t�]�s�2���d&���>�������K���V��Z�2"[UO��C�O_߯i���*�� �{uIUb�^���8)�h���!��H�S���4��n�\��:�4��S����W,�Aux�������)G�q[�-_i����_k̦�W&���t:���8x2�W@b��;��'ĨsA?���ͺ9^o�;ĝw�oj�Lr�"7�Dn�g�zZ���(�,z](ԛ֥�k"H#i��􅑴����!,��-ץߛͤ���@���J+Tׅ����(�{g���[�1޹�>��M7���>�'�����Ki�SP,��������'�Ղm��ߨ��X�a�̯:��S��%cj#Qܬ����4��71aӵ_����6E����0D��|��;���ފU��j��6���ȶ�'�x�?��x7�M�Ⱦ�g�l8�����Xv���}d�w�ǲPZk���֣7��d~{~��}����O?�����
��k���(��F'�+һ+��t|���s���p
��Y�����jV���uHf{;@�����]Y�1$}ʴZQ�Uy>�J4n�Mgl�i���۴�({�^���l�S����|�=ХE;���Fe�Y�	��<��%7}��kq�\���rmWDMt\������EQ�.�������ʕr���\ �S��Έ�ά�Z�m��:2���=fʋ�Ġ9E`ҕ�+�i��_ӣ"�\"e�XxD����MGD�ߨk�am[����E��|������XX���x�i��;��[������n|i�Yܣ����<*��S�����1E�k��>��xSd�	EӶ't�kR9+� 6ɀn�i���	���ԥ��V&���:��u�W��ț�
�o��Ț���G@�{�k���m��D�������{����ݐ�(�`�h1z*��Ѫk�	z�K�qND�F�bD�P#fGЬַ��'�V��PKc��#t)%�0��m2	�Q��'���a�|�Ƨ?]�_{��z?�7���Z����F�vϮi7�8L����<6bC/��E���>���8���X����}��eE�ra��(� mJ!��rSn6�m�6��Qz��I��%�K<GW�ܥ�j�h.X#�e�D��,�����x�>���Ѣ�nyU�B��[�k��rq�����g����x�7����F��3Hcŷ��u>v��}�N�7�{F���}_���?�s^��ԗ���j��5�$��Y%�?~����ϧ�ɤ�R׵����\�����˴�?�� ��%�*���h�A��[��7�M�zQ}�_�6ә�-�����}�yR��(���@�H@E��Ƨ9k��I��o�)���w˱����t��f���-�0KI%�? D+\ﴙ).8�H$|Q;��x0p����'����o���g�UZ	[�������Mi!��뎎Oo/��/�����j�ot�~�[}�n�g�~��@gFF��It�sfc{.W��6Ϭc��q4�]]	��W����BUZ��E�.��U��	��]�"Z]aޕ"�/�V뛛��T�/���^���_�6_�e�{
�[�n7�:����8fVW5-AM	:�I�@ktFı�s�g�(�q�;0�{pg>-Z�}���|�2"a��Iܯ<��j_a�Fϴ�ؾ��qПT|G_����M��|�������Z���,^���nu���֛w���ѽ���-c�_��߽'ަJKFF�T-��l����r�dm&/X���VE�5��ѬǶ�~�H�{ꪺF�C�����✊R��us�i7�t�^��vS������V|h���Y�6�Cf���8��͕~��Lʒ	�=��|S?��4C}�	�Vid"<M+�ܻ��m�x���o���/�=f����l�'bZ�c֪�(Jݶ�;Z|�c���K��m�X�5W��N��%
�o�h|���W��=�қG'�_������o԰�����R�Gcd5�S,_�W,F�G�TY/i�֛�[ߣ�zќ�Y}��o�VM�����kEW�u�#������v�y��������7�~+k����U�Z4��m�Y1�U!zY�Sq�����zR��}?�ZS���EA���_�����e�b'�0-���nܸ�����Y����z�u��e�@	a�N!thq��M������{����GO���D'���^]�����Wˣ{w�f��7#c<(t���Gz�N� �"�v8�t+4�h�<q���Q��O?�ϖ''wh���������B�"�S����D���_����Y��/�l��d��� +F�S}3����]�*�Q#����.
4��u�\  $#IDAT�+�q]��~�g#�O�q�����&��q�����}��E�yŅ��������x�;����2)���z1�Ȱ4$�$L��օ��1�{�9��)>��@J��_�X�M�T���a���o�t:��:I ��(��*{t���ES4��H�p�K��m�eo�0�A�N���w!H8=Yu\���UJ��C@@@rIa��\���YBJ���k%w�ZJX@����NiPx������|���9gΙ��y�Kh�e��JeF����m�Vi,(:M���n�ﰴ�#C~Z⯩�l��%���6:9��Y�°NC ���J�pJ���7� <�Qɰ�����8{ƭ�ZČl�[.�O�_����u�!mN8pNrE_�Rpƾ�%wpZ^J�]��p��o>,��q��OR5|��L��X�In���g���
Y�C�g��Y$<�'m1=4�����U��s�3���*�eɌ����}6wf�d�0|?#Xҙ��ܮ�Ga[r�D?�.h���z�Uȋ��aV_�`�%�I��;����hy����ټ5�$2�̂x�a��_��3�S�=�,gOnv������������!�{���J�=�;�Xҿ� î�}T]Zd�TWj������.��|Cl�"|*����x�	������S8���*%�m�RjƎy-�������Ə$�
{�q�wVؖ�����-�p[ ���<�ӆlS�%��nk"*��$�Y"9 ?��V����d'{�(f�<�{߱�g/��%6}ElA֦ǺR&*��
��פ�Q�e�,n�dV��M�10"������J);���;���x����ѿ���,"��.�S�i r�>%�Rw���x��Jt�:��Pa}?U+p�j�Ç֭��<�!�>	�.�4<;����\��b�=l�(�iP��U���|����b��֢�%�/O�5���_W�7W'z,Fjl4��{V��k8<��.�ɣ4*b Z���ɷ"��
E�^�$}�������ۧ���q����O1_�g�d���=�	v�c�8�N��`��e���6�O�@���V��(Iz.�wӚ��Z	��|,�҃��я�[�߬|�P}J/��3�j�d2M�z:��H�8�W
W�h���O��%�>�e�w����>ȡ}�=�ԵI*mP�������`o/�$����N6��ߺ_�x�P�W����"e�=dC9E�@�*�8Z�f����i�? h������M�����A�Sm�����qSݨ�&�jy�]14��1�t��]�*G)T���io�^���o����f��3"E�:�k-t*Ⱥ�� ��5j�!�g^i�ʡ�֚f�y/�Z~5�"��λg�#?����x� ���~E��<��RZO�g��r�<�����S�X�r�d���8��G>^��͛�CL��"!5?���ed��d�l���f&����t[��C������w
$�)�1S?�CG�X��Z}�^�0$���6�}$���[���Է׳��Ș�X��'�hm��Փ~v/[�ɚT�����f���C�+�L�_U<;��BR'�R?��52�p�^��d��IdCz�ͻ����!���Qi�L�A|���"T�X���a3M�&�'��X��>^� ���>
��#ɪ�[�Ȃ�_a�.�W�9��[-5�ɮ@B'7����xe�ro�.3_ i��ܔsX�z�D&{@M���$�j��8�ش�1�M	>�c���1Z4j�|��5��0n��cUI�6���k䮽��!�7�#�7�!��+�N��\G]3�]����U=O�wǎ�.h0uYo"m� ~BC�5*�"h���-1�[6�\N5�k";#��M�����eUώ-�\="��B��%�j�U�Uf�% GN77D�	ih��>�d�A{��j2�i=�X�y��!���k��_z� _����'�l�*�\Z���CX��<���}���2A�a&�l`�2�������{��p2�V�Ϊ i4�B%â��8qI/N��_K��(��D$1[�}G�uon^�k|��6;ʱ�%��/�|�-;�Pq���	�<"ΪF*wy�Y�*@G�?"u��B
��6�Y(&J�J~��_�(k^�7�D�0*/Z1ȢQ]��n�5���~���9�FB��T�k�X,�/+J.�����[ ��n�9&t_:���Ïa�i���g�5Q�0ߎM!�wߐ�\���B���/�]��/p�B�>�P|Oz�?����/����i�N�� ���We7#i�g�xR��h��>nȱ��k�<ΐ��㋐�2��0M�W&������q3�;Z�����h1�d³a�
-<Ղ萬�QۺݾVￌ.��e�-��>��|��1n���w�w�V�������7
U4�Ll��w��M�Y,?S�l�6����P���[�&.�]%��u\$�A��=G$/7
�K13�;i���A�Π�J��L똻+1F�.z���:�����G�+h����j���F�3��+����l!� ���W��̃2���٠�rU�칏�D\�ι`{�d?n�[z��5~�ީ���~�~� #y����M/�$s�u��MyXˉ-�w�X&�=(V	l��}]�j�qvVVT�W�x��`�F�EpyQ�:,{����gР)�9�'��;�lЎ�rU�7���Úѷ�wE��-\y��n�;f�u<�w��N��P5��)}�����Y�d�|��y� �1�ᵈ�&Dm�Vm?��%��(�Z�;�N4Y��T�";C�u�C�E��MAf�1�?��aI�p�ɬ2wu�װ9V�4p�+|�_Ev����A�iugy,ߛ��_�]n�m_�HZ^��,d�lN������<���ӵ̃�����!p��.ܚQ=���dEWh�
�y��%�<��}�D<�^����f��"<%E$6?R����X�m�!�!��*��2�ZJ-�L$tq�aοo�n����(��#rhT6��.ZJK�{>���I�i���q��ܞ��Ԃ}��(�c������Ѩl�|M-O�y�Lk;()q̦���ǅs�9�j�^���7*6��e.Q�������Q|���I�l+0�bp��n�{i�8�HFm�f��p4<qq4���8����MS��mv�<���k�Y�:�U�#�-�I�?���!P߅���7�����O��=�(,_�ͷ�SY���ꍫC@C����M��i�rs9�z�{	�2�P~3�z�Q��:�X��!���fh�^����a�Etoi�.�/Ue�$n� `!�J��+���|-q$��6"�[�e�����#ccr=v���Dn�`��w��N��` pBO�q����	 ��o���U�q-��|�Fh�!���j@]w]�ŏ�'h$���	�
��)��/W�)�*�;%���k3��i�"p�WOU��f���iUR�Y��+��J˶$ζ� �3_J�"7R����a�8Y	�V��P8d5�P�����g5-��|oR<�汔&�.��ZGn�Y4���}�����VUw�������Y���Kv����|͐dY�I�S7��a7��%m�s a���m�D��qK���H���YW�X2ـkv<�80�-�@��dۉ�s}����"��%�ԉ�5�����=� �m�I���,�=�5����Z2���D��y�#՝��X^�	�냅Mg˥N�Y��I��y�>d�VgFS<� w,혍G��X��3$���Iۭ�����p�.���%�
=!���8[�_����Q0��t��VLAt�뵧a���L�L�Ϣ��N�A���I_��ǰP�v����H���FHタ��.�_��
�~$��T�5�#��� x�K�D庝��<�x��K��)�ص|/�ShM)g��Ek�M��o~"4~�)���m7t�{�gXD�-��j%�%��Oi��WΎ���O���]�5���7A�nB����y�������E��,�ڶ��x,O��x�dZH:*����#���Tr`�Zw�b�g?}�r*5ҙ�}��|��jL�ZhV��`[4�⪙�w��l'��I�Y^z�d u����2��Rj~����Q-Q���ZJP�F��A�鿌<.�`��߷��-
ܥ�����m�*[���g�M�vi(����5!�N���}p�}�lnv^���fl]R���n���ݓrH�b��uG�mۨ��M����O�j�|�]z����rX�c̳ _]\)�?���rL�$!��@�0U��
���:TW���Z��5��=e�5mj�+�0�������LlL*U��|�w�:]D��/'ڹ�<��*�aH(lN�l�%��$LG�N��s��������I=׊|�����W�	E�(6��J�zis|����b������ńVDP��,雗���T?1y��fP�1Y��v*��%��N�Φ!�/{X�	ί��|�4�󜶟_�ۘ[.���0��}��e�,z,�c��VU�����iGQf)J{��ʈ�Y�f�]��C��$�b��:"|���U��l©��{lZ�Z���^���2*Ǿ����aF�C�����~?��iIuS=��('���ѹ�N,�{�r��s竍U
�/��x�8���DH���p�+��ū�1��
)�&+��o���K�n�u�w
$���G ��� �ڬAC���|<�\G䫼D�ߜ�)��+�N�<ڋJ�+pcTg������`��I���|$�`n�k.H�4}��o5����L�0���FoT�%T^ԥ�E{������K�b��������&��~w� L9Y�]�5��Un�����D6m�9o��4/;�D��)�R�/p�;F��q|'â<9��bϣ'��E�{��҉����c��m<y,�;S�U�ٞvE���o��f��&��-
ۮ�(��eR'_	[��������|őֶ�����e�X�p��Դ�R*63÷,�.Є�|n�S� NË$�Q�it��c����*mO�W�4(����+0�Jm�я�a�tA�^��kkg��92��ʳ�5si��X�IO�nvQH�R���?�%߄���ϖ;[Zo9��U>�i�=��-L$��<̤���:�O���ES����c9YȤu����a��+��T���s�W�?�T�+o��Ǡ2rZ� ���=����P���"�%,��Cu:AJ�U��6�&��5��r�h���*@����{G����
����׮���&Z���)�d曗��5;�����<6�H�|�d\�u5r��r*˞���܈e���2���.��wV��Vw�a������\VƆ%*�7�0�2�o��LI�U��U䖌���
	O��Q��a�ۑ8_=����Y>Q��x�$\M��ET͸@�~^��z.o����Fmud��&�!�0�H(�d�c�S*-h���pMQ�7��+�,���ה������0���Ί�D����)���l���õ����&V�k3��Al���A���ϱ¿��܁��6��>:��c3�w|R�(���xYո���W�P�-'mÒ����O+�eq�U��.~,�����n��a��c~���X��4�bLYq*�DB\�o�t�K�k1_�yRt�"_��6M�%�-oI~��Tp��$)��������&)$��JeCú������Z�5EU�,"V|qO�u�����Ά�U�#w��0�(��������>�����Ѿn~a��O!U� ?{��\��i�G�S�5hN���O�J��=yn)����?I����#�Y�L�0�y"�tț����b��v(��v���~Y���:��aT�d!*Q��������~�~O��^��}X7[o#��1�j��4!7��#���Z!��p�#��ĝ=9r�剛��/��3��q���7��f,�b�O���DU�fM}(�7t�3\H><E��+��Wl���@~DiR�P4�Q��6�G�yi�ሙ��AGS���A�*��@���lzYf��yʂ��W��Byiq�3OJ��� ��V��#<�>�ڢ�������OŨ�i�N$+��]~��VQƓ\���((�M��\�%�2nA�����/��fM�[�h�Z�^.t��M��"�#�n��ӫU�Hm;ׅ*P(j���L���>�ȲӺ6���ˌ��Oݔ7/I���(T
02���`�[�O�O���	�u�u?f�}�C/������DX��N>\Z��v�/��lCA�.�+6%	���0�ޭ��>� 9�y^-N4��V&��ޤ<U��6+Px��A�Q-\�7KV�9mcp-�����K�H�I��t���W���v<2-��e�A�A�RW*�n�/V�.�sz����0J8�HB|70���]E����̸��9���5w!ww�+4�����`��<h�p���{����0����K��{�e����M߽;m\(OvsW{~�{!�O��\l@K=�2�bՈXFBt�Ҋ�k�33�'DW 8��b�����Ɍ�b�︎fV�a}�	%�a�ȶ��Ul���v\|�Z:z�	����� ��3�D��i�E�b�z��T��d��Z3�U8�gۛ��M����W/�~ͥj��k���ކ�i���o1������>�4���Y��I�)2Ɂ`}��x�(�$\��A�[�E�H��ǤDS��D�HB�2��$����/(��+�j��jNP�3�[e�4E�I�SS:����h�U�6c���:���JQ 	M�wE߻+K%�,Z��0Q��UEP�;⠵J�f�Y9v��BGF �!lB��2�]!C���b��C�M�WεN���ў`r��Ue3��s�d���K�1��>R��BXӓ.�:�ҋ�,X�Zu����]c�h�"�s��r8��DR3\8�=*WI���
cJz;�'r﫠�eH�u����A�83��,^㮢���\Y����u��ws�Nt�i����Q���U	Pn�P��1)�.��D��mY���B�#�.Xm,�q�.A�4�ڟY�SLJ��K^fK>8�r+BrP�AB��K���5�1�S�O4_
۳�=��ًt����m= {bX^�.� ��rH}\�uwf��z�a�[:%䪯�[RJe�KǀU�jVǵ��\g�X�bbCrk '�)�
`���	~�kC���n\
�+��ִ
�⃘:7�&�V��t���	,��V.x&cOra����s��;9.�W�C�� N�Ò��U�5�'`,�G�x�9��E��B0\�=B �|id�G<m��D�l�&1}�Ze%T�F���N��!�FR��3Ol}����f�H	/:~=;c��PY�_K8}Ѡi�y�㓈x�oƶ���@�ǴL��21�ꂣϞɴg���9mT^Y��{=�m���t����(<�2���ڑF�;L�}�L��g�o&�����g�d<����EGw��ΰ���0iA��8Hb��6��J���dE���=��_mBrS4� |M\M��n|0�*?fG�W��@1�z�9�̶�I��*��e��� G%�@-}�t�V�[f���4S����7)���������g��t�zt6}�L�O�
�w� 'ۂ���y\(/�d���l��D]l{n�gЖ��(��ڛ?g�\[|�{�G*bO��v�}��t���c�J��z�^Lsj����D,��}|���-���a�����kj�mG�	9�S�HVxl��"}(�iM�g{�A�QC &$�]����͟[3u=<�ؐs��?g;j��G�j��N�(&��a�Pqn�o���C'Oi
04%ck�3���ĭ�_�F����Ť��sď�W�jA .�T��Mb�k�~'�����g{��4/��o��			�
�g��&N_I� �d�^�fB�_�$��Es�#ݘ�3L�t��4�帀Ƚ�}U�q����f2Qʹ
��-���u��=Z[OJC3�= P�8���:������ͯ�����K���V>�~���w�]K&+y؊~���O�?H/+m����D�1-�� �C*��h"XL����r|�B=���CyY�zW;�&�8jU���1�Qb��|�*���������Y>� �ͨ/5�Vt%�ʙ��cd��QmtO$��s�+:A�Wcb|�����Y�aϲ7��)s���`L&�̠�ީ��r	J/��+�8�1Ɔ9��QW[�}�666��I�Y��/�H�FX#)ӻ��sI���Y��k���<T̽�m����V�&�������B3�`$��B@���`�>�}��x1����{�ݕ��Z}��襰N�����NC�u�y��<c�M{fbM��6'ޙ|ʹ�Z��ϯ��ٗ0R}�_�,�#�q|�����}�����a���>tѯ�.]�j^����p���v��[@oD2�vVG�{��u��^YM��QǙ�cGἀ��N���'[�LBow��!{��Wm?gH=��6,�E�Uם^��E�"����V;�{�ȭN�u�n>Mt�9sW���� g��&�bh����7�jn4��>^>?;{�\���w��N~����d�[��y��ǣN�P�f��I��t�&�z��(rr^?1��� �p��������H�l���7mk9ޛ�����O�[I�4�R"sߖ�:;�s4s��ϱ �}�j�;�t����v��֒���3?�gq�h����7�W�=R�%�&�������GS)T5��!K�'E�ܖ2*����޾�d�А��QN�J�����L��:1-��:������\M6�ͪ_����T���~�߮OV_}
�S@8���~�a�?��Y��j��k�<���_���EE���G��Ⱦ����߭vԡ��������1�	�烷�����v���s�es0�����3?[�ߵ��G��Ȉ[��Be�~�3�gm����Uq�7wuD��A�i6w�%95 R���� PK   l�X��� � /   images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.png���o&�����[��ֶm�v��ֶm۶m����U������I^�y'g&gf2'BQ^  �KI�*  �Y4��յ�?��^R�	 @����� � ??R�B���W=������+�O��O[���6Y��0�I��I^a����8�S���{@e�ΖxuV6Q�޸q��Mr�X�$l���$҄����vsba[!��_���%�{�����~s�ύ38������$������bz�m��x	�������^������<ý;d�ȝ�7a�����$��?$��Nu����h�Ɗ|45���IX��ˊ��>m��='*���'�_?^��<r�|��p�q@O�������f�����n����O��}P}ʯ#��y7d=t,�dE:�K~���!�����%�� �������)��q|�J&+��VKyri@]�����uQR�c�|5�{�I��au�t���Ԏ;��X.�h������K"��`�כ}e�kq�:�ŏ����a��Q��?V�~�~<Y�?
�Z�~kzH#����yZ�; ��_���������n��6���L�u���m�����DH��	�����)^J0�P8�8�cȅ;�r��y��0��o����L���{P��?<��笔���(�i���?���\r��խ�R�H9���\O	V1<���+�*�h�JY��]�6��0z[C��5�%�c�������sN�1��e��.��P��o���'e�����"������v���p
lqVh����m�[K���/��7���u�G�T&m�骦���WBԷ&��b����3Ǵ�{��^�>��	^rh-n���Ǘl��'/ė����5��C��D��@��x���"�}!���֭%�܋�el��l�J��=EQ|/�sGo�D�I%�s��� �]�+����3p~B��5�#9{^=�	�����[T΁�O�~��9Ρ���_Y��Q��$���0V̑1ˆ��M(5% x� �p�/N�,/w�@���{yDXoW�N�^��|�� =1"� ����Xª]�|uECf��O�v�)�Ȅ���
i�'
8#���P�1v���9�ٺ��͕�1y:����%��e7��5�y`��H]ݠ��LN�9�j!�ᣳҭ�V�A���t��l8ط��`��ڳ�p�����������o��' \(���P�����^���κ�����w�?��A6�iu~�Q�l��<*+�����"<��X��I�I�"������ΜR�{�^����ƭh���^l��8��3���V$_��ı��q�����k�Ke�2	�/׿e�jtO��ʅZ��D�����*oD�n)�ɉ�M��9����[/��|�W'�����N�O����e��|�s�q���!uO�U,C����a۱��\܇�c��}s��rs$$ط�A��l�,:|���;�A�Ě9�c�M����7�����tx���Uw��[m�ω�3� �^�3��Ðr(d^-dA��b�ܰ,��n�����#]���b�_V�Cn�&�V��W4 ,���J`���a�5P�R���0��/�d�o ��آ�K�Jiw5a��Y��*��)X�m���U�ZH�W���J��̇����J��g�q�j0f��E�] ��0��}�eD�	ߦ)��m`�L�xʭ&'�d��j����]\���\���[���0�t�܇����x(0ˡSC�g5�B1�V�U�f������!,����4��O$e�[���	sk�s_�"p����r�̙���|�}�`�o���]�>�gs,f�����[��n�p�GK+M��K���֞�
�E��Ɔ�Ϩ����,����`�5�y����D�Q���]�^���\��E�����H{Y�F!K�e��|���%�\)�ٵ�v� ��,?8���fK=��R!�Z��Ci��^~q����R��$��C��E����������_�l��-�df��� �S��)MG�l'� ��1�k��d{J0���������󑌽�,�X�����b���]-sg������6�Z�	b�93���n5���A}���O��2x9��%:����g*a�z��:��?�r��?�w��� �0f$�gއ��٪��
���S-����b,�#��W��Kl�����E��L������șxhV}!:�2��[��3�Tus�ke��oV���6f�(S۰���-�P�С^�$Qxy��ngp�s�>Z:�,dX�1ۧ�g��ޥ��Oa4���y���3�m���YsImS����x�sãY�
�+NJ��5�4W�q����wAyۛ����+_��q��GZ��s�#���Ǯ�'�6�J��c��P�X$��nЮO%�-���L�1��1V8�?\,�&�{W�D�ӕ�P��t��i0�3J0f�t�b
�i�p���H�R�����
ϴҭ�:v�^��֨�o,�4� ����<>l���'?���wt�=��^�����o��[��?�8g���Y/T����w��b�Gp{�������U��Y~�x�U���1|"3�AA1��d�~~*��Я��hQ���M�MpA�zY  XT~�2KR	t@�f�
��y�x�'�"���QdAn�@S6��f�����|��}QBR�ҸBN��3���ZNZ[�����S %$K�cE�_ns�x��x�X���iv���N�Mc�؋z�)���h�zA�=**.�_����K�AQ��i��pP3s�^$d��.��H}�B�ֹ���o_�@�To��!��a�h E�@L�����J�K���uL�D�<��UJ�_d�Ou@ڞ�f�H';��$�@�N�<ۺ}��no�~.gv�0Iv0��z�^m�E��"'�2PW��\oq=�<BR�ת$�u�[���p�(���6�m~Y�\�� �ʎ�(3XIo#&y[������)a�+Z(nh�qn*n@���t�Uw�B6�M���,H-,����AS�;�rc��V�o=-������1Q��&9G��w�*��i����b+%��;_�X�7>a-P��lja
a��ÂJ?G��Vro͡�l�FE�������"�=�c�[@C��Y�����Ivl�X�f�(ѡ�_�Hk�����peL)�������������Y\�h�-�x��JNF��YZ��5vx\@����^�
�F��=��������AA���Q��Q����0�^��`X<Q�[�t� ��Lk �^ސ���p�U����^��C7bZ������6���'�m�bQ	�A�l4,�@��Dq���S�t���ܶ��z�r�9��O�Û�|u�?~�>�?3~oU�X�� �|zjS���Uf�l6�]���;
It����/���E������q�1aN��շ�X�:;�%񒕞�Y�~�VcbE_�e���aGx6L�a#g�u�i�a����Be��6,���7������ਃ�j�D�Ҟ�L�����ieA*�0�Q>����a��^e�*:,��2��2�^$?���^��*3;�z����s�ky�1����r7��dB�p��q�� �@PCb�~&d <ȭ���6 �C�H&�1o�*
������~O���*(ӕ|�����>���:��̛�7�P�<}Ōi��A�v>�;d��iN�bsc������.���d!��1���K���օ��V�����=wOܼ��`��n_�h��mx����u��\=݆��w�5��댼<1]�'c��6��a��wN���+O?4܂�J�c~.����Q8N�����8�=�w�Ҵ�H��R�=\���!l[q��;��}ۑ�����ZT������H�=)4�]ؒ�����d$O�V:>�l7��V�р�@�T��A변+oǍ~Ƣ<J��T�L�R�i�A��z�R��>GI��8�� C�r PW��;t�v�~������F@�S��4�U��p��/`"c�Px���<���Xd�3�:�7�<�WTYa���}�q�����R��[L�k�*vP7/������H�S�h$��lݺ��9�^�t���b�^��
E�U5�z'�1s3b���O�g��
636o'��q^���RE�1Fo4�#V���}��'�Aq`�-�ñ��	�ev�{�78!��k#E@�L�Tp�? �b|(��q�٢��ҷ�L���b�?z�[�Y�n���v���ue[�qk�#���$9�d�����,8�T���!D��s)y��h`��V|'��6��÷���i�ZB�z�0��gW�H�3p����WV/���x*��h81���"�2�x�~�NJ�W�vg`���`����C���N1c��&/x�A��|�iRf4n�ZLvL��5��)qА�5Z39wĨ�G��;6��O�h4�J[^^��374��PPu=$n���Da�����h��� %������g͡!�����2��]�ܸ�/;�(��}Lak������_�Q&�n���R��\�~��;��y~�������4m=id� D/��,g���Ӻl�ji�]�0 ��("�.����TO�m����A�/!Zʸ�.B�J��3��X욻d�-��f�88|Vƌ�`ʹ�0�a~ݚY6�j�Eh���<vVsʫ�?�B%|Q�ЏW�e�dQ����Ʈ`ÁUXS���4* ������)� AE�P�J�tT���,�!צ=�kd�x��>��M��ӧ�Z?4�NM���r��!�,7���Vv�y*�t �����"U1�P�+���Px�,�8Y:�{,�X��c�d�W��Q��n0��E����T�����K?{u���A���B�J�p��pj�wG�r)��P[��I+9�!z��u.Zk��-A�,O,DS'���*;D77��N�(AQ@��{��H��BAV�"Φ���݊��z�?���l�b�:��U�}�#=x��0T?�1��������$�6���I��7������mlm�=T�W��)AA<4��?f���{�~�=�$.�w��n�]�eteL?�BE��&C�k8�H�ղ��5��s���"6y~��V=��[��F;{�m��|��ʘ�`�%�1�pzw�J�b>hY;D�X��!_�l̧w����hO����(N�`�XʰI�����Ȉ�7c��Z�f���#[U?����d����ǹ���n<]���5&����.굘s�7�K��_ ����Us�-.?e�e]u���]�抋bL�I&C�p�I��a�$��+��K�t���0�-��yf]� ��?#-J�]�2{�.��SI��UuЮ�(�)��z~����)�\��h�����i����,*�ܐ�e���*�~"���%XPj�U����8|�=u:#\�]�CQ{�����X��ݢ;3j���h��1��p,�h�.X�l�G@����t:Sh�`���V��2ĉ�A@C	�u�=.��B���7<��(q��2ޖ�����2��5��8�6�d��Q`�2Ŧś�̐DTһ��% 
�ڲ�tj(���d5#}kKl�J��M怣�M��A��ޝO�`�hF�t7j��;3{RÂ���(8��o�k3ғ��+����MW�z6!\�^��
u��U2�����A���x��&3��h֥?u����D��� qG�e}�9��JJ��f�ep�Dguw��0D�93�-Ջ5C��vA�~�V��4]qrw&�M^'e�Õ1��]�s���1�V�G��3����csGL[��=�o�U�Ʈxv&�R�5��g��Q��x�/��P�a+�3'9]�hlc�p�ʬQ7oؽ��ل~�֋8�5c ��E��w��[��Yq��#��v�
�:�׬�!�g�Պ��%Ng}�_b������I��+���ĺT�ߞI�qfZ��� �M
���D���j����&�J��̉I�6s��Ӓ`-ՈU]�eh��H��wĆ�5���?b88�꜕lђ;]."���"Ma�ۙu�Q���	�3���mdFc|�\c�L�y��כ�	1���,�o�m-#�S��7�ǘe�s�jCHѐ7�FA��+ơ D�Mw�=��;ѧ�Y�v�k06�������#݌�
OL�*) �F���v����Q𩇟������j��W����}Kw�'U��@���f۽�+������t�H	���Fc�$�lM�I�j��K\���o�^�e���A�}�@�3x.6�+�.7"j%� �ڭ�Et4-�Vx�UJ1唲�f�T}���#7�E5� ��l����Թ����_�Z˕%_?	�M% �q���<P9:�5:1��4m�������c���xRh|4M���|�\b$�N��>!;�����4�BZ���t,��Yg��)Ԗ̢�� �5J���f]wC�qr����T���Yʶs
�N��Z�ģ�
?)gr�s栞��[������#���"�ݖ ��D*��s�ڲh��J���/	��IL6�b4�� �!�E� b 7.CƢ��	��,~斣�#x��/�sr�Dn��#��w�w�{�
¡�8=>s�k�&�K�3ԧ��Z)��P���k����"�x�������#1�R
�+D����}L+ݾ,�ɼ��D��>���@f�wO�}�:'��~?_�1��w���U�	m3�fd i)���Ǚ����;j�%�oڧ�f��GzS�S�	m�,Ze�6��6H]sQ�c��%Nݿ�Qf-M�t�I�PU�C,?'O�?$|������W�)���"d�&:[n�9�5��#��ӀW�gQVL�1���;����-��BP���N��jJ1�ȉ�j���pǌ�������h7G��N��ȹ��U��M����)��H�t���!-�z��Kc�Lb�w��>OX�`6��O�{�V��	
٫�}��݌7��	ĸq�/> ���g���Ƕ:>�Ѝњ�_�]m�nN�b�.�� ����\���d�
<
8�:M�< X@�
#m�1QE�*#e��^�v}B B3���d����Ev��Fb�tw'l$|*��r�M9ŦR�9H�`��������2t�7WE�{��c�w0��`3�������m��:��*5?	���5�3�I�;�p,qB���{�q������ܱ[���=�Q?ٔ�_����"g�3GA���lKt�Ѻ~�-��Sxb�)��6��:.��z~�MƢd�3�]�{@oܰ_&x�%p��j�$u��G��,]�0��u|����1�H6����Vc%�����R)NΎ8���(8~���R�L�;��4�p�=lZ;觋+��S�K{�L���ʽpz@ a��~�x4Te(���C�N���Ke�r�4}�J���Q���s$J��wv@���=����:�=p��U��`��A�����!����qb�̞��U�F�x�8����˲~��җ� ��cjSŵu�b�I��X�9l�)�x���ܙ�"�ã�z�	+#���>��˼�!��2/��+q`�������H��:Z,��	%������p��yf�,�Dr����~�1�w�4GC��������%��+��X����j�E�D7����g��Ì6�5�sM³$}���I��x��8+*-�K<Ǡtɶ��	{����;�@�k��p�hH�/��B�H]
�I*�_�N��{��]߮ɑx&���x�J��]�s��R\v�ӷ�`��=!9�[�����O��A��J�����3�^��}����XK�l:��֊���B�T���t'~ą��rۙ~4��yncߥ���g�q�c�fM]�_њ�����kV���n���:K�8�Sm���e��c+���2b�\%8�[.T�GR��}^~���*��e�⢐��S�JI��S�x�\�.]�6Ӄ�ja���l)������~phQ��R���$�^=�]�*
�+*�NLI�]��z5U�F���C0�&��/�DG�RכmG��.:Q'`�Q���8��H*���F1|���:am��.ݩ��v/S�b��C;���v%gy�	��G'|��O���+�sJ�����üdn�'�e�Ry�P�Z�7N�9�80:o`�a��]�	��ICDp�m m��kW�ٖܲ��̥A�z��:�&XYMN�u����Eg}���4F\\���S�t]I��t��qI���+�C��w����"$�.ņ����[�n^�kӂSuF@zQ�Ӽ����j=�Қ�T�0.䮧@H<�ގ��_�� ����SY�C�EB��U��a�ٯ8��Z��J].�h]�,���ە}��Dӡ/�1g�E饚���Km�y�J4�5٣�4dK�rZ�y�j6sdz��a��Ԁ���
���� ���j8�o�L73�s�Y�3���i
R�g�ȥ�r����L����F(N�lx�
�����^��8�	�<���A����y�%�x1bz2l���S�5e��|R�� l�"D\���h@y�� y�RF��sSJ�H\B��lA�O/����rz^G6���>�!�����I�\Q*�@�B5Eh6�; Kˆ&�I�#��%@Q����[�s2xW�rKB-0y%���!����#�X��!#n���T�#y?%8a��6zT;��l�.��0+�#wZe9�a3G��G~N�}l%OŞ�3�w����tP5aj�.]�2$K��cˤ�=�uc�6HC�����5\�����m�F���u~JŲ3�ܢ�`��^XC..  |K[�.«�lD?��-��Z�z.W���p;�}${Tsk�ƺQ�P��{��qgV�����Ҏ��H�w1u/�g$hŖ�AܩC	��p�&vW��A}QkZ'D���d�%�a�LV��:���������iW���_���%���]$�N$�y넳 ŧ+�u����Q[��^󞠦��=�Y�˗!�bQ�d��8��z�֢%M"	O��˷j���z� ��?GSELg,�h��V���Y�-��X��5�ݳ�FU��Y�SUW�-4c�����0p�!3V_T	�!�fu�0�4Q^��g�?��/)��B�1���֛��P\���P]IOgN9d�A�Y�:i����,5� ���gw�%c�{Ư)<u�b��ψ���lf|�f��$ ���ꃄ�R�<����g���3=s�Lq)T��D<�k�l|�O��ˍsiF�c�t)b9��ԑ,����CO��a@W���l�4q$՞^���M��5�][ЬJ����������I(T�.D�'ڑ1{��qIg)�/A/G��
��B¿X7�?��w�;�o�����T�"�1^�� �n4Jg��/�~�U
�A�@?�[�JO�*��{������e��\�x/w�q!�~<=-��X�E���qCb�\Mg�m�<R:�|�ˬ��[�K�[��i��xO�᝹'Vq��������[}����UO��5�ꃘn���� ���_��nEfj4]χt�{m'�}��D���?>���հ`��S%�V$]W|��B�����[��H��_��iYO��H�_+��|#���ɕΓV�A�i��W�I��h��k���9��v�Ӄ�t6Sj�08� .i���I�9�ܢ���t��n����."d�]Tg��<�jK
���\�/F��yJJъ,Vy���+2%���oD'W4�h��f��2�l�>p�R|���9�L.��x�/Λ{�:(05�����S�qeG�Rl����iHo,����7��ϱI�i�m�����#�9uPz��>�c�O��n��G�@>J�E�ʴ�]�R�2R/jU@k��ƌ+��:07=�|�]�@�R�N������~		OLٴ�WYUu��S/W�a�JLnRxg�$��;d^�U�J�x�;�,�vBi��7ٖVw��i�O(Sbcۢ��}n��E�Ol���������u��>�վ[�0�Uk��&I��\�ZBMe�&WS�rbY��Kn?Ş�����#8�%Mn�O$��<BR&��wU�$���lG�
T�%|u �����*{`�\`�w�^ S�G�J+�
|�����G�l�d���ʜ�
z�&��ɷ�!�i��B�qztG~�U��w��x����\vߥ?�j|�X�|n;��� M#�&FT�I�`B}5;��Wgh{`�p���Y��?��wv���Tip��j*�CA�xPS��?������������|�bg䱡�V	����9�;�p:�9i_9�����I<�>�9'��(���4��N%|�V��s?Olo��61����1��2����*�rN�X�Ӫ�@�:N���M�|_�=)Q�$nu
�A��O4w9ĉF����P��|ϴ�V�׹��ҋָڶ��Ͻ(�*�9�ҜK��ʭe\m�����'W]�J�F\����>d�!�T(!��`��A��b���I��JoeH8k�q��N����-�����ԍ<��NB��-�E����yt0��Ի�+��;ӄ"e�0y*Nd#�3����>ꗾ�l� v�;i�?D�����T�3��9	h�xB���9�:'�d^�4���b�~`�~����j�GD�p,
�j\���]&����Ԣ�x�{����%�y'�Y�ypf�Y<R��@��
��:t%#L��j�L�\)�u�(��V߶
���c٢�>�ME�e�jFV� �
��y��tJ���B�!� Mg�h�X�bMe->0d�a��c��%?����I^ �$[�ǃ86�ڙ%<��{r*�be|�H?�O����6VT
��;���Y6[����c�*���B��fk9J&�pp�@>ߋ\�q(��>�*W�Sr�c�s���r�7���L�/�@g�,ŕ����6��[�Oe&���A��hNM+��V-f���A,���QRV�_?�cY�
��
�#��y�]	�x��-2M�w��F�p��0�}�JP�R)�B���&�xP񨡧���}E+p��l�pvT�.L���Lǆ�b�n[v�����!'=�p���N�޻Yr0a��,,��lvs��i�޾f��i6H��b���3��h`�p=�]zZ.v�6���:Z���=dB��4�4��4���r����q�j��s֐k�eZ��0'kh�>���YG*W����?\��l.b5�H~�:+;&:S����yG;*@B�_A����V�8mK�5
�@C�K�����ۯ;�rF��i��+��Y�#��3������=C����84�Ą|
�Y���:<Mi�+������`��o�	�u�E{5��+n�g��	A�L(��v��+�;�� .�����-M�ݦkI=shra�9�^�(x�;i�2P'�y��Rt����;�W�cC��K�,��{�ƚ4�X5
�>�Y|Dh\�'X􅙆�s��s|���i�|�����x�����VFH�
��c�㎪���1F� n��ͩ���V��OYV��{x�2
���L��y����_��G�@|<�GZ���&a{�rv�=��6G�o�&�*�[�m鱰X��[^�Ld��!���js��{�" ���5��W��͐����4�ر�rf�f�O<�����O'�}�� ��D|�l����Ee�scg�\C��S��.�YAI��I�i���c;��p�RZ0���ɕ��z��~
M�1�u�#�b��w�"�Q$;^M�L�l����S�����BD�Yު�$B�;��E^�1��O�4���.�q
G����Ɂ��8�y��EL��O�4SO�z��%�Z�LI�	�'*ln3gR���S�S�6�=Ň �a��rTIF���Q~��"� >���'���r���QcˁX���S�sc�y�v�����UcAex2�	2�_y�h��Mf�������Sb��&�����6Kx��6�9g�Kґ�%`��؆m���.5sR�L�D x������7���Qb骭��b���*<�����V)�9����Ԓ�	���Y��1���.�/1(,f�p�U�Z��ջ��@!���3s��P{1��'rf�w}�)o�&����3��u7ϝ��#w]<�]Z��1¦�O)m-Km���+�� �.�p�!�\���;ݠ17��@�0�A��ܒ�9aXy�dA9�w��4?�!�#�v�_+vGkudt��I�ۤ-�&=eޣ�Z���2B5M�j+x��V�%�C��U�� ɠ^1KS;h��ϧ��F���G2�ss���N�Q�{�s�Y�f����ȺÄ����k�Mt'e36���6	pg ޮ�Z��"<�1����:�_��1���9���}�ETM���o2��GE���:	N)��_�e@䝾���`;<����(0���hqQ��T[����>���')U�'����d<\��K���}��R���fm������qL*j|&ZX��ie̸
���p�~Y��I�w-�O�`N u�I�Gu�uװ��h�ȗZr
�Q�/�j��u�
�VT����gt-h������p������=.ܡRQ�Y�k��G��f5~P�	�U�����4F�x���5��H��n���v����kt-T��u��5���݋@���cy|�wa��G���v�.D�'��� �����W��ιּ�=�޺ؠق����77Ej�Ts��ϱ6ȅDΡ���rlȷt�y�e��d�X��RyO$W�,�q5�%������������� ��7�ŏw9�}�z=���j����`+I�B���~�3ԧ2�x�~���K@��u[s�?�2Tuy�|^�8S�$����u>���a���:ņ�i�
�-��U�tj�,()�]O8����唎㪣��L��M��ִ���;D�69��>O6�5fm/�4�?c�H��`�oħ`fg�<k0��~�l	����jfiA���հ>��L�2��VS�J�����ݖ�=�*�Pwt��QU�'=�
�r��(qqf��-��H(�m
�a�ENS[wt}L�A�%B��Y4v,����8�O�K΅�a�.u�ЀoI�>�j�v�ky�F chލVTx��2RoW��D��d�߮N���oi�圎ow�6D���2��� K��I�S+8+� %� =��T�{I_ڛ�]���z�}_#��b�5&?��h�Q1窛5(�;v���։M���Y�>qّ��h��l��r�^l�c�g'�Fٞ��ZX
��Y�߮�?��U���A*@��=f�H��Hlƈ�����\=8�w���txj��D3��p�(B'�$��Q�S�,iE"���T�ČM7/�A�ƴ�f��8�u(j<w�5%9يE�#��u�9,�7�e���Q��ׂ�����@�*=��i����C�:@���>�Ǭ;�������Ҙ�x�N�}��E�ّ2<s�=�s-��q��]��ܫ멏ut�%E�5i��vU�������SI����h4������Mh�%{J"�7�Y*�\bs'� ��7$��b�;��*^J}0[����WP>� ˶k"�vy�j�x�A��m��GG��_+m�����I�s#!�ƞ��~�E��1��ZvxA��O1�9��fN�B'�Jn�z���M,?s���AR~u����0�-C���M��x*Ӱp\�Aq�E0������c^y�r$�9i\~��p�zdEJyܾ�>�ء5���G}?�#<JO.�����:�.4c��t�Q������yɹ���ޤ�;��KM�6/+��Wz�IUZ��)lѐ���o�I�x���l�=��L���#��n�ڂ�^�9O��QDL�Axv��u��2�d��R��0&ri�O�.sjí�������<������F����gL�̲�!E[O֮l���U�HEA�Cp�
oIͳ�t��!� ���jW���.V[p��h�߿�3�KrV����f���$��7Ym��[�nɭe�W���XQLcCt�Cc��A��sU�jK�@�Ƽ�]Oק����P{O�n+����Z9��B��r��0�ӧOT�����闚4F�]#P��G��Rʠq���r�k	�EW� �Om�*��j�Z�~������7Y{�%��q׏�h�N/y���r���[{ڕ��5Z�ŀpFe�s�UQ��^�2��N���� N�N��)z�-�0e��>7'{��ST�qZ�߱E��X�J��x���"7?�ْ���rC�d�C�ٹNa�#0M��}�,3��Q�T�Rr��]Fl�-��pl1��Z��0���X��<��ؙz{� ]��VT����GE�������T(��bH�C���?�ۯ��?U�=���׈U���q npp���4��:����I$_��΅?�w�q?s,�Q�� 8����c�x�r�{͉Hn��[4*�ϻ�퓄r����{��M{};�*`ls������ă �y.��qIZ�ҍϳ�I	���C�Ͱ��ZX��;(�
�~����C�Ϭ�@�ܩB����N:��?K]@���g�Ɲnŉ�b�F܆�El�o�A���b�S��ܣ���ΰ(:mQg�����y�����2t�h���Kzy�T��5>S�b"���c
+t�:G��p�������0�(I-/)�Ė;�6Ab\5�Ś�oNg�B��%W3e,4�8->� �� ��όƒ�?y������c[�k�7T�;D�k��V�� �E.H�!!�Ǩ�� r]��~�~z�|Xi8�`���Kk3��l��Q�{��Kkm3�]J/�
�~�+������u*�a0�J�����T/�3�H۲w�~�Q�ZZ����^����+ͺ�4�0�Nh �Ǘx�r�w{�ʯ���N��ǧq�Qly�])�wm���ޝ<&��$""b-�Ji��n}���sѝn'��u���F�w����Gn�6�(�K�k�������WB�z�W����?��D����JY����1��)w�s���	�6�#�~~�G�p�\��Ž8��X�X��W�������p�b�E��w J����^/;T]R��C���'�j/�T�7M��e�g�y��;���O��-����B���>q[��v͙n`+OP��[����yS���Ļ��,�y�D�:����7�T��G��S���t�����}m��&�0{��+�2������$Ojc9dj��	U���w)�V�K�&7��;�^�6ւ�)t�9w�AQI"���y��s���\�-L��P~359�k�<�hwч��N�^PM�d��S��z5�r0"�'��y��
_6yל�ڜ0��p_�%6��3�L|�lO4��^@�I��]ă�+�xyz,dV	�
0,3�����&C/'>��^߿U��>����"Xe��XNKC4V��87�����V�>˶��ϑ֦훐j7�Ԉ��<y�s���|��c���͖n�,�++��y����j���!�3��_k���15�-7K�d�x����Ŀ�sVܖ9�fZysQ"��d��5/u0�'�M�mqef"��� �<H�.4�z\h�뤰� s#�z���"��bF�qA��;S������d�g-���|<�)\9%H����V�ёK� <:�r��s����iDr��@�l����k���r'"<ۀ#��'� ����:��dnb�ǟ�+�ȃ$I�j�"}�rb����>�)ጯ�F�m��b��Xu�G�}� (�R	�7�G7�9��!=���at�>��(3���I���*w�9r�2I���7�4HSՅ�J����p����j��[E���ֻ�2�A�kh�2jN�ZB�m�1�Ě	��N������7)q���4^L���I��$���Q/4:�����:�:�W(����9]�/��m���w<�@c5���sh�ʎ߯�h�	�M�L�ɷ��lz\d�������O�w�~+Zm�FX1\�j{��:�]))Z�]�t�|z7�6/幕�ਝ���:$2A!U�,���eL��.��E�N�l�(��MZ���?0����v~�R�Lp#mn^��t���Zsݠ����Z8:�N����%��*|�'|���9�����H�#D�p3^-S��ra[��{��%g�~F[��=xA��}���X�~bzR�}��I<ࡢ&����6�s/�V�Mn��|�X�uR�$]�͖�zy�`�9K�����h�:Iʜ�	�)_1B�+�7o�T�������?b�O�>X$m�����T��VT��g=�� �&	��_ɒ�>�l� f���ˉ������:~��ǝ���<�?���:�k7�!b\����U��� @���!\��A��w��΁풉xkevp+��"	��dq�^��5.��4�����NÍ���D���~������8n���O�C����e� ��yB�/���n�j����V��a ;f}�+y<Y�TVQS�GZ�`5�:�y���vε��	�Y@̑�{]_ �<��qM�W��I�:"�_�s��أ�m_&�il�g("�CϮҳ���<��%f2�abSc*�ɂ+��bKn֍���	ٻ��N�!#�jebW&v�,Ԗ�@���R6��}��`S4g�sy����٘�g@o��S�lOV�,���^��R]�������k�Pt��[g�8t� `n�.���h;�a��p�����֮�<TJ��i����{a��(�n�u�a���I�͝T���C�H�����G]D`��\$"���*`�Jt�CnR_\�W�pE/89�]�y���߫��(��i�s���;G&Ғ��^�uG[K��u��)���8����JJ.�xz<��ǌn0�G�V��l�����fm�e�D�bϋ�����Q�0�qR�j��`�ώ5�ʒ&gj�.�%�Y,���ȏ
Z`m`Sh�cԍ��w?�ɪ�[eV
>�Q1&L��

a
\��:�A����� �ӍQ������J�'�G|Lz����
E߶6xi����`_m6���������w-#<��Χk5�?��ɕ���z�{5T���qi��C�i� [�OV���K�m�3����_߭��g���bśU�Q���'����J��V�B:�A�Yf���eS~e/�����/���a����h,�5�b����}���2��2��LfV��z�iU�fk���o��-���`����:�o_KӞ��Z�cg�\l������k��l�����A�i{��{�U^u�x��@�9JUC���O�M�M�-V��tFc?� �e�#.c�72H��<����0����+���^�2e��X%td݊�ZX���oq�S��l�T?�.@n�\_��`j��eǈ�>�-�^@-����c������*)��da�٫Z���|ر���X0>�5z��"�*	���L8Bz�l�
���}k'��UW�G�@�����Χ멆���Z��e�kem��\�Ϗ؎R��L�;�0�����>��;�k7�F��;3���لm�{��7�	����Y,P\��G�m��]�)�ޯϤ�l1�۰0^�VSj���XuiƊ����u�T��6݇�R-�ՈM�ثP�l�qh�o&̈́���*w?��Ƕ�=�.j�g�s�n��:Uk����¢(�������jKO������:��j�o��jK�0�7��1�ꨖ�>[�=��AU�k�:Z+0,V&(�A+��i���z܏LC6h��s��UYbZȂ՗�L��Y��9[k+@b
z�n���\���w��k@�Y�cfQ���L�
��6��]*s�֜���+<�T��gU�L��Zb<�
e	���q72�[+$�0Ȋq�r��vKA4�	n%7��������:�I�{��XL}2�9�pŻѓ��}��\^�3S��*D�^�	�R!�����k�b�wZ��$f�	�k���>C8 U@�d�e���bw�V ���T:���;u�w5Sx��C+mJ��yE����G�ڨ�e�w�_c֘�mF�D �^=�eRF�.�w��{�Ge�[7L��n]���	ƍ�?����!m@��|�GQ�IuO5�Yg����=l;O��0B�1gcb�{����*O$׀�=*�+{a�m�[�$ �2A�D�녺��=��o�zcPZ��!Z�W 2�Io�>��h�4�8¨GK"b��V����G٩ׄD51����s�v�g�jb�3�xգ;׸W6}M��AZY\:�.;�V0�	��ES@&����@,�%8����
��I�=�z˰�o��x�%[A�҃�u�e�$��͘�D����}����O�Qp ���~e%4X�p�	"����o��Z������+���Q'>bheBbOh~2ʷCYl�19B.�a��_���^�rr1W�E�Ƴɕ2�'���d�@>_ks�ҤVR{븢�{1:�;���h�u�K̶��;��1>�L�
��`�mQ{z�0;���"��l�g�Gl�`;��?>2��V��`���^��;�#X��+�`�2�����c6�Z���Ⱦ�Q8 �սC��3v;t��p^�;��9QN��@�e݌�J�*�<���~j�	5�keL�bRl��؀�^��F@�n�>� ��s,�៬�1���1/&#J��e3�F�֩���2��Z6ױ�V��3�l�ِ�5�F�w�Y�V��Mq<�Mc��P]�� -YSX&:��+���k��>p�a��[5�����d���w����4<^�an��_�-�L�Lk6I"���� 
�1ȯ�0����ٽ5���kNNU��n-bn!�:i����]6
�=sڗ���eX+��{���`�������~�V�b�X��?��I���Ý�_�ɍ�����-�Y���D���lw�^_˭�c6����MV1���t73�\�
r�� ��o{Z�DVcT���.�g}�Y'-+�C�z���b��
l�������(C��XSP�Q;�b��H����I�O��]T ���-dpV|���������0���:�6�s=X1�^ �.{� ��>����-�`(q��g\#���0E����}c��F�^�����B���W��K�@�花�d�#�7��3)�\_I_X�+3>hSZ2�m^�B�
H�H���tc�60p� �����(�-U;ۖd�K<�����XOr����0�/�/��S��|���5W:t��d���o=�^St��B�b�G
*�Ω$
��@6�6�*#>9�����!&�� �Ί�4)6z��F�vf'�2;;e<���Z~ү��v�=xH��k=���#-��R����-v;�4�J�صn�([��1���%���[$���"�ϟ`d5ݵle�v��ǁ2 �w~앵5�6�l98�g2����t4��єeIY�b���?�I�ƅ>��W�
���P�[��K̯���h������)m��3cR`�c0E�p)���1"���2�d���a�(�ؓ�7��1#+BaX��� ?3�Њ�� ��e�<��2`F��D�)�u��fw��K{�A7k����E��i��ى���Q�G���ʬ,�X���4�`��J��+�+`l��Y���HCjT��j�'��Gv�I ��-6+i�E�1�_%�5e��on��D'��ϲ�����٘�F����� do���?�z몂�~ce�����,w�~��4��e<���"��]�"�|q�*�@˚*���(c��K�� Y�&յF�/�s��K��t��5�Tй�w����,�zez��ɜ�F��x���FxV8%��4J`����ۿ����{�V���F�ʺ��n��"�%2l�H�$n����lp{�^��6q�8TA�˧�c�5X9<���t^�<CE���>���gv/-����l�y�mVr�md�*6>�� �bM����|�:�8�v����n9U-��L�v���<�}T�")����@wL �:2&�{�X���šNq�^���������K$<!�=&�Xti
�Р�ި<j"���M,h��[Ϟ�!���`0J�P$>g�B��aѰ)8��Y*�����5v�j�����~#��s� Ys��;��z:ޯ՘,��^�-�7�� �Ǖ�j�s �h>�s5:(����Fb�Fw�8.�lF����R�o�~��(�:�cPɲ�Y�׼�k�[�vDGcS6b+	,�;?�hu<��0ϏS&ǌkhQ%O	�q����^��:�w������k�_��hp/J�"���챋3��k��g��`-�N������S�H��h���y�F�������V����浯.e����d#��a����zA7`3e�1t?S��ÿ�W)����OV���<yX��P?;A�A�61�ٽ��`}���l����El���QۦoX#c�ɇ�bA��\���^F�6��Ɔ���0X�t��e�<\ 
!"Ļ�K;�""��m����4��J� ��ũ衵��x�i�v�'���䢗z�=�D��am��<��Q$s�R`���{��!V֌����욲� ����(BM�6�x=?gK%�ù��374!�+�0/g�0 �Ѽx������ ��N��FY���ZCun��PU#�^m���d��e�ǥ��s����n��<���j���!X!`q�ݵM�`u;}�eS���H!r���d�,��$R2���uU{�#�� �Jr�[�����d��$��>q�v�Th<���y�k���]���d+�3-X�o��%ť��������:��a����� P���:�ҧ���Bqy] �Y�V��j���[3�N	4`�(�����|��������3$Iӥ25�(� ���|����'}�����?���Q�l�f�K�*�EH�7\T���z��)�Gl�n��<�ҏ:6��jŅ)!���ʉ��7��\���}xJ>��9����8&R؞��U<@t� e�(�fg*jL����т���t7L-�&��H-̫J�ji���?�n���քV���B��KtQ�8B\����k��:Y��Gl����y7���R�Fj��o~V�7o��)�� Gd_��tq�ȶA��]I�ݖ.P��6xQ��z���� �V,�B��;�~�K}�_|�+�[pX��Z[�)$xnɌFM��cRBB�u�
2(}S&�s����jbٿ�	�����)R� ���e}{'�?����(�z��3t����[�Z+��(��~��Z�k�3
��~yJA(�	{%B_:~x�<�]�Anp�^Z�8X�u	��a۶s�c�c�F��k�}�ƈF��'�E���G��5��ve�ʑZ�c����'��
��N.[M����7����Q+�1���+#-��<H�Ǿ&�}�t��~�4�c�<j�Jr���6����O����p/?-��z�����ѹ��[�&C�(��b�u�
�	m��<��3lL~�u���*��V�FK��*���*��S�|����@'���`�=�:+9Q�YיԶ���MZ�1pmq)<zX$0t:=�6���zγ�>H8���>��C��Q! �BݫW������v�x�/.�"n�]����Z?����J~���'�@��p Nv�P��%X�m­yL�Y=ȏ�k�_<�d7e���s�j�����֛�/tQ���R��F�TA���yzfȖj]7	�Bk9W�6����X�%��ۡŵZӇՒɓY�����1�n���q�Gs��a�y��t7z���@�\�R�����:P�ʐ�+�Sp���w���c?0E0�ӳ�\���D�[E�)b3�Ģ��Q��lD�&�L��I�秮P�s��Q`�RZ��Z���>�Lg��ց�d0!��Y	�C��{�"�~�x.̔�K\vZ��kǔ�$�ŷ	�&�+\�d:�x=�mc���"v'E�]ڞ��-��ҳ���R�������1���vk;�A�./�F�H��Kit�L�n�B���	�&�6D�[l�������N�'�cc솪7���ӡ�go�&�<n�ֱ����h��uN�^R���T�y*�V`�r?(�p+$eo`(R�B��!�sR� T@��}�M��n �>P5[��Ko8�O��CA�T�h���!�l�Ԗ4�z�ߨ�y�	5z���阌�Zj���v�L`���!�c���������e�t�3lBw��y�l�����ޭ�����h��.Vo.��:�3Jg�e�
���v)�o:l�Tw��N#�]=��pe����e�uFb��ny/WՅ���%v�X�
j+����L@kne�jPv��ѫ�e���Ο1�7�����㹮���Vr���앭)J)��Xneį�^�]>Ah�k3�W̙����umn���ѥB��!י���y�0>��k.�C��:	���.�~��k. �,o��.�����~�zH��8�\:��m�$�V�K>�}9���i<͈D: �'��4�g�6�m��lL�9�L�������j��� ��s�H�RvZ�܂�qk�PX#��nа,:c�#�妎Buek�f�m�0b��VΘ�Z=�'���f�(0�Ȥ��E�-嘸�u�9m4W�p_|v9<l��/{S���{�vj*1��D2u��u=�B*ix��P"�Q%���U����Ԏ������zA��o��m'�O��Z(!pK������k.(D����t�bU��G��[((���a�Hw,��]=��U
x�_��r1�31f}E�R:~����o>Ȼ�k�е#��J�x��) ���.zkI`;n��*[�̏�G��F�x�o�R7/}d���w�brn�f�߅/<�k�4�w�������J���J����V'c8?��nAa�XeV+<zC�����-������ K�E�g�\���l��2�tMQP{�����ה��ul�ܚ�Ȝ�Ţd���L.�����G��~T�Hٜ��[�1���٫+�Q���$��dG�S��?��޽��C���U���^܍�74.,셉?'�Ltp����.�'�XWa��1�y��woso�țk��%��HK�L���R�1㙅t	��]�q�m�i�=tF�o�E�L�z'�U�u�)���_J�FVŰ� ��s	�%�H@԰a�0{��;��۟L/�����r2��(�?m���K�-���-=��9���A$<��[ñ�:(̓�&{�e�
}��=��a���C7k�Z��w��rC
d:�yă���H2�@�%0 Pe0��oj7����ڞ?�Y*����?Y��L�M���ƁUAl�M�ƞ�ȧ�[@~Z?��v,
��MJ��td�%;J���
,�4��%ܕ���7�NG���K�����wj!�=���D���ƑUm�F����Uw#�-.��FhI�����ݘ�����,t�vˁ��xʓ�w���A�z�`��}�p8�NX������+�T0��çz-���}�����o�g/�Ե�W�����R�x���B8�~Q���~���q�E�D�N�;�'��O����������%�H)1��1<Tz�!co�>]oMܻ^��+�h��]�!AV�,�gB�J��.p��|V�c&g���Z��۟2�!.:�Is�{O�0=S�FK�lA� �y�<�fе%EVH�`S�d�Z�*6i�M��W6�8�V�s�̟�w<l�o�Lp��� �_��_���毕����|Jŏ�p������taC�a�X	(�Q<XUn<��K�+��,���tf�L�-�؈	'Q� �(�x�1�=�#�^F
tu����%`���VL��{U���{{�gL��]�
4+n,����C�:���xE���mh�'�u:�S��*Y�F�#۠�h��ܮ�V�Q�#�� l�v���� ~ j5����^��kT|�4V[���AA�����P��­�����]�$iQ���'|>��/� M�����B�Z#��.��2&6eޭ�hnt��,�zP�C��͛��g�|-/�.����{���S�0�\N`�8��7�d:��K}�m,�r��bAp[+�@�b5S�=�eM{siNr 67�GI��6[&C_��B�<�Q��֖0���B8*O���ۓ)O��8ؕ�ĝ�Q���䰙uʶv:�=(�r��xy��~P����|٫���'��? SgI#�m5�Hbw��Ƥf�A��:� ��}���'�gC��&�G�Ŷ촦�ѓ:>g�ťG�c�Xu���榈�z��)_ 5��Q»%;5�[�bI0���S�]�=L�
%�nY=r�7�/yѴ�u'5���[� �5���C 8��N�=i�L��V�O$Zra�	Bϸ[�]�馘� �����G�㞺2
}Q]��h�>���CG4�h�lE�;��5kSˋ�Q��ޢz]yL����"�O�+�f��2(�v�@�bg�b���LV�>�z��(cfJ��_��l ��^�CR`Y�)�����h�^� x���eG$h
��Υ��o^��+lw��[�����[�*H�WV����VX��3�v�楌fc��d\�56�QV�]��z��2�Ll|�XK����`s˥�!�w�M.�F�0]6�ʳ���h��5z2�Oſ�3�1�S�2��{����x�o��r~��D�$��g��O�'絏�59(J6(���ڴ>o���h�i�E�Nx4�ʰf�}����{��0?�;\��SMR{� ���]$̊�_v?c���U�kz����;򘙢Xט��'<N���3���,��f)����q&K��:۟n�~צ'J���`L����$.d=�/�w�[��Y��)�"-V��Pp�P���2�U6���E�
�f�#Q�HԔ끥+,zG�$���u�`�q���{ۼ:�n�=��:Y ��{c�;�>�Is����6QM�m��C��L��z#���Z�l�F�a�2����hx��|�:LP4E����.�N�Bn���YT��J����pn��Yt���ɍ׭^}�F�&{l\2;���٠�Aߋ,t��E52�*gj%�k�$/K)f�0�c���U	���D���N���\��g0�*Ȯ3c�,��Tdx�Y�Q/�%��:��Nr.��m#e���U��ak"�{�����j�X_M��P$ds����$ْk1�!Rg�VG�̅�A3����_��v��F#`����Ӣt���k�{DVc`�6C�P}��"#���|��>�T���a�,�"����p]�a�����ɠ�ԗ�V6ޝ�=zoqi|J��w�o��� $��or���6�-�!�kF*�/�g27�9�:�V����҆���},Fw+R�O� &��
g�[� ,{;V�?�I��W6$ۈei�ś�v]�϶͛/�X��4���v���`"��{�/B�#o�J{���;�7b�']a�w�_��jz7�6�Z##�{,ͣ��� �[�lWX�3�hH��}��Ҩa�kL���Aeaw�nS����dq|�#}p��{k}�*�*�#�XJ4?�puH��B4����|A,��~'��7�kx*MO������������>��k�/hW���gTm�4���"����#E�E�h�M��5!ѝ�0�N� �W�c�cd1B�%ڊtAbF��a�W�]���~�?���F//{a���"
����K,.�}��/Ch��#����x�w�-�S�n� pQ��#�ʍ����E�#���K㢲���H�:|�!�б|�떉��V��P@��!��4����O/Ӑ�_T3��d��e�t}�`�|9R.���"�9�*���=V_��p�YFŁ�	��+\a��e_�م���3���\I"�P��
ύ�\e_̽m*z5b���!m#" ?�|}�L
sϋ�
�il����<޶�R��4�$�X�\I���ޫ�jh~VS�j���
w��'>�[�/B�Sa�h�b��<t4<@���im(]�G�����G���r�R�g5h5X[�j�{���%I�4pA]�\�V��-��*����
����v;�])�&*�Ɇ�(@�a�b�Ë�����I6T��{�i��/��g�π7�>���q�B��<��|��x�L#�)��K/`0�2��k���4���5�r<�f�(%�\���nD��ҟ �o���@,ئ��j�;QJIh�5�Y��֠�Vz�4���ʍz�L��RIѱ\CX�z��^�F���r'��,rYJ5`��� >Y��_]/;K�F��KL��Y��V�Q��1.wɽ���hÈ@�EI'����dA��;�Qc�7q,����<n����,��:�XPё�:�����d~��)�3 ���EO�K�ɇ�qPx��ֿ�Ȉ��=��r���Y��2^b�4�	0��&u4�eQ	�q˝g�c�o�X��|e/?r�;��EA��*CX{I����?�t9���ٌ�B�h.U���gA
Fs��@�Uf��Z�i��}VC�6�f�i1�uY���Q��y����xo찖�kw���#�ɈpJ�9�β�<�|N�H��^�p�<Y@)}�lȁ���P3n�U�ٽ9dU��>����>�H��(�J������}���	��x�	�:�R�SK�J�H����nT?�iܻCgk#yBEB�6�����������v�?c��`%��N���h������&�L]��Sķ��1,s�#����0��(��{)@�S0j$|�0�����x�v�o�d'	O���4���}u�	�°�����d�P�&�'%qV�:Y��ul �Xlx �p@ �2�<�9�n����� �F趘�s�FD(ނ���J�����d�A
R���9�$Q��<����P�a��X�1�����9
�Oۍ��g:Ѓ��E�����q�t��̃C�3�����ŔY94x���vd�jP�]�r�6YAKFH�%8ܳ���4�&��A�;SFqx���i��1DK=�5��V��̰
��n�҅�������0r�e1���\�R��aL�UC����e3�*�i4�)l}��G��[2y.b�>�����°�H������.��0�����L��t&�O#�)����vŖ��fK3��M��p>����:|��3nu��\���[Y3c��ʦ�]�������)��&�y�9�lr,��	����g+y'���O��q��Q���:�����M�M����P�h����@҅.�D%�E�PFȆ���#H���w�>��7��|���$v�c�|�{ �˭�\ch��^�;�^�3Oʳanĸ9�> �!̈��syؗ�K��4���C������v���f{�O��G�Mz3H=�zjHB�5��P���L�maMC����d�X�P����޷���Qs��^��*7X���<g)(��4Q����qϵ�q|>:5!��^���ŃnNvwε�b�������r���e�Ww� #8"�HHr�\�?ֽM��<'{kC{�%�x��f�y���1�Ҽa+x�~Ș���#��]&*��4���u#�ӻq�'(�k���q�A�1*� ���㘺�Mj#���&㦳
����qS3��������|�/�Y2k.2��uI9����d��j�%n ���s���牏q��c����1��˿+"Tͣ��%hٯұ�x�>�K� ��
�X`�JisR�����|g� r�.�P�H~�.�,#�_�7��Z�9O?@���K�b�z�N^��n�[�?�`�Ы!�ACb��'KY]]�Ww��n��|$�g�ɠ_�(���\����~�7�?pfЏt�;�z�����"6C�\;�����y=V���4��2��Ƭu���)!����}��/�U�����;�ƍS�|HZ��k7I$\��{�b��r�bT���A��u�b/��"L�.ݔ<ꡎ[ʞ�3/1�ђo������XL�\H[���{(�в�>��W(����;�p�zb��M�#�-
ީ~�S�N���R����$Bp��S� �)g�'
�����+eT\�|��Ќ�����h����04�ga؊"�c�i��>�΋���t�'�k�ׯ��q�<������m��1�|z�0f�y�l,�e�<&[\8����f��4�u��2ϙ�kg����ć��Ê�wQ�C��Kc=�����i���Z�ٮ$^���h�� H��[�I�u�z	}|��ۙ,���y�R2~��;��wW�g�렶qZ���[��_��V�;l��兒�������b|G�f��͇g�,;��J����j�A��W�]W*�j6�nZrY��>*m������ׇl���u��d��H��3�f��`CÝ<���ݠٿ�+�a�AɌh��=�A�k���o*�������=��A�ϻtN"�[��SHlm4�P�F$����;���C�pѵ�Ѹu=TAt�~u���r"�cX�����i8��[r��Et8�^dH�j�E�b�����5]��b\�A,[i�M�4�v�x:�ߛ��?u���j���ar6o���q`�F��L
�� g7%R-֟;��a���r�8c��I��'�1EHM�a����#����5�<̻x�j�"L�Le��LV+�=�������;Y/�r;����kzzO��8A�K���w�Ï?����F�W�,пx��_�����%hI��	T`gSv\?�
E؅�2s�
���xd#L�!kF���6�T9��LJ�iΫ��LB89m��l^rU�����:�}�l4���9������<�9��W	��ܚ�c��:�!}�s7�_|Syeڨ[����	�_h���E5J����evx�W��u-L���
x����p/�Vg���a"��Tm8]W��ߩ�������iM\:ϕ�6�-���tÿc�.������)Ӏbą^��_����&�� ***���gj'yش�������w�Vɠ���%3�Y�聫����
��H�3���g����ϖ��t:��dO�~(�d-�Sr�/��2��^��1I!G���a��0���h�G��B����R�˕��n�"���Y�HqS��z�A��Tn~x+G$N�L�0���O��ݭ\ݼ�]n��w�ϟ��>��;������Y�f���u��k�l�«��\�"���[�aa�,?�&�����B�����v̸)ޑ),f���@ǱRK�����i�]�̚�>N:�^��ü�������0�[���x|�, OTx�0PYҨ���}�����zv�y��q�r��:>{��ݸ�6#�6�y��h��˺{	y���d���շ��j�6�\��NW�'3���uq!3�nx��6��$>J�q�a���H�Q�$ٯ�����߯��i�F\�J���0��F4����541�;`�'Y�(b�F��h8�y�8!Q?
yn�d�A�5�+Ak�ܜx�l��F�����)D~�$ǋ� wx�\��p��b!=?f��Y�/y-�F��6�.9�=�������^��f�~���j����ie��7K?���@W	� P	��~�����N����_��G����l(�3�^�q��Q��ƞϞ�8�f�s.�H�k�mM����V����Vs�=a1�j�,=�� Fi�n�|rhƼ�J?���~��.W��6{倭��p3"'�[�k�L4�k��9鼶��$�!vHڔ�
>G�+^ms��D�S�̥a�e4��#i8��q�&Cb)�Ƥ.MN��RG�9�Q_��HY`?ϭ.��,�Hw��^z.v�F{��Ɂ(׺�rxm>(1H~�����\<����	�?��!�2����&a�V��������<S�_��xJz>��TE8����dtL������nԫ�i^�H��+=�dV�iᡕ���\D���aUx���0��E�f+y,c�mm�5�C+C?չ�iX*�����/w��5�{���(�k���@M�/w���dj�lX��Q^��>??���_�|�_�R��zsK��j9�����(%��-K���)�ea���J�� Xr��%�Q����ҙnP��f�ַӊ����X�g��%�� \ЋB�_|�z7���G �������(($h�i��<SxD8�����%lx�2��N����Ȁ�����=J��qZB��%BP�;.���#��6�+�:�Lc'�Va�E�<~���V<_�r�_��&�V�Z����]D^��r1�EX�� %N��V�W�G�'�CQ����?^���{K�[���W�j�S���&��|:$�d� p�u������<|N$��h�g�r4>їr:�m�3O*�O�3��hM�q�h��[��_��>b��(m���$��z���1���Sk�c�^`v���T2���7O����T}��D���J^���&WW��r>�Y	��կcùJ&��,�ޒ,P9AU%�ݙ_g��SG����\da�j�Y�o�UQJw�=hm
�«A�$��TA��B�"�b�'RT����osg�#cPG8^Tg�2�֖0��l1�k0���=�2uxY<�`t���C/����xI����qK�A{�55�1�浡b �l�I:�s�q ��z4t�-�|��͆�qX�s��2zi����vT I�� ^Za*�qH�����������-,�a���0��C�0VA��-m��qaY(ֿ2��C�"]`7��H&D���3t��~�@9��ھ�.���ōn�p����uC5$�㳼���dJ�(�����!����Bi48�j��P�_���]��+���ƸN���l��`�ċs�1�J���!������DQ ��H}��1g���q�v��!Q�\�A�75Ps�~��� �ܪpi)5vF�md���sxU�=��=g(��a�xf�����y�¨���P1�`�60E�����m=��[	K�8o�*[���̮]�f%��RL�v���XK� b���'6�*��M�WKI���B�5�!�3f�+�x��ۡ_Y�߄���$Wϵ�vxsֳĈ��`0l�v<��L{�T���9e��8��O��ŐA����8|�c���M�!���J���iJ��p�\T��
�Y�P�꿣禋8!�7��"^Q�.�q�m`�<n>�n}��~C
Ɔ��P��D���͸���vd�F�.B��<���OD96R��XC8��w1�sO�������h+V�����Jօ)�M���~8�MUD���5ngj����n�X�޳7QS��}F�n�]��uC��0��üE����2����9�>�]x���A�,��`�C���do�a�3�徑)2�A]�{].�$3n%��d�c�g�04"�W�&ǄA���Y�D3rn�9�;K�V���{�H��S�z�%v/�r84��UE��Əʳ�WR����?S�~6�29��жe~�lT#\���ʥ��h=�	�"��������:7VѰ	�HER��Ll��C��>!�������b��I���g~}��K°8�W
矇ia�W�C����<�
!�wNR�����o2nM:�̌�����͜dld5����!��{�1(y���'#a�d���S.��WY�ˁ��ϣ����W�0f��p
�����\��C����,0ʃ�^.?o�v��bɗ3M���p�U�O�/�YZ<�o�s����W"��#\�6�ĐJ��g�
n�*��fir;x���W<��ys�{��������IYy��n"�
�F�a���^�¢�ݳ�n�ck���bcR���~^c���!є���zHJ���X��<�r~����t����g7�+y�n͎i�ɂE���{ު����([����;;��ᓤՌ\��%]x$��L����<��<�ތ�u�3�8�PB�F���ލ{f�G�/�l�@n��p	�� G#%j~�u���R�Hn���dې-��{�v��~ˬ>/8��!a����86)��u���Q��:�_���\D
ظb}��ES���5,���&N$�a�H.��L.5�?�{�3p9��:����$�&�^[�]N���;$�-��8�}��CB�Q��5e���;-�~� Y6�r`=�H�)*�˽$���F�D���O$2d�4�g��o�(M맹��R1x��4B�4��dPK��j5��p�����P6N�Q�����|�D8)����
!�[,Y�vq�W{��U��Q���������������B��=�B7|�=J��"��'���ܨg���[����߽�Q�^_��0&S9�'GY&��Ѹ���Y�7��_�g��_?�g@y��%(-�2������&� ���m�S�����Ρ���+
�
��C �3�ǗA�/����̨�ƹ��e���v&C�Dҧ���uԈ�����<�1,m�u�x����͞�,���LP��t� #]Y�����D)_�� f2��|�Δ^2��U���ԏ�[x�"� 9`fn�x�H`'� @鿿�w�����^%=J�u-�v�]�'[������&i�y<�<�������i��C�T����AW2<4��h� �����̀�.�Co��
I*q�
���+3R�m��yF����W�C��7/5 ��u�)�p������/�c��\�(�NFi�U�!�g�0@�k!J�r�ҔQx��Ϛʱf�3[� ċ�Lw�+��CU�1R/���,�Ӌ�ۓ�N�������������7+�n��z�B?������NGyz�#I�_?}���_���^����<��4������c�,�7����pt�B�����7��
��N"��R�c�(1���N �\��pY����Z���5�[�-a2��K�i���J��h�;��UZ��~(��?�a9Q�"������!�Pߩ)3^��̓Rm�\�|�a���O��������D^�����E� �� exp�q�u)'U�r�M_�������]lg��w�V6jJ+�w�f�n���<Lo=����J�N�'m�),`0-�%�VR^a+��q��P��S�Q:tA$�.��0l(��^�ΐ1n�l�a��0��P��/X�̓��J�"kZ9�"��Pz�$�v^�$�\yP��.c������Z�)֑{k2�Hq{�+�P�ڟ�y�H���u�����?��[��~����r[�%mO��ye8�Ԑ���^��IZh�:�~����������/��i����@��~s+�Ŕк=uN"7W�*P��u��l� �er��m�(�b�#��(�&��F3nT=α7l��2������mq�<'�Z�T�PE��zuu����Z;��u��/����$cȥ�)y����+�H�u"d���3��!k"���#ri���<^z�����2���v��̏�\�y4>q��J㤉�N�!���չ"��jx~#4{��7���w�Uf��1ݟ�/+N0�zQ�!(D'E!g
$",�=��g8E�iH%Q��N���W�Ie=em8��=(&�B����}�Ѱ����=J��r@��fh hZ!zg$�T��M�I^�}�,��ʚ*�Q]�l�tgWo͔��6}C
�v"QdwBjP6��2�ټl%?�d�F�7�~����'����gy�\�����v���e}Y6�9@:l+�q.�:eo8�(n4D����ӽ4z�\�9'��R������o�,��vuB����0<��rZ?����C"f�CqBI)�J�;[��J�NT�z|.�i�9���6�ͱnz�Vmc������փ٣7�͎��9%#����%�Tx�b]�V��� ���ɸM,���6�����i�b]����ݼYZd�}v�.]>���Uv˚Қv�hL��S7��5��H������Y�/|x$�hj��(1�ώ��5�Vr���c$i�?��gC}�<z$��.���x6�3�l���{��	 `��No���Yi�zϧ�z[���O��~ ��٭��e _�����(&Et��U拾�JO�=o=Nmo����K�+l�b̈[7�D���b�3D<G6�s��h���l�K5��Y`8�n��5�c�?�q淪����ҲX/ZD�5c"A����0�m]�����@}����k+y������/��������[~���}'6�Y,Wl�]�W���cɊ��r�_�56C�X���3���qK��j���֬�r,[�5l-�����^��������5�f��`�lU2,�s����z�e�/04���B��h����Sم�$��R�_]k�d�ȀAG�c͕�D���{Y�*��A��}�j�	1�����̿�q�Ӝ�mW0�m���x�C��)�<��w7�sq�x���R@♕X|"޼䫐½��t������]�{�bT8-�SR؉ǲ�&.H���R��8F�0�)&�;��R���j��;�t���� bc�#�D��2�b���w���{'x��dy�_LjYe3`��eW� �A�8��Fb��Z�!�gY�m�����b���Nu��Y� ��I'�ֆ!�0�����Q��aa��g�kا{�����kK�|�O1N�	B]Xқ�}��XGs�d ��I��b�N//�gA���o��� k݀�W�����35X'����VL٥˕y�8�ը�ԫ{�\���A�P���ey��s�s�# ]j�
x��;�I�*�z��֤eԷ��4��0�j+�
a�DI��zb�p���'/��P���Cq��T�a�0�Xc�𜖩F����D��w��K��׎bxYԣ�¡�b��8����zT� T���ϠzY�{@؟}[�T�e0��>���66$۵��X��C��eb��.N�������J^P,�\j�e\���,> -�j��Lo�+� U:�;#Z2S��G��ش\P�T�N�Z��tF���Rb?�&Eax���P/�؇X��e�j����G��r���L7����4���]MW|>�B�O�X�
f}Ox��Bd�9uf�I�<Y+D���a��s�o��C��<S�S^�M#�b9K<�����L�A+��k���4�׽+3��m3�$��%���ϱ��&���!�=�N ��{�8� �h%x��E���������r�0���^�ܩ'V�&{�����T3T��޶��r��e�X]��������1W=;}=�d_�h�Ax�KfųeD�lj��S�z�<�0�:WS��Oe�0P�9���X����}���]��o�o`Tz�q"�8��pbW��~���TO��FKT|�zr	T��ƭ,Gޫ��(�O+q<� �L.��=av���鉱��5�J��1�t��6��a��0���8������@1�s��RFn������z�!�a����T��5���H]��A����3�{���QaA �D���`f-����uk�	��K�qd|N��dYT����2��N�+�D��.�����7���.iA;���xtX��������~l���;��N��?=�[�g84Gك�_Mt�ZC]���ݤ(�b,���1��L���r����<{�O|9��s���5�.�;��G�B�ƉU4@6�1���>יִ;��0_os޻�����*R�O��0�h:��To�������3族����G6�.��rVCUV6�,{s�¹�ɋ����� /�O��������_�Goqx�v)B��R&�! �g��(��i��`m�g�)�[�P�*�?b>�RQx1���-���:�gCh/Y�3T�Ѵ�p��h�[*��������c�׈_7:W�W���hh���5��&*���skm*��v �0'op������7�s�!F4ϖ�'#9�ج�[�!��+�o�+�8�r4,�@`�M�@��a
/�Y�lӋ
O�!a��������l[Y���|���x�-��ϵE_���*	�L�G��8��s`�R>����.2:!g���r�a�ՉB{����~��%
�j/4T�/
�7��X����,L<�͒��g�͉�����Y8������%i�"��rv�FL�� {+�v%���(��u�;]���$r�,|E�Z�3맵u����E+����'0�j����P6�nx�Ȁ�PK���x�$ �44�Iv�`�'����mN��1|LrlQ�n����0"B�	G k�Ѓ}�������z���/��t� O�찅g�A���//�j|��
���&�_�y||��v+��Gyy���n��|2��0�eMl��s�[� 19�a�����`U���ߗF��W2;�d�׻��&NV����0PC����/�#��*�Z�)�r*�xV%d�Y׆����N����n���N@��ݔ�9���?���A/�6��p��N[o)�g�S&=�Zjhߑ,��]7x�}_v-X����
�m����^��1X�z ���M����^Y0��4���l�3JyR���Qv��UX�d$�8.��ƹ�4��,�B��-V���c��9�P��x��!���Y�����w�k5<�<=<����7Ǔ�2���l&+]0t���O_�><(ƂZPN����s>S�N�M�Ps���3O��`�!��U���O�6��F
'��M���x�0��}�PR�I��vl|�]���l�֙]|��k����@���L*m����K�z4�-�G�gHK�{������������*\�y�(��C�L��=�/z��<�N�1-ۖ^5����>��&��3����٤{���i8��^]��vC�����OT����j�Ow�l�Sc`��ӂ�f�^�a��F���Rm�Q#��s�����-Ԭ,�F)U�6�ֹ��6�1�wF�.#��,�YN@�d�X����0�,��W��ګ��Dn�n��Uo�H�� ��T�d�����Ŝɔ���E�{�Px�>'��P���?6�ӼIOi�G88�G�Xo6f�k۟�sn���6��r��8GC1��C�=�i y��͐ѴT�Ճi�xd%/�8�2U�ޕ+��1:1��?~�M�c���λ�D���ٔ�DÏTz+3��]!�xĀdlT(F�a�.��zd�\�Q�W˻\�ݞt�\�Gp{s#+��u�Vr��E�h'�uCSl��ޛy ���i����Ȭ7U	|>z��'�4i����
�zv�tj]p����I���5�Ȓ�@�!��M�}S/���V���=��9��
%h��EP7�gq�q��$��J�q�lDh��]P����,�*j����r��+HX���ʊ�"�
 ,-�@� ���0�=SW8�2㑹G���/��77�H=����9�N  ��ڂ"����M��p�Ǐ�~oƭo�k�`�тg
B�Վ6rF�
��z���J'$���S,Q�J��&+�Yզ��^�z�U�]��ӓ�u>n��]�4T]���Z���TKf��Hb^z�䣪0�7�������i�O���7[9?��cY����!��:���D&�%�C�l*�r*��Z�~�J���������6lMY��N[���˚�[R�I��;bnM��l��F.[�9�R~�ʞ`�N��6=�y �YO+
��W'2��8��<Q�f7�KO=�����m��b���h���t���� O^Z�p�Z��u�Kw�?�-�j(�򮜳����ZOW����Lx��#p��ky׻�H�A��XS6�$,pF3EȤF�N�����׃.�s��N l��r�1t��x5�/��ł �8�4Ԃ���B��bv��z.�l!��E}䓾w�F�<:<xt�ֳ��[��Д�$��hԯ��G��`��ֿ���;dI�k�ޢ/8����VYay��q�%�|�6גX����γ��񿽾ᚂ��A7eRc߮^ޛ)�Z���>5`8�`���u��A�Q���ƷfL�0��	��`U gf­-��/Be�^;�|������	N�U�>��:�lW��v������պ����2J��L�Vk�J`�������ck�=�w����Eԃ^�����˞��roQ4�F+Dqaܦ���5;_/��>Qe��!��1��Yg�YW2�l�V���̔��2.�M�R��ɸM�sӍ��	�r]�Õ�݀k�^"r0#�W̋+Bƨ	��7$.,c(R1���$6��Z����oo����
�#{[�xQ��%��$������	�N-�#���ɰ�ڱ�����漗+5P�+y_��'��ޖ˘u�V^	�F��'4ew�﵅��r1�`a ��u�x�A=h��F߷��gѱ�*��uwE�M�;��W��)�,�_?�V�[F�w]���	��∧!�9gy;Y�Y��;��~#O�QO{.�F+h0~4X���2fz�������%�p��u�;Y���xo���k����%��� f�P�aiL�c��r����&��ï��ԏU1�ߝA:	jjDw��ul�h�	� ��'P�R7-����pX�p4�}V�W�����0���Ğ�.H�`E	��#15T��Jƙ��<B�$5& �= w�C�*�W�dB!���:��'�����3?�x,Aҹ\�gr��(s��!T��oNj���=���L(� krA�{�k���볍щ^�u==���P=���C|5Wc:���odv�RCw%|_�t�u�*3�O$i��	��U� a�y�Fo;��7.�#�� M"O+OYG?Ğ"{�u�� ��βq�Ntv<n���?���R-E�<��{����a0c�驐$��7�%h�Zy�P���!�غ��x �R_�NW,�B��_zk��J��;��`��M԰���t8�����%�r`D���ú��L0�x,��-���xsE�EPK7��A�r��2��lʽ1��vt�(0?��FNj6�'�����ƛ',�)u=�Y	c�뵞�����G����r�A���I>nɶ��[D�w.�� �AR���<z�:� �D���A���������ȼGf�;;�B�"�e+19�����;��;&D�Fױ✕~��C+��qA�V=��z=���������x�޼�poI��^C������n�G�<롱�ɗ�/���d�|��'O��馅aQ����D	�&4�F��2���Jㄤ�̂zB��*n��ab�0O0T$HN�.�����:,i��!�B-�#����~���=��0�<5z���w|�����c�er"��Uc��ګǷ���9Jq�Qȍ>�#DB����������T��HpI������"{1��nMW��� ��(u��h�̺[�e�L�E�g貅�J��1fK��A+���<}���L��`��،O�1\�5�h졃��?~�v�_d�*Ȯ����.�4\y��B��F�~����J����j!K��ۃdu�'�^"������G���e9���
��3߽^�4�a���{֌�\>YDd-l0<+�q)y�٣��:3�B��1�5�������	�RÍ�����^�=y�]�/�72��|P���A�'0JZ�� �p��^2e�3F�3�`? � ��� T;]�����6Ι%f�0,a�}�ec��@SW��`�C����hkw	j0Md�4U�~^i8�d�����blZ��0L�@>]7�5�ww��net�O����B��/Q��u�!d�J�,�&�h���O�Dbמ���g]�B7�jL&�(2=:Te�� �Y0����{$ԒZ�Y
Qc5���H"a}��OP`rR8�d�[�_��V�9-V��i�uOL�L�k5����h)&��6zg��(;���{����X�����t�!,.����*`��
���+�)e��l,9,䡟@��b��F`_���b�4�O9�%b��^��^%H��wS����W���b��+]P��[6-��q�g�~�^�9�SG���a�Эe@=-��亞�[���M�n2W�6#�C��I���8�@�}��<�
�Kr`�5�a�+��U�dL�.����~����� 𰢹K��;�AC� ���!�4bXQO�������k=I�f�` {���T7�n���?J	=�7k����zl+]��^�<�pdQ4՝ #
��0�ʏ{u��/4�tl���J�Y�P1C���	ei�g{�&�����d���ьĺ���Bћ���{��Vu,47/x��pu2�{����]
��4�0n�x���a���6[9��̎�0w�y��A�l�C^��(�9S������z�$�j@�ׂ�]Y5B[����@�	�]���'��ٌ0b�6�6i~��bJ������)�l�7��{/��$��%+�����dD*�����%���P��e�E��W5�}�ެ"��Yߋ�G�V<'����\z���3nxQ�!W9�0!���Q�Q���[�S`�ul�^Y�G	Lz��Do�*!xOa�"qAc*𰄡#�rpB�uS,�p,Q梋e�%Z�z_�]-������]�����'=��v/�A&(�4:e��z0j0n��n���0Y��vM�����x2����J�.ƥ�~:1� �$J�BޚY��y|�n�������ɾ����X3��7���� ���[�YHK=�s�K�"=[�m���x�d���lj�ԺU��Z
�@�b�&'������_�{|�+}���R�\�%w���}�,/H8 \�{@�~�/���쬔
O��"@��'fq;��^@>�k��dU�VI=;����Aui�����m��:�H�ueee����ذ� fx,UM�8*�b�������W�x6�*ɘ3�&8l�y�r"x���
���q/�s=\?��\�����C!z�k��;���M��e�������<Y��Z^�um$5�(�_p��>��AL���=��t�����:z�a��p*]W���%6�·�D�d&�
����U��M� ;�������'��\u4jp���O���;Oz]?�j�����O���qs�κ�?[��c��"����z�W_���xS`T7Jf��i0�T�,�i����[5,0D��k��w��	
��������J'o

�n�Jnr-W
�����ƫ�'%�޷��ota"};[�B�zх|��"LR�6���4�n���jmiw�Rb�_�`�0!�'7|c�� Wh|�w��)@�I�%4 ���� �֍��ނ�tE^��A���Ga|�s=���B��?���Y6�ϒk]�7�z27r�C\ȾT�Zy��cj��%�U*L��X��D6���4�e�ĺ>	,�l�D� =���ES���eWz�Sr�v#�f���;[m%_������$��J~�}'ǻG9������ֈ�E�1ʳu�F�6�!߲NX������5�oO�Cޚ��lFϘ�x $�|��0F���4�p��{��+��6�S6�:nb��Z#��u�!�pF�"��h*/��u#"x�Cz��+ԡ����g�a���vZ�p�� �|=G낉Ʃ��s�n�N�op�@'���L&'�A��> o<��z�hE�n���h�tse���JjHȧQBh|J7ݭ.�ܡ9'(���j�F���X��L�V%�G��z-�� E���D�J͇�J~Ұ�.�_�ߒ��fE�~~#t����:��n�y���ڲK3� �iQ�:!3<ǒ�\���a��NI���9��[�Y}������I_�^(1�l���y!х�ԅ�N�%;���5�Z��>ox$�L�rx���1)�W�xk������ E,ks��4E���[]��Q�%]�E6Y�L!�i:I�v��@�\�d}{-�j��ۻo�j ����Rr�B{s�ӻ��<0//�<���H,��Jf��I'��:�X=�B�%_���ŀs�<.HF\����{,��Ի6�l�[B�H��a��_c���3���k8'�O���͛e�؛�gL�S_��:cO���=���
�':7v�\�5�[���<zA�B�{���,f�r���|�C|YMI���\5�l�c�ըmv�LO�T�z�v�����T����FB�u�0v�U㋵ Fő���q�� #�_��B8���&IUÛ'�sFCo{�m�j�ɘG*S��}���
�֍}�
�1����<[V��l)�h؂������Z�o�Gg���ʡiG4�Eh���;xna�_�H��3C�w:��Q��7�ky���;���8��=��]x���yB�w��`q��n��u���}z�\2�`3n���U�԰��m���*&�j�g�N\�"����߁��G6IM	�A0Ҡz1��-ԃ��F��g��a��A���LtN��g����J7�X�(Ga70S�b!�ą���x���5�Ԑ��n�`�����nʵn�:^��-c�U;݌��[��c�IA]4��E��s#����$���F�i�v��/,��P����^"6�T,�f�oK01��u�2�IÒ�'�����P����T%���!)ݜ�l��"*���ѹУ~ޕ����`\��Xo�������1�5��A���s�؞axO��3,F	�J�jH�nO�L��k����Z��!s�^�kV��L�J?��!�#��%�l����C�f�;����P���NwP~�x�	ɢ��ǭ���t"��߽�!p���Y��#1ɉ���A��w�`�4s�p�"=�%�V�Ђ��G�*��/���m���y΍�_z�a�"W�';	��Lo�w�-���_�~�)�i��
\��xNNzBr�Ϧ����),)���9p��cT����
Lq��?��/�@~@���3`9̚B���|rz�� X���J�	�X���Yo�7t�H§�r/'6.�ՠ�'?u�
�	-�y�.d=	�Gè��wd��!;7�`�����Jne�F����ozWเ5_V�U��(9>4�q\ϓV]�4����0-A�t�ql>l��zq�Ylܛa��'�P�dψ,S}���$�_�(�z�7K=X��{�dyX�t�'�ھ]^� �|��L��5��X�ٛZ�΢��ܻN7�n,$O,I�0C�P���2�-Ў 8�d;������J-�����:?۳\���I��O��j�xD����`�4���[�?�m�5D��E!a�]� ��)u�&f����u�W�NM(ݪ�f�_�[�����jDO��^��UT��iy�D�FG�Y�Éa�kx>�e	�L�ª@Ͳz�S��+�wY�bp����U�%�S(�Ld?��a�p^Q���8U#�A��m�Pb⇆�g@b	 �|��j�#Z`��ut�L�D���0NM����A�	���3��w��^���������+ݠ�u��8�1����C�$�dV���d�OP�d*�0~�ۼEp�\ZǺ;Y�}��_�<�9BJ���.�Z7�l��I�j�L�� gѵ<��RO��.p��B����
�0(����N �_�]+X,\��ɣv-�~CCgN�g6�&`,Z��7���E�������s���}h��L
���h����D�R��$�]/�D�«p��.C�'O�ǀ������,A�7;����H#+
�ڌ0
Y.�;6aƺ@#�0�s}���Nvj0�@��P�v�!?/�|�ֽ |��B5�A��䰈+�yZR��%/�/)�m�9�	J�����R=�j#wꝽ�Y4�}e�B�`���VȽ'�]s:�Q/�5�"����q�Z��A�-�����'�?!d=譟ڣe��_�ԋ6�a�֍x'�B�AwS�FC�	�i��:Z��?�\�պ���0Cb__�u�)�:ڽ�7�UA¨E�
4�3��B�gJr);fqX.�p���i43e�0p<�T�8B%��[��1��bz��J�6���>�����an�t�O���-慑o�00���Wt7��]�4X-EϮ8��[�y��<���0�=>���2E��p��ܳNH��6��}y~${�˗/�j��^���ݏ����,2�
��F��F	KE������o/��PL|�#{3/jL����&(	um�R�0��Q lB-�i!�X��A�Bh����P��
/���z0P�<Of2>��R26L��f4��
�5��Pǅ6Yi�E#�,ױ_���@���d���F[5�z��:޿�~�k�s/����"PM4,d�p���
Y���-m�(l��z^Qd�r�'-�b�eHM�?yØD/ tB�CK�YG0�W���,y�Њ�>�~f�gk�E��n������:���)V#	���,�Ʈ4t���p�ko����������y��Kb�E�#�{fn�T͂{]{�/|e&�ڂj"	�7Q��2���F~�{G&�"T�9x��"�7V��R+�(@�R�g�d�vf�V�����V��-�h?�OБX΃�AS��="��fFi�Yߐ=ab˴�ʚs:N}mN�����8� ˦��}��gsY|Ǆ�,��l�Ɩh��R^[L�|��'�ӡq���T��E�B`C�D���$�B�.�:.%�r�b$W2�&E�2���,t=���@���a�Dnn�X�7�5���͌�`?�$3���q�(������Z7d�A�Xܨ��&�G��fOp٠0hfZ�R��,W��[�ή�l~\�����qg�R'|ރ����є9�7��j8����G����X�cy�<5:~���µ�!��o++�A�������e�R$a���1��=���^G��2?���F�<[�:���xfu.Xĭ����(W7k�R����>��L�H̺��pHӳLk;�ȳ�Ȇ?�@��Y�V^L���LO�e����O%��f���E�.Rjq����>�Y�\�D�wI�@���D�����Nc���Χ��YQ�c�o=�Ԙ�:�' Pu�����|�nHZ�<���� <'�Kr-u�Y*G���~@��~{v�V��^�1*�j����O����[�|` ��t<z��Jz��)P�Vsd�W\S3]X�3�\ջCV}��g$��Q����{�U�_�T��L�?۸�s�ꏡb����T��Ȃ�@cj���Z'��Ȃ��ɳ�0t<��z�̲X����ΐ�a�V26>i��P�Z��4��~����I=�B>���굮`b�Pm���0 9��:�i��ߐ؈&�gd� ��0���9� ����0�˚��rC�1Jq �c�������&,E�$�������JSsF����5a�B�(�t�͓�[eQ�[iH���f�<�i�J�u=���1�ձ����7����~w-���Z��y;Ȑ�jy��}EM.��� ��'�s~ܐ=����
U�3�̌���\2��H�agR�-8h=[�;�G��{~��%|����lW�ި�R{UJ�9B�D|�g�<0�G����j���GHA�Q�,���p���SgeR��&�d��7��B�Wy�i
�b��)k ��ÞXqw6܎
"��jIN�w�m����`�a� w��ek�����![�'9�Fϒ��@���O�aqO�w;#Л�ߙU/Viҩ�WoU<�/EȈ���h�H�ݹ,�%Q�����	㻘�y����`�Y��Q�L���b"8�R8a�h�����6n�~5 �)�������`��ehXI�o�샞�X{px��H��^Ð�5���9s0Q�UO�]Q���Y*��d����9,"�BX������1غ?R���^�Y�S��j	(*��}~��:MO���¤c`dq*1s���:�ZP�x�M�!"i$���@��b�o����4f�9��"g8����www����%�In�􋅈争X���$>��u���,)B��~>�3��w8����	�����::��0$��?������^�R���X�Kc@�y���S!n����w�|�{����]�)/g/�kf�9ƺ�q+�d;_��Ê��W�/n�.Z(!:s�p��F5`�T%t�RE�* t��: Ƴ��5��#�� �b��Vg��Om:dSB#��
}N*�h ʀ�m��l)1t���'k���?�Ia�cPY��m�,-s�L�0��O�Ճ|ɮ�b:o��B��Ϊ|��j�@��a>�a���Z�1o�gSn����J+��qQ,]|��[_���-bu��=u�?��X:۞=�������3Fa)z������L%�n�݌�4��N2���N+1�Y�B�V� xD�Qț�r�'bdDM����`�׺�����P��p������G��<k�#���ŀ����(�����/���͵K�$6Å��f��	��.�3�����z��T ��zƙ��-��G5�,��yV����0d�|��1�*�c�։.�3|����===9�h;xnы��L��x8���p��>�(.���!�$��˙��{%C^�|��@O��d����:���@M~[$t���T~X_�1o5������zS�-ʞ�B���b��y̯��V7)���O�mxo�ct��0u�^��#@l ��v09l�PK�������'T> <M�93�s��z�;)�]����1<����9�h��$�q�"!p:�xh�ڢ�~�IB�I��	y��]��[G�CXZs%xJ��:v�!b= Q�5TGD�l>��U9�$f�䚗(�������0�	Z�L?��f䭖���.�ɲ��AeY�@AR'�{T��qa�k�L��a~�g��[����S��{��O���
�	��
���P�x';��
�Xɍ��g֘Lt��湯=\��^^�S�e6Y�z;���a��t1 �8S\7г�d	�g�H�L��'���.4����O?I9]qcn5��[�\�	���[�uN@s�)t�6�����V(������4�=5�s�1E�Y\�RèA��-��w��e�"�V��u�K��K��0zq��]�u� �6���G�߽Q���eCc�Ul�քI(���\k�Z=_R�ꊌ�)3|-�n�i~X_�T~O{�FQ���ck��'�m4��ֶY��\�����o������ѷjH�T��)��C���P"������Ǌ���|�<���S��\v^��R�4ަ
#���ai`ΕU? ���ۂ${:�tֵ>�V�ޙ��l�,��E��a��ؘ��
�E�9��$:(M�`��6AAJ!�a���u�35n��\7�mVԎ{�k�����Iu�d,�|�M���snd��m�:����õTY��\5�z˺^"��Hq�>FL�]h��zi��h59Y.\�	�y����Q��?Ӹu�\?r3l�x���-'-U0l������S%t=,�߻VH�dK�\����zV�T����B�k������	�̾�g=�����N>t�N�޾�w�ox�H��\���)�ȁL�^*�ۡe+}A%�e+{k��4�]�g����ֲZ�N����x{�v�����pzY��gݐ0l��"��v,�j�S��-�>jW损�X��l�ˑ$	#�ր�ya}29��	�4�H��x��>�!Ah5s�]X��V#�<B��S_m��g��T3V�d"��t�͐`I�%^�T=�:O�������`�%��uޯW���ݿ�� �ݪ�TO��w?�R��TVV�o�������&��N�e�+sbҿ�͊5��A[��	�R�8�I�N�\{���X_��ԆvOSc��O��`3�̨sqM���2i�[��o���4Ww��23Ľ	W��$c�gu�/ڐRH�^]ɭ�,�̚%n��В=;е�:�>�9���B��K�K��L,0����-�p�	�'JY�\���Z�_�!g�7˴`��9H!�6=<c�W���R$�/>�Ÿ۷�_�.Ov��#��5 K��F��3E�6���|^��t ��y��:ܥ�^����!ˁ�?�":%c�����>\���N��~���~��(���1@Tԁ.�ؼ���%�Y�&
4���&@U��U=x-�2z�r>�6����s9�����5�@��Qc$���q���yi�c�b��*jD�REAe ������y4���po����$�l֩�9� �IG0j�����!ݪ�"�ίË�g�AWkf�9�V�V�0�(�nu��	2J'�\�w�`�Q�tN<c��R����g)���!�P���O&���V�'T;9���l�y<b�Cc	,R~F�sMb_l��t��ܘy�c�s�7i/Jp!z���u�lO}���]T3��?AB���=q�U=e�-;��RQ�MQ�pN�l/�klz驅�;Cs!}�B����^��ǫI�A�5웬g�������Y�[s�޷�����afY��3�z��jY��ST��y�wv�.$������L�M$�p�!�X���]��N99u��Y
'����sWKS�R�m翽�T�[�n|���Ԩ��46�e�<[=57���ڤ��Aʮ�b�[�U��m?�L��ڵ�t�����蕞��x>��8AfH�r�$���Iz���ݫ�k=�:fY����'`.�9��"]q}  ��Z�`� ����F�]5j0hu�>.�mہ���~~���ɂ ��KS ��0T�P�Ǥ������|����^e鵽��A:�;q���,DĂ#�Kl�7�Bw�'wl���:[��
 @�C��!B"��uCLuu�c�$������Go|�#��{�����롪��ՍՀ̐}�k��?���}��j��s��Ut\7F<��'�t!+����%���e�:�s� |j�l��e�3�FxEԂ5�=ꀖL�dkx6�ɕ!S�H4��.��0h��R���#Ja�u�lE��a�Zx�ꡡl��9Vsyw���+=��3�RϸZN��r�a��߁��ʲ�$��,�G��~w��8`���F>=>�="�ѐ�nFm>���I��Hc�:��+�����nt/^���"���Y:�d��y�dk�#�9�#�����Ը(�j;*<���FxP����]�)o����G������7����m��K�z#�V�i�A[��H�L�ٽ�N��L�1��,�_D�V��ga��:	/��_�<�O?�d}���=�p³.(��t	��<3�Il��3�q��_�k{f�Gd���QC8�-�O�d6�`+���?�L���ȟ��㢶2 ��	�������;z�q�,�tx2���H$4.,:�r2&p'��7TM�^�X���4Q��F�����@2���T��KD2�t�\��2eKAh�]��E��t5��n��|���@/#dw��ҰQr9���� ��>��O4Vg4qy4���q"nC1�r�p	J$_���dYY�k�J�k8p���=)A���Q]��s����UN ��0���y�M�����~�}AR;�R����r���J��(4h�b��q �O��YrӲڢ4�t��%�%�[����3�*�o��<����nK�B�[k�5�sb}���P}w�߿<?���Z/O�q� ����@��։�p��G[�r����2a��$`z�����~�ð��4��[2���b��ɸM�7�FH�Y��'�"��S���>�8iw�A6�HS<�,B�K1+�^. O�wd�[a�e`��NQJ��t�uZ�+V��<�{:Hu����� T� �i�t��ǭ�yײ̈,j4e����c	ӧAg�jYM�X�e�0�����nff��`<#Dzx�Q�|�ʱ�����P�����_�CZ�:�٧�BLzi���΂2���H�qCb�T��`�{]jH���
E�{`q~- �xsܿ�����O�)��  'P��0��w����q��������r}=��zۛbG�Z�[�6��Ywh*S���B�e��,�ߟ��-�<��{�8��?�����;�ײZ_Y�]î#MKW�g��]�kU��N�k�!���E�u*��h�ބH�6j�1]�y8JeV����s��I����-{��Z"J�~pL�ɸdb2鬿��=.����~����=t�ZθO`�kd~Y!P0�����ߘT�}i�J�=����v��|�kL6��t9:�ف%z�"�=9��:ƱRG�s����WbB�hۊ�Ԝ/�,-���ξ�{�&���y�m�����!N,8_����	��a�~<N�G; ��Vj�G��1�t��"m��M��l�[x/+���f՘qk�wRw��B�:!���K}ӄ�mL�Ck'*?Y\/^�l�z���Pl�ݱ�
7-�DI]�0j���
��FL$������*���+[���VZ�Ɏp�5���֥�q?��� ��ˆ>��O��P��ᆘ_j��2��z{D!�m��xꂣTٸQ��x������n@�A6��p,�t��nٝn��)[�y*5����u)
2 �� �wA;�ȠGm(�n��O�~���&ơ����i�C�� �8�J��e�j�ݚA�c�vX��50l�5�yZm�;㣣β�umz�����6[)N�y]Ty4��)����3�P�َ�W�ǠNW,�Hg"X�NV��zg;}��H����Z����fR�`Ѓ��5VyU:�-O�/@	������X[��P~����GO�����J>�X{q:II%d@<0�(G��	�0x�\���VLф^{a�A��E��m����:�6��|?�N]�l�~���g�/�io2�"2~�������A0�e_Z�%���ϐ=�-�ș)k���λʎ�$�&GS߅N�Lm:5�b��f��'�|��wo?ȇ�7o�I�FL�V�N�L&$i5��f:�\0���p�3�D��y���@d�w�X�� ;��^v�����?ȧO��ݾ�齮��)zA��j��#v��p�2��&�v���}�ԕ�)u�D!c�cw�FUC��WYX��$t������u[�ۖ��i)�κ�SC���d.�J{��z�P�`�G�b��b%VȺn����k�`���Uz'K5�� >}�J���=0 w5���E��o(�OyG6��7����t�α�a�,�Op�!�� ټ-4j�����Y�2��T�S�7�<�A/�k��4[o��;u%E/	�ª�Q/�\O|���������{�
��O�+�K��~I�EeʪX��G*X�u�7=n�4r�A�M`�����{��Ǿ0�HfsY�g�εXH��4ͤҽs�{���T?O��5Y�$�K�Ӧ��i��d��`}�q[�Q{VK��q�2g5����I:�-��:n��z#��\v�z�z��8�u�4���Y�P䨨��^01E���LY3���?�8vtp�,\���;������w�����������uf�z+%Ib[(M��Æ�io��A�Y�F�����Ef��(]��g`l�����p��JLC@{�|�{ʶ{=���������W�5��
�U�}0>rA�q�7c��l���`�b	ɮ���3�j�L[�#9�%�+3�bU�[T�t"���8�"����d+;��S#��r�	 �N7g�vo�y颈h��S��� ��Ԕ�QO�9ORx�1���T�Qʑ��3[6`�qo�</p����|a����tgR̬5�u�,Qo��O���Y
��Em5���~��C�I�-��
 ��ࢉ'fr����t6sr4��+aM(
�Q�pD�&��)�U�Ƥ�� �un2�Ǯa/T���v�P�s�QV�2�^̰y��'y�):�fx��d�0~X?�:���7�"���&B)�r���t$������.Y��t;��}� ' 4e	��̊5j(M��c��8Z�c{��/�T�����z{u��֛��i� ��)x�7O:d�fݸg��.z�e�ă�<,.��80�AZ�^�o��7������F��Wj8����V����񧟙Uv��D��U����cbqƊ?��Y�3�];�\x*�Սܨ�>��tN��`�A��	��?r�FV]��Q�������lY�޷�	i�+��#�#@� ��'�yA#� B��������k҇�c�~�Z�Dd����F!qo��s��k/����No�MA1b�B����O��xd�,�ǝzW�h>��m���)�u#)��=�y/���˼���}Fw�J�=k���D;<���/ǂ΄�*�6Sj��%˕|:�q2ңKd	*c�D�m>�ƶ~��\��������ɢ�䥖7ɸ��>h�k��9�Z$o�K�yH�О���B���M���٦K2��*�DXFX0+[O^D�j���$����:�H�$nu�0�����3i��V� �y�M�C�>�V���v�2/	ܻN�m����=z�ʔR�w<k��w�er�E�AabY�Ģ�8Ⱦ�-�,P&�y���wV�C��B�I���'�F95t��XB}�O
qY�9k�*"��޸�K +�)��(����g�E��Y�pYxK q�����v��n�22in�<�U_)s���`闼D��z�R5������+e.�����>�����"S�u�:O35�>����M��3�k>����6}�<�Ϗ_Dw���ח�t�����������Nȱ2�~�!�{�N�I�#�Gm�rj��m6<'�����&c꫐��f�eh*:V��{FIa�3��ϖm�3yzq�T0�΋+yV����9+�b�ZGƤ,�i�dC~7Rl=�뜭eX��Z02�a�bK�s,�X���jѪ�L[�ѹ�SӜ����:WW)����\n�ȥz���s�%f�e��A��7}1��i�_Z��c���sjP��]�Õ��j�<*x�L�&�8��5��ѯa:{�����{��c��f%8˔�7���@��e����Û�����l@��!�E&/RX�Йޙ����������;x���(�	%aϸ�r^��	�ۅ�s�Vi�Շy_A�״�PGS-�8�.�Y��ϬV��f'0u���)������L� ��lHm�N��ѯ��$�"�LY�������Ȱ�tB1D�6�j�{�P&0����j�y���}��6�����OG�x�A��w�7�tg������Twm���b�(�6pKbZ3���v�Ho/���ޥK;M�|J���]��v�fp�W� �V>n^���Jo~�&]�b����(~��ߥ�}2�V4�G��l�p:w�F}e��G�[+E����ӓJ�I�	�/6�"��bX�k;����_��FcwRD.> "��\L�M�D�^K�K�}���O����F}��,�(]s�̀����B�̇�$9���J����W�̳�5�a��?��?>C�δ!��/���5�'Y�vT�c����W`%���u*�c�f��I�=��r3��;�>\��j!g��������}�d� ܭ���rfe��^o����@+w�N3j]@�)�yϒr�
HP&8#���}ɑe��L�"��G���g����g�Iw�]��n�]1l��>'X�:k�dNĄl�,���*�S��k�,������u�w�H?�Q�|!���{ჹ:��>���b>;�;���Rib��%b��u��y52�*̣S�>�҅ ?��x�3��B�,B@�:�h4$�$���oӇ��� i<X�%�^�P�,@8F��f~%#�o�n�;+]��$Yd��;j�z�=���>V��e1����������I���eXY5���n��A�RE����'Һ��4���:�#3ğ*L
���?���h�M�RQ�(k�tʏL�����Ґm�Z���E�s��]7�U������y ������6TfŬ��4v;����/VB��3f��9��<����l��t!���CArC]#f����>�<�'Tf�z��{��ש����>�Ab\��LyB�{�-��҂\=u��gp���ەL�V
�no4Y�y�����Y�Y�A<WAs^T
ݗ�=�!�����0=����rQ0��U�CIW��"G���wqOa�����s��k@�u�|Xs&�������R[p<��I�|���o\��>�!J��t��1�|I���~`��џ�0��T1�g���|�FIܫQ�@�4E�^�+'��5�g�H���,����G��ܾ��tm�(��"����ǩ�G��� я���m:���l	�Nm&ZPGf�&�`��e���[��������H(�RX�I1U�xXl���J�{+�Oi|{!�	8��r����,�n/nR��r��B�f�+Ed����$Z��|Q_�L D���tuycY���|&�đ�c�K�ԃ�e��� D��n��!H�R��^��yum��|k��9p�S ���\�w�s�0��d�A#yFFc[ezs�=�Tr��,]�a���G�(��f�ń���s ؈�RE���~�g¾����-�$G���������.Mn��\��%��_"�4���|l���>7v �$�d�괹���ݧ;e﷨RX����U�u��d�yVI�)@��y�ON>��v�:�$JZ�Iަ  �	?�����=*8H�ߍF��|�d1���Y�]Z�$�YL�'Y��ݑˌkY ąOm�v�=מ����h��_m? 3���S�΍���z�d�Ay�Q� :��V������v��uh�iB��6�L��"��R}Ad��#�-aU5.����W���6��ͦ���wN�q�">D𐁁h��cGYi����ǅ-(����en7�\�E�l��v��\���tm_<7��ŕD��'5�8q����(�K�~�J��zds��N*`r�A���S9���<�b>�Q�-�r�Ȝ��J���$5X��p��L��)��I�rC�`!�"�d��ܷ������呕tٰ�"G���v���e��W~�K�B���4�}%m^/����� %e�����g_3,�7gv�g����^�}�FK�<�j�b(�l�Ц�Œ� �_6��U��`V��ӟ�\�"I�]���o�h��`����Y�b�TdM�~*�e�����U?��d��D��G�~��R�������~-9����p�d�W<�i(�hT;A�ʀ���=�bM��,;�*��e��r�Lo�`}w}�?��_ν�S��lhF�6U�������}�❢�J�Zp�h��Ad�/�2@�L�q�OS�|�%��:�a�~]��K�J[��m�i{}�sM!Ћ���Z�l�C�ݧO�����ܺ8]*ɫ���Ԑ\*�F
]�4 -�������Q�i4M�(&O�ĳ�۬�yH?=}�bZ�Z����ΐJ^����
��SX�d�"j|:�i�SQ'j��;Ґ�G#R7�CWV���|��K��u�8��xO9�pq��UM������el�B�P��z"@�=���x6	��6�x� �;�|Å"�M�G�s�}�1�l��ѿyp��I���+i#�W1S�(c<a?'(C��SY���	DL9U�Y�K��v��&u�\��-B��@)���E��(���e���`�����rI�e��y+�vsi��r��k�����+��lr�<�MA|t���ʳ�7�j��Ѷ_>��x��EF�׷�����\>��^�J�����{�8ɒ�9}J2��Wt��wr%j��&}����!�}i�Ke�F��0�>�_��tx `gvPJ�LU�|�)���>c��/�O^d����WO@��I��On�+`�./,����j+��g�_O���(<�R��:�n�ұ9��m���;"	B��w�`>��|W[�Q1� �������Ϻo�����V��\�yE5�y�>��F Ք���G���e���2 R�no.���O���yI���~z��>�_t��'�\�vͦ���o���2��3�bN�k�>?�l��q��5�P��9E8�l�!'.	#;���6�M�#`6u˾t�z��蚉y��ǡ�E//�g n�QR�M���|�^dW���H�/�~��<MZs��e�$b��,�?���9��_z�9O�3��]�����5�ػa[���)C��n�g���Z�W�u��@΍+ܒq�~_�l�ٽ�ܦѲ�K�X�Ȁ�A�ݹth���V�$S��7���=�_t��Yp� �k���/��j>�C�A��N�0�����
��٪���ݧƧ��3O�ѷ,�Vn[��P���E��
ư.f㴰̔��x&�LY�S���0��Nٍxؘ9s���4^��=a�v��Ǥ��q���ah�����F�2�&7Ԏh�^�[c Wr���>���ПӾ��2��(2o�g�~��3��'z���-RI��yn!��E  ��D$�����?3L�vd)�چS�����e��Y
<=ֻ<
 өP[�W���Ս��i�����C�M��H��c+!�-�{ss+�r�:_v��[	�[:>���(��%#�����{a�� ¯�a�5����<��>e(T�F(�I:XzN����1}���5{���<�<m줲M��,����%$�A�CǢ���9#��Y����0] �5�������QX�Ss��$���gI������nP���4 ��I��������DM�&�CT����8�2͝��b��'C����W_��w)F���*}�����KQ�����(�-`0��F��g�d��R�,n�[; �>6�������©1���IĢ� V�T����3�'�@D�Ү��p;d�N���o�M��S:~yR�!���J���%@�G�1@����ɟ|fJ����-�ݯvy_&V6Zp~�{N���q6S��;_W���ɴ�l�W�R�pL��%�Qa�F�V϶酇[�<QY#ǅ�*�l��2���>d��l�4�hG�n8��~��8��;F�Vϝ�B��X;��̝��maYx5�ZPt����� ��ƭm��-��]�d<2p�m�E_�^���w�+zT�rl瘥���+���kO�{�*pЫU��a�j����x�>�.��EZ�fRcpw��y��O1���Yf�ڸ�v�g�����i��}ƻ����K*.U����a/����/O�⼔i#�ʯw� H�r��jXș͐U@��r.ys��Y��p!�=g|}VQ�~���H���X5��������͇��yv��I���vVEx>L���a�]YФ%qX��@�2�B��ͦC�ݫ!�ngj� l�D8=8K�4�`����TЛ,;G�˵cd[31�|N_��`kBs'<�.��I�w�xן�����t �X{��m����}h�@Z`#C,�!KZ�[�dlG{}��ݞ�:&1i��JbA8�T���t;�6�:�,�g"��҂�8],3��[b�m�lݺ�Vzn]�춍X[��j�:����ލcrp��:d�}x�g�u��0{��d����Bz�`��G@����Ӭ�un婵��bY��_ZL-�.oJ�z�_�-ل�)�.��Si�r��H~�L��Q�����Ý�_X�L�Pz�k6��\�O#��R\���<��5hn*;� ��}��G�L����<�)��Ǆ����$��3_�՛�_�M||N��Oµ1�lm�L���+����#b�GD@&�]��Uy�y��v'������Yw�MHjO>7�郓s"5�\�+C�F�Y�����N]��	����\�����*�vM���S	�:�ڇ~��L6k��ళl�͂i@OJ�D��3ɶ
N��þ�$z��m���+1=����͡w:V�2���(%&>Wӷ��F���=J��5|e����Q���j}��G�'W[1
�[]��)���&���H��)d}[O���v�is��Ȃ��t۝�RU(�d~){�܉I2t
��h%�=�@g�v¤��2Ԑ�$�� �����ԓ��q*�^Ӯ;O���v���~���h�S���ߣ.A��ն@�x�K��F�GɈ�u�,Ȏhg�ч��+ڮ��!�thG��2����ùI��@uT}��[y�e	�k��S�ą@6����(�>�*8gm̵����	T?�N���ʰ�X� �0��υ�T�٥�`�*�)Y^ 2qn<=#�Z�0FJ����U�L�N����T)i-�v����?����?�!=��e,�8��d�������K��3�gQX�P)��!�y����!��b�=S"(e��sw,�j�������9oT�KuB���t}�޿�{�I�t�	���s�O�9h�99����JX�g+l;�EoC-��:J ;���malW������l-����Ӛ8	�A�ƭ�dCɰ�썍I���l��m�d-��Z{.iA�|gȵJx���t�����g5�a��a�~X��+�~w���ƲL,c"\=YPK�l�����M����,�Da^>`�  ��AY���C�H%��ﴆ��o��ihZ��sL��d6���ɥ��h1qhʒ/��撫�>�Y�*?h�a����D;��_M\H�
':p��>���#A	 s��37[�V�7=��
��G-��Q�Ue���m���2=W�3���}�̋�W+�"dn�r�P�.�B/�3J3�����9�z�Ʊߟ��A��n��ۻ�R*2́�l^�?�ot�p���z���,���L� t������A9��@c�x�!R���q�	��M�Sԉ��A$�
QbR�t!C�YS+�ma�Ɠ�|��4�3 ��!pe*V�g�d���A/�\�fX�лKΦ@�k0� 
�FL��x�q=���ӕ?WU� �:�
�l��#pgd,��م�{����8���5��Z@P��\���Ɩq�6����}�!M1*%��/��e�o��JZϓT��\,�5O��Q�6�g�鬡G���C���z	�0���*���Ԛ��hj���~��y�J��8X��&n�M���?e�6���ڊS��JC�j�R	�B�W
v2j�k	��G;ZSp+�`(8�<N�Q[�
�:�*;Y�A�j��D��ZA�{IH�YJ�yT�E"�_>�5v�'v]��D��{ݹ%L� �W��ZA�h���1�������7�޻�ޤ]P��]��ұ-�pLY����.���7�-h�U�n��8�pHQ|���~��}���J.n�5#�By6O#/�	b��8[�'���#��7m�4���x��Qv	`Z�*�G�2ĩVV3����Uv�ޞ������S��AGjvͰ�s�JF�2�8au=#���*/SF�ZT=�<-c��ӿ�	m�|�߯c��
��ɛ�Ǚ\Ƥ�|�z��9���}�Y��_�'�Ge���I��K�b(d��32ZĴ�ı_�L��NϏ��(�]|9���F��'�|�&��/�J�X߿��(��c�R6:�{=��5��gv8�I�v���E�b,B��~�M/�i��Z��ϢC�bp}T�:��5#�g�9Jf	����l@î�� '5�&d��]�Q�.Y
pjwVQII'L�x]�6�9��A騁��`��"�2Lb�s���n1��Ժ��hZ����a�����IHŵ��6ɨJ��H�|�{`@�L�b)��Wj�IO~�~��[��dne��MyJF�Yz�\7�v l�%+'A7n���)��:�z~������J�;|H	\��"ρ��ڳ���FP ����̂�7�&�R����qw�*
��QC��43�U=[ֶY�h��aB���}�F�� % %.�?�������^Y[�['MK���\
	�Hʩo�pST5��Ќ!H�B�S�j�J�����^�W�z]���� �{P��$��=f��\���9�y��M0��7��mA������^�d쥛E���U&�F�\ؑM�>4�AΡ�#��F%�u�"ZG���u������^vO��~<��	B���b���bV6'�3�����M���7�ߥk��w/ϒ>��B���0�e�\vW���ػ�%�	�.F�V�Y㪁z�V��ə$TI�K ��QL��r���f�2��~ѿ�{  �҂ǒ����*�;�1,�,`�,�b<T-�ow���vr�o�����[3��ǳ�_��{k��L�?���U]�y���%�Z�?�s��8���"gLi��(0��о�l�����lK�B
�R�P��q�R4rb��}q�&.ox����%"�2�v+˵�O����Y%)��)\>)�2��RI����y��ҁ�>*n�"����O@�G;wm�OD����W�Oߕ� ��&f�N�pK�<?=��~�I��}���f��QZlC��<�:�Րiz�V�
(��ޅW��d�^����G�,i|fS�X ��)�_e��2��0�z��9��V�́�1t�L��ɟ�����!#���>�'9+~�^a�Z�c��3.Om�I!B��\T:���ٚ����Nk#ː�/�R�]�����S��������7�ٮ,ȝ+K�2Ⱥ��t����5,���Š�'���,��D�r��3�@Y�p��|x�NY�>�^\��WV�XV�����J_�F�r����	�K]�$\j�8fA��d���%A���tR+ �~`b�Ϭ�e�d6��\�O���ݡs�Jl�1X�}D4�B��i�w�2���������5������.��(R��L��7vK�3v���}��^pk7�N�Lhwq�P�d#H?zT��٭$O�s�JGw�s'�Hyn D��XP���OOǝ����:�R	EＺ+]y^q�Py�����GRr+e�nhl���� $I6��p�����KܻL'^�]��pQ��?z�?��s���:���Wui ��.��$��Xd 7����p츳>$�r��S�A=�(U�g�d��[��'�U��n�Ȯ^��Ԅ2��3'�l��Z���C	���� j6���+��+\�U	�#,PJ��d	�ᔞ���s�
�!}T�����u{YW�(����.{��{��[o^�<��P�_�A���њ�ؒ�OSe��p��^V�4ۼI��.қ�����%�1��lh>u�2���4�*d��|�}��e�:����С 3���wmZ\X�j ��m��TZ%��������6!`�ǋIzo��?�����U$��sZ_^��gX�1Y,�a������>*A��?2Z�c� ����0/ҷoo���WK
��M�˂5>-b������aׇ����]{|jw�3����y�hrl�l}t�2:�7�b� ��P�����yR~)��9t����q:G��RfI�@M'��8;Ț������6�P؜@��n")'������}ɷ�����mh'1������dA���6T�1�㴴sy}ez��v���˟e����D� 7s�Lf?�J�ESR�e��
G�3���I�gq��짘L/��##��g��Eߏ����jI���Wy���V挊�R.sphuWMw2��"�$�T�a(��
<��~3dG93�qyq=pM]�n��|���e�����Q^���b���0\,�Gb�՜�d� W;ç䞙e��iЃ�}T9�5��-�[\+2^�ͧ���� x��V������.�lwO۴�%0;lţ�ܿ�uyP�F#^�t����X�cuV.-8�pl�
Ң��b��	Ӗ����������v�jm��b*�R ���\k&ˢC�ͻZZ� �h�Ii}ܹP%�$�NsA|FQ:7R�A��+M����L�������&A�L�d�C���s��v�����"�k�:��j����%��p��*gD��ӴG�6e���vN���2������=�Y.:�'GT�k �{z|��
p���F�qiY��]����܊���h�PDvo򍻴�t}y�Ϳ}y��.#d�X�	��(Mil�0���ςI�E���:�O��y�O㶓�Li���L%�����.���GsR��f�V�
���ġ|��b�M-W-���T�>�EY��I��}I��GPxU22�\��م|�Fv� ��B����s����F2�A���~���p�z{���U���u5c���M���H���k�{l���3ȸ� �ϰQoo���d{�>��:�-��y3�5k�	�;���J�)>c6��B�@sPV0�}�K��k��r��������{I_[
��Mske���B������xP �A蓸�-��げ�����R�s���/�(g�'R�U���V���2*h�޽MvS���-��~)� �#u��1^�Ā-q��͇���ٳ��n˅��
!��K��#�?���݉�?b�S+Y��YB��a��ϓ!��Uw%fya���^V�����-_�/��Bo.*��P�]�w��U~��:C�3�h ����;�<w���|�0)ި�>����$��	��WǪ�>-�̭,kVG���=��"I�u���[+	��V�O�����/O�0�(��շn6@(Jw�i�=�E~�gBˋ	Sod�]�l��d��+SJϼ�IF���J8��*Nn�L�Hi������!Y��3�/56+ЏC蚱�x�c�7`s&2`�β7�犻}d<y��1f93�P�s���\��L��L��m�W�O̐�����à�N]Ri��d�N�lAR��,��I�T���&�^V�wח��Oݹ$S��d��>`/.jp���{�f�>h[}TtMA�Ogi�ڲ�[��"L��l�ҋ��[+wn�{].�e1kb�l��K�����>�	�ni�T�B;t7�/is�(E�_���E�����:�����Rk?�Z�G���2eA#I�2�S}�����@�Ͱ^tPr`�./�"��T2�]��ut��M��Jj4ܮ�.�Ȅ�s�T�����% ��/��a~PaG���X@!�y�����fgAm���YL��P��CR"�d�~�=-�@8i���̙���3�Ãk��C��Ju gb
�s��[5�/�M��2���q��Ke���<>Hl^�| y��5���'�����q>�$�,��d�i�+i<�iJ���Nb��t���]���|�|��S�A:]��	���p\��2��0kQ�$w)�&�p��_Ʀfa����g����W &�]����8�i�Ut��Z� T$��\W.6�Q��(r�)�4ٹ	sT1�Y��-W�I=X��޳�����7�a����)g��O9u��VkϨ�"y3��ʿ{�>U�H��!�e���|9(����U���P���N�b��I ���b�m��V^�i2N�0*$��k/��i1N/�v_>��l���*ɖ�;���O~��S�:�k� B��]�����˜ϖi7�u�vAR����C�qp.m��Y\��Y��0�/8��\��jUa��0��^��*�\�rXg]�C
��P2p�,�M+| ,���G�v�G�$ie�7eZ*|�o��~7P�T�zkS�n��9v~5a���\/�	��S�DTA���3�f��[+�/��mv�./��>&�Y`��6��k@?C` �`�Tr@�i�������ʣLp}�r0#���5�8e�ѷ�鐾֥xj���ɠ8�A	����^٢��0��{�yZj��Q̭�<�E٩���F'9���Ƃ�U)O첏湴�8�h��0����/ه�p������"c�	�I���� ��+۽Q5���S�������|�y�Ƒ����M'@&��2� 7X�@�:���{<�Yf������zdbdB<..��Xdݶzb2e��e0��|ڛ��~����}�����<?}�sm{<Y�IW��t�����:��<�ɏ�>[ ZK��|i�u-<Ze����Y
�
`Clf�#ê�n�uSI�K���p(˰����2j
��3�c�y�>�ւ|�S9�2���%W[I$�P�v��[��<�N���٭+��\8�X�R��N $���A)e\�{��ZKUy�
p��麆�j�}���>�J�=t!��}�I��m�|��������A��E	�k��|����c)12�oV�6d���;�ٕ͟��?mӯ|��̭�Z�Ȍ=�/;Ep�#�v�;��V��=byr�ƞ�l����S��G{��ЏSY
����lT*�=����b;{�	���2KG�K�h�UOp4>hQo�<�¢���f�H�.J�w�v�3�������-��/^ɡ�=��?@����r�SO���O)4#��P�������D46<�� A���߳2,?��:r�v^V�@<+*�,� ��We�̒k�4kw�Q��>�93�ku.x����E�t�-�.�������Bb��Go�dN�t�����\ۼ^�����6w*�����8]�ޤw��=�>�d�O/�e�����K���Щ�^��j���w�> K��g��j�~_��U0�wi{���l�ʂ`����û�ʬã�����zC=��e`dNR2�z$(H��F?�d�.T�g���w�T+�q��;)�tM����E,]�<d̳@��Z��EE�g�P��lX):�cY�ŝ{�R���f�9����SR&՗K���}(HJ/e�c�>N�@������3~������'����������2V���V�#�"�-B�K^#ƺ��8��*�q0\;�d�^H��"M^]^{�8 �.�5�\'0��v�.X�t5�--N�E	C�~W�S'onWڤ>�:�d��gJ���bcCP�[���l��!XfZIބ�QT��_yZX�L,�2F����ܗ��u���E��(�٫��E/����}��rN���:p'Y$�^��C���Y�){����9��������KH�9DP����SS�!�qv#�vS�9��I�)Lf��M�@�DnWV�q��p?!�_��N����ߨ�����=�Dմ  ��IDAT����V
!e��sK�c\��Zzr`6k+E�[��|4���7�
Ȼ;�D6�Ւ�A��R�!�]���X��a�0�����HT��llh_ @�GUNi}(�� S�{r�]�Ve�up�{2�^��֤ۮ�x���7a��%�\�?}��?��P���>������H�j%�D/���M$�ϫ����c�8f
�E,
���5�W$��;���Z�pA�0�'��U���m���r�m��$Ⱦ�(7��+��"y'�8�T��gy3K����\1�.̎`�M_紖�;EY8�{�-2���+ 1N��%��!Ӏ�޸����{'cS��-���&�H�<�tŏ?��'�1�*N\�S	���w��9�)0\M��뭞_����@}g��u��� c��¥б����(�(�L��3�̓L�,7��% �"�I��@���T+@�`�����$}1��u}*b|R]FpMC����\��du�8�k��x~Ѱ���8jޕ�k�<��`a�B��B���5�c��v��'��o�'�����xg�(H��J��^sz~1v`z�Z����+m�>���R=I��C�ru}�൵�0�ѩs�\&(���jJ�d��j���䛰Ɗ�ь�rV�?	��=5thQR��N�Af�F7rҺb�������)��l�~S�wI��¶/���%׼��,;�iS*����nh��&l��Z�
����9/l�ҳ�8�*'"�!	n���r�P�����(�~�ߥ��L��1��*H/E�x{M��>��έ�Dx�g"5RW�~�EӔ�m�z�1	}�K�M�_��4=�S����-`S,��r�B.��S��}��L�둸��/
$®Un�A����.t�#�i��zG��ɟ~��M_>�,$zO�*._^hڔ�`)�����{@�l�Qߜ�.�/����2;�<��~9��u3f��:G���`R����/7����=����!1�d \�yh�C��� pb���B���x��l�=��Ͻ�|m~�X;K;ܖ��6�9�	�j����ݠkН��y�f�=��
�J����R�C������H�,�[N�8/S�{�y��cz��`���;e}b�*eF�Ui��� �_�~- �����OS�A�*D�S_6<I�=dx978@i8�T���상ѵ�<)]�&�(],C�v�Q����S�K�H��)�BA�"�zfB��+�:I�ڹBuU���g�ItF��TV�QQ���G�� 	������s4.��F��1��ށ����[0�N{
�ĩ������ wί�:��)RC/5Z7�/�
'�^�U~�#�1j���f���F���C���LB����T8e %��ΐO����E�wrk�r<��ce��6\#��L8��}T9�A���.\�M��sa?�}����m�G,�����m4_=�sG"�A�zV���v�s�fCZ��8�����O9LjVP�����RD�p e6��i�C�z!! z	�A�@��P>sΆ2ؘ����{I���JϷz�P�:7�FJ�(����gPjxE� eTD^V;R>��!)����U"��Tw��d-��[73q��.˥K�H�iK{��Yښ򰚏��[��ӯw�U�>[ư�H���޼fܦ����أ�\9g�2�Z�GD���M���$���JO`"��i��f���	��c�{
.m�y�JPi/�F$Ƣ����R�Po�hv��Ҟ�N:��h�t�{�G*2��%���sG��!!KEw�d��� y�5ѯ| ����:�¨�d�n{�X����X���AG�p��+Q_A;q2�� �,���1���z��]Y��mQG0z8�,����`$iw�Bkaa����}fW��y{�;��Z�Y	Z�.wbA���2�l��,�ny��B��S3|����+��2'�1<3����;W�̆�=�IQ��P�xfdD��&�}�]�������Ч:W�8F/���id,DJM~/{�ff�����`b��2�V�<���OI����JA���ݦx�u��nvqJ�_z)d�q�����x>���g�6ׯ8)�d��4�������1iG�����/���)]]�{��uA ��#+��U��$�ͭ��|ӡ���K0*�y<��6\�*�Q���F�4�lD�ڂ��6�̟����鰲�a1IWdy�3#�b�Դ����jy�,�����.�l��Y�Cu�̔���#�Ry��#�pvm��0 a�W�Ր�l<���&�[��R�vV����� G%�l�=1OJw��Δ^�5�HS:l.�Є脘'��eLl���Č�D#Y![-��\,����r�ꂛ�=�W��2��:{p�׌�6���{.r@�^U$�P:6����W�����ƣ�]@���u���\)6xN�<ꝡ�M�7z]�f-)�7�l�j�s�-��4ѿ���h���|,\uޏˊ茉^����G��U���߹ЀUi�6�B}����D��\�L�d|��;I`����h:dA��L\S��+7��9v�b���+��
�l�㤆1��-G�/T*��4H�0j�1ܺ������+#�	��"�����i���3���[rI���<�)B������ ��=���Qӧ����I=��y���6(��e�vbH�)��[
 �<^Ǵ]��7��DV9�/�dd���m?��, �3ʗ�2���ez�@�~���2]֓����Z���tc��ś�����RL�̏�����{X!kE�< ɮSk�j}p+[���n)X�s�#�����S�?���8���������G�Ŵ;�N��l㚉9@�� �x��ߝ&�!k�D��V9�A�ރ����+r�d�͈v�T�x2Ӏpj���������)�|��t<VЇ®�]�M��hJW�C���X֎`
�n2{/�Au�>{��J��� %�N.�r�;oXk�!
��[lݶu:�#�E�v�L3�v������\�o�n&���9��`i������.����m��C/lKW��B��l=>�ۃ��u�e�V��,�M�6x��ѽ��G�-c�������(_{�����������s9���0W�i�n�,�j�Kmf����9ϱx�=�o��##̘3����NeiƤ��ʺo!d�N�&cs�։Y#��:W/�b:|>1��W>�eP�������uUk�W�D��1qS��t�שt/��-wz�֒2/��4m�/�i�|A#0��R)׻b�
�KJ���n�s�<�);��4�����=�ϖB�C��6��ڮ��&uv(τķ`3�:eǍ �U�!�x�{4�'T�ۃW;ɝ��v:�
�5�:'�I��T�4p�Qx��P��Npܤv�)��Ҵu��"�����&�D1B|5y�IS�ҡ+������d�L��H�پ�-ӷ�_+ʠ���%|2j;�n�\�w�v�!Ǵ�ؾ�Z�����٫�?��p}Ⱦ`|��[�¾ȃPo��&�DقE�'K���n,�q��d�*o�iR�����[���R�SkFdG�.��!N��Ӆ}R<Ke��s�>�X9+�k�#0f�RT���j�'D�v��)�V&��AQ�=2��\�	Xػ��γ�}�vYH�3�J���D�`�<U���v��^�qI�D�-7��#�^^�
:��~wԬ�Ѓˁ(����|o���E��:��� 0���~�!��୚�dp�f��\Y�w}kϽ�;�el6kW@ə�h:h��\i��~�yY�ۮH��4�|
���ʝj$(�K��['�saPB����(�ki����Ȣӛ�\�S������w��<Pg�s�=�GM9�R/zj�gzL/G�@�0�$�W���ޱtOR?��ʱx�J*��)���Vb6���mI3��Zr*�"#�̖�^:&��\���gyH?�1��W���Q�Z�!���Z��ԓso]I���r����]�pg��v��h[i�����>���&]��~��V�o	0�Eid#�H���y���_��J���8iW����'nQ�@�#g���L-;s�x6�{X����S:�uH�����,�FJ�v*ӣx|N��wi�?�+[D㢎f|�Sp,?��2��nn��x�V�&n�FD6�Mח.��ޮ>2����MB��s�k������O͌�:)�z?o�o`�r���<]��q����$��9Ȁ�"�䩤~7�O�Du~'CpCL ��O��+-|zZ�̨,��:��hW��>4���Nߛ�b���=V�5��d<��p&��%�n%˓�+I�c�'��� ɥ����!s�OP�?��z�� ���a7R�[=����w���>O�XV�N�?���S{�+�,����u���
Hw��>m>������lm�uY�r]�Rm̄,�]�z����Ծ���⺞I�g_�CO���g
��:q�\h��)dr�v%%Yߥ�&<Z�#�!Q�xj��(`U���&������u�8'�@!�~O�ʅ�ݪ�V�:��[1�1P�J5d��,��PT!��y��W�}E��5z�닐��]�-,��'n3��}���|����2�Cs��_p�Z7��--��Rc�sU�D<u-�J�r�H'i�<�9<H���&��SL��c�����kMGi�S��8#���	`lz ��N]�J�/�;�%����AS�4�
,���y�&��[���J��/>2�y0�B��3��=�����y]
���P�-}*�l�Ϥpl��"4k��ɲ��V��ߥ�\^.$��ͻ��ρêPA��f���n/��:K�7l���&��G�,� ����f<}��=^��}uc���r�
u��I�A�凲H2w.�������O �Bq�}��j��>%�޼7�gU,������Kr2{�Yji��|�V��,qt��S5�<KA���k�dz���c�&zo����������Ó������>�tU�ڳ�����`J�}��E����By�Oo~�!���R��?TP�saJ��aIDW)�����ߡۧ쉪âO���ó��ݫ:)T��SL<���&$T��%%���E&@7짪p�tl���/W΍`���,i�o��QwV���1㹆���i�ؿ=���3�*�zv��VE+<��J��؛�'���>��
n�ΒpK��k�i#�jK]�ߤO�'	��B�6�)�%}
�a�;�%Oq��V�Ӈ|6��&�q���F��b���|/��2��O~��H��۟����@#F�S��Mg�Te9x/Ҝ��@�E�&u��V�
[�W����z�%��s%��!@���"�\ʊ�e�6pM�s���Qf+��!o���$p�l����M2���� ��`�c7�����
FC�>��x t�{���֚�z��\B�¼yg奦�![Ł7�Ϯ�Bteb�%���_�28��T��z��-B�qR�4{�]ZНK;���.g�ց���^;���C�%��9ey�K-�z��ve�Ƈ�2��|��Y^�s�}�F@�߼��ǟ-�AtG�`��=>�d���,Ó8�ŉ���>�+�/��ot�0Y n�Q4Dn}`���`%+�vE��.��g�,��7�M�^e�	h�C�}�,�^d��3���2`^�'t���p��Ku>�uK�� ��LECn=���YT��t�b���ge�����nRFpw-U�J���~;��:�ѹ{�itͩHLo�n������f��(���<��BË�|�{i�1u�w��'�'��Fo���N9�!y#�r�)�sY�Q�9��%c�+�G�Y�k<�Ԭ�ք
Hw�y�YX&�g����`��-c�����@.�8�y���;�y��p)_^)��Kx�f��lڥ��,��E���Btdr}�x�ȸ�>@�y �� �ȡ�p�b�YFQfg�G�x�B��͟?� ���ˠ���t��ǗiV��A��wi|���yc��բ��m�L��!�� �������$K߯�o�����_���̷����}�M��ǔ��ͭ&�?|�>�łڿ���:��?���כo��7�l��{����m��5��괾	�oy���vR}�V����I���Ł�(#q�QIA-�y�8��\T8�#�k@�_�C��eq�3s]��R�Lz6�qfH1`"3���X�沸�L��y��͕����V�-,9XX%��C��N���j�'���﷝_݉��+/(H~tQ�k����"z�YJ�x'G+dW�����O�[�4!(��@Jg�5�2�{V^�ϛ�a�H���A�����}U��̿�"I�{TI��w�۠;L_?�-]S���2DKv�4�_?/���ya�k������}2�W�*�g���E��Me���t���}�����A6����̸<-ʶ{���`�E��RH�X�ʍ}�KO��D����Y����w���cy�z�'N�tⲎ���R4Ι����=G[C�& �H�(x����-X�p�M㗭�۷�;�X��0������*}��[������J�o���%���$���M�|{�^VOiG���`�}�/?�����af�=�9�ʽ��Њ�<� )���ý���i���=߿���2��[B����4=��{���0=������.N�x��Q�9c��[�I:��@�D
* ��~8߿�n���v=��*=����5����<�z��C������Ĺ�G��m����~����ZM:'\αX�q����鉜��GG�����E�BR}Nk�h�T��$��0��E�%���9Ť�+V6��([�㰙��y��9� ��c�p`��D�ss_�Q���a���� g��\z�LrF���'k"��'?���/��ֻw�`���U����y��Yj����� �����grӐJ��Tus���-��!�8��ӳ�d����rj�s�7Z��P��lO�(��@7�Z)>�C�^s��>Gm����?�Ò�eAeoץ_�sUv���F&��l�u`����ҿ���g�<���3onoӷ���.��: �`�a=p(Q�M�|��6�]�}�F�xD>���3L1�� �!��@��`'z��}��÷��ͻQ�'�bѾ��"\.EOY�~l{� ����-R�W/;�֡)�k�'����mg��O���6u���e���$�̅o޽OWon-�&-�ޤڮ�
�ƞ�uq
2oJ>0�žm~i^�#��G�6��ߪCitu�lErMuɆ���S�p�ڕ��I׏�^u==�iii���Q�`�2 �m�1m��b*���gQl A3����@��b��m�Ep;F��G랁�bE΢�Q�b�(���T4����2����!j3U� r��e9��s�Ld���mϰd����$�	7�=�ɼX��8sh�K=�����4��D2�U6�	�A�����T��L]�l�Y��N.[^>�5>응�e�/	~��N6��\�읚_��v�g.]��v��׵��a�]8��h[�u_]�P*�@p��/��FF���^��ÿ�W�:�����H?Z)�����M�����(�d����4������i� ��ڴ��Y`�?<��2֏]��C�i�t01�`�ﯡYHZB)��<�ɓ��v��<�sn��8�kD����b��59#�)?���sc���L.n��g�c06��A��e�ǡ���u�H�����9t?|�]�}�6��C��JX
h����ҨKY�w�Ԥ*�-X��W4e.��8l�"Y��P}T-�*�v��1���7~�]`C����
�i[�K8��Y���p���讗���_>i�;7���oE�B9k�ehĠ��"��k���//k��t��'��<e�A ��ڜ�S>o�
q��m.{3u+o��G�t
K�ܟ�٬JT��Ǝ�r���� ����9�<���s��uz�N4d'b89������d��=g��2�y����~��=� ���'ף��+�����r��������+^]�|Hd|`��br�#��{8� M�Nl1D�ޘ�wdQzA�6&�PWV:��β�"]�!B����?h�:��}������������SK>s�NTo"U~m�5Ss��0��Ʊ��*?U?���*ع��
��^��;�}�z�YS�FG,@{?` �-��N��o�5~�$ãZ�:Y){�,>(;�R��g_���!�F=�\�OC8��cO./��w����������	R��ԋ���hI	U1!z��G���Y�v�����kfn��*��}xIi��Φm��� 3�	�i��J$��Н$�I����Y�޼Q�\%������������m<���;+5�@{�]I��z�|�4.JIm�t*�^I�ŀ��F#|�UeU�O�";H	���ƕ4F��Й�X��}��4��?�⹴�c|F�S~�ſ�;��t�f ĝLX���9�g����Z��x�MЦ����>y�%0��\:+���p#2g=_���M�L�<���ʌ��a�r���}�s�Ã��O�&�3����n��`�3���l=�\J�����Z?��w��O�mzy~I����/u��^��U���"�'��)4���t=�I������Yغ�B�ٲ�FRݍ�����[0e8��1��Z� ���ϫgeoE� n�EТ@��mde~���0p|�]�뗂4�\��<����2L�a!'�h�ں�JW�}��Dd��B�>�lJ�T.�EX�Kd*�$��A2�\�
{�o\��\Y����.�L����qQ5>��X�����x�c۴V�*��JO2���d0 ��߻v��(����T9i�Ҿ.&����ϣ?�/S���n����X�W��t��o(Ղ���������]�OJ�!���$4��dQ��KÉ���O>������VϮ-��z��2F��Ep���M|>L��`�s<-�У�]eQH~^V��?��g�8�~���L��$��̌`�z (���7��g���A6�����b1{�� ��� u�x����R�oS��f�G��f��LCa$k��2����M���u��Vpñ�6:��f��v�N��"�y��h��<�0�&kl�1p"H�����O�������l|0�?���gA7���~0u����s 2�qn��I���HY �5�"sc�A0�y�V/��������!RNm�q��M�T���/�{m
h���ץ'�+W�
h�uڳ��K/�B�>g�j�F3\?X���@���!�%�F�71J����̋�����C�е�ߵ�H��㜑S�۳3I~���8���}�P�e���9O]ʨT^pab����A��9f�^F]r3\N5��(6 l6b�"r�c�,�sqЮ*\OJR�evti!�\�ϡӫw�U�ؚ��~�ͪMs��E�6��N����1cꆅB:eS^�ƍl`�aŹ��95����!��{ή>�{�}��{����`���)����a�ܝ5��!�����}���2=�������3M�G΢�1ȟ㗰�,F�?k.����^�������X�α�\4t�' ���Rw��m����1��?�>����a=	?t�Ni�ݯ�2P2��j��4�C�f�~	\�f�1ד:=�a`F���v�u'����jYT2`��Mҭ]��ȧ�H�H��x%}J/	�Z@���+�l�"�h?�U$�s'��fw��9��zw>�rKI	$TαF1���ڭ;��?4�z�a��P:�C��?�A�gvq)OY�F%Z��Ӈ����t��v��R�R]��I����v#�z����(��x��=�N����t��� _�S�Dzg�0�E�D�9a��)hvƂ�� 7{ܫ9���L
��m����B�7m�0}����'��
N=ɽ0ό�r/�Ap^�����נc߼�)5݉������EFf���͞-�r�JfA� ��r��Ƃ%����X�j�����!��DÒޯO���A;���y�p � _^V��t�H�]A�:wi`q��8��(��4�_^��U1[�M*�Ԑ��x�Q���tT�~X�'���d˼?��9M�/wV�>�z��i��;o4���W#�Y+l�3����f�L/�Ijոa8ЕqN_�������\[��9TY����q�n�����.�o��5i�W����Qv7���� �$@����dù��V�۝L}�i������&�<�R���d�}`�N@�s����Jnr�\�=�-/��w�����?Π/<ڮ���}�奪b(�P�uz? �3�!�������n��Q��6�|⅒C�;:j�*o�B�%3���đ��`YD1�� ��-�� ��տƞy	뙁��!����i]�A�����04���&�T����WO?�`R(SiNnV�����Ϟ�;
��C&Gvu�V�
���)/g��<ਪSV��$iH�@P)
���"�rz���\��QR��������?c�>�r����B �D��C�se���~nk�2����{t]h��|��ޣJ�f�jf����G��*���Y)����Et�欜c3m-4�$-�*�MP��G^�=��̚V�#�(im�^_,u�Q�������:���}���kJ[�dw�7�����ORߠ�Ep����Y�{��.r�aLֶ����%��p�5�8U��zy��L��]|�غ�T�����(�_�~7�8x�V]��d^�]��0��J���h ���3d��Y�ӮV��eh[�H�G����qK-E�֊~�B� K��3�e^b�GbW��.`m?3a!N���_�7:�HBh�c}����縗>���B�9N��/�拃6 c����u~��YO������v�%ET������ǖN�J�q54�	�R��NVz�P���P_X��˔,���&~H����R{_U�R���#AU��R���qVn��D)�N���/I�s�-6L���F6�s>����š��2�-��d�ݓ�C���N��\��,���g� sP�V4�ޞ�~R�
��cQ�z�ǖ�YǬ�	 #^~>@��?��[/qe��ej�[t�{'�
�UiU�*,�5��c��B����$��Ҳ��8|0�������>=�׳�zgV�.�Wj=ЄFwzdk����p&	yW�����M��m�y���&�l�����\d�����e�M�L�j�]��6DH�� �c�٪������0qe �kLgS�� �����az��72r����9�&��G�W!�G��^=Ma^��Fc>�xS��n�-�]\0��u�"��߻S�냰�3?"h"��(a�^��z���,�f����c��Jt�3^���1�,<%?�W$�6RR��TU�F}��<R���ofӶCz}�-���sy����cX;~O�ȡ��5[.;��w��`�L'�X�K�\^<��r��&ͯ�w��M%��``��5�)e�\
SBe��kf� k��� ��_��N�9��5�p���O��!5��d��L�������{�ꮣ�"�RYP*�)�t��!xqM	B≾,�C�{K�c���rk-9�-(��p��P5;���j��C��e�pv�t�µ}^��$3c��ĞI8<�[��(
�E���2 �b�#b��4���Y\_j���޸�>�o���8�@\>'���v��r�]!��hh���Z��%9	ZJ<�qni�^%"��rW7���w�*�y\�����E5�V�m�w�)�\Գ,܏#`���]����!y4���xo��;d��j)Pʩ(�N�W0��@�!��y`�X8�
�UvG�&&/;�pZ���LYB���/7�ʝ���r�!�G3[�QR8��N?��a�h�pUo��c�|0��l~?��Z�������T�S�y�0o`NnM����;?�|��r�VԖ�x�R3{s#��<���&|ؙ6�2��4Q��:ASa��r��$�j_�dD�iI8e�I�/�W�0�1�sI���r��K���ڏ��@ہR4�3�" ��K��)����{��pG��1����X�i�+!@֤�ת�z�g���G����J�>~�ݠ&��A�3q_HIfl3t�N��]����z�/fi��HW�E����s�^�U��);P"c��7�*U?a��+=�ևjEd�#Ih]+�GM��Q;��q��9�I��ڃ'(�XL^�!���{BF~
d��֮�\�o���>|󍾏�*�
��ɪ�:��>��}�<��{���w�;ږ_1�M,E�hj�H!?7� .�����*M
���p)�l|Xw�� �2&bdn���C���0���)�޻���IWKm��NNF�0S��x�%b�6Qu*Ks�4:n�E�'݅V���<r�t����,�2����4�:��>��ՃRI3l��q}��(pF����\�� ��>Qݜm1� �y����+�/�d:�h��z����^/hN�E�����5s�+U��*���/iN.�SC��f��9��G��!.�F�C�H���E[�C���XƁ����\���ļen��6tA�J��3�+e:��V�����@�Re�=���BK�+$կ WO�Q�3<��P����	���t��u�M;�E��8`	����M�T@/�3���ނr�p��+�WXGڡ�����
Ҫ�+�8�"�^,ԣ���]۽����^%��׶�T�����2.Z������0vF� ��l��I�f�>hr���SZ�!��N �B� �����f�%>���v��ґ���|��V͎@u�"Ø,���']�
C'CV�� XW��~h݃`���9�=j�A'�(���pB�:���$РUy�<��P��C���̓Y/�^&�;g���Do_%@�����ǁ�7T���j�P�t1w	8 �q����_�E1�E��K����b^0�F���l�m�4�gZ
�\rŗ+�T
��Ǧۉ��Je���v۽�ʳ@�8ZMe���r5����n�ݗWɵ�^k�ʔ�-qV�'��v�q"��y�(�"D�tp��B�[�q�F����g��>U_�&�12�l�d'���J�ɴ��JW~�P�r����Nr�XvQ��=�����F���q�:�c�g,x��zm[(H�.�^,��h�-S��C��U��l���>޾�6͖3��ia�b4����R*��ܼG�[��i�%v��ϳ�u/�.T6e�e0&�0jP<&	����Ź��Z��^@OcbkjAp����x�dl�_J��(�Wr����{[��V*
����攓(� ��W�����@�=_ٺ�3������WT�SÊ�4�l��F���J>��>=�ߥ�>'"�`�X\]㡓c�v�v�ۣJ[x�����9k�2�ɨ���W��l��~�w6�D
�þ�L+�̩��E��z0t���E�l5�h]ŕ��S����R�5r�+n.�(��bS2!̈yS����l�];^^��(3��:���׸$_�2�Nђi0��ǖaè:���y�	`H���{9@d3f�G�F}yRiȽ�\�e7)��G��,R5�d���2lf�2&�L���7/*���e�s�,���ZI�d̼��(&�F�����sw�;+k��k�jǤ�r�}Ջ́=��#�����3�Gˢ���$�۩�����a+�{!�����
����x�˰��1��a����j��֮=$VK̤Ǭ�N��²���\L|=F/�q/f��f���!m��$1����:� Tʄx_콍c����, ��7x�SX��eR�J��cZi��Bm;s:.D%C{�!	��c(��,Czg���+�v/ie�cMVb�|�n��E���×����w��J
:���7�e�K_>~J�_�|]ۺ�Y�����+�5���(��n-�R6�>����G_\;����Z���
7lYx6�nZN`O^��X�ەx�,�L���
C���nU���q[rl�A�	�{>���_h�X)������F#�V*�J"ج�v�4�s�5&G�h����~x��}�r�"�2���T �B����0kY����!#�0�� L��48 J��F�lG��)�i��g�	��@c��l7�*��� c�td%8s�!h[Y/OH������p���VJ S�_8�yz�Keqh;��Eu6��|Q'o��e�t�\|�Q����<���=qZCхaҽp.AoC��>�l\.Ǯ�q �w�.t�7�K�jn[�>+/1'X��-�6�1DW�����eS�d�H>|�b�:�|����eV��hm��#|�r>�S��-����T%dpvOX�{.(]W��:�>I}y�OO��hAy#5����C�VNC��e%�^�Rb��\�}���<][���Pݻ�8�����Ez���e��7[��a��*�e������BU��ͻ��?�'�8�Xn����C��ǟӝݧ�w_4��=�l��/��~����!��؇2�ܡ2�|]���n������qK����u����QLG�`(h�����O*�E'g @1���P��\܉�������w\} _��0J|e���ǧ����j�#I�5�Y�H EzzfeE�qE���!��d���p��5��~�nY�9�2#<��Ԕn�����i�%&t���<�T�r�6���&����?N��&��J��>�ӆ����"5���P��\0FiӦ�?�Q�R����gt�T�
qN��x9D%�M`?<x��q��L¦�ߨ��|5f������L��9Mc���G���?H��3RG��A=JY�K�2�O*O��1"Z�{�v!��B�y����s�e%�i(:vS�XgwגW�-�cJd������+7F�<hGj�d���L�_<QWse6 ��TS��f��'�˹��"�lMQIl�0L��݂ȵӫ�e�Ȣx�5�?�-�(Iw*A�&�����qj߻��Ke}hXゟ��~њ����{�LP{!3�|}���*p��ệ�\8E���>Soo���Y�4�2����w���Q���f�+C��V�%"@�~�;�<XYS�Z�p`90k�Ѫ�h��z�El�ap;5��7�Ӭ��}p H�E��=)������� �-|t, ��>�؛­�"6��B�a���Y������Α�Q)e%���m�>l�/7��I�Z�����c,�)#t'z�ޏ��X�Q{L��m���G2��@(&��`�J������iX��(ި�X���b���`�Ա�vu�$ݞ����$M��\�R��{� ��S�N��K��r6�9ȃ)��ij�������>|�둹�$&Z��;�k�D4cp��v0{A[b�<���w��a�b�?U��{��K|j���"d�<;��G��Tu.w&~�)�&��dU+ی�cٳ�#��yR
�Z#S�}���Jӳ~6��2��kˀ�oT�e�{a�hݲ���e�8��,��P�����T��ޝ�8��0-��_�����k��=�?��?�\�f� �u��Ђ����A��k%p���d�>Ђ ��`����va�}?��5�g�_������
M��n}���-�9[`�>��><�3�-c;j���ɂ��(l���S}	|�Y�QL�=�Dc�3��Я��/�����_��|��v�����H@�r�8�` ��M�X�~� �����N�~P�,Fu]u�Y}��CP��2��;`��jt��$Z��}��n�ևP��)D��[�v���8@��;N�xc����n��#1Rƕ&��k\�*k+�*��?�1!�/�~lz��n͈����{�}���A��;J��?#�I�_!�������|I2�sa�&e	l���B�z��W��G�4��d�ҽI������,3�Ч>�ϛv*u9$4���}f����}��:(3�0�4�3�Edp�0�8QN�C.���f�bmY���mZ�6��t��+FG�;8D��e�XY��ϧ�*zf��(g�FX5$��;LL%��=�^� X��O8�X ;�Tۂ ��*t;�:���Y�l��������ZmRkA9S��~~u%x	,�|�.ˎ��� i�<-,��J������͵�I���F���l�(-�T���F^�TU�I&6̫��ìP6���r�� ��z��%	�a!�uoe�*�,W���C^�~��u��+_�rp��L�/�㬇_*|Z!7�VÅp�T���;&B�D,��?m?�=L?:Q�?�Pj���JYʃ�W��)��B�r��`��zQ���f݅����l�u�� ��+�v*|rX�P%_yԲ?�ͤlc�df����=Sy��+|9k1��)IA�x<�6{W��K���_$����d}�Lmx���<T������ @�SM�4��V�T�I-�}��){���N!)}4�P�*@��A�`��"�Ɣ(p����lxv)�$���8}�Ё4���P%2�,p�m�0c�ԟ�Ϛ��ԁ+��E{'ї�w��K��v�){�������^� �$d�	,���9}�d�Ű� V��$����dzLU'�$Y�W凫��e��-���0y��a��B"0��^݄+�}�Z
��WS�ثO�^��=�ϟ­e����<����,�� ��iRd(��r�����Y����0�q�.�z'
;xv���,��^�_W�i<������5,��ۅ�+���}���vhN���__,�ެ����6���[����\��ެЦ+=@��{�Rb!H*�n��N�<@���R�G�r�',�8}��a�Q���!nzA<"�4$�ge��=g������2��n�
�����	�_SAd���������6e�˥����krRM��"���4�����!�N*��cF"L$��W���T����e �l8��̍㵤�Z�Ƣ����� (Nٛ4��� �t��U1�r����\ק��ņn�SݶI�[��Hh�Ah׾��j^���9D��|h凃�/��dl��ښ�Xִ�u8���Զ ���p����d�3%ך��W�T��<����5�R�\m'E	@>}z����ު	��שs�)�V�M�@�U!���>���,p�({��7��ւςv��I��{�
P�)NV���ꇁ��=�X:�YT�����^k�ծ}7����ýl9���0��J���xN�a�vY!��J {��J�(��(c���p��h{��~���b���1��˖��UN&���-e��;]���rM�D�m�d�jS���F%6lCx;dۦ!���K�{U��/� '�8�z��)$�'�)&*�F!�>�����N��	�N�v���	�tM �A*mA�i��?+cF�Wɒ��l�'��&�O�XB�bতSi:����r����EH���;�4|i�'�d�x� ��xj�����9��P�'�����f=�I�Sf�I���au��P&��� /�A�A���T�s���"�i�vv^��G�� ���Β*IS�{�G)x�QQVC��Z �L��ͥ�b��U��/ �:wR�9MV}>�}�4�5e��@� ���|=l-�e2o�Hن�YY�XJв�X��0_�i��?�^��v^���e�=I�l���aysnn�5�[���\����r��e�V�pw˩ ꫻+���Nx3�y.6�5�+Z$p�V3e�G��L�7�e'����,�927����Mk���fn�re�i���
p(v����ˢAL/��������\��jtŇ�{��M��E�2�
5{�+���H1յ{>��ǖ�rn�߿r@�n>E��\�W�.����7:��Y1c�L#r���2�1�9����Wj�[ �C���p.��5h(�w꼧�Ʋ��yl�;r��|�iڒ�	$l���I����*S�����m6��5��M|�n^1%N�NAM�vP�Є�{�{OR������qok^#��8�K���6bG�i�qq$�e�zʂ�����j��|�t�["��ݔ�&XI��5�G�����9ǓӁ����.NN�#�]H1e��49&t�X���׮%�:zA1�5c�î�;j��ρ<!���a�z����)x�,i��
��*�tZZ�xG��+o�}Y��ܮT�Χ�z�0
�d>i�i$���6b���觩�;��R���t�Cm�P��\5�K��,�)��\��B��͚2�Vp�	6�y�և8�7�a���u���xK�>s٨����XRh���ǘ�5�J
݋&���}�W̜$��7�������J�Ub�Ѯ�up_����n3�/���7��&s�$[5Ժ�q��"a���8ѽ��R�Z�T��ezN(80�$��i� �3O���}� [M3]͂��Cz"�m�Ž��71nN�$�OLX+"�g>`�laN$�h)�-��n+5]�W�Fƾ!AY�Y�&wt������b��5�y� ����P�����EKn���
*����,pk�}�.��.F)����:Ġ�^	x��CI��ې�M��h�<P2��E�Hte�Nq�F�X,S��O��>C�|��Jx�&I�߯>�Ѳw��m:�N�g�jf��港UZ?nh��� C��0��i".���e��/�	�ʨ�Eğ�!�����u���eQ�5dm���oa�������9���A�{����&M9&��Pz\D���ǅ������2�l����_8�q*�C�����	ٕ��dVJ.�w��%<�l�Y�z}ş��<鵧�"�R��n���Na�̠a}ڊm���x��6jd���1���JX0�a���,VL-J�e�voN�}�a�=��/��v_�%+� ���!P���!#�P���^ۿܬ�КO^�l�"�cֻ�a[؃����J�Z2+�lՂJ��ݰ8I���b�������D�����l��!�f�j'���)�&�לک&'��m;��i�2x 8,8&[�n�J#��VV�SJ�>�G�.N��F��@G���KE�N��]�r4e)�{��y���2"���(��w^�?�}�_?�7/��d�D��e=L;ǎ]�<��$���2/���Ã�gu�9��w��B���ݧ�3}�4�}���M4@H�ht��iZ�͍V��S��f�d�Y�R�d��R6��T.�1��U+(˒�&s�W��u��4��l�2+\yWX�\H�'jǗ��W3�t��LV�Z�6���[L�<�Z������_��K\N]s�F;{M~���4��e�G����S>٥���Ɛ�_�j-7VN�*��^��v�Z}�i�{$PN:���?��|>��s8l�E3��:,��tD� t��D�`#�(������7싼�E��Y6�����p#��t�'J��I����+�V4����� p]V��?>+�C��D늻�*i��v
��g�[�}��;ys9Ջ����N�+}��8au<����dh� o�u���%��I����,fpq��s0J�*A�#�����9�p/���bMHc$;�.�M��L��x�����Q�2�IXxo�"�2�ޕ�_
r1X��Oٓ8|���bF,��rȎ����Etʚ�;M]@n�"7DO���g����D�-��R M[��!B
F)�6��P��^�2��1�h����v��R5w�z#�1����:Ѹ�r@5������l��"���2}V�Ip��M1��7�{��ܒ����ʮ��K7z@���Ca��\�\�UE�k�_&�R����Z�fv?��S��޵�����>�XP��)P �\
*|0"��>�����W�>�����	�B4�%``A�����Yk�~���&���~�t�쿁L��Z��6����V�	2<MFKetMa�ik��=J&o/�:WK;Xڕ�bȰ&�B�7�WL����o.ȕl|vi���k�qb4� ��aK++w�o��;%s0G_���	��������߇���_�|�U��j�^�B�yX %˳O;g�pE[����{�=�[[�_-���/�%|�W+K__�^,��l 1���ˮ���Xt�r���P
������6<[��B9�w�ċ�EF(8�GB�[��8�+�6܅'��^���-v�d�b&�4�8��w���WM��$�5k�v�zx�tNM�15��tM�F��:2d[qg��%}�>^G�^����Ɯ�1�M������K��{��v�(��]��ߗF�#ń�?��h]����ġ�?_�L�,�c�"JPy� ��B��̣�[�:V��� N���ҿ����v��}��p���]�֨�BP+gh�Ep6ki%�v�g�7
�2G�1� �=L�'��\�\�2��V����j�	�e����d�7P�,˻����x� U��ug{�(~�n��avs��]kc	��zp�g��4U�3�\����+p���5��ƫ��U�Y�鿉��9SB�Q��#�$�pc�RW��ӷS��^�6�� I.Q�4*��t��U�>1��,���-{�X�	L�`,�!�k�j��g5�2�=��S��F��wϛ���5T�;��^�L�dtzK��v��aM�7J��&wy�rE�}.��K��{7Oa�iSEs��-��?r3�����A���C�'`7��5�T��R��
����������Qf�\I��|��dz��b�CIV(\��	���i�0�.~��|%���d��M=�DɢTM%6@P��d�Oa�ĈHS�Tަ���-2/X/I;.1Y�5\T1�t0��.��S�����H�E�g!����#�:��K�`�)gʱ׃�������U$;0K���0��'����=7L������6ac���u�oX ���w����"Њ���{�o[�v������-W��M���4\UI�%-����R�(��e�����}a�W���vX�zG@aj?_�矐 ����wYyi�f���2���+��:V�<h����5ؒlYy�d͝z R=��K��.^Д�D��nڭ�>г��p�V�o��u�$����Ӳ�ӧ���uqm8����}���p3[*�ܜ�a���ʻv�ْ
[+Ѐ�0�̍�]��YP��_���T�?g_�as؇_�=���{�vڄ����f��e+�a����E#W�xXi�蘩�7Q�=y��D��wهT���Xu6a�T����{�^���^����-٠}	t<�#�F�Oh0�.�ǅTQ��Y��G	NƚTC>/A�.)�$6A¦��u�Aύ���hА �cVF1���r.
����ڧl1���a����zp'�JN���I}֓8���-�]LC� ���?x\zI@X��c�7��FT��U�Ŋ�^�� L
��Ðk�yGjAPSg��lV���ts[w\��}|ܲ�PC�]������`�j\�ső��J�+[��:���y�2�V߷��1�b&�J�9�����ҡ����u���
C��E�8'Y��·l��a@ �P���;�6SZ�m�~�ɑL�x��r��.�B�}���j�9!_����{J\+���D6���!�,���F=m���9�k�a��~ƹpZ�F�(�-R�"d'ٗ�~�ߗ��,�R����N�b���~z�j�LQ��!��W���^n�E���R,��Y�U�Kf"?F�ix�2>f��'�p�Z��Mj�o�R�h;[8>��WY�v%�a�ng�H2�&E��)R5u|��8�1YS�Y!��s�����v�,R��
������ٚ����v}ԺBZ���Ó|v�.���N�/�,�w;[Beƛu� X<#9�E����C�F�@�*�Qb���}����i���s����5-O���2	�ީD�f1����3w.�`n���pjS
��{+�^�M���6*�n� �-2���- �p���^����m�{�-��7�hDeB�d���c8���"o���0�R�,H�Cj�S����^�RU�"~����>W�����K���װ9���k����7�˿Z��e��۰�	�'�fd�e�}l�nf�>���l�س�6���&���>�Ҫ#��wV�gK�s1���ʶ���dfdb�v�n,-���a��2�e>�_��f�Rxb�?�@8� ��i�I�O�q�;�V���+qS����"6�L��2������E�?Z�v+ua &��5d�wN'��@O��!Y!P��Ϛ>+6�2�����Y����4�}�Tv)�8���:��43�p�n���52���e�|����l�l/�!�ώ4'PM� 3��A1e�x&{PȰ<я��]���������VDx����ټ���0hpn�oJ���lz��ϟ?+�	��9�����Ի�����ڔՌ}F�ߦ����+ʭ"J6�r`��1��ƴ+�Lcjeo.�t�d��'%&}�ΠYK�ấ�{:ǌ˱p*�,����&���S���q��Ol����+{�&p��](���x��϶qNVvrMy�����$FSe$��Uՠ3����$����K'���߭w������}ƫ���|��e6T$��8갰ףW�y8��bY�u���=�q��d�!�ˍJT��gm@�����T�A圬�U�����}�H���a#��Vx;w~+��A���0���ءA��$
IL� )�>�*TM��P�����qys#&
*>��O
i� ��2�������ߙi��������e� <�)e�X	�"*xQ�K��ު ׅۄy�;%C��ڐ�I��%��D�>�/�F�Y{9[�ޯ�����<�⽻��Rބ�|�������aj���x~�m4��?sR��3;-�m�C��Us�M�<y��`�L�+�v��l����� �t��ZyF	��-p���N����-��v��z[��ɮ�t�ؔՉ�P�wB
n��P8�z:!�������hCY��H�&�p*g��_�h�4X�䩠l+��C��K�C���0�Lד�L�gMdh���T�7~N&���^��a���.��=����S�p���oK�nr���,4�2��U�>@*�9�ɓ���mX#�h�Y���el7�B��q�%O�?�u���0���LӉeʀU7˔7V�j�m��Ls(�B�:�EL�$�Z�#?W�a�3��u�U�2¦��٪�Z{��1���N?[�_�ﮎ�[�#��c�K�Tp����ͦ��܈�	j""�d���|(���1[�$x��B�X�����R��cya8�l�ĵ�.ןe�d�gy�?��:(��,ͼ��cտN�b$���}:N]M���PQ��}8��~il�=��xN�5�����J���'�<H)�N�����Qe'�f�U[HH�,M���)gO��x:�����r���<�E`��v���I�V��s�en@!��~��'��G]�8a�N.~	Q}#m��X�^9~��Xc}��>������x��(G��R��^7����2~/W�͇29��LS�~��Z
�)0�I�6Mi���.=;)��m�)��|D�KC�!@ƒZ��ާ�L����[�3��a*��5����6$e�b��C�v͠)�Y���U%�1d����J���:���������2���Lu�)�Ic�m}�^������ޝ��J�,{!��rO	\�Or�����/ANe�Nj�=�>�5w'���e�䝸lSYF-ĠRzg����^�^��ִ'���{��~'?O���i�O������詜c+�j�ue �}�b�������x3p�O�CVA��w�����������g��8��>�=Q���Q�+(����K)j��A¢\^֊3�t0�NY�w��[��Yq���>6�{tх#�;_�S��82�g̲I��/�t��y���U�n?��|���ѝJ����F��Χ�>|)���Iyު\��Kٟ��&�;�Ξ7��� G�Y	��UX�v}B)� �>~�Ӣ�EջJ�����@��c�.\)0xp��R��#/ճ�0��9�ӿ'��X�'�n�_���H�OA.)	��%�Jt��I��+��Vxa+$5�$��N�{���++�S�9�ռ_�fc8hƟ_��!A�n�<��Q���$���%��.ݻ�U����6(W�>Ŭ�>ؒx��mg�am����E�"��n>�+k+��D���@ H6k]��¼d4��6sljY���V�~}z�/knvo-�'�<0kF�T��b�����Ƃ�֓����{��ڕ/�Nʿ?~��k{�:�³p���죈����3Z/��!Tdm��VH��
��Q�ł�q�Z���B�sp_&�$����b���E�z��ăe� �9� L`#����p�!M���K�{�$��I"�G��5�D㦾�KU���$Pn��h�:#�Q�i�#O$�B�� ESs
����0�����M>����V�åC���\0ONF���]O,��M�?����|��]}6�x]fY�P�ZDw�AHK'�`(������߻��}�@��&�����S�������fr�[ҥ�iTŠz1�M�N�:�뻥��y�JR7���-ϧ 6e������2�sރ	s*Y	��,�;�M4�!���]z_�Q;���� ���ןJ�t-E\���i/��uhq00ȉ�� !	���&-�	���l��>�vSJn��U�*�{�M�]]KJ��em'[�G+��p���8E�7j%(����4�OHl�|z�����Q펒�MJ�v=v��b�O�i��7���&���g�/=;��6�}�u^�~�<���=+Q��
*�t�+ǣ1��YVH�֪�R���ޘE<�P�f>��$�'-�+�l�DJQ+e�����<+�Z�h�e��=Τ�g�V�*01x�Y��#�C�I���ic��챣�AI��wé��C��vP}�s"6��SJQ�y��y�
�0i�۰���|e�עu�&�O!��5�Dgp�O���l��ra�f����׍�Юfǰ����JM䲦-�j�oy���C)N��gR����]�=W'�t�7��� ���*�p��Y>���Ωm"��ٺ�����pOD����F:'���z�p��lM$o�jQ^N�.D����3,ʩL�}��� �d`r�cS?����s��PQ�')%;~��
�}>?z�-��K�+epcAM�<��ķ�R�:��:���
�������-�p7��>�S ��8�)R���ʂSi��:|���O{�H}�@��&�X��no��~��óZ�JS�L�-='�3��`}�,ck��e�__���.�m�x�i�^1����7-����Sk�į�Yٟ��ѽ��`HTO�a�r�&��Ӗ���,m�B�V��ճ� |�
E8X0$x,��m�:�R�OP<��������Q��H� ��
qX�l��*�γ�7�\ٝ��3�p�1�s�;6���b&ī� )��D et�RRc�c�{Ez�S��<~T�S��vt�s���lH�5R�Q�P�H�P9�֭��w���oD0�QI ����zk�����敝��� d��_^��/�����-|�oCe%��n&y����k�>`�I��DƁ�/�ē�ߥiaR�er�p��ZDHol�c	P��]����h���&z�����zl)�KƷ��J��B�;e|�Kٞ�u�D�U�%\Y�0J���9�t�2�Ϩ�͋A9E��ډ��vj@0��V���$�{�)�H�ү�<>�B�2���n��b�/�do2Pf�ù�@fzI�~�1\g��%d��8�x���%�uw�-c��ބ\�?�j	�lN^OYG#(Y�TÅ���ųel�����3~}�yCo�4����6��B!_}��	뗝��v�5�<xJ�L7�B�O�m��L�7[�t'd��8 �ΰ8P�Ҷ�ן�FC	�(f�W�� ��"�:#�y/�#qU��=�4����K�2�^��bZ���0���2L���=q� ��̠&��t�w�>?~K��|:��S_K�� i���	�)-��W��}��܇�j>�����LZ�����ׯ��5�#!���Y��$��Y���߶��y
���Sϔֶ1��� ^Z�P֮9/����
؀�f`��)��y��d
�ӟ���$;�J��A8�X���cƐ������W6�]�	*P�&�!P�BxףK&ݳTB���F����I�2����-��	��&�i���}����	�w����5��We�C$�W�KpK/�� �d+qT��D����hf�`��m�\HpQh���&&S���땤�����`��B�eFP��w�a��See�x�����1k�fɲ˨��;ze�%������ڦ�h��X����q�T9]Y����fZ*�{��:�dY���[x||�5���&����y�L����J���=`=���R�-$+w����XF <���_��Y3�c TIA��bs�b�������I�pU�P��3t��q�5;��o���R�z2�F���ت�O9?�7+���� @���ĵ2w���p�����I���^��+@�[7zn��٢�x*^�u��_4rQܬ,�#��[�@����}���*�,_�|������?�i�V�BJ�@�����}*J��@2�]cA�zi�r+OY���2Y9Da<&�խz�|�/��[=(N/~��F�	�~^F�?����_��/1��(��x$x��1�i,�=.��W�x���1�s���h>�����_{x���3e||��̇
�?d~)�%~k
�!�822W2	ț^����4�wחsz��樓V�`r��d䓘��R�O��l S�os}
���0d�������p���&T��;a�Og�ѧ�6�F��]�aK+�,�uʴ��xV>h���W���2.^[�x��Y[p��ms6�%+�Ky9��B, ��*F��&|���>��7+k�R��z�Z>I!ׁ���}�W@��^��DR�r����(c���맗��k[Ъ`�XpG�G��"
����47J���( �<�S�&v�Ww����'�u{�����Vi���ab+��		W�oW\�2@>�	FԶe�+q�Nh�u��-��Źw|��nH��&� \O5Nr7�6����"��j�Y�xs���Q���uù���χu��˗������0Fu�J�</|
����"|�=�d��[\�'�a# �Pa@�x�('��}قc���d���AL����e���d/�X��� @5�Ӿ� ��(`JN3;?O���I�"5߅�A��eY�x��+k�rZ���-܄M���$84�4�E�m�p�"���L��˟������&C�?�������Ȏ &���-q�u�ʢ�����t�K�&1�$�\�x����2��F3=�;�/�ql}�o��;��}Evg�{9W�v�K���}-�SK=c�he�Ag9�w����X3}K֞@эz�I"_rH��(��`�~����֣Ŵ�l���΂*2G�<�<��15�,�<�'�ښ�Ͳ�/pP��"��U��´v�>W&u>nãUk���.�ځN+跊���į��/__4��w?��}3�,��lxx��ӛ\�Vfc���^�B���Bwk�n���>s�ihQ�qb�R=[���;)/�!F�a9qͿ �#�y���ݨ��l�L�'�|V��W��{:2;A�.҃RM,XW�
�r3Y�ϫ��ek��o�'n��JM߷�6<[i��=�_�ïۗ�n���Fګ2�Qz�$q��LQ1�!.in�w{@�m��e&SavX\�3�8��U�F+{�����l���l:������m��G)U(ë3mt~W�Tn�{fcX�8sI},6o�Z&���[H�L���u`6�1@� &����s\�nZ��/�����
��:�|I�<y�&ǮK�6eW��*��4�F^��Mާ�WWw�0{5=�:Ρ-��mndA9�>|���Cm��6���Pm�%��S$�l=�&8���<�ۻp������7Q�%sp����CȐ1��<ׁB���<��z#��� �	��"����XS[�k�X&��>١�� q��VL�N
�����3d�_-{������~�gkM��>�q�C�fl*6}�ק��X>I�Trk���ٖ���b��<��p_�ng�$���	�x��٣퉎�B6��6�6�E$��Lb%u�Ro�Q(	WQ�����2�`��@�*�_ݬ­e�w�7v��<��_n}9ɻ�v�G?���u��*<,�ß>~�����݃2"1АW++���[�ۗ����5l�S�I�ص���D �:l�
{3�\@]J�v�꺧L��'K�1���a�K$��D�4�ɒ�$'�Oq"��d-���>��TC��w\R0	���n�h�fp��,��i)P�	����o�T�2-m���$ƃ�ԔO��k�;@P.��1l ���>d�Ț'�_
~�5��<{/6YD"�����QYT���(mӡ ���$j@ ���(��G I�&��C�4t�	eD��n�gO��8���23��Gs�ޗ�1@�/��Y-����2j$E_�Ŕ)��-�G�� �͚�Q��mO���Ꝡ���Q-!�R�lEx��~ѡ��ކ�	���O�:�jk�� ��~���߿Z�C_��KD�B̨�+Z+M�Wm���@ہ�<���G�F%}�Y��y�ځ�=h�@��$-=먢,<!�⹋���ۇނ�|z����[칃}��_4ʑ�F��Q9h��Bn��ad}�v�n8+3,8�����
n��EM{񯲨���,z%�-���[w45��v؅�^��ߟ��_ޞ���N;-کSUv��� ����eY�"\�9��I�R/x� �O���)P	]��@k�Mr>]$��Z&�
�����Y^YD*?>}��썌e���4^��Z8�o�1����n� %|�����{���Ca�?K�0��ܑJ��9�q���l���G�?�b
�L%�����o6(Ӎ4�"f�`������j���r��󚦶Mr��`��O�uo�����WOgu�~�!�\;�J��lsˈ� �~���w�v��r�9�	7>]�l�u�L��������JA&��9�x�Y �҉K��Ԭ'�e!����oည4�{�C�o��P�N27�>�k?�ϾZ����/���g�v�"]=?�N�?)����R�J��m-�#g�d�}��#i�e�>%�ڂ��U���f����=��鰣G��Q}d5PrJޫ]k�B���zvn�֮�J"3��0YDa�@'\�={&ǈ^Hb��`֮� 8�mm��]|����4�tE��s[(�6�H�����fJ[|g�Z�����翅�6�b.�s0b܈�Ng��Ɖ�PvD������'���5S9�J\�'��`�g�z�z���9���ᔶ�I�FOMp�ب&�q���
���3�d��|u�#�,Z��I1�]�A�2��#w�#�7�"�s��B��28��`V�`C�^���u���wC`��n���"x�A���Ka���I�Ә6��7ey��L�=�es/&�� ���!��)���99�^T+��ħՑ�,��<�I�+����fY��Dx������2��i8O\}��Y�1h�iCu(��@Wn[�D5I��Q�MY�7�@�0��Tx�$�@�B9s�zr>%a*$-�����'GpS9�Z	�?cM3��^��/�O���S�'��O1��>�
"�ezO/o�=vךf�1	޴m�m'3�����5 ����r��kVI�+��赶���)5q¯��,�b^�A)tY~�`����0���l��� �Zv*�7)��^�j�3L���=,����*���!TV��h~�F�2
[(;t��x<�E<�巟�_���h�RYav��r�egRPf]�q�JNգ}��"��݌�z�$�:�]J���'���*3��5�A�*�M�����e���n��ܔ�zE_A�ç�>�;�.��A������z���t聥Lk�+��&Q���N'm���SS]��)��2�=A���5�fY������X��䵽Ov��$�aʺ�n"�t��CĽ)k�.3�Y�b���Ir��Y��0D�d���-����}
�����>�,{|����V�p�k#ww&ʼs�Snт�fX���l����s��,��0x�vб��J�.����]�L)�.b�2�����
χi(
��Oڨ�{T��ޕr�;�p�n�,��[fAQ,��}$����W�^c6U)��ߓ�[�`�:h�8�uu$�����y�;9��~�C><��s�����q�Æ8�d<��d���@� �U1�l?��[��v��#k$�X����{jP�Qѩ~�T�v�\U\Kɀ-x�J�*�bb�X;��ap�˼=w�I�4w@�� ]��[��8qV�+	CΧ�z1��lľ��]�������e�>���-���?BO�O��)J�Hs���O^^v�q�W����R��2.h�l�=uj���o��I� M=2���N��~G�H?|?*N�D��R�M��P����n�q	4��J�-���R��	uT���"���Os�$�#��]�Y%i�be�8�G�UUC��AT���SoNzY�4:7w�ulT�2[Am�������Ƭt+=&�(�d�м#A�s^(qP��Qr�O&������h���ZO�� ��!XPf����{j�p���"��I;\���Y�Ķ�[B:�<f���M�A�:e``���(���d�N���W;��K� ��p��������:8��^%ӛ��s�i**vd��� ��n1 ����t����ǚ~Թ� �ğ:�+�N{�O��;�[� <W�بq�8o��Y��n�ۣ%��Y��oO�0�b���Wk��?­���XB[������׵�CxZ�Z�f�e�`S˄7��s���kKvH.a4s�ׁ��ݓ�l�������
8���6l_]��<��
��I&� =S�� [Nm;��a����V剓��wiU�F&'
a���R�t�k���ٿڃ�H�in�A��,�B���=dD��v�R���A\A���v�߶��o�C�qˉ�@3�}6vrT�\�7w���m�ia�I���5M����3$�{_�B>~�o����+z`��t8�K� {�2��U'�	m+y1�m�$�А��� ���3��Y�m�6�='���ߖ���Z�w�D�v秔!�'W��g(�Z{ax	�_�iB�^�k�/�����&L| �J��q)xp�˨+G�F)U�ݠY��k��4̿���YߋIh�W��n+�d =��䳍}�,"��6GS���T.~��,جM�ʁ*@ԁh:��Di�k�I���8i��+��l�ɫd�r��b/�w�ָ ��f#�^2Ν�7��S4ꥉ��Ȼo���_��Ƃ���vy�p������V��e�Vt����@�Hv۫'@�"ך�|�bY=@���qʒѪ��y�QԝC=�Y'��ثI�B\M��.�_�Cٸ�Ϛk��K*�38���X*s���-�J�^�n=��9�A-��z.US��Bm�'���"��ʆ��N2�	S��{��w�p�/ ��U5����������º9�����<nvk�� � ����i����\B�3�&�v#Q���E5׉ǔ�G�*��r��N�����Ox�������LAN"��m	~���_�9�����Y4����w��]v���Fʰ���ęJk]g��T�(y<�Ig3��ܹS� �>��.=7��]̏u���E�'�t�~����i���W����A��g:����J%�D$Ŵ�3M�话U6��0:��G�^���H!O�Y�s�\�Ų4�r2���CY�J&dm��P��p���a5*E�j}�'T�l>-�/�8N�E-D�D�`l�6r��3����y^㬌�����_��W��Շ>�{eҴ��l� �k�����w�:Wzϔ��]�Y� C[Q���ε��9&��c�zɺq��Ji
,��j:X�iu��s��5���������`�^��"����ǗW�E��ѭ���]x���i�]������:A87`��\i���������W��?�|s[6��<|�DO�ח������Z��E��@�on�������'Q���X^ڝ|K���=!���F���T��c��v �.��D��4�L�'驱8�F����l���iSP�7zpd���656t*q�K��S����Ry�8�*%'�qy���C�
4H�x�4�L��R|(/?��AA�yK��!�M~���!�A�k����J���Er�
I���{�� ���I�a:#���=���@��H�n���h�8�Q�X�C���^�3�)�Q�I��)@�@������B�EqY
Ǉ�k	F�gĕ��R��Z�կ���l2����yJ'�)f�yn�v��P�A����$��u��ugU1�̘�VM�z�I�Ɏ }�W��<D^ZH�t==�_���禗BU"@���]t^���X0_Z@�E��C?
��E�řU0�R�|�s�d"'�G\GgAPJ�r%m��Q �(v�۬(Y��j|AC���cҡ @��:�����.��z_�����{���~z�Ug;�&(X8a��>]�[�[�[+����(C|�.��+�G����F�W�r"�6��[����2���֘Vjs�ַ�E0pa��T���Û=��v��ŕ&��݀"�Oc�&#�=���r�`��Tds�,?S7��V�BA�f ʯ����9����fwq�� !����UXo�WSU鸴N�D���,���:L��8��̋�L.�,$a��s(���M
$ɔ�&y���)�@EJ� ��T�0r�����i8r���eG��Nz\A�y�+{�W���u��A�A�����)�=�]nk������6�A�ž`�Y�EO^� ���b�_f%�Wb+�c��(+2���˟ס�Bq�%a�Ԟ�Kv}Y6��G�,�����c�ҧ��c֣�T8�|6��%␅�V}�� +'Z3|�@"�"��r�}^��g9�嚸RZI�{� ������-����� ��9余�Hf�!Nl1��zi���:�޲:+�Eq����,��֓f��P$�#�N�V琗V�z���+�d�ә�Q/��<Bw��β���7$�W}��Fp�t"�%\ْ����p܇�ۗP~�r��M��t;_��l���\�������ه�pu�����p{/B9�+7B�oo��o?�~}~{� �z%�1ѕ�Ej�6-s����86����`ԜC���h�c[6�͖1a �/�hD�S]�a4���@K�>(����*���篏44J�Ё.��S�t�;(�҂�P#y��˼1�]E����1_S�^��.���O;���R�&E��
FY�T����E��EqN��ٺU�!����;��wp��Z�K��m�d�S�4e����5� a��b��aHe���sIf��wrNe���/�OѪ ������,C������	���X3�����Z�;M��F9n�(��fP5�&	�}�½��YK8NnF!�k�*�\�A��|��36wku8��6x�YRk�-��{.��� =9�f�J&��8�;��@�S}A�F����Z�,^[FG�Ũ�쾿j;������8�W;��(ap���,�@Y(��ZL�5F?T}@@1��2���⡓� c��̈��*��)kk��$޹>����vP�fEv���W�����a���Β�uXb�z�Q}K0��ve��흝����5<n�$U�z����`�ݡC�
���MC�ˢk�\���i���{Cd�i�,͵����1��\`�{su�����L��,=��� �&�>�~w��Q8�Ǘ'Q�$�5`��.6C@YΧ�>��i�U�qxW!����kǒAi�$aK�2�:*ݎ �c*X
�}	~z����i6�^zIRG9�����(�����KV�5��,�4�琽ϧWe����H3<�{^�
�1�8
�������Tm���_ځy�����3&���)+�l>�tϒϮ��~�f:X���k8}}	��&�N�&��z��	���ʲ�X�
3�_<5 r�@�
�����N����W�d�d��w�ƞT��3>˰����FL)��(����C/�;����	y>�RJꭡ�Q�.t�{�M�cj^��##��O���O���f� ���YZRR�7�z�!$|��q�uI-�i�5�;��V������p�R��ԝ� ����ȸ��~�cv�����{M�k���#���)&U[=���YV�5�PXz?�4�LY���^�҅�q��ܼ�
����%l�{���sB]����s�[1�=��l��T7~M��p�rx�l {�R�kKza��a-�!w%�l iX�CA�?1���_���Ls��1e�+*�:kܗ8˲�&�|M#iw��閜�\Om�܏�NeU'�m%.+������x�p�2��wK^¯]�_4�T/���]��!��T0��ˤZ|�j���1S��}q��)�;�*G�X��; �`�^]���.ј�A�6�3X�j��BnP�Ct�&��>꾌2���K��-��������$32�����p����ˤp���C�"�>n�kx���<�����#�_�:�R����]���}i	���Á`�;L$s2/e���6mL�-����.n~�eH]&[N\��e5��o(P�|~~�=>Y�;���)PM�tdm���Ya�ϸ7tF�xI���CS��{��\��y�QA�iv=�0 ��܀ay+��To��!��=�S�q�Cʴ	4�����A5u�S�����R�=7��cX�b��\��AS�eh���L},��y��������ihW.�L�����Y"�mr��W��)N���J>��!�b�t
��㐘�Y��g�v��<y`bQV�f���u��2��7��!�����u>�e�=�ݫT���Z�aDZg#	�U��۪j����IT)>E�T��y�\�$��&ҼNR�I��v�H������.,�1D��!��?y�� $���I�+;ܶ����B�w{6x���P� e��	Ы�C;-��ݡ9�I����aa����*�ȋe��E(�֗��N�_��.�X�3Rf�G�wHEi��h%�XՃm	L�ȴDh����ص��]d�d�ݸ��'�{�;D%� ��l�
����։������i}h!����'����NQ�����n#�KXo����ԕ�\\�<�t�M}�,�(� �s������ڒ��F��^9��3v�P�n���=k-�#QxS�q��/5�c
)U˭UP��=�Mxۼ���]x���,�)a_{}���TM�<�e��bc�~C(HYvy��bHc�6�4+UTe�]Y�i7z.�4|�]�n�H�t�tRFh�؜iB�Ol���޲���ߔj;
�:��H�a(\��D�?�u9N ���&w0Rߟ`�ɩ�d�@�1g����Rp���� �S���p]lN�Ys{ �.�ݫ�\?>>���d,=�=2ѭ�(u��!|�A;�t�$�c]�@f�*K��j4�����,�����ep�J��?dޣ7����G��#�%���Qooyu5x?$e�wS��j I�h�C`ui����)���r�>v��a�ԣ��pb������-l�����^�d}d%S�&���o�E��["��/PL[�&�쵯,���׭��
e��W��: D�_TY��HYv:+$1_R����lW�;5%O"��3<d��?�G�����;W���,R�
����'NO�ޟu�� '���]F5Rk�M'3i��S�XH����%z�������e��t��[=6��`�XM#y(`=dn������:jr�hR�+�@l�W=)�7nU���lo�˱��Z�\4U?�j�!�!b�a���ˠ~���ҍeN��4J��`ԲpQ��|s���l����[��^m��44�+��.[�̨�SG-��#��b�{?���[��#i�\���t�T!UЎ� 0���)<�fa�����B��c��E*� �8����no����N�ۻ����?��wW�E^���2Q
�� Ǔ?'�Av���Zܛ��iX�""(w,���.S���q�6ejͥ���A���E��oޤ�{���.FP��Ր�x�t��@��=���*�gT ���P��M�ļ����5q8�: K)�C+��dNl�	��.BI��JQz��嘤�P#QO6����`b�{{fӥ%��(�U�ѷU�j�6ZS�=,�(����7�� >��~�t�=���m�|9Z�cZ���a�@ǋ�3�O�"�-z��Y�+���G���`��0�@�T�T�=SR��5;��l�~�h����'�����R��Dy}(a;�_���a�
�da��h{��oU�5�7�`0l�#LD��r�|�>�������������H�O.����)!#vW�E�|}���?��3�nȖB#����Z���Uq��\geYb��ۛ0��_�p޾��V�ި��]�4ki>G�g��K5���(
D�T�D9
�x���,s�e--�/Y�y�~�dR����}J(�T������ p�A��������#�H'OIj��� ��b�ɣbEe2��vcSv�T_T���ܒ��!��w��o�4Dh�1!��Lk���C�&rt{ٰ����Lê���wx�&i�������U�6̣墸�t�-�'�	�F�_-�PNU�g��<j�P8�]"�� ��Q�j��J��룊p&�t�Gn����Cx��.e*A�G��o�.���/�w(ŔQ`K>$��R/4�ݾұ�����q{ �tO�x�2�v����'�������q���@ok�Z=	:��dD~:J���󎲳��~����r*qm��e��4աM�L�J�����Qy�#p1H,h-� ��C���? ?Zb�7n]!�"�;�a!�aD)n��5��Z���6�x�1|� ��-�ۆ��j��Ɔ']�2�
�۫��M�@2���WJ�t&�����l7h+3�Ȁ�A�t�2�2�^�[�!9��s+��d��&m���o�X��pc"�;ᏽh[:�#h�;���<�_��
O/�x08Ee�N�,
��(U	�X� �O&�>T�}C9/�����;(*Y����w9x6�r��->I7����,�����a*�h�Č��: ��K;��?��ݐ�)ifm^�C���]��W���eػ�t�ʖ�]�1�f�}ꁌ��?�-x%,�W��J���o�sɇK��Hlȧ^`����������v��$�,��X����@���ޠ�!mD�,Q��E�[�ķ�gbc �Y)n����)�\~ۃE�7������Et��ʳ�\����T;ʵgY�"���R��!v�>h)����B���j���M�zO"�o��9�B���ͽ��2F�TxZ}�}�����g#)��{k�(Gg0Qh��������m8�&3[D�d�m�]���b��G� �����~X^���*W���NJ�������G���B(��N�۰�����]�����J��+�W�a~{�O�/?[�l��R�IP0xI7��f�l!_N ��B�DG�SG���6�����в���?�c�'u���C^2ש�cϋEΐ �}@���I���\k�*���q*�kR�MAC�B��l��1�TH�_Reo�Ҕ�'�w2V�5q8J�����������좢ˡ�����.�Gi`�x>ꋤ��6F��-�l���bI,y"���綦��P��X0�=�������P�JW�p�ę	��P��z�l�W"ӦԷ �d1-�� wG�5� �����,�m��h�,٠��%�1��W���gC0S��8VO+%�+~��͇3�_4�)�{d�����@�ӿ��;�5�?��gRvRJ�dw�_�szN���V B���$��ϧ�@i��&X����ry�S���2�I�\�JmG�{�����	�nyQ���<���W�XZ���	�����~x�~\�;E�ٞ�5�*�O����HSѺ�-�U�*�@����J�o>�b�
��~��8��odM/�OX0��S�\��Ne)&�2�s�����hg���X�iQ,�f/,S c���!|��ѧ���K��t�S����	륖O%9�XD��V.�IY���Rϯ��*{�%���|��3UB}{�4)�*bɓN޴໨���	������w�I�lk;�޴r��[Y��$����C/*�����O�R4��_L�9�
��x
}H@C���\	���,��ώ �.�pc�w���G��S�\��U&b�q�sԫ-$�K��K�L8�3���N[�L%\���A�����HRPnUS����9y=m���ɴ�R·�ArފnU��#��9�`�8;F��_�M��8i�i����y�z2�j�$��QE�u_��4�i@�����&I�Z���`#27z�P7�^8<T�0�o1y/=��b����#�2s������ۿ��ڍ)��9p��4���+�&�--�w_۵��y}
?Yp�g�;���=I�t)r���>L� �M`ѮW��S��|�?J������~q�t��)���;%�Si����� a��n�s����F�����׏@{��؇�v����TZ��ցļ&oܶ��fSzh��zP����.ڗ������5�]�݋;�e��N&W�6\z]���>�K�R:�Ԫ��L,����w6�nV��qFy;�b�gE�/��\�K��#�@�	�!��H�k��p�k�ӟ$���y{RP8#V��go5�����ܾ��2
��G�RJ��'�L�'��ڝ;�k��-u�U�!�15
�m�]	�3���A+���
�g.]ފ�Xk"�.Um�0�q��|��� ɒ�{�<߹U9w��2�'�dВZ�z����UG%bLǽ����-{�΃�l�=ۨ��(O���V����D�����P����O��d�B����A̐d�������;���d�~�bտ���E_��Dn3'��E'��a��~/'��o$ ��j��Z$lP/�����nBѶj��H�j?�z~���+��O-<ZM�Xx��>=����)��u� ����\���s�##fp���Q��Y-�#��3zlL�l��6oZU�Z�z2]�	Äԋ�����S�H�;�<�+{��2%pSyTc�ʪ�"�Mam�B�H����`�Iy�d��0�[�����s���WYyp9C$n�y��<�ŢpdYE�o&� �!�$^�,�E�U*����U�{1��\C��Zzf�
x�n��έDZ��XL�6qu��m����0%�vvX�8��|�aI��������!C<Ἃ
,�ot�a�-��B!�L�6)�������j���S�|!~�;�O����q�٪�V9x��s.sf���d�Ro�(p}����Q^*!	�,�����2\������hBk��Cye��C�f\�,S��(e^E6�=��b&޸�h|�^�]}�Kb���)����@����o_ �����|q-����iqM\����_��(���^M��{C�y���-��lW;�v��9���E��No�]��"��X���_�Gt��g�V�.sW0)	�7�k�(˒�
��}H�\��O��ۄ/����n�L�<u�I��޿�/�:���qc`-?�1�Y�j�fV�Hf��7�3l�7���g ךXFm6ъ�Fq*Ejc����;E�:eNg���g���
�2���D�u+�;�ɝN5cE�/����k+�s}�|���40w�����RJ���q��`v�>���"
��ԋb�e���t������2e2_����{��N�!��m#��l�� ;�ҳ6��Ь(��!��WM���&x	C0��&�J��VbU�����ڏ�=˜�|�Yz-�����3%0��za\�Q�WY+������;C��2�:7���� ­-U�/#� <�0w�9�ץ����Q(��C�~ԃʽZ�$�5|�u��Y,�`��F�������@|]d>`T��5�H��A�	9��O%����Gqݷ
�z��j��z�kV)̪��hk���ev�/6���տ��72��8�gG|j�g��E��9��|9�B�b%�I���wGJ�	���7j��gz���[A�Fo/����xޅ���=�}w
��6�Y�B��k���Hե��N%j�{~���_j�ίV:=x����Yׄ�( �H�����j�P�,�e�����!���8�V'^�b:u<^l�Xp�������)y]��z%%�N�|)�D�3�X��NB�����X,v�8��[�rs{����$J���c�B-�I��_�������{]��)j*3S�3�Hmw��x��/vG�����Qr[:h� ܥed�el�}Nzh��'�F��J�`(q��6���ԃ}���2XMꢹN:hryL�/���C%�/��(H�
([���K1T��22���1�.���t3b2k*�J����.B���\�5Y�3�=���O&��"�݂e�&V.�U{�6��-�X����͑@zm�'QEG��R���.jEժ,f_��Ƃ�l�b�e��5'���:�gy�!KJ�[m�x>�k��HF����E�9��𸆼��}�
}V��$�X�؉UrS2Q�g��Je�>�O�b�HӘ �I.�T�:��է@����l�%��B�C�D�ݜ��'7��rH�%�#oz:P5D�z=+��AUp"��J*�>��$LIР*Ji���xpB�'R��(�tќ�r�$�9��\�����(����J2�Rt�p2uz�b�mqB+����HcqS��V�ci���az�~�n��Uݐ�i�EJW➦�8��M��tq����q�B��xm�=,�P��o���2�S0�DMu5�Kg��p�gB)�>��<�j���>E�Ĵ�����٦L>���؀~L,�#ր�'	���|�FA%lpY�8Y澒��N�Ke�Dx��^"	���%��	�el�k�:���9��duM����H2VY̺��ԹC?�Y�:p��)�yxN������m�/�C�(k��������(k��F�g�� ��,�=�d�h��,	���6��F��2��g�{=d��yUQ�W�g7Ϭ�M��[7ZHv'���m�v%���C;�6j�V*op�.�n7 �,C$�Z!�}g2��9[���μt9�^���Ȣx�d`�1�G�G9}2�X:H��Q��3�꺰f�������n��A��X1ݱ�1//�{��x���T��͌�����!����]�Ud���.�Z��<d7��F�9�W²������P�-, �?<8��>%!���@-jM�r-���nqr�z�
����6�%��8xӬ���Tj��E�&m,֬SƧ-�D-S�}�Qy"��<�J�����3 �?1(p�M�G��`>$_�ʧ�*K��(}LTk�����RF�ŬU�IeXA�+�K��d�K�v���R(��$/\X	�֛���uU4���v�^���T�Ƚ��1�̕��u�C�t����G�(�^fF�!x	o��~g_���d�xO��EHӴ�F��\Y[*�%��r��,e��.�Kz ��U=�r����9z �Ş�����fK�$I�����GF�uuuw�l/0���+�'�?��3?| �@�ݝ�9������������"jٵ��E�^����fj�",�,�f�[����4�H��H�r�������������#x
ɬ�x��`��[o&)z�Ӊ327������Sms�ŉ�s/�&�RHk0����ԙ���,�	n�]T	�^��jS�M"���x���"��ߜ�,��r� `|I�-�Y�Ӫ"�ɋt���w�grZD�A�����sެ��{#se@qN�Ɂ\~&���]�/��4�4�6v}�\͌�������j���\ �T�K�@:�fK���m����K\Q6�2[w[h�8���ЫW��&�혌�.#o��gt�0�Ux�&2����:Nv��X�*h��>��ls�TCOP�B��?���F<��j};�G7��Ӗ�y���[����V3m�I�ѓKWt�����&Ɇ�f��hu�ud-��z����m�E\K�G�RA�����ߺ.n޽�E��}#�>��p��5H>\MX`5�\r> �I����5��9�,�b�u+�V�YN�xoťs\7�e9`Kϑ�y<}�̍�ԧ��B; v�L��qr�0��c��0��H�K������u��iΨ֍$~LW�2gP���Gvl�$��0����gP|],��yNl*Ljb$a���ğ6��������S ��}�]=&PE��`�B���3��R��Ր�����5��L�p�`s�e���2����1��]�(k$��44��������ܝ�2:�1}]Y���Osɒe�c����������$C#�1�2�R��t���Y��z��1��D�����P� �Z�xD�7�;�b��@���	^��ѡ��5�6�3�W�p�A�� ap�`n�紣����f�;�ED���r�ԏ̌��7LV5��B�
!�Jt�b'֟�	�w���j63�pՑ�=��1<�t,rV��x������L�ח�Y4/_��߱��T���$<�04���-�~&���d3%)LO�y_I>5٩�d�����3�b4bܣ�޾�[)�jY�I�D����u^又���Е�mj:�%��fk�vv�,t�,.�ث@�ט�Y�1#[���� 쉤�A>n�͘N��W46)
��D�!��
�x��3C����\?)�+��!��j5r��S��*Q�h�`�wu~a�Ƃ�z��+��\�sr�'�go���! ��8jM��{��'��s��8��L�k�t_��e��ޟX������dn9ͳL�t���W�������gk�9�0��������@�GOx _l�9�|�V�8�^���gAPY�j(o���o���U�� ��j��=����4�7'�as��%iۻ�{5�<`�M[�A.(g��*)w:���E:��^�w���Y��rv�%i2�q1����??��t*���</��"?w��6���	�1&�����$u-��M�)�����=�\O� �4pU:� ����ؼB��Q�<�Lj���s\�jN{2=�$Y��~��J�/��tU�֑CT�55zeR��ܕ�#���a�ꍹˢ']ü[%:���Ibj3�y"EM��0�$n]�1��T�%�\�QȎ��6.�1�lp��Qt��Y�G�-;�%i�X!�V
&('��J��10��T<aS}�;��(�V�;�3ag�hݞ:�w��}p.'r{@�Y	]0��=�:6�nn^kZF��w�ʤL/Ks�$�51�R\=丙d!g��&�a��u����Q��=���hu�g�L�Y:� C]��'����B�N����L�mw����Lm�avR,�G�Qa!�\/J>��b[���e\S��sV��2�I��I%>��H�;�;�t(�����D�#�~��j�+2&eG���ɓZ�^p�_��� ʉox�]fe��>|Y_���h4@�^�>����78�u3dfxy��AvO�zb� a���i�A�I�z�����/.��������M���l8A�(Xx�cǡ��
����2_*?|v�����
�q�Z:�08Y�Q�:0���fj��v1s��R�h�̗��ƻ�~s�>AcG%w�+NH.�4R���Ld�Tk����c�يgySKU�@k������W7���3��tG�2ʃ��n���.�q�h[�h��۩.@��B�C�9�'��9W�|�w@:��y�L�$�;�V�y<���`5��x��P�M��,��?�YӨ�d��,�۸^�E��hf�����/
�-�����A�~�]}��Z\;��EP+1�$�D*�5g˭�N/�):}���
X����󨮵y�Dj��^�a�f	,��V�=�F�'M,,0}$T�t�p&q��1#��V}{���ϙ����(�D��;\�34���؃zl�����Dk�%%�m;2E_N���>=Cd�+���8��� u#~����]��o��M���4r�aäw,ϱo�=�[9<2N��[�&c�����9P���B��M�-�����Ϲ�����f<��֦��ʭ������]���\���ٖi�2sk��gr�.��̡���GP�6�jK��o��=�i��	Ǖ�8:���T�'(�lB��`�-jtZ��pz����1�,������"�L�Zwp����D�����v�0(^�&�֬5,�����6#{s�Xl�t�\̸e|�2V�KM]��u��#��Įga)/Q6��U��C5rO3n�}�l�cjA	�!۟I7o
z@j���+�f'	mV"k�i,M�IL��Ɓ��!s�#-�N����;�e�M�e&��=á>�>e+e(u~.zJ�0e���לv&u�T�5��o1���\�~{� ����mjN~BI}�յ�"�
]��3��ֿå���TJ�*B�%w�Ǽf�ܚ�p|�n�X��.���U�Z�^@��G���롑��X_O��A����w�i���@A��p\����r��cb�|{v�  -6��i<�;� �O?�r�B>&�K�*��J��h�7�����I�ғ��ȝ�P��]ۍ�Ѻ��yA>�S�=�(�Y��F�EK�x`uZ�uRP����i=PQ����G�s�Bٗ��%�Z�3�%6�B��"�']U`95�n V�[g*5�E��dZ���1�������P�|i�n�@5E�6<����Ʊ|����|<�I=C�ct�%(�PQt����;oSozȢ�9���$�v���°r+#�x2���H�0E��L�/��\h�y�p@}�LQ���@q&q��������5��:�|h���	�8fL��$z�捎��,Ae]-�)ɺ�Kƭ����}�]�(��Բ�����`B��_�� �=itaw�1ˢEz�簃��#�O��A+���q����+��IAR7��[)�fa��^��Paj8+�S�J��X�ԫ^&|Τٺ�sJ{�;!%���;����� zV�}�=@�s��.3�s:Mc����a9[��� 3;��6�bxqnc~��Me$ybVZ�~T�a��X<c��0/q�f�^�(q>Τc����I� �Xpe5*��!ȖP0�����9�	J�����27^b{���� ��Zd���'���鯘�y}��{- y:���g���22,��/?�Z\]sVkQ���f�=��<P�]ߚ��&��8�� e(��h��4�.H��L%��r�;UI��	sM*Ki�ǻ�Sn:���ȶ8r���وQsO�o�C�ה�Gh[��!���X gK�0��=�;у˯�ԟ�TE	�!)p�%���P�}�Ӫy�on���yd��Y)[��>�ߜq���Y�{{��F3m������Wp3T�z��Я4O�.��̌;SҺr�f���D���Q�<����;�4� k�y88��gord&�k4.���z��T�Z����G _���~6Ӂk��_���!�4�k�S�3�B!�.�~�)-���d2�7�(�®Z;F�S�w{J����xf�����n�2�
U�\d�X�'/Gr���i}�N��f��f@}�NmY`E$��5�T �\���*3�w�E�'	�"���@�ĂA��SY u��8K�p+wD�F\���ܸs���!�25��.(ɿ�?g�VE��Nn� ���ȵ�����fAG��D`C�;�
F�; �j�S�I�	�lf�@������^ѫ�Ό-�fd>{41���g��ѧ&Ѿ���93tgrq��tx�#�(k�����H�����W�*��I�ا��$	PE];�A@�����Y�p?�ĥu&Hտ�{{��Ng_��V[t:W�ϝ8��^�#>c�k�|�^v�n�������^o�bk�MlG���5{�I�t8��cs$������	l�}�6�\���f;l7pzd[���l���C�A��H	��:ql`Iɵ�
+�?��xn���qMr��L�&�8v�(�#�x7nt���%}靕��D��Ŏ���+Ǖ,nltKp9��*@��#��F��v1��l���t�t�"a��F_�Q�kq�A�H�+o�uA��5;��2G��y7�P2�=c�����k�(������En�Ef�3.�ˡ��w�8����O�˜\���@t7�(��Ʌ��&eV̤Pz�>F�b﵂�y�Ɍt��Kc?o6�}���Fy��Md�tA���/w2翕�?
���������	.�"�*��QY2]y�fd�|����Q<�����;��v4WD��k���Rq8�8��J�(��X�+�Np��)i�2�=�t{����p�٦��እYv��	�x1��t"�Ou	�6�ݠ/ޮ�lظ����{&\�ܢ�Np6��B�9�M��
A�P����|��]a�v�MQ��4	��v�;	�dO�D�
��s{#����������z.vRj�0�K3�^UO��ni5��+o3+��AD� �0TA��;��,�^G�D��ͥZrp�k�YD��??N)�l�eI��Sͥ�q\�T�t��L����V� 2� 1�!7(=pӣ���4dN�+(��`ef�F�����5�wS�.pL�8q�SoΒ���ٌ#i*A,@� ޅ����#B�gi��䛡�͉D*P>2P�ə${�h
c~]�3�.�919dR�8�Y]�.��7��;6��Ғ�6Bބ��7�BÂ~4�t \���)�~B[�v�F4j@w�H�2��ˍl!�yZ�w��L�<��2%�9�/	�?	�P�Y�?6:�����vG<Q^z������05wр���=f�d �c�'���&�yP�}��|��%���#���q���f�R0�	Z��Sm����H���7����� �9����l�0@	�_�E=����k��b�0�Iڣt�|�=�J��/���@�Lz��0tJ���A|1�u��lTL��č�F�ٯ��ėB�sH�V4��s8�z��2O���xl�AF����q���^q̫8�.lO��7fO)��AxOk���(+C&��[E�۝'����N򫓨)G���v��7�I��l@��x��f�?X�d��#ٌܱ�o:�\���� ����n��&��S��T�;�OY��t�nXv
��B��໒��K�)�m`���*aW��`P��s��Q:��J������`��;2s�2�Ǎ�a�Bk:Nr�.^��q�#�I��ߒ��Qjdb����(0��F�4�.i��i�AB���Ժ���%x��\�^���t����V�-�5��s�$�
��I�Q�
�cl*]O��vg7��k-��F���_=bF���햍��80g9 C>��>�M��;.P�v���A6V[f��t��=s��XF��I�%d�p��0�U���]l.��⑝]>�#��0��5�g�L���X���'�$��4"5�X�m��hrG�M�Q ަroi����/ &�SI�ZĂ�i�e���9d=��D~A���s2oZ0�$֣�8��tD���]U��Щ��c�E]G����PL��QG��M
n��*N`��-do�`uF!5��A����NA]�u'���ɛ�n�}����)�O��<���.i��'�����z���z*��'��
!�b�}r:Lav�cQ�k<�$�6#�w�'��hn�ML���]��E�ɑX���,g���d��3DGs�g�s5a̐��e��V&'ň�E�n��vu(��� fH:����푧��x���7i���ܹ��hL��&��n�M��9 ^���9q� ��h~\��6���k{{s����F�nO,�;�a<���α�pI	�B���՚�+��)���*j�N�a@��[Y��2C.8��ĵ��AY%Z;�>@���W؞���qn
����y�z�	��۪�x������Ā��^���#uk�B�����F���7�YNa�����.߅�Z�o�u+s�1ج�����%��x�,���%pJ�]�xq���rr>�e�=(1�4���vr���@]�����	J%������,�Eo,�8W ����9���Qr�^��Ar_z�����������i ܙB8�cv��#Ae��Q�(����("$��h�x�;h������2��_z��T�,� ;w�1�5���K��Ι�y�t{ח�q��:Q�	,�0pp��藇�b��TԌ D:���.��L,N��2m�7zO�x�M�M���2��:��$���-�����o޲K�Ƥ$�fZ�m�yP]�'�3�i8�U��	�3X���}�~�H`�NK!�á����f�RNJU��n�����ʅ�����P\���p�a95�=�f+�s�H8?Nui.�͝;^�4�G肺�>1��w|k�������M�������5�5����E�4��[���e�w���`sn2KNJ�-�9��+��ZS�Q��8W��{V��D,4��z&��:����m��=���!�$�Fc�(I��f���E�:W�3l��y�L:����b�B0���4Ռ��N�S\Y�ͤw�� @��N�x�%�T�3�����9gg�� p��<������$��bS#��Ӕ6�5��O��*
|'a>f�3�,������=;�:eΒ Z�8����+!��T,��Y8�ʇaGw:6}�LP2ǚ����m��	�Q�Av��'�rV���y}�������.n i�XB�C���%z��c9'�Y����Ɇ�S<O�̊�
hy{v�7�5�>�42H��7�L]4�Ҡ �j�C�;A&0�<���f��'��A�0��nI�]�<��e���Ew&vf���gk��9Q�˸V��/-�E�(nGzUb�ql��Kfn�0=8x>�(o��[��o
^67\[G�k� �	�
��|�*gp��W���ѐ�&��ÃLAn6 �c����\��1�iu�K�_��ьVH�%.fN��ݲ���%��"�jz`����Z���u��f��2+W��ۺ>7�TY�g��{ސP�U�[��6g�{�X��#��s��ś�آý���Ϭ����Xl�x_��w��2���t�&��C�Kl8Rߘw�KSZ转���l��Z��\�;娡.75S���j_�5��s���=<��p���$�{Z�'�U1Ώ`c��^ꑓ��2N�N�؄QY�9
�dlX80��Y^taJ��&�1&��h  (�L��º��v��\j��C!��s*j�����en�?EY��Z��.�>��1IzTA/2��?���̓f�:��:�2cP|�B�\����5����������ˍy�L.K�:kA��%��ݲK�X��Z̩�7)�gS�$���0��Y񛬸�K8^M�᧸Ɩ���?�ò���(��iej�+q�C���B�
@�s��V��k�����AZ����7)1�L�(;]Wf�B����V]n��iQd�h! �i"כك��(�J:(�F��9���Ö��ճ.��s{�0�4�}Sd�E� l��2��6[]��:Q�Ĝ�N��Kkv,���؍rk8բ�	+p�2X����9g"fٳK{�.�qֆO�F�	��.��6�w��Ъo��a���e��]_(v����nO$4�#/g�2Ct#V|%��-UH��~�Y�G���QW�.cY��@��'��_�t}��M��w1�5b5��@����j&�zŹ�`O&'���R{6���習�XK���	ѣLN��$edʬ�\���<����4��,]}�uo����t!��۱X�ytbq�2E���.�-�W��rO�_���2߳��K��Hʜ%�T�e/)���|�`�:�ϋ��0;bd�I3=	x׭U3�-n�;@r7h7p�鄓�c�2(���rȳ?ZO��H_q�-�X���u"�Z5�	AEy�,���b\A$��6j��yƀy"��8�D�v-�S��y�J�������}�v�]+O�k�R�$,	�V�X�#дf`.��P�]�=�L�ur8�����ɟ����p/Y����;ȹ�d�ZQ��-���!�Z65j&|�B�*��um���g6Gc˽��6��n��_�di��^�d5mnPL>����]-�{N�;E-���W��?ą�����09Z�4�7�.�ì���g�'�����A�e���y7�1�����2�wq�'��у#|��l�wY,��xY4��-Kϼ�]������g���%uGy{�&�uR��)��dE��M �:�35_���8��iY�|��ܪi66ȑݦ���c�b`S�v���nGo8�Ynw���.�5�xb۫K{����@6�a%hxt�|��YK�q��YA��ڻ�<����C[ĺ�}�n* �4�L�Rv��z�Ex��b>���D��GQ�D�620ȱ�J��]}�?���c�zJf-�L4�a��)��	s�)�Sklu�MG�d%b9)��jv5W"y����d����C3%f�whB�ƴ�bA�^5()��9#x]LF�B������J�5ЈXq�G/�v�m��䃻���t�j0��j�7���ۗ�>����!7���_��g�a��%�D4��ǔ_��O��"�h�.���N���3�1���R�d�bmW����1��n�E��qϜD���?�E)���q\��F�	�R�H8�ytB)1��J�R�����hx�G�g���c����&ޚ\��f���$8�O���q����E������C��let�$���	"�1�('t�A���ݛw��>��䃶��g���(.ף�OX�"C�_�����jH�'	�GΖն@���[���QcȄR$繩$\�DH���V&;��+R��[YPj�.~��ɚ���l]%�V=�=�</}c'Ԝ[7	�Jd�EʸQ�,'�Nf�b|����(YN0�jZ!��� ��sJ�,����Ӡ�8�ʝO�C���Q֙�t�g�4�L���)�Fr�E�����]���;ylF`D�9;���S@���$#��� '�1�浩χ%(gѺc�+��׷w��n�?޾�{��^,�9���^�6������$��&��3��e)��*�R�cE�ˁM���7��+'�a����Uf��2	zF��D��|G�Y�b�N����D���E�?�̇Sb�W�ʝ���y�ſ��KzA���4S@V�(Q��}�F~ˎ��Ϡ�����A������W�^�c敞�P�ת�~���v��2�s=nH�1�tg��?�ͳ+{|qi�Zfܲsz�����[XeY�/��!3�z��k�N�ƞ��<�dP<`Lb�s�N�6��y�y)ȍ�
�cTQgw�1��(S�=��J���I��T�n�!�g�!Gbk,Y��6&��A���Z�k�X���p�,�'|6H��N����w?� v���lM���4�!� ��斢}Ƞ:W�f))\M���k�n|����\d���t�}B\���{���5kCc����>�vU��NE%8���I����:����_�����s _�3r��z�	��`�:��gX ��ym�Lm�xIZ�	/��9�#��w��/��4S"�3yB�� �'	\����o^���⹣�r\� x��*�(�`��MH'a�z1���;���������U��f2��`�Զ4/��^�b�G���L��1����ѡ�eFi����h���>�%����v~��L�Xw�p=��{&�'��A �%6?K.�ʍ�f���$��L	�(�U�
Idc@�*p����R��w�d?E[!H�(n?6�!ƥ�҉�'���{�i���)��dۖUS`���?,�9���O���mv��7��Ec��i�M�i-+�&Y�p<8�H�Ѣ�Яxn�;eu��n�o�vwǌ%<�adn4(&������~S3y�%N�]�3��k8jsSv
��x��1nǓ�����(�!���=n=�L���Y�6�JV]7�W�<�O<~�7����#�X`j�sf^X��v�w��#-�Լ���#k�M7nP�F)��-2��%z[pю���Y��o!�E=��Bх����� b��h�L�e���0t!��!:�:�f%���M-�:ny���n�jP�{S�3��@q�����F� ��ʈp���ڃ����s���&����i�	Lǀ��j~?-2!�S뚦F�%v��F)��i��^��#�Y�� t�$R�<p��D�ۚu �ƹ9��o�v���>��G��3��	z G���w/}�� �!`T�f���nr:��+�g�IVs�-6��Y[����2�R[��<L]ɖ�2�,��'�W)aO�u�L��z/yG�w��'�q:����Xs?f��@@���a���2��
3�uQ@�Ae�,�Q���tSK��~�.���rp�z<pN��]=��g�W����ʴ�&�����y��t�-sZ�0ˋԲ)��Z��6Fw��%2�$��M���"�"���{�آ�ѳk7L���G�h
V3\/�e��sr�1�KT���='�ꈳ�y��|��
�:�-�ظN�7�2̥We1(�?��	�R��WE�q66:}���)Z�j�������yH
�(�'� �i"I�6NSG�v���4�gsqs��r�l��U�CF��wM��?7 ��D�Q��$�z �Aꎋ�sE����zc��aep5�C��8I���/�q�y��h���'�:�)���E�g�İ3��4��E%�y+lNsmy���_��y���_v)�,԰ˈ��-_�Hmz�����U/�O�O���|�bD#8I�Z����L�����O���܌l�xl2_�XǾ۲;��খ�����k�]=��
я��yU����g..l=$f۷����������@����:�>c)-	��v�x$�R�*�O�A����f�_/��d��ȎP"���R~�P���x�� :J7��
0Fw��Xl67K�����;��Klf�r�QS���F,�ZY��6I�b�-�����D��an.t�u���H�x�n8f3ѺxCWB�99.VB ��؂�3�q�P� �y)ۜ��F�י��aoID��Z�,����4�S0y^��-v�����&w5sĈ���;�z�a#���X]N���u�3��<^>z��X�;:���n1"��=�^i(c��i�q>�UŨA3�8,��F��9�:p6��ۍs�v�XZ�X���+Q�$[T9O�r6��`��Y��25�[]��p����s"��R����E'�P96�sAr��P~���l�����o�vĵ8���Y`�܍�Eb��	kt�^y��`|Ju��x
�R��R�Uk*���i���]�S��ġ́o\dlKR�dKn'��N�{�e���WmǗ����[������O)X�&�~��M 'K�Ԩ���~a�g�lM��$��r��0$J�x �%�Y�H�-z;F~u��X(eBn;=7dY�C�M]z�e�Ԡ�OeE�e��˫+��	�~&L�Z�� e�fm_������^'n4)� �U�g�U�X�]�� �;a�CL��	�_�j��E�V�#x�|�G.�eS�2k�� p��<	���"�Y`�p)�z��>o����	Ƕ��I�A	��8i;a;_��)̜�(�*�s�/$Y�R~�C2�<�U�V����_�،�%�HJ��X��s��Gk2�yTcx��hs�4"��:kͲ�,���I��4L�l�gGuB=����ڦ�{��w|����S-G/�mS�odv}�4���D�x�:��+�Ts}�!叧P�}��'U �(��k�48��l���$��V��ejI�N��,����s�0�j����)�4-K�(s����2�99}�wT�ɱ)�|E&�ٳ6b�%h(Ss6a���ɢ�G�=bf6�;��J`=�Jc�����|7~~+~��p���7���gU=�7�n���ϷW
t��N��������=}\3�z����iL�-�g7&Y��6���������n��Q`w�a=����	W�'���E �����3X��(-�yTS��K2虙%o/ӡ0=�fk��P�6���s~�}92/�GCGqTF�=�(�l��I8�1{�0i�@ީ�f�����NC�a��N~�U����������tk�ULSVxse
L/6�<k�S`��!��M��<�$�v��l�vh�{(,��B�T�I�94�����U����3c�}��I���s�P���R��Zr���z8�[̗ ��]� �@֭����8וVfd�?�{c�H��`OVΡ)K�P˦�_��n3.X"�We����<�L(	B�C⟦J/O>5v��#�O�Cq�[s�]��,s��|1�C+���O�����4Mad�Y%~�x���w!����֗U%h�ŝ�6��|���;���uA)���!�o8j,Љ8�Z��0�Pm6=�F )�E:�t��U�����|yE��������/�ps���gϞ�_|a���K���y󓬬�yrI�v}V�n~m��ojF�&��l�e�)��G�Q��KL�´�ܐ1"����m��e�oeJ�� ����9���D�e6(|��U#&G[,��݃�7
�߰�2I��G��a�))��9`s�Nta	_
������~AY��H`�����_Mĩn���k�k�/�D�Y����I��ޥh6Es)��+)��`�u�]���-;$����q����6�&ŝNj�С���C�3�2�8Aua��a�ߛO ����0gu�l��Φ~��{� ^��a���-K�R���qgW�>:�{E������/��t�d# N�(�[��##�_>O4��D�P��9�߬>h���^|��V�H����n	/�y����>x�"\$EG��<%� �4��Cb���m��M`>�d����O;�Lٹff��������,Kiit�끘I���t|Pe�1���El�24��k����r����İG��~6� �Q3��_|f�]-(j�&���ɓ'���3{�♽���fh7�_�b������8r6uY?�ӫg4*D�z�ּ�>�7�}Mu��ol7쭬4	������k3�\�yᳮ�:�h��C�h�$l����BʱE���d��Fq,߾}˹���A��S[�(��TGn��HAE	U���C�2�!^��{���?6�����Ĝ�L%1ob4h�̳z#�kY<��!Op��Q�n(���)3$�4j�y�M�C�BR�@.3=lR��#6��A�j�V_��D~&Ec�68W�zn���&�C��z͸�X�1�`��/n�d��8=z�pS�Q|r�����	ds�"�[�d������˟�Ϛ�H�H����@�xF���v^�bY���<�#.B�F�ſM�tsU�k�-�lz���D��*�� ,Jj�\F�g�� ���l���I�a���ɃhLKi~=,���%�4^j���\<���^>{n��/�q1�!ѹv�����w�={�)��N���G{smk:�${���>��S{���Q�vY���v��fP�;z�_^�	�i�f���.�o����k.��AȷG����N"�, �]l����N��>��7�;ن��7)�lr<TMNR��Ѱ[�`2�U<<szH��=)�@Hj��V���'���N�5�$��s�������Om?s ��jYܣ%����d�nZ�q+.�{��G��~��;0Xah����l�ڐ�v]��K�O��{�3m�2s
=g��>ZY���Ʈ;�7f�1ss&O�B��!0d\ ��k�8���|b��nKǀx,w;��݃�-�⇏�XZ�pX�^J��-;l�� ��E����(�37,�ز,đ�a��:�7K��2��8���/r���������x����菶��y�42��:�D�v�i1���=
O���K��W_�W_�Ʈ�����ٛ7�i}=֓�zK�����~�?�[����<޿�Og�^���4._�o~�[��~gO��p��-Agd�׵<yQ����}c������J?9{l����������|�h���ǌ���k�C=6�5�ã��Z�)2}mZ����� Ph&q�����t��i;/ͩ܌���&�ʣ0ǝ�g\�pF��}��^*���������o�c�
j�5�ȗ��5T*��<��g�)��6����ȩ��(Ɠ?����!�#$�9�O� �y��ʕ6w<Z^4�6*Ա[�ȿhbQ��Mt?0���Kؚ0�n�����'����|@L�1���Y�w	9-i\���j�<�Z��py��҇�j;���F2��(�#�u�������."���M�s���ғ������M��=w��|�R<���i-#��#6�r��M�\B<��q,��v���jC�=(�8k��2�$΂J鉊C[��P��g_|������y�.Wޮ�8�����>����_֒t��o~2{_3��~��W��_����/mU��,�.�0E|y~Uˑ�����Lv8�Wg��뗟�W���~��S��r��ښ�&���k;�Y�y����7�d��sW�fwk��}kp�!�d���Nx���Q���0���;�=���˨����p=a���u�%ů�s;q�V���4���6f�l(H^E� ɘLRg���H�5��y@N�E߮��u�4NSi��f�����g��H�#i�a$i{'��,Փ${6~�\����DH\ŉ�1 S���t����Y��� ���_<66�V���i7o����8�m�;��4�*.���r\/Yc��Y�|D�������2���4�7qr�}�A6�n��A��5'�x)#��<�Y�>�,���}z��{W��^Wȯ���l���o쬥9�]��q�������D�osPO^�S�]B�ё�GRѼP��nR��E���,9���?:�S������20�D+�����Zo/jp�w����.jv^�Dկz|m��������?�3�m.���_ٯ?�ܞ�]���X��M����<Y���v���y���f�I���z7�r���[Nu�h$��n�Y�j�]�ff�E���,�GCb����Q���wZK���͝o�gl�܍�Ԣ)5�u��@��yR�|F�y�1�:��߂_��pݤ9AG�%D4�A�F�q&�6J�F6Qr°6[Y�OĭL�AR�F��K>g�m�@19p�FFwON9?}v���󏿜
�^Mi����SK�gJ�'Or#�^�@�-�P�Ohy f��&2��ެA`)Q�x�An�{����+��Sxk�
� ���A��S�)*Sr�ߎ�4�?^RC7��X���<m<hM���^�XgLL3N�m6��z��e?���/"�&e
��q^�Q&99�/Ή���es����Hp3Ԓ��,8d9��x�G--_>������Ok������}�����1=��G5��=���}bO�<�����%���}��}��3{V۩�~��^�\3��PS����vQSK�GWW���{_��qw#���\hXʴ�\��� ���{0d:�G.^�	Na|�`?��iSY6�q�>���b�n��t}�R�Φ�?)CS��`��}=S���<�|a9[_�)��������,��\�d �_C�`=Ff�?���j=�Qd�'��'t�k�9��s��r�h`�����']��@�0��8���9����6�o<~Q�4��F��e��\�}px2���4h٥Y>?2�ef[<���������]�~wٔ�����xh�=Т����k�)vUCӟ����1��J��<8���(�3��#�QJ
*K|���l��<��ڰj� ����a.�:����k+�VM�Ґeʳ��l���Yً����ӧvwoo��ۿ������y����K;����դ2������LnS�b�1�f��ym�}�ʾy���twM[%�`������?��\K��� �,澾<�[	 ������O���JǢS��F3"��Ș�d]s},�J���~�)����u�4���DmA�=Wfy�����u>�/:���<`4����Tfj��
Pr⹎�[ 4<����̝H����[�˓rn��I��N�P�� �4`h���ᚡI���$�Kj�{�%��\|���g���/�7��aL�0�(�f����66�nh��;��&^#^��v �O?�Q�}�U��4�����JX�9^�4���.���o<���L�����>�{?n�f2�L� ��I�ߐL�Я��ÐՅeT�����V^sߛ��1�s��i� ���;JS���|,A]�X"ao���a���`����颊�[�f�ٜ�5�P��F�-�Md��5}S3���������������~S���OH+�����Ћ�����������������Ԓ���l�v��ô�g��������7�?~ϛ�ef�W�<`����R
�5y�A`6�N�KE��`�'����p��"F7h��˕���Ѹ
��?t��1��2�õF��l`�%>_hV��Q�#�k�����q��UB���<W�e��4��IW�pƅg��::Ǭ$��I�p4\�G�<�i����-
�� 	)�Pe�����T�m8;;������?���	nkݵU�
/d,�N��eP����J$�i��[R<�[�����X��K|آc�}���9�E
�SPZN��.�Ω�&�@(�{�U��9W�?��@�i��J��,��~\�.��@[aȁ�{�U��;} ����Tn��_�����[�,�����՝���[����Y�Al�#E�rn��t�����9������ˏ0,v��(��D��6\����!�����]w�o��d��}����}����I�,�4`i�#,s������G;{�31`5l"$�̾f$�bty� �\fy���:�M����0���8��UD�4N5�����1O���ݜ�k�+�]ώ̥6'�uC�F���"c���4W�h]���ZyhO��47������Y�YkjpL�W�.�K�5GXr������u>�����u*� :�d�fn��>���*��$�dq��`���9��VP�	�)J3鵔?>�X1V��_��A����SPN�n�|��� ���r��� �-�W�w�Mid��f\5���gՁ�Z�.�\,���7�%��t�gw`��mN�����\�$��(�e��/� ���	��,�v6�zF������k�vz�����9���G�Wg��
_�"Ge|������z��2��i5Յ����t�����.����)K|`1谁�^p�l4�i��S�������G+7oT�ۮ�V�l�s�Zo�b���}F]��y��2�g�)�&es��Sc�(�zE���f[e����6��t�kD��BB�c�Q���@Yj�;eP�2��Nr�Qe�k��ꛣ&�͔�1T�6qC���F΍���	�e�3W��w��N��;��L�_�g�LJ�B���6g���aN&��?���R��a��=��#}9�!��E$_\t�L�u[�������{�e�\GD�>�(C{�iQ�-�c,�F�}��c򡾱[�܋ں�� ��E)�H�Ś����-�T�K�q� ׿����(�����7��1p9|��l�Rɳ_�Z�s`/��K�9��nr2��������J��41?�����'�r��r� !�c��$T̀�IL��a��|č��͊%+V��.��Ef��4+ |I�H�ԑ3?�Rx�.θ.>�q�F�^qU�ڌbm��j8LN��~,�/-�P�t�P��n)�w���e��]Θ�+C5����S��E�l߇?�jfX�pj��� r�p,���靻Řh52��٣��)$�_��q�`��k*�\�~�m�Q.��S�c[`��÷o׏�n���_dVY?xʬ���N��)|o!�'os�Ʌi�;���s��ٖ���A��(|�k�[Yۻ��/���̙�t~
��Ǵi4E J��ͳ?S 3/�G/�3�&�lP��2�8[�A�ۙ�f�����1biI��Ì�w�E�G�N���H���_��x��F�Q�ܮ�.�q�:����=���QW��\��ʧ�p���7����C?|��k���MN��9w}��(�L�VNǅ[�`��`PɲӃ���I��D$_��s������$4O����a�8: ?�L!����3-�N�ڊ�͔���4�*����&+�'9c�6uN?��[�ײ1�A7P�1��O3J��EuZǸ�g��pɋ�i�1ɘ��I!}r��ٗ�Ϗk��>*��[!��;�m��la��	���������/��~z�3e���UN���O�S���7P8�*EH3�,m�d�����`g��g?�k/�ݥ��ߴ�g`����h�8_h��=v��ٌ�Cy��q\�M�,vn��d:N���"��_�D��?���{�Ŧ���v^b���_��^Q�ĿSPm��V>��D]����,�u����|ˁ���ޞ=N���Ǵ���̩G��y�~g��[;����>q 2�	�$@����Q$�����t�I���D��}�g�zsi�n�T���<J2
=/;�@�GI�>����� ��� �+^r��Ѱ*E�7���8�Ǥv�j~>a���f����?���Z�^^ɢ��o�h��pԌ���2���6~���{�b�(��r��oY���AA��r����1�p�{�36�ɂ�x��9�e�J�����nW{���=��J�;l�^�g׻;q�^��l��4d�>����NR ��'���dK������ Sj���.���.J�e# �H~s������Rf,`�f"���28���3�����!z��>s<��n��c������IS ���1`d&�]�z�4�l���πA���9���`6.��b��:�>�-9����
�Xx�E�����u׽�#m����~����~���x����~���٧���]4����1!��=���k�����ڤ���;��OMF��4�x�{ =c������^6:�(z9�cq��y��%69B?��lps� �D�5���T|S�	���7��\xC�|m��,&��y�LN��k�}��m�I͈֡�Z�����_ՍDλcs,Ä́i`���,��y),,��ْ��:�ͮ����T�~�l�.y>�X�n������k��'�g�v^����̮>��^߼g��nwO�ȃ��oV�IU���2�&����9��M�&�\��Kf10�)�VfH���b��ϖ��i��V�xP�I�������9޲x�ۍ�C�}�P� Ω{�1�</(x�%�ھ��^
r��l��c-߯�B�!D� �8�L�$[i.��|k�e�/a��f��r�m+�Y\v�	��*�R]�w���;{���/���%ʳ�����?������7���6����x`h�k%���G6�o��x��v�\���]]��	�[���r�J`Q�hmQ��z'bzO�-<��S�%�}�#���⚜ʢ���)@~��$Bga��&�"���XB��{Q7����A��\���?�����b�]EнĽ�T�O.Lg����v�As���`�7��Q��=ۦQf�3�p��g�a�#/?�\�,�Fj��%k���<yCe;yrIі�Y�ל[LvF�pOx����!b�Y�zsN� �dn'A f�t}m?�yMũw�ޣX����G����Ο~|N�> tY�N�z�O�!�r�O�\i�,M�O���8�XH�wm.;��#�ˎ�J�����Y�������kE��rctF�(�9,����%�/���W �R��s��3��SDi���ֱ5tm���_�F��I��=�""'�6{��޵�Ke�t�������a���Q�J��4��X=��5H|����u�]~�؞����_|eO�s{{��
��/�ԯ���<����}��[{u����E-9?�7���=�zl���K۾c��T;�� 7�/>�\Z�zc�����]��`]��w�7���v{so��{���En_}��]�xj��VJ�8���+RO8�􈛳�zP�dw�p���t$���"�zR�,�7LHi����Y��E�v����zN7��yd�8����D�6ɘ:���2�o��q�Ê���<���ļQ��x8�[�ݾ��C�W����t�|&�@o9ē�Ș�q�$A;��ʇK�o̪�䘝V�6�u�lhʮ���?���nV���O��Cg�gu���y?�{c���ov{{���L�������nz5x���,��4;���I8���mx��_PZ�w��c����"�.�Z��`���e���D&�M�V��'����Zf��O,�r����bW��Nǽ�}��s�#���7���j��֓��i���:zz�.Zɞj%�
[AGԖ��_�Yo�s46� �Ew4�����~;��V��Er�Wp4��a�]o�SMY�@�xr�Ȯj �|�E���E�y�� @c����ξ}�������[�2�8\��{�9�4�w(ek0�������=�����5S;������~�֎�����?�xd_<{I�ilD�=���������/��Փ˺�jY���^_��>�_m���L�s���-a�96��������L[2��I�a^���#V�� ��S�:6�,p�'AXw��jgӝ�������V�JxrN�S����4V�sϐ`�YN'��d��Y�g�ڊ�O�X���v�u�}�E���8I�jS�T�o��X�1\�xF��M-YߝvT�`�zN`vzB�	� }�r�����=���T���S���˗/����_ܺ��-jl�ٛV�Z��l.	Fv�Ǜ�Xk&��21yf�?�Y���{�F�������b��X����^r�F��_����x:��;��90�[�j�<��s��T��Lh��E�*�g�sT�t,��)N�s�Y#����$m�7�(�u�����%v𜖥<:�a�7"+T��1hQÀ��n��W?�P��z��L���?����k��S���pk�T������^Y��	���ƣm��|��~=(���n���lun;�s�������k�co޼a����W�$F��'��||���=���g'�������kp��+'x{�!�I�u*����$�K^���R�K�h�>�������2=R���mcg5��5p�AfpG_:��g^x�S�ٮ��,�0�����2���	I��y�x�8X�D\ead ��HV�J�A�nZ����X+��t?9�����r����X��E4�2=׎:��v�%�76*���9�M� v5�?�?�H�A��=�C���?O��맪�����O��\��>z�25����IHv����r<C?ͅ�'"�Ĵв�vs�����L02�|>c�E'�g�p��/<f�x� �w�ܰf����o����<1k �)K���H���|<�h���1�%��<��ϋ ��f��!o1�׽�)�E�/���ْnyI�Y7t͋������,����Օ_wQ�~��S���5������������y���?�1{�{����=~�=���|�� �����rc�0���޾�W�Gw�2�z̯_�fy��I���j���n�"<���ܿ����`���ݼy� �Q��;��mfa�j�P7e�����W�.n��s��xTW4��=f}!��������3�&�s,A}9�ן��ک��W$���T�c����}9D#A��J�_5'8wxd��*ɧv�wV���,�hp�7�f�\]e�u�A&f�
�f�v��uq[�_�ogo����u����=";,YkA\TبN���c�a%�����'���a��ʇ��2SX
�'Os��4�� 6Ef��f�C��d���7ϋ@D���ED�yd)���\T�	2��n���Dg�<P�G�X��&e�1{y]ڽ��w�<HM<O'� 3{���Ε�Z�����]�Ls�V�`���ZV�G������kz-���Qn�W���;�zHmJ������?����g�߾��b���=U�޽#�����dgn��"�>�@�2���޽~c?���Y27p� �T�Ⳬ��Ȃ�bt�(��лag?�������~z���I 'K"Z����D ���pm<��ܕ�����O�Mn��ǹn����(��\w�Fֆ�M�D��X7�㬆>#6l�0��˲��y#�#�>�]4":k^E���B�j>�È0��D��� k��tPe!衂Y3�9!,]���٢W�2�|�-8tJ;g:���L�_�09M	$�f�ʪ���ΆU=�^N+�z���vKw|����p w��q���o>��
s���f�byӫS�J �gP�ϰ�b���,�Y��v�1��T�#�K��/�����,4��n`a����=v�8��,P�{��b7��,cX��=ǿyr
o��r�%�)5�*�K-	�s�?:d��r�Mn��x��\-]��Qv��v�
��[���=�$�$G�et*��$<b'�f��������}��'��/[k���������3w�����3�������g�r�ן�p������L���q_3�oT`3��{bm�Z��v>�`�4�T3�׻[�����ﾶۻ��o���Ԕ  ��IDAT{:�+��\�9�}�D�q�[����@��-���\��2(d;�(�Y����b��ۮ2��<|�mFi�o59�h�'�nd�������(�~gA5a� k�46���ҿ��&X�j�o#�ztd]%O��!�} @쿳�ט&�Yۢ(�,��S����0�3�q�Nj�P��fH�c'xxkL��=��9f`�8ֵ�0fql�����GaA�g6<�r�-1jY���+>n���J�J���|�̅��e���"x���u�A`BP��C;Nn�U��8���9��������Ǡ�+�~�MS G�h����8wrwS`&%e:����i�rtn�|D7�ߕA��]��&��ߛ"�:�'~F-!^��g�@��̥w�o6-e�b�8���pm��H<6C��y_m׵�<Ыm�Fê���zo�߳�8�_����X�3�V������n#g�����\da[��#ŠS&x]��o����5�]�s3�ٹp��I�p�����}pvٲ�Ǯ
-Ӂ'�e#�s�I���y�]g	)P���H2��0D���{^��o�U;\\�=xQ�3��w�i|&�?}��=�zj;�IMm=�I�Kil�}b�+�Fc�%Ν5|�/a�!S �Z-?O�N�=�e�e-���M�fc��1����{3�͚�2ϒ��f�(�$:����Ȧ^�� $��4��Q���G��Jk�X���`�������QAF�JSL��n�V�.~� dA�����w�M��^���&S/��BV�c�̒3�s?GnR'���< wy�&P����Hcz;�ó����]|���)�#�Co懚'z.]�T���0�I'�|ɉ�97�%f�&��3 &-�p����>Sx�[d[��ye!�A�����>�뼮�{ˠJ*K�mN����1�7߱�{�F�`F���48���"�fU�I�����r[k��c��Zj�����A"����Ԟ�6��1�f;���O���@��3�׾^��?�`�w��z@�
Ru]��>�δ�42qR[9rБ�׍aE� ��AWx�9�Gg��.�e�\:�QD� ��~q(��Nן��Ts���,�"��˫�Qn8�����ގ5#=��^�C'�ų�v������Q&t\��@�	��S�6���/C[���FrBp]S�A��'ev�oj��O]��L/���~�m�Ѹ?�J�qu��m�ĽH�-g��a�	U%,����A��p�����{��'�=yl���R3<5�4S�������y�9'Ǜ7��q��F���V��돿����JǱ�zqʭ����$�����"w�51���� b�)8	�p�	��L�ewӱ+�<���vXhJ�xH���|�'b�;I>p�D�e�EV��;u��8����bb����6��QB���L���u8N^DdWuA����h���8�nTyq��ûeG���]�6*;?�T�� d��S��V�;4�,'Y�#8��7�r�^`��[;�v_of|^t!�<v��k�����
�q�eu�֟oEK(=&�k�:�[�nj������p�������ѱ�1D�o-���ݶz,c�K����� R_c���^�r�Ck��
�4����{��X��YoD4;j���5 2�;�N7'/F�<zL����]�{��i�T��}]Gh�L��-g��v#�޸?����1�	�����#��>������� ������f/?���������Ξ��������i��suyi���̞��nj�����b�~��`�']o�ݑ���^�i^֬	�	�=�$����=��P��'��̱fpw7�\��x�O����b#;�\%96E�a��dtďww
Z�z��5ڝ����Ҟ������M=ȭn��y�:�q�0ȉԣc���}����
���d�H��;�aZ���.��'s'�ق�����9؝D�P�ݽ�)���v�D�a�4�S�aс�ɛ<ͣ��5�j��fB�Mɧ��4���`�1ℯ�{T3�#>%ŒW��d���QM�d�W!�P�P��u��0	'
V��)����V3����'B����;����ʐ��j���z�s����M������Kj�	���|���z�<�ֿ��L� �b͉�42��M��k�V��'�N��>�7�xe�G���Ȉo�F�Ǒ�ӷ�k+�f���k�/d9�	G���9��9��������n��ynq�������7���[��̍�����.p�zs!�u�.j��!hj��8�Ma�#I-�kP�k���{{�����3:�؀@ƭ˩�r`_���R���3�tN�Y��\1���S���/�t��6��IL��V�\Ё����F��6�Q�78b��������/_|��}������M���r�A�F����~� !y����6�z�϶@���3{��irg����rj�YG{��qM���;�^����PM#��X��:��J!����ʤ~��'Wv������M}���n���7��bm��)��SV�N��x��O�z�����}���l:��Φ�RPA�DXR+B#� �b�\���륹�����d�!���� U�5|�N��b�8ک��;ʱ	d�B�ku������O����FQqG��[9��q�5�0/P���Dϣ+!�T`ţ9�lm�;�̀J
8h��M�����0�=���G{\���9o�c-���K|��Xք�M50M��%-�W��\���j]Iy_o&�D�Φ�cBV�F����� �R3&�}$�3X3?�H�zNj��;���[;���q�fC ���\o.d<��7�Aϳ'O�~�a@� e�-�L�D[�driB;v�Q�r�/<5hC���f�Q�:,��R�&n�+(n�q���n���C��[�x�]��w�0�5���K���yR�[h���8�;�&�5�N�O�僲�ŗ����\Šk|��޼fS���+�z��~�o~W3�������d�~���:ȿ��z6u�U���Wpx����s>}�	��o~z�n4�/dl�j)zV�'����;����z�_���
�����Φ�k��9��3�GJ�a��S-���^��;���Fϩ�E�2��zC���v���f������Z_�Hͱ�j�0�^��QZW*gR
s���y����ҝ��ރ7Xfim���ܦrK����Ж��]=e}>�"�r}*Q#���Gv)��$o1�{x���� l����ko�e���X�ǒp�#ސE�]�w����U%o�y����2�Wu�j�!�/�(//`a�'rh�ۅm���<�������]M��~S��T?�����������u-%k �wi ���_<f���Dݽb�g๯�v�n��f:�]��T3��Pb��ԃy��{ਸ਼�Z��j)�nwGg�u}��~�D	���!�C�U���O�l����m�D^]�R<�����X���
O(��odŞ�;�޾~��n� �K�<��(��8Aj���{��-�BÎ���9��(1��^�L�Vg��K�Ս.���)C�~����$y���o�F���~-u��.9|�������ԑ}��`y}Y3���u\כ�# �ۚQc=b-��^m/�/~��2x��ġ7a\���O�ۛ��MV���O��Z&�#x8���w���H�(`���̾���w S�^7�=�4�Jt����c5p!�����9���P7�}]���o�����z�j�p���}���)6�g�9����<��"�t�T���{p;!��p�g^���f��KAm�)m�Ut@#�,���fzB�$X2�b�(9h�y͞�"���m���T���f$���Ҫx�#�d���{�M	��G7@T6�)>��E�c�����a��D���"x�L��_554�A�M2hQ[����^��컛����{�����גv]��N����^K��>�E�z}]4j@@�G

�F������7%)Z���Qʠ���rcRG ��P� ��c�-3��|`w�v�!�?�rWe1剮�<kЃ�a}�D	�w����qo�:��_]���[�e�u6�\�}9�\�NUWW�I��E��� �K� ��+O�[ �� ��&��@~�	؀� B� �H�\mI�%Z"�쮮:u����5��Ƙk�jKNS�:2�=���u��k�˜c��7�O���R����*��'(��ҵd;I�O4��wf��ԠNi�#�i5_�[dȍ���<gxqh�g�>����z:�wr������_�7Vm��i^V�_H����J�g9o��,�
6��x^�MK�����0�xZ-��R��b���F��*sO�N9Wo.�8��F���#�ã"�gr�i^�ӧO���c������/����F�~t���=v��#w49f���\��ժ!�#�\C��Px��+����:��ј.=�r+�7�l��b�C�z�ܓ#V��ZtN��
�(ͩ�3�N��HگtU&"�]���n�FȌO�[#%Qk���Y�<>[�ϒՀحĴ
v�x��q�O�w�) 5�����;j*d�$�t�Ho������ܓU��آ7�y�bŇ`8*$�����p��o,�|fm[���ܖ����,�9�#	;��v���_\�R��T������|����%��X�ky�	l�+ԣ�mʞ*�<!��Ut�%�9>`��K1��a�9&����<12SٱW��,�zkY�h�O�Ȱ��s(��xJh��Q������(m���*7��,��]c�y.��Ն��`�1����G�[�y�ڞ���[V3&փx���|N�s�V�������)C.Xf�u���m��ܭ1�����22׼��pc���*�P���vc8���ӭ 8m�)�:�%,2��ps���ວ�5!?}J�uw7uc��p��bLz)`�~�ï�P�h��`��h��)�#p;�q?z����O,�c�2���ZO���q����F�����Be#ψ@�d1�ݭlXhtG�d�Q�;8
6h�bJ$UHׯ:3���k��L�4�C�-�ׁ^��qv�����-61�7����{{��f������,�E�)K�F�I�È��֔��?j�-PjG�N	<�Ukg!�A������H���)Ȩ7��ǲ���q|q������+��C㖢���p;õŶ(�����8�[���f�Q�pS61���3		+�o�5	a�97,F�P�_�v���4R{bB>�P�Bb>�b��7�F�����t:��*�x�d�K���V)^<�SH�(�!0����p�آ�-Ž�ʀ�6�n�s�)X���&�ð���)Ƒx��+O���
h!+g��s���SڿQ��jӺ����Z�����jv{���j@��W�e�;V�K%�Hݖӌ��y�?�|��o��������D����*�C]�}�0j��w-��#����]\]1��8��5J�2@!d. !$��L6����^Q*s���˅�uBQ(��G�X��}�.��C�sΨ���Y��j��Ĝ�.���������rZ��^!#�e��ԩ���g��k��mdW�?�?y7����rן�b`�؏!c���uF��5��KR�Fx:�3�sg�Ʊy^���1��ab����A?鶉|��lVՌ� e�p40m�a;F�x�u��@ZS�R�K˰,@�C����,�^�zJu�(w�!,ù`� �C�-y*����
�]��!.X*�	��u}��y	E�b�ɤ�u�x $7�=�j��}l�ǙxMHR��&Ӥ�a���y���]Є8(�����x��)�<��;-�`2��)���
�k`��dw�@*Bp[���u��p�k�F�*#�� �)0p�E������2ŴZi�����*0��,�
�~ʊ�K�
�J���n�Ua0k�/��J�/����#2�r$��<,n,֖�yV�̴	0�"�}$%(+R@�SN�f`�A^����+�3�@�80V���;���kߧN����yt���{_����������Tn�6��&����8�z\IΞx�Ԕ��E�=�~x�ȋ��p�����ڑ�G�8���d��\Z R�(ęqõPu>���+uF�չ���xeyf�d䂷]ߜ �T�a�AHD(Zkh���`Ɨ��"C�&ޅ	�!���WB��,*��1*\�ڣấ;��q�^c7��yr��#F47ԯ��Gī��c��Ҝ�d��*\����oMގR}-�Q�
�X�?5�Ͷ��@��(�BM\�&�?�5��CZ�7AoL>r,ǜ#TAn
�a�]�2���"�X����]]]�Ջ��D�1��K8�b�p��j��HK�b�V0)�l*�Dg���B�%�D�V*!�����F�B~��=�22�Eʊdkx>��:	O��r�-��P�W.2m�Au.F��6�r߱9 ?vtr�a��ً�8��z���m䂄o�\��(@3���(f������):8<C��)�%rg���FTy8��S)�Gۈ�Na�x��gh�P����l2 4���4i���4�p������T��b�'jw����i�QC���g/�k6��BBTGxϓ�Cw2<p_;��r� ���̠k!s���2(T�%e��Us���'t-�=��a��D�<Jv"H� d��(2�N=(����z�U��N�����W*7�E������H9J�l*-D���Zl��"}G97y$�����P�E�(��io���צ묈@��q��yCE <@	���;=y잝>!��#�=\�ܹWw�n-�/}N��ñ���S�lr��R�n�V�Vy���������2�z�����w���BT�|�lr�*]�����+�����X�0��xS�g�z�NF��"�e� `��b0 �:�\^�t��T]H�W��`�V͟ X�I�.Q�Oܩ\�q6�=D~gLsEZ����9}�085�0`�@N���F��H��>΅���Z	������=z������ƽ�z���$�pDm�¦Y*�"ճ���%Q��9�Q�����b�@|��
P8�����Qb��Sk	k�kbQ6=6�C��2�^[��&��K�y��"���ޕ�sE�/1~�4V��@i�Kc_i��\k�G3��Ad��h�5�n��<�h@G z���29>&�v��.^�܁�Dm)!��+ِ�S�L>|8����n3�+VN<�,l���f�ٝ�u`s>�+*�e��`TF5�_��YC nF���/�EV��!O����F����TDdi�y���jm�^���(&�W�Ż1n�B�P�d���7�������5XH��5�iQ���"��P�e�?����=s_}��v>8v��k7XW�j='6r��C�dt�"���G���<��cj6A)�����4&��f�~Փɡ;#�����nO����0}&^�d>!Ɍ^���'��~�=�s���m$�C��g��&�O>�������kF�I%����X���!�Ä^CN%{�=�G.��,�	���-�0H��t1�-��~G�ia�L���4
���w��8.�$P�B�&*N�P#y9�	P�����l=R!P?cuh��<S wD.LW�xy�����Wǉ,flH#,T��G5q���6��!�ɢ�*��i]dakLo�]d��^� �k���#Qy9�t���t�AG��3�(���"�p%#Lu�Cϔ���N�8P�+�c<۱l��a�c BɗCn*CTy�K���O��[3�v_#�&���~$�W��~]��345(�q�����:��[�d�����J0��SꢠQ�^�9b�&��U�H�hϵFw�oST�CGt�6�5ۑ���Qu��n8�	n�zA
�l�>������ФǱ����G�'?J�Q �S��N/2��ad�D�,(�>��K���X=�N�$���`�N�w �>�w��� �P\n@FĜb���!7�Q�0;�_�Z����4�C���{t<t��_z�C7�V�$�s���ʹ�����q`;�F�+�}M��\�(������.�kư���n��?���@{��A��Za	eӳ���
�V� ��*^L9[����ъ�^�z@)&8�<�!)�3z�!_C�-h�L:,��r�R�������aZ���7zD�>wZ�o���p�	�]%�[�v ���sy/���������r=w�{�ђU��H���HQ�B�*XOn41畁KN�s$��BD_'s=��$*}�l4��%*����gggntp��� ��$T��&��r��䆛��C����IP����ͽ\�rN\�)�bE	T��VF��øW𴀇{��=^6_��E���`��1� ��zْ�y�L���x��!����1G�<�M����̓��j���)�:Q��A��Y�v�k���c�=�9b�*QfcJ%aM����dS^O��P��d��ݏ?p.�Ç�wi�v��,�g�2�۶$�x!���"#WȂ�����}���10����VƂ@��`x�GC���̽��t���]��]y;���
�{:cs�Px���4�Gm���zEQ�W/_���̝H����S���_w>/��? �L@�|���B�[`$F�ā��h`?M�P��t�x>X�`�H��#0Y�j,�W=y�U�U����-�d������ڡ��x���jY�G*�N&$�!�	5�d�j[�a�a?�4�a�^�e2�3Y''G���p���J�,�HN����Yq�~F����;:;uA��������j�]<`��V�(��I�t�~]���C�da���'��i����Ʃ�z��:<<p�����ch��-��#7�0^��,rL�Ūg� �#(�::؂��f��1�nke�%[J�e-:�6�#��rw|z➼�T�Ł �3D�ڐ^��������:���fc�
jm`խmӖ�娆�x�%��z����t�U�^Ο�|��p���"�lgSzq�����Zx��>�fU��E���IC���C*�zT�n��!F����c� z��>�\�(p���jg�(<0��� t=�^�#ò&��*�.$�7������Vϟ'���l}Kn=Z�O1^^Aƅ�5��VS+&腰��	�	�ؓ��}��3�	E�&���	M*'�������yK)��x�7�\ hFN
���VN4/S�7�����K�e�pW�{z$0�>r>}�=���S���%<�2���D������^^Y��(2t�(�Ra`FrK+�� ����gt�u�B+�|�X�ͳ����Um�F����-��KO&�蝆
|Hr\�]�zG�X+-�9�g;1�i��Q�H&�x8Rqcm��}�@����D�#$��V���bHL���-�ۓ'O��~�Ξ��5e���ҽ���T �ٮ�@H�/����'	����&�I�u(=v��ɁQW�0���`������X	��4�x�f�u��V�: �dգ�,�v���IOt��a,�N�ʦ3��O�����؝����=)�dC�9ӭek6[��|��d�*c��ԑ�=�_��g����|���Pƒ����|��)L��l��x�����SLݪg�9�6CO;dک����&&ƻ����+dޏ�AE��] �[����ab�2��Lq���Y��."�a7��R�R����o�����t_ʰqݸ�a���[wc��O�P7��_�P��C��b��F��ЍT��D&�������ռ7>uc�ײ��J��i�Xn�!a��cW�u/�����?u׋)�*���3:�HP�P+��z�^JH��_|���q/��u�@<��=��}���{�O��2�VwS�`��n9�c==>3l\'�ͽ��d@9h���W≡H1[��0������}�+_��3N5�.�!����F�Ў�g����ݠp^^9�0�)rO�gs�0Ia�p�3�R��AC41Q�K �2R��MDE�pT������B&3�һ�{zl��'O�#�珤1&ށ�g�	��QX�%�<���C�vNO�zc��ěш!u�,���V>(�ȎN��o:�� �Jwz�4Jˍ;9��(E&̏���0S��
��ш�/hY���v�3,TEk# ��:e|ּ����-p��D[�x���Z�=��L���L��^��7�fSI``ۈ3D�}c�߱\?�r�iwx�PM��^!)/�֭��F(�������)ӵ<&�iY�:�7��j��,� z"�Y[�����8	<9-�;k�^h���B�N�4�j(�4}��ËN�yi8�ƺ��h��~R�Up���G�`ݍe�M��J��49z��7�[���c��ol��F2t@2C�\%|9�)U��^&ӱH=̄!���켲szx6	�}��9�h�Ah(�_��I���({#�9=>q�b�@?��t��ҽ��g���e�==gy�p0v���T��Lރ	}�������wk�Hj�'b Eb`d�Ioz#�Bd�,[�bY��G�Ne8�n�
�,ؼM"����k� A�mU�ؼ12�`p�'M,'����O� ��ʇ�<z
)!��UٴJֹ�W�xO�P�>:wK	1c�U5+�^���g��Ξu%&�ݖ�`(����������RBC���h	hw`�_���5���x1Ђ�Z֖��IR[(pS����S��.�B�3��oYŋ9���@�A��\H8<�T� �F���DKU�ЌǠfz�g�� ����'�z9�]�g<�s�'5C�������I8B�9�Yl�b��F>��Ǟ�C0t�_�v���
C�����1?�~�e:(�����1�՘V ��6���9}�^	�Y��� C�ԅ|Ϛd�����s�a+Αs�{�JG�����1s�����&��j/mzy~���~6�6X%^�yI~�:܇7�c��o���K���Y��)�c�jV����P�i��0��
�C'���QA�(!T!aM������%LIĽ��Q���|����ӫdRV1��������-�7��Zj�6�9�>��Г�;�\�Z��"�\0@e��R^��G�5�Tڴ\)�sϯk=�rM���\W�RИ�W\'���k5<�RC��8puX3���^�
���_7�Ұ����F��������he��p�Ԝ6<�Z�r6��c���t�$�?���wqqAl"&*{nb�J�k"��,�t�p��������������1��y ^�Ce��%�Z��6�mIC�`P�8U�+z����[c?�7h�SF��#0Ի^���TW��Aߪ�:Dr�MK�t"�e�7��j.�؎o'#������KH!�Z��Za9r\��ԬX�{�?٨HוAY��b�L�o��_.$
��3��o����eB�����o$D=�,�d�`j0#�L#�B�sL$�J��&}�<��Ǐ��i̦��]\�t\��ߛ�e_p�����D`̸�[q^=��:9C�FL�ຣG�1*��X���Z\����k��sM�"M��o߸U�\�ktbA��g8���#j�_��7�E��)�ෟ�BZ���t�̠M�<���YMT*~��^kw��F1т��+��"o�S�[`uBg4�ѳ�`�@s�xޘdg��gl���/nH���M�S���
T G�d���f=%�[����F��"�I��l{�Z�+�m�v[,qKpsGHL���F7L\z��!�WI|��J�r��<P�(h�BC8	0�Ĕ��կ.��]H��$>
�=�𘔘�vf���h���*�8'x� ���8q�j��_�R'a-�-�>�Vv�IdP57}$�yV4�c3Z.�U��P�c1i�q�tmU��a�>x�)'��V.?���g��<[|OS�ݰ�p(�<Z�ؾ���A���gb�h�Z����h)���T?�`�UZ��>ov?�ڃ�1���Y�{����B-����H�t\�\.���C��\��lg����;��3E�� ̽k��к��3���@�y�r�/�GT˗�kD������)vz(Y��c`���`"ψ�!��9D6��+����܆�*����=3;� ���j�wi���Hۖ"p��r��#�M�pc�`���ؼK7�H�v�����t����]O��	�Uf<�G�5�3X2y�0n(@ �7z>Ф.�1#ʹ�1�B����Q�ǁ���$��Ujs�L/�oϜ
����@��U�H'TCd;�T}�@��&dd���pF���&4d��)�D���;'�s����e0�^	
p�N��݉glx8&����H/�����a�.&|[GA���H�V�,��5,�A>d���o��hi�Z�P���m`!c�Ad�E�yT���h6=w�WW�����uƬѼA���.h�=�x�����BK�S@�o7����E�8�$4��Pq�F{��G���ح���1|E�61k���E<dc�s�2�\k���{*�zT;��;���qw]|���M7+'A�9�����x����[�ŝ��W4�h�|
��[w��%I���N�bz�b��wl[C��g�Z�F��1Mر���OgJ`�D ��Q;����Z����(�jR�N�'5��&���Bǂ�YL��w�~�b�6$�1g�v�%m�-�x�p��D��Sc�x�E�&ǃ�F����sQtl�r�f�A���cX"�7���0Y��~=;MS�����שo)l��&�t�F�,wc��ap|K,�J� �5C�V>�IRȤjY���g!`�0��Q�S�ēE�c���}���	��*+�פq�%����7O��5���*O���k&������k����Jt}۰�O����s1���oi^O�e��Ϟ-�#
�y�.��}L��	��I5$�B�&��7��kL�!Pm�U�ơ�Jwh%�g�p#���<=>$������r��bn�P�Ԙu��ځl�����$��c��y��#���xS�jƫs�h�k��a���=�g���b(=�_d��9����M9e~��(3f4_~$�'<�/��uIOo��s��P῿v�@�j$4���X��f�p��#X���Z�k���q�Z���r�.>��ymlP�De�P����Ѕ���&�1�=��긮���45+H�`}Aov"��D�!�@׳�ҫ�#��\<X�%:� �>��y_9�S[��vAm�߶q� �L�������C·~��6�A\4j;ƍkfܺ�A�T	ʜ�+e��Bw	12��V�V0ꑄ8L�w�����^�c$�w���S}r^�\�ƾi�G����4� F�)���J:���H<		�d� �O�%	���dr��ǿ����  *pf�5�kQ l�k1�k0�&S=�tp�9q�b̳�t5�U'*!���!*����b�n���ߐm[��ᭊ�
%23��� ����g�����`0bEl�0E�*?��O$\(ငs�p�5�!'ј��#|A&2x��뇧X�%VM#<�ƱSwP�>
l�(�L�'��c�X�)�g��������� ���6�N��C��C�����}T�f��� ��Y$V��:�{�ț���k��>�s~~N�m(�4�\�]�����2Wb����;��У�R�s���E)sJ"��B;p�r�n�nXd!~<۸��!���[+Q@*�>'��#u��S7}%^��k~��j��ǳ��+���'�	�w%�=)���à�0dd(����c<��
l�s����k�����p���lHz��q�����
(���#.�o��wҡ�lwۭ�o��E��L�vp;qrj�h�m@Ψ�Y��W^5��/aE*�yx�?~�)���M�&�D8?;g%	�*YW���U�~�5�%&B7p��r������=W
ptX(��$`�!d���~�'���T`A�xvp���r�2�S�e?l�|g��(H!aG��@�����p�?ǰ٧��wʎ��o����&d��)��	�5f ��3�a}�4,� �DER|��ڈYGxQ̍��Qiw	rF'�>;잞=f���z.�>��*�����+�5�1ȁ6A�z��ɺ:�'�f 
l����FJ�`�|ϗ�1�w�1�	C������b@N��ɱ�����\���D�{N�2�,9 ��3U����V��.Q�5o��NN��'�2���ўEqRC���y<РGg'�=�<{�g�|6��34E������"�A�V̈�9����c߮�+��;(��w(�b��pmLCFaceN�AF!��d+C���@��?b1���o�W�D:�t@R�)��;��Ӊ�������䇄�]c,!	[ɕ����Ȳ�������G(١��C=�"��l^�'g�@� ��>��[>�� ��}R�޾qk�M�$Q�n�<u��gV��$*��{�M%��D263ËB�0m��;**��N%��Z�ܫՔ�PLPٙ���b�5wc/�ƭQ:�����Y�9�����Ų�"��ۂw�閌�_���Q��IV\P!����X>��԰��!;R6��C�x��P-�G!s�a��8<&EJF��y��V����A�]�� 9�@�}Y0K٩���h"�!�L\W���6��-�h��F�i$�<��Ew��ȽE�ę��X�r~'G����M�ʦm���v=���6%�NŘƊz�C�CFy?�i�5+���84x|A=Mxe��Oݓ�S*�#�I���D��:o�W�=w���{yy���P����9��zLSxN��gܠ)�Z����Q��<�LÚ�U��@վ�<%�)�����7���4V��>}���o�?��'�5�;�6pm,X�;i����팻.��f6��5�b�
����k���k��4ݶ�re�T7��(�`8�q�}�yP�n�p@H�v2ə#˜IKғvD�V�kO2R5=.�oC}� 2�-[�$�#TO���b4�	��o]�!OqDʧT)�M�B����,�	+�啦�I�Ǫ��7WaA)��RLu���)�"���3��R1��&�,l�������J;�p�a2��m��ޛ߶k$���"���p��>5%�d�iddP߿�Pm*x�2hU ���F�;�X=��YΗ	��V�h��� \@� 	�à��<�MV�G�.�v�	�c�3*�Bi���xϊ�Ōy��f��!?$;4r[��&��uL�G�C+�n��
Ԑ�
Q��00-c��:5:��%ｧW�N�Ǡ��,�
�䪹Pm�,$�F|TA1.��:~�/�R����
׳�V�R;4'��X�S�/z�VG/^����NO����Z�~A�VV��X �M�>x�=:�q�������g�tD����a�u�&t�SO�a^�e�� 5����d C����RO�К�����lϋ}�!�b�k��^���ZY�Y�h����94�;��[�c�|U�Y�Pl� h�"�������$nEnӫk�o�uԳm5����k3�$��]��3m�Y���M� +M�J_�V�P%G
|F(���z�X~���q�φ�_���3��#q��s�$O�TV�r�S���ᤐ+��8 �݊ Uc�8�	$��kǕ���(�?�FN
7�2��m3Y�����cVm:w�9T��]Tqǣ��*� >2O�һ�`��U9: Vrp��kG9A�]���F�\9���dҶ�ވg�m���O�]A��'�w�Oܑ��:j@�0�)J#�r�>�y�SM���^j�>�
[��5:��S��,bfhfƽs����*`	զb��ޱ,x�n�Yb��hyE�%w�d�������'�<86L�R��,dTIs��)LdS*&����"I��R�cP?A���^��mо��@J�3#s� O�g��bˆÄF2���Z�G����Y���0H8K̟x�E�zom^
J�~D�ƾ"JRR�0���Gޤ�Mo)ϧ���3�������K��A+�RbOg}�lM�(�<���#7�
�E�p߀�k��
�n0��f.�r�+/L�b���R�P��}1$TEi4S1n���KdN�BK2M�c�����g���l7K�2��J-�ҕ��-��!!	��u��:��g��Vs��x��!���C����A�6H�I�"r� 2�5�٪�&�U��u�&^��������*jF��xR� 7����H��u�Z�
!�m�=j�� �t���=�^J��1��a @5s)u�b��B#�2 1ޏi��*]%�4њ���0�)�4�ct�m�c�'�mtl�c۶m۶m�v:��������Y�V��W��n}rX�=u�Z$�΁��-�s=c7��"}(D���'�Ή����M�z�!�y������'[i殻{i���{B0^l׈r�&�F�6��\S�Nh�T)j�F�`�(-���ʉ��� |w�Y�X6�r������c:y�uI$��1mF����y'R�e*��l��A���T��Jf!���
�>vw%Փ�� �Jw��gbFX��Kt�.i�0���2H`���2N>�z��dWq� �D�U�-�*�A͕���ç�`�8�Kڟh����6x#(�e��ty��_ڰݞwR	��}!f)�C$ĳP󗵾_V��x��PrZ�7Zp�б9������n��M|����u6�`�`�!�����ɇ/獢��WE�����<���m���Po���7�cuj���Le`�D������-���dV�d�'���tzΑiZG��`���>[�7�Io��5��c^��/���B�f,Z4,���o,�.,�C�7��`�n��aI�g���1є�jG�d��O��C��5P�"kJ�1����9��@�Z�����@��w��h����C��#��6?B��p�
�5C��}\Ļi ��:�# ���h-z҅'�Sn����28�;���	�k��~h���� �N�<�KY�r��}V;-EO�N@�؈BtsͲx��r���M��2�;g=>b4�FL|�z�_���5��� �^���x#��3b�#4|01#��;7w����m*W߉���U�Zb:�P�NJ���X���O�^Pi{RB�W^`")����3�|�vQ��y�/Hj���K��+��-�E��)x074�
�;�mbX�G���1�x�%	��4����r/�}:�����V<�/�ll�a��R*�Qr��WH�i���E�(&�0�������7�ӄ�Q�u�v�q8;��X������2���Y�㑣z�||��5��u\�#'���|^����<Q\���N+��F�l�m\�{���X��)h�(񖏏M���Fn�����Se�&���(����M��I=d�Dxy�	�@޿]5w��ڐi�U<';	`�<G*@m}<��)1��\��gD���GǛ�vr'7ڭ��ʤ�����G��v+m�zī=x�1u:����,I�#L��b2�C�Ea��EgӑuU�y��*'�H5�aL�3�6�u�;��{^����"o�Rw2u�����H��.ĸ�ѹ���B:���C��S���X�0� S���h��o�� ��nd�� �&4��"�spB��W<m �W���?���"�������s�<H:�\c0������)x.����a�[�jv�J7<�e������b�vť�E�t��U궥��u-=-j����~O�]L| @��鷤!�
��XYp�X�����"{燴-� �!����Z�"��IAYW.�O�n������]���}���4���M�>�t�~͑$#���bg�$�F������!V���~d�s$��3�.��8h�;X,n�'��w!炕O%��ZHK��G��&�4¼~f��`�}?խ�c��*_����V��y6���-S�Nť_��e�]%�M_ԃ�4�Y�*e��|�Y���g��{���0q�Kˍ����3O�~{0sz��%�������M�5x2f����s���Ef ���b�l5l��������k$��tg�&1(_�J�?F�t����'Ý��V�/w��e�>�h�_����PD7�A27}X(�����jhPU���!�O9P�Z��*sD�r\[��NfR��2O��G-�}���aw/��I�A�Bp��
'���)�xMѯ��������z��&Y��$�nN�ļ|4@�G'��CAB���o"�Z�
�nL���}��E^�$�v�|�l���6�����ÜTǜ�ţ��!״�]=�>W��I�m������j88BG���o�x��[�L�-6�Z8�1���tb=R2x��/Sn/D�7\�|ŭ;c�A
�9\9�*��<���$'`�*��$��E��m�M@|o�lݽ/������9$y#9�ڪ���#x�rZ��:Uu� ��]�۝������D/�����8����L�qF=m@�A���2)ј��Du/n���L�zq�k���&)�l�H�#���b�t���ֳ��"�e��j���u�fe9��5�-v���o����f�b�1��X�j�>�Te��1}Ϫ)�T��K��A�&�]ļRD�SE�����O�l�\Έ|�Ouoq�`@�gޯ�_I�#l�4Z�W�%�O4P�Y�����OOM��nD�D''&'���/s�J����eq�Le�ڝe(�T�v*U{D&hm�=*��Br���85�1��B۲����@�n�����x%Uz�q��G�Ke=x�*��LYLV|)���W%���Fl^14�1Z+� G�� �u���H"���a��Z��(}c�o����#�I�S7ȓ�(��q�ܹ��Fz�x��>�P;d�gm��t�M5�q�@Ցv�ܓ+�!�]HF����v��P#|�]&��D$Vw0iUT��P��6���Є�@��)<0Q|BZ���y��*��PQ�"�9���c�������em������%��'!Cأ-c�8B�`L{'�v��"'�1+�/����`�k�(1)z !9��F�q�R��l�;RKA�7J�6оjc[#a>>^�h��b���j$���~���<}�Eu���+��1�TRA�y��V��r,&�g2-U��],N���j��K���g:�q�;��Ȫ�����Lx6"�G�T��ԛ���%� ������Jwh"leeR~�sg��tm�5h�Y�k��#a��_|��H(�P�ʏ�j�@kXܹ���
s('��~@A�K����V��V����^�����XIH����IR^8�{���k(��a����@ͺ8$t����q)�{�l�b'������yԐq�&�G��.�A�F7�!��C���,�l�":��BR�5�Qx�|q��`�1�0����+�jA	1�#O�s���G�����;����#�d:gX���J� F�}���1)�眊�?n��*����UxM#�ۢ���ፑ ����e�%@�//Jn.���]���I�?�����MW�@!`?��%qQ�����]|:[����}�}�a�3�v������m����XW �OAr19B��#o��a��9�u�G�:;J�j�ي�����!V�S�Cc�*��W�)�X�zf���0�Ub��t�uۮ�.#�̐|��Ky�+�˨gI�'Bw����&d���+�wQ��u� R.5~�6_9��Mz�{$�&�#;�Uj������J�~y�@��� ox�Q"���ۼ��@;� ,xL/#�E<Y��e�Ĉ��o�Ӷb	�R_�0��i�Г�X�%dP��k���Z��O��c�6H���׈���г�'4E��Rd&�u�8��!-���)��D��`��`ZTq>8�d��B Iy��$�Ǆ�U#���wO��!�MI��\rE<��c�� b���� ��Ȍ`?zF"��5��%ܜ��!b�N�#`_zq�DF�Y��b����0�雋��y{tO�z��lȈ�a��|��-���t�k��={�y�}�俍�6Uc�4�\^�e0K1[s��L���#
��<�	[�!S0B�2S���CZAa����'�>��m����I��I�y�'Y�E��v��v��o5P>�(6S+��\��qYZh�5�U�{�2;�ŹI���,[�*#�Y^Q�&,I���E����"���;~��������h��-��F?4Z�z57��4*�`�k�0'�	���=+^�'Ƙ(�.#�ã�#��
=��t�݁c����,�ϑ<C��K��7?�
�r�PnҼ��wZ�Q ��iӬ��w������7��pbe͸��V���T%&�0F�����8WZ�8��Z���'#b����Bq��}�2WEp��݀�{�B�Q�x%_�p��P;�In6l)���Ҙ�i~HwS"Qm�_�ge�x�q�O0�5�T�M�@�3e89�8e�����?�Y5V�����0�'���	�����!;���:������@�����*��#n��R���>`
2x��	��E�S_��l�"̚c�' �oW<I��C� ɀ��t}PH�X,α��Q�Q���lMa"�!�l9>O`�p��F����v���D|# �������K1�z��tܽ^e� j$�Mv$%Q�7"�Z���P���+ .>�R�o�V�4މ~A3Z�x����vJ+D�Լ�����
�!���AQ&�]�`^���@�7���z�a�O}#��-4��>�k6v!(���Ч�R;y`�-Lt��m�_P���䰗�?L�@��U��v���X��)d�p�\���ӄJΉ4{n���J%��U��t77+,oPɶ>WrG2.J���l��$[;��W���U���=q�R��_��Aoȩ)�r��~��{�l�{�Xc�c�IS���!�� �5ґ�~bz�q� �����cDƁ�,`��{�
�@����U�0]u>Z���N��B?���,|Y���W�|[��k4> ���̘4�/��G\�<`Z�9P(�<��V����E����ϓ���U��&# ���ZLAw/D��Eض�G�B˧F,�|C����"��;šR�i��e*�(�"G�=����o��
I2�k ݎ'Y���aLm�����.@/묩�5�V��SXh:�����&�&Zê�*�X�����b�(X�W�$e;�����U�\��dEI$(ߌ�����q*J�R�I���/�Z���۠�Rk����mЩ��d�T��۔NC!,8fQ��/0��kJBh��"����z���fi���'�[,�^�?-ީG{�*��<ҷq��G�����2T�9¨�X���4�*��T9��x֡�fY3x���� 5����e�Xɫ��8������v�U�Br��PD�~	>κ�k�����/yjv\�����9����z��b����r�|�������6v��GڌFY��hdT*?�*�(�XX���+�;��;��&��Br%���l�l��JO����� F����X��R§�A»�����8������x�Lw����;�4X�Ҟ9��\B�w%n?�AE-T�^G�?���h;�nA
��_�.��F��,IrfY��؅e:l������������T ����mĸ�pxnu���ߺh�Z���Ǫ��ǫ�v�xs��UËM����3��7%�
��
�P�����!�6ȔR�c���%�.å��^�i��
�T��0A��m%�*d�|f�0�^��D�7�d&{Je�Rv�W��� �X���]ү��+��kΉ>X���ս�?�/K����'��Y#�5�B֐���ks�l����}�s��gw��9�v�e�)H�f!��Y�T�D�E�Pa2�ƫf�뱜�t���;}���Z$�q����3}�iw�(C�2]��<+?�'�;���h�cT0���l��A��IK���/���D�]�pFI�y7��i��ܸ��H;��D�(!��)���ё�!�����:�Ĥ��EY,�M
n]N��q8#�3_*��%2zPH��.�lb�N^0P���@�Q"�T]�N3��+j�G�����t�p��&����e�&�ٞ.�)�wZΌ��M�LC�h��a�7��>W����h�C;�C6B\+���MpG�.5�v���SЋ���n��V�n�GE�.�rl"Wb�|�����&?9צ�.0g	4�&�q��������i|�!�dY�b��4;�	�n�x�(Ŧw�����b��f^�yy��}�d����6�,�RJ�O����R��|%9y⥵ZOs.�D�X��`POH�W.�x
I��N6�6�+\f�	6ot�jY�����!��Ӹ��tX@;��W;K�¥�Y{��Y9h�k�[�u��j۴��a[VW�m���n�x��D'q7�)_���ǋ�]��bp|���=ޑ�^�hve��#���Bh�O���W	�1�}��|0��"�/�9}L���z�.�E��N���4"N2ľ���QT�<t��{���l*��K@��1�-(���i2���o��x��<;���Pߑ�a�'�)ޤ�t����T��Ԙ��_�=���a�QL���8����f�BB(�ݕ�P�Z�v���#�	q��{��-B	�5Wg��ĳX��c�beR�h	�]�\�t˩�����5!%�7�V*4t��&�� ��&�p���<ZwRo_�r{�]aM:9�i�0�j+��q�k '�-3B�/{��5g��(U�y	�؂�?�bA�zߛP0��6�QE����[��g*'d�D1�~6iN�W�@Kej�J��,��H���P0G-���,����U������6Ht |�AnaX�HTf���@��?WOZ� ���]߷͟G��[18�W��G>$P���|J������*nt`�opv�W�6�e�9U��SJ�W	�xĬ�Vs�Z���ri��e4��զ�9[
��b)会�����+Җ�ӿT"f�~�fKl�͌A�g�R	��J��H�d��՛Lr��n�=��(�G�8����+7���f��a��A�`Yk�-� _��R������~蠴��1���0�11�2�]c-�q�o�ȫ��g\2��j]�����d��7q�$Г~���]_� ��Hs���/a��̾nu�2H���:�[z�bU�rne��
6��`��I���/bU3�R�������;�#���l�i�G�&���b�
o�i�i�� HQ9O���b���$Y��{9�td|� BH]�u��V*��J�4F]匧zE�%5崛=,Ⱦ�a�$�����G�*[n���f�~L9��&����m���F�H���v�}�xr��AΤr�_�`���b�����]���g��&7�k|��b���2�j>�cpFj���.F�N���7�*�dzSݮ3��WX�	^� ����j|�h��$�W���l^���|v��;�[���(.�[�I@��S&U�D�.�ai�C��3�CY����y�%� �y��eM��E��Uu�~�;ب9LWe���M�3�; �S���mY�������s|��]m�RM�<]DZH-R"}�rP�l1�͉�` ��
��{�ciE���P�����wq�η����~�F�G�$qTԾ��[�2˳Ɛԩ19���=�++-��̳Ty�lo���
�!S榵-��I�F�<� [���%f��"R;�rXQS��M��$���^4�$:�>pE`&�%�����N��4�l�.-�[&�7Zf���'�b�%���D]�X��s�aPٳ�����b�@XaTk�>Є��l�� 1&�bZ]��7Vܨ(�7;b4O}?}U��]WH.M�>���`̿8)��!x�� #�9���i�i87��o�\R��&��
�p9o�����[{�����';������VM�g�ȕ�@ֻ��C�1 �T,5�����rϐ�F�(�u�V8aN�T=����d�������H�L.[�j���k������3W�~�7ic���} Y���D��"�@��/��j�6���|��$qma�
3�YIMB�
�F��ԨX��d�7Qq-mt������5��b��r

�Ds�oI�]���-f���Ӄ;tJ�E9D�����\����,ǷV��1�Z�5��ꡂBNe�ㅈ�UH"��;f5���<���~�=�ƌ<��^6m���Ϛ�v�4iHOJ�|���%x����:T�^m�j��M�8�Wޖ0��e�Wh�UP俰ίb�ێ���.x�P��W�jA��x #*�3���C�+��+�(�^�]�~�A?Wo�A���NU�t�sy,��u1f|��䷾�Q���!b%̶Cp@1�Ə�N���4��p�!�̽��u�#�S;1ʭ���J�F�Y�����[������5Gф��lج��K[��6��J�����b���G-�m[^nt �7�����w�g�q߷��?Oޞi��Si��qe�Hv��椕F�;�kaԄf*i�k�wՀ�A=N��f#�40�E쑊��`�¦�La����F.���8���(��NPT�	�"P����X��i�P�>V�x���a�HH�y���M��;*�-�&��>�?@̭(h�ᗰTx^���.�tϡ��Q�!�����":�X4V��ͪ3M���L���.+Cgn��4L�	0qR��,*X���ieҢ]�'�� ��r�e�A����`�c�\f��yk6T���]�;��<�>e�K�v��I����=�=GT���'=1�M�ab����h���O3�'��+�En���xgr���:��������SD��P�����籸�4P7���X�]Z'�E(���R����Y���:b�k�x�I퓠A���%P����z�˨4eL��	�o}���<D0�iT�vcg��q�dڻ���ғs7�&�7qrE ib
R5�)������1s�;B�K�?��ɷ'4 Y��� ��_t4�ڇ�p<�q,����z6[�j�M/����ʕv8��mAuHXZ�Y�a�9�qw�:��;��-A܈|?��=\l�㕍<fަ��Y�g��{^�!����J-�Us'��%-3�T��1���d�(�>��J�J	Z ��p��0��6v��V3����C�@�S5�JZu�Q�0m�_��U�����9L�#�J Nȍ1&Vi����i�I2fŅ#�[w)&���b�<��5ssca�7�R14 s�/E��A��w^D󺧌����:={j�J���3���� ����izq"��L-��3]���=�P#�.L|��׆w�����:e+�^�U�9
 ��'���5��a�������ŪSv9�ѡ���b�H-΢I�f!�����^��d�Lz`Cs�Ą�hg:6=��X+���D��<Y�f�&I�t@,��⠄��\cJF���I���#���A�V�)��<))��,E3��Q+�c�͋G(d|�z
>f�H��Qָ�-?u��/!D� ��.v�Ř���ԅ�&;В�%b(�)(�=�N����V��rRBIV�q5UD��R�L�0�e���V�
ycy�hV>c'���B�;���ո��jt@[p���
ue�g~���{?��LOm5���t7��=
Ԉ*�6����4�o䁰������uq*��N���7]�c5S��#�׊�}ӯ�k��%h�����c�����k����� ;�9������!�wr֞?,�]��c�%��m0*Jn����+E�-%g0sp��-���s���m�6�����˘*���A�8�S�A�n��� -����pL���^��C^�`W:����	U`f(�h��O4Y���N�t�����L�4(�(V���8|��3?��u��>6�N2e<�d�M8ҝ��1�81D��m�aBvlWM�.O�����ȑ0�"=���M"Y���T��p��J�T��2 �������*nV�}z\�8E��OI�L!�1�g��V�)F�E�j�& ��ԣ9=�l�;�4�\#!�R�5��,����v�oC>�Yd5l�UQ�H�ٜ8Lo���8��Mh5 �����5�
����3��8ր�I�.�.�����p�~۫Q��=<��E�	���=ng8������a��S빍\�DY����?lߎ�{���Ld�:�
=ј�G�,�U��;����RJ�$���~���;M �,;w|;{��%i�3Q�F�}� ��k��!�{��+��a�����j�od�������0�g����ȅ����.:�������V�a�T�([|q����a����v�A=|��^&l�e���i����������cǯ���/~�L�� ;fcp)�x6�X�n�hW7ԵZ�'f�J�$�C���c:�(W*|��i� F���Ya�&�S�J8_�OY�\?��Dd�����Q��^��w��ܙ�K_W:�����8���[�'h;,,M��&X��a�ݜb�������{��rj�v\h��[�l�4�W��hD_��!�N�}B���Ƣ���}]�ɧF�*?���V@�ʿ��-��dѹy¼���~A�����tr0�x˂Y��R�-��Fj�I���u� \���jAc�˾��g��;�ױV_���M�(�	U%��-��4�@�)J7;�����vdz�^����%�~����r�F�q}��pԇ��1Ch�kOԚ���6X+�J�#���k��Τ�~͸I��D�j>?��}W���>s��C�<�7*�����շF����x`��n[��c����z���l34'}s�R�]��=��eN�%q��	6N<���YȬ��n���e����>`�dՆ�}j�A��U�|f��4\TΘ�6 ����ϝ7�G]y2�_iw8p"n��U}��+���7̇��oZ��ēRȄ�]����귭&35~��=��|���_}/c��8_3�b��Y�>[��C��t�5�����ٱ�r���Xo�K~�������������������D؏��-X<�I��y�@*�mŔ����3X��rn���Ա)���uxh�������'S;��ň*�]R�=�%dBw��N#�J��ty[U�䯉�����2��d�'�����<�ڷ`T��*��a!��xu(걑zr�+@�d9rK��$?8��&�+�]��w����}v�B1±���'���ߕUW�W��Fb*ɽ��c�:1�$�e{,�~�#$�����c>.��Q� `����Q=#��:ִ�xC�����g�D�#'��t��֘j�΂F�/�����\��qi���Rr;ɀ�{�l
��b�5�����s!�!nbǊj<~��쫲m�x฿���x��a�n��3����*� +TY薑>�[�z��17����-P��QA�$�H�K9 M4��w��om��khJD�D�����u<Fr<�?Dq��p�ߓ�R�P�C����3��!�H/����&*+��e�QY��O�q��N.w�J.����
��ǎF� BB
���Y�{e40��	�qdNc%��3j��.��Ook2k$�c��Q��7�b��hL�߱�Q��9�?�h����ǈ�dƿ3�b{�s����ο>mxgdw1��"�{'��cP�;s-FQ#E���P��Ȳ|��u���];s��P((q��`�2��a�O� �F.�U���f��tܸ)��g��uR��a�"�T�)�HW�o�M�,�mg������t��kP���E�8�����@�Hy8�n<�#6����+|�v��	���o*�����`z�!��+N����������Ԁ�����D�Y�,p�n��vᵡ�������87���t��c�H��e_}�G���+i��0Cp�u���f�]�ң��X��j]�ĺ���?"ۃC'�����E��E��������}d@�gW���Vr�>D9�'�}���3�Q���g��z� �8q�?]��T�:����i�H��bc�dU|�s>�EY�����N�a�����f	�*�uAb+>7��S0��TW�Ji
��y��PQ��G.���hwl.�b)��q���#�V�%X@�=ڵY�V��(J�	t�R�i�y٨��Q��#�<@�4��*C�; =�C��V_A*d�B����,�����6�Ō�.��~y�5�/`Ѹe[�`��Z���"a�&&��w��;mW�a ��SQj~��T�c��AV�%�z��&D��!�p�J��ʂ@�����F<(2��~=4HBR<8���ؚ�JN�0Ƥ��7��Agd��j�SP( ��J�#��\M
]-�9�nk��Lnڹ	�'v�cCz���J�pH� �h{K�*V��OȖ��z�ݪ��Jp�}��kO�����J9NH�\��_�iO�^��I^��P�h'7��x�4Z��X�q'i�G0��fSF�ޱj{�"�C��0a�R�����~�?+)���L���]R,um�[���0�|T��=����[��V+���1�AZ�;z���Q�U\�ukk��0ij<.�ǠD��G�Tt.[�\�� 2��Dc���Ѹ�j���h�y���t����#S�l�t�76>������6=~w'��vrl��n�Lu�[����^s���Q(���
[9?v�O�k�#dTf+^���``�/��w��|�>h�O��O9˂i-c��L��ȘyB�{c�=�oq3�`�e���@�W�-��H�?�u�A�����'	�m�Ҏ3�	{7�"�� +,ZJ.��Gf�[&�A����T_�$b�v� �|	 �c��jit��_���!K3d#�],Vh6G�v�0���{����x��⸲��(�W
k����^�w/*�'�|�=rI�Їd��(�aY�����~�o�S=ϐI�V9�@ݢ�u�؎@ͭ���o|���|���l���q?G��O蚤o�˲k�R�9U�R����������d6y6m���gŋ�Fb
-��v�$5���J؟�"3���8����K�0���`F��J��R��@�3Z\���%<|�� �́_BaB�漬�;�A=P"yx �d#�>�?�?��N��>���=��hB�&��|����TZdL�JL����Gp�{:�1� ���6U�!"�;R��f�åxa�e�J<)�� 0�,fF�=���xG�kN���'5?�BYy����[[f��~�{a�#!7����������%v����A]�N�1.F�="���#�����ы��$���
�1�˩��(�q��q�l�t=�Z���I5��9EuH��}��}�no���Y�Ì��g`����=���UD�L1�fl�<k^�f�t��e̛�Ⱦ�����q�����ma��B��w3(s����'-�:��A�5T���8L�恌�l}
�R=/�7�eh���,�����<�ˇ�.�=�u�F���W=��j�V��3�u��Z3�|��n]#o���_�h�C*�o81آ:��a.N6_����=��sO0
f�o�e\�jd�W��QR�q�a��D5��b���N`�KZ9�lפ���|3�)#2-�=H�-�V�^�3I��w3��R�Eq�����V��]ԨZ_FQ�+WrC��Q���?��G�Z-$T������}�L� �b�/��.AR��m������o��=��{ ���vs�س�$'ԇ�ҁ��x���~�"�	�IE�0Č�e�c>���2j�wC��cm.
�f�	/�g�x�g���s���7�G��M6пw�Ax�����ST��?�.۬�kJ4H�$��ȸt
o___At�\6q#��T۶�l~��`�����I]�3~��+_��S����ȭ��Ն�A|I?�Ӆ�5�v��O����G�C>2�;_���}�]������z�-P���7Q?�{%	�:F� ��1�f���a�/P�%��=U��z�ŵ|���W)����7�o'�#�.�UB�5�'4Rc����ט�3����0n^H�k(x������&�]3�̜ӝ>���<�`Wj99Z�=���lr�ޓ��3�{���/��c?x�3zO[��������"�_f姅s�F=�ăA�zσW�̽���@�OJ4a�n����T�~zz
�J�M�1��\	��g��\dD�a�ڡ=�)Å�Uq����y2p��������7�߂�H�<���7���y�϶�^�Wӗ��C��
���0�U	�CaA/�fBE�6�>bB ���(���1E����$B�s��w�l���-��}�iz��\s�,�SV�X}U]t�,�,��Y]5��E�9����v�ϐ�f%�����V���Dr����~�vL������J;=Z[�����j�P(�D禍���;��=��tXX�b�+�m��f�N5p��?�갡ͪw</��~	9c���ɡ T�N�9��"��`y�������r�}7JU�����D=ح���|j�mW� �-���ui����'��@K&������{Fu��#?a�������v�����gGV�j��\��VN:�����M���CQ�`ۺ�5DVX�I^�ԕ 'gl�T�Vk� �JM�7V����WO�z�oA�s�hQ^�M�UP���!|�E��j���4ￏ(3A�lB����Ũm�%���o����w�4bh����Էұno���N�&nTpD�Ɓ��O��A����ҋx�	<ad�4c��|�����PH�3��t�/(�o�&F�>��umL,Uʲh����؅��� �͔gw	n��j���3��W	'�ͣ	��xE������^�!H��h��_o���kn��z�]a�.��P$yT�"�f�Ig����� ���l}�T�1�Uut�f��15�26ʇ�������(��)U���XLk�_w�g��S�y
�967��m}Ё^�ok`�Qi�(�l)K���]]]�DE���`�0�Jl�J��U�A�im�ଆ-V�K�5׽ٴ����D�mKo�^��Rl�Gh����� J��XM;v�E�Y�&^�(t�����@C�s�6���(�������d��(]`��T2n�K;�pb����rD�6�M�V���5�m��'�TA�-���Ҥ;�d[��i)i�낽�Z{{�	��E夣nS����>L�o{LH�c�`��~�.b���8���Y�\��n��n�0!rj�L��!����G�<-l�f�2�X�%��h'����o�����k�"(�8����j�SH��XmZ��c)���{(����D澄���S	Q�r�S��ݦU���zI����dS�h.��f6z��t0�o�C����6�+n����H4�x��c��!q4A�e��"�@�擓3XFJ��	�qC+N�E�\�fE����͕��7/=	��U��$M�/�:�vu"a��Na)��=t�M��I��� ]4��b�? 	v�0�%uu�q������tk3�"�	7F].x��}���.����?\
�$���j��D�+��}���p[C"���^6ONZuɝf�p�$�Ռ�
�w02u�A7�T�X욞�B�����W��T"��r�14��71�ǖ���XQ��pk�iC��B=��M�=�!P�.��-A
��OJ����m�F��ȚX���%^�i�ʩq�'�~�enrc�嶒v��(8�@��\����2�M������5t��S]K�t�g��ؕ�c�hMb���ԏ#�;���kR���"��S����U�a�?���W7j��#8�dY������'ŷ$�1���y�-�ʽ^��l��*Y��^|)���8�=�D!xv��q���p�p_^����O'��ͷ��YI�ʶ�U._g��Y
��lgt	k֨�X>-^�k����'��E�笑E���?��5��
Wh�K�l�Ң��C�j
���$����J�b>>�DPY��.�ǆ@�r�Ǹz8ʹ���r�ЀCH�0��@��udg'�ߗr嶅aw0�۹����U��N}n=Zx�D"�`���"�b�>|ܯ��)j�[ɤ5�yx�L�z|���|OC��_�O�y<�����5��2Lכ�.ţ�r����tG��2��
�8�P�k$$٥	��5C>ep���ӭ7���[���o�;a|�s�WRt��v��}�0����ʩ�������;���a �\qd�[t��F����7����tU�,_RNW~��p��P���lU��ѨBY�|U�5�_��R��TP�����d����d��o�����x���촶�mΩ�i=02�icQ�J4���;Yr���jE��ow����U��1�=:�f��#e�.�u��X���:1�YƩ��L�rݟo�s�Y%��] ��$�y�����s�;ۭ<�J�7V���ݔ���i�s8�X�K�V��n)�6u2��W�E: �7�Vyy�E�!�HJ���>mZ �,�2	�Y��Y��J��܁��7,Ld�s���� �E�6�˟��2LX^R����ժM�z)<���tÎE%P5��Ā����s�]��300�2<�$�{�tX7�TR�d���>Fk<fr����_���k�V��F�C��Sg��3��q���:�4�Q��`v�riB�K1��j�%�s�/C����4����b��$%Ͱ�Kr��=���������������|ߟ��v� ��PEW�aJ��xs�B#��s���� �ED;���r���WH5��yo8Z⡫S�We�/�p�m�l�eQȜ;?�	���mǀ{G����?�\����l]�y4�kʋF�j�~O|��mV<р�mO�Lِ�d-?�uy�o�1mEʑ��f�E����Ӎ��{ �
Be�{�k@�M��4��k��O����o7�~�N��ŭ"ۖJ�F��o%[��6�a軸��z�bSOtr�\�r�����F-3����XìԻ�=�������ɐ������̨�Xizȯ���N��b״[�4*�Ս8�[ȓ�ٻ{��{h-)ܓ5�q0x�9�f����:�37�y��3ﭚ���ZPM��i�5���a0[�:9�!��IU�5ə�I�^���c�Lx�$5a�m����{���\�ܵ�B�����!8��r	��ۗ`��#���!�Ꞥj`B�&	�	oU5P�����G�H��`�iL]�a�,���s���d�,RT��s�W-kn���5X��`��,�YX`oH��[i��%����-FԠ4�a�PZqH�Y�����Z5]*맱_9G`^��h��jV��e7���"%�!�N���e$��d��ܫ٬k�SP��3X�vC���O��*>��5��)$X�M�9���=�9{�۫"N�_zd�G��,��	uRL�ꁸ@�Tb%�r��4I=�ˉ>渪߈�p5���*K��������M�U)r���~����6��=��T$�#~1���z�J�=�����:)G�Zr�6e���=������8v?�"n�`uT`	uT�Wz���B�HB���ڔcb5V\A&���5)/�?H��ˉ2Ϥ��N�Ey�
�Q��l�H_Ҧ&b�0W(��$��¯�a��w���h$ش^Y׋?���>���>i�}�֥��d.�')>�X����l���_-s�'�䅍s����.
H�<x�D��|�����=d�����Xl^�2i�H��e���֞�w��ܩ�Wg����cEC�J���O�J9�C���|m����\����dr:`�T���2�m�G�ȁ��<�(;���B?����j�l@\:OqgN��֐G`|������SI��')���V�n/y_����kDs�
܇�f'Q��Z�"NV��AW�����M�C�K9$��R�w3�"c�Krp,Y�gDφu�e*��n��XqF��3]��q�a?��Um�5�ˮ��w���v��k.�� G(���	��z� u�nƗ�,qە:g�'wU'�}��z�������.AA-�0c�o)qn��_'ԅn��F22�'I��|��<�%��d[|	7v3K��ߙ��x�
���{qyd���-��Q1����K�T����!c���o��Q�?�aD�v��[eJw��d��3���������\㒁�0�p��t�G���=��։fѿ$�Xހ�ߟ.x�[(6��ݺgϋCaO��0��~��n'N@緶h��[!(�k�,��i�͎�kG����tO�{���>�F,~}B'/���
Z�z��Lw�*�������±�Ʊ'��b�U9����\��>�Ǽ �$�!}�m�Je+�c�^�#�l���ZNxWs-`V5��r����2y�����K�3 X��V~8���GDݟ���p8���կ[�[�� ~و����nnG�D��Y��C�0��3
+��8m7��P=ҕŅ5�u�?Z�������ھ��{�ŝ��ѩЩ�d˥��<pzh��l��p�U�d:�8����h��~X��	�����&/_O}�$/��͆D���^ع쨄e�S34&�-,��?O�y_UKxy����7wr'ؼ��h��6�vSd~qz� ��;�+̊�x9֏�y"��^s���h���H"lG������i3=<�0��"�0��
����H���u�����%��۟��P"�h�Pv��>�D"&
�>
	��5[�����PK   ��Xq�q�  i�  /   images/963eb574-430e-4d09-a29d-074ae2ef552b.png4zcte]�퉝�m۶m�<�m�c��$��m�Îm�7�{Ƿ������Z���=V���$,,  @��S�^�  4���Q�u���")���; � �b�j��]P�9�n��O�F�<B ��roLit���������ANNjڏö�6qw�=37実)RѹbW�XF�!�rW�o� ��Y�E;:YͿ�3���x;ҋPE
+Ã�.1�i�uW�kTj_:h�om`�Ue�&f&�lO��>�R$WV���`���jk%����|d�`[�cnV�~yk.��R�f�\Qpx�bRj�['���OWs�$�ZN]�]U��"����S�9���D�! `뮎�蟯�"lحt��+wK��� �pX��V�ar��W�"�����|�~M����kYù ���Ϊ��+f��?SN�&ٺ%��G#��W�S���}�{q��fS�Tt�󓬄�*e��z1��?ą��k��'�.a}2��+��KW�n���#A[���._���c��(�����Μs�e��´�tI������r  ��)ո��`���vi�3\oy��v��A�4��h�'6QPG]=�#�&�@w�v6��͸�v_�lVi�~g����-."Wa�Ŷ����y�ǀi�77�ez��/A9N�r1u�P�
��r(��{��2�=m�����#�yB���A�������SQ|�U�7��o17�C���v��v���槇\_��e�J5�4)9��z�������Y%QIͭ���S�4qu����E�����}!���87��E�:p���ֿ� i��n��4�o�/W_q:<X^6�A����y�N��7����+�ܯ%2��0�j|�x-<�Olj��z��h�.�U�6_3ER�.�.�K���=4C�`��}��	"��g�Y����+Z��zn�9�	��ٞ�c�����τ�y�W�&��J������Q>l8�lŋ���5��=h��݇�JG�;s;���K���Ե��o��5s���?�W�=�s��f!qx�?ٴ�M]`��ی����>.O��՝�����׵����#
UJH�� g�H�R�I�זKKh�c�>K�p6��;���`�v����y����{|���ή�OMC~Y��k���jd��,�r|���p��G>�9����V�ʫ�����7�J��z�O33{b$Ls��U�T*K�L��N��wD��^���_GzP�v��]_�-��*5g� ����|ojl8�����O�����h��˓Gwяu�[3a�-�tf+�����uJن�	��-��)-�G+�T�T�N�I^Z�t<��mU�]	�4�n��Ǆ(��c�>�Y-��ܸ�9�o�V��s�<�:���f��7�4�3u{�yOo�^/G��ǎ;D�q��Ī��;8x�#vX�`֤�R�H�������C������O�� ���(`�мZc�×w��tE(DR^WbĲ;7r�iߙ[��v�W��?�*Hb�^,_�۪ɪ��t��5��1�B��d�G���f���%fBi�G�jaP������
����cؙB���uY��}�{p��_��9*��;�w�$T<7u�6������{�ǌ�XOC�4u�U���s������xe����5F����s�tE8���o������� T�&_�m¯���J�����%,	\������I@�a:}�׫�̩$�C]>�_��aU����� �AjG�f֓@���i�Nb�h��ϝE�+�F��tUUY��$ԟg��J�j�Y彽�����7�溤���f��q���u�E�_|��:d���ȆO%:����o���/w��o���o����~��H�3�o͕�_Ą��gPSs	M���a��g_W�N�P�B��ع����[:*�_nTl���b�����=?̴R�����"��AՇ��Wy�CsJ��?u�"׽#���ܦ
h����35wK�����Y�zQf���d��EU��ۓ;�KϷ/nՙ$;��ICíx��	q��\x^555�,��>U�OA<�����:-|�z2a�
��H�(3��dusZ����k� �H{�\�{&Ξ
��өm�ګ��.�}��<ߧ|ҝ�lx�cy����iUg� �+�C�Y#T�b�R�5ۿ�����P������l94MT!��]���Uv���L/��/.��"���b�Ʈ0��4L���!�m�|��{��]����r?���%�hWlǅ����ݣJ�S��99�Ro�ڥ�ˇ���Sю��Gӭ��#A���ה����f���o�DpX⒨��tg�f�� �*�]��Ny����r�X��}���Wm)�T>�{ta2�U;���o,oݤ���͝���TE,.'d�)�Mˡx�:�;��7'%�������G]�Ms�J��8��鬕kT�W���|12���-A��'��&3�Ͼ�^&�ݸM���#/��٥�aǖ%]Ί�L�汸@�ϸx�����GYt@�?B�\h}W�i.K�E(��q=Ц7�Wj�(�=�N�<���VF�@�j��&�dȐk��+Ѥr��<�������q=���r7,���������ܿ�}:U
����A-C�����/�E|w5�R�����[�������6�I#Q<�59=�Ň@N
ƾ�1%��ަS{M,Y��dW�������&h{>��Ͽ!XYU�N�VU�j�S����T]��P���BQ�Y̯�������&HH��چ����{�.{;i١��v,��g'�|7�{���o�?<���̸����1%""�����dJ� ��ӗu�w'���x}���&S�55�G�2���449�J���(��%����nϤ3JW��kT��j�*�����i���N���~� ���������ՓBd^۽�f
w�{���9&75
��=���A����+F��ӤFS{�=΅i)�mWU���WVF�sLٰ��4����+�r�̠M�H�׌-�+~,L���0ЅO���Jzb� D�A0?�CF�%+7���.�9UVV�tos줒pfz� �n���}U������s�?�k��k0ߋ�������۝�RW#�N TD
5�Cqz:���JWC�3m��w�����[6>���Nn��ET�b�4�y\o)����������C 6l�������._>--��((;��͉ӵ[��)4x�)A�����i"X�DyW��Z :�]8������?ZA������kS_f@�HrV�캧��^�ҡ�Cz4Q+��وB�7F�=N������}�"�j�[����]�h�7?�CzP/]��^���b{e���d3>�
��#�k����-�&�"�8ܑ��v����9fؙ��Z�.��Ӄ3Y�W�ݷ��bFJ�1��	q{�!E|���ڥ�^I�o)~3B�΋��|�M̒]Cj�T�ot1nG��N������?[�b0~�������N��/�t��Tz�[ķR�[$x'X��/��������%+���aU���9�r��� G�h�`����ͶrI]��m��Գ���eG�hGTr[Q�����lI_y>-{3��ͻ# ��-�{��n�̑K�{_o�8؄�D\v�J��[ͼuS�q��v�D��r|;[:�tiRe�L_<.�=��2�Ӿ'�Wut\4�}N��c��;�de��8�;�M��.{�|t�ݡ���T���hhhF�-�6�mO�|yV�y=����uq��s|q����T��~�k�Y�춡T	�/����R��	l޽�w���=���.T*���A���NGo|�O.N���	�
��ާ����,�<�믛���刋Lic�كBk�t=����S)h���]ww|*"���J�:����T�������PYYY�	h��H��{�WR�@������{��$FE2e�A��Ƈ���a���Y�}�KY�ݖ�a�~�;R�kqqq�E�_+�*1�B}�\�6�f�der��R>�X;��D)2�L9Ȱd/s�ty3V�0� �	/kGu�R�қ�#T�Z�0R|4Xq�b7oH^��~�ՋY�u��U�v�Ʀ��[�}Z�q����egg�C2����:�~�Dsbe+�N�)�:3�z��c.O��G��B�"�Փ�.jZ���U&yla�CЪj&Y$�C�<�֫T$S�:E;N#Y�R�M'v�d
(}��.& I���c̆���S��P���)�ܺ��K�]==�����5P��'_Β�ȓ�R�]�C]2H6�����F��I��b��C� ��`eK�(+/�L�*܄Y�.�<)��Q$Ѷd�/dU��38��/bf���s8V�>�N�6|�.T�&�"�O�������Դ�t�þܕg�����aaeE_�"�5�f�:�P�[�Zǔ��5��߯��{*��5�0����SUJ�ËS�>>����1㟗j���D�<�E�{�y)�#"���hǌ���
%�HH[���-�,��t���R^� k��K�����͕���Y0,���;\��e��O]^6���2�7���{��S���Z=�`
��F�j��Q;pB0��g̺�ɋ��5���s9�vp��naoo�v|���u��Y�|���71FLvD��i�����T�LiEGGv�r5D�4��s��^�TyF��M�x��Ac�Z�/���Kg�La��@"�g�#F��Wh?Aj�*[���s������q�����q��S����Q���u�Y�H���S4�����4���n��һ�YW�+.^�$,��*��E��<JZ�MLN���EK���,D�-��;��ח�e��>�B.XD��Jgco|���G'��T�Ԕ<��H�) ���9"��F3vIL��:�3	 r3��A#?����wڠͩgp)��gm�z����w�"jEee�ֈ�ϔ�:<!,�y�$P��y��\x<�W� C���	�5i{n�͂im?ؽ�/� ������l�o6��:�_|����G|>ϟÔڜ\�
9;d�˲���P��&
�H<P_k���&�������F��Q��3���L�g��Z�Sz_�A| �v�
4Lb�H�����	Z)1NQT󒛺�z'��]��;G��i�~>��1�z���񍖮����d'���q��fUU�T3��[Ǻ!���Ѓ�|��t�����}�'Kۘ�����Ǉ��5,dH�Y���N�8���!ZKG��L*%V��\�@���i�q�h�#��&.��wT�o� ��W�v�\r�!0��r�W{6ș�~�O^̺I�k�9oz�]�:���HΨ���������.���8
9Jf\>fJKc8�I�5#��Ê�_���.pD�FA�o�	��q�-��~7)xeg8���������s�Ζ�%8�w�qŒH;�C�!��N�Ӂ�759ym�Ԍ3��Y�W�_,%��6Us|c4+$�2�@��(�s'��~`��gd�L�
�&�'���zlU��W13!�\vV��d���E����Rvn���C�wt8iʸ�'i������3G�>�ޚ	�C3�݋�Y{�Vk��R=��ڿ���b�M2Vk�Ɵ�
�F�LLL�<Ң�.)d4�8H�E�� *:�u0x�`9#@Xv�R&[%:�ؠ:E�j�I�����5�q��xߒ<�("��s���YbĄ=�]Q+c�^��`<���排"��
8��S(G1�{�_6�ni��)X���,�J��K`v`�dvVv��֛�|���xP�!.�-9��19o�Ș����2c�яW[���yd�"SSSf-Z�UYp�Бp��0~�L���0�{"asʗ�㪢��ީ�=�M�1G}%��S;ƃkvSNy�x�祖,	�PI�cb�^B�B]����w�:��aU��E������!�����K�㠇Z>�R��}���5{Q�F�ql������ޫ4�M�(�`_!F"��ߠ������U�HoF��q�_�1�Ԣ��<�qLd����+������+����f��,(��S�jأ�u�V�O٦y�L*B�
����������+Ϡ�B"�_����I�@���0�6s1c���c0lK�B&
�(P��Ĭt��Vl�X��Ѩչ9|E�����ܭ�z��;:�ާt�*��x��D��/!!���"?�jƂ;z�����P��-=1f1��a�s�u���� ;��<����\�f(?��!_�bN�,��y�������DV��&��:]k���A�:8~��ب�#ћB8B�&�I�b�n�W�����[�kx����Y��l!��+�5k�M�֨}F���8x�sU.�d�(ny����h�>Ǣ�-B�b�av.O����^FYN�?�� d��o� L]�qvv��W[W*|Q��d)R���<.1�˲Y��$�Qsg�@Ca`�@{L�!���U9�X��"i��)�<wb��S�8?!��[^�
lHd�^�"�#w� ��=�ي�ʮkh��r�5���P�H=��S�|��e �H�^�����Y]�a_�����(�^ʻ�
p�5Y�;�Hm@�<��c?����/����9� m�6G�<#!��`Ì��'f���<,�N���@�@z9����CF�t����K�8Ux�I��x����R4��Rf�Yt,?*��H��-d�*"�_ߤ��'Ӧ}��w(;6��~Q[�,��vk�j�S�����1����R���d�y��-�&���{�u�6p�^��1�n�]�{#���hy���Z�zim�x���w2t��t��<�Tq��E�4]F��*[���N!�\7�*�A\p�}�Fɂ>
�ύdL Q����T�j*0��a��*�� .@{��R2�+�5�J�VX�	��AL�c���:��vG������x�	�������7c3����N/�@�q����R���7SN~����p� ����<�SE��~8'�g���@��� w� �;
x�(O���p���$8�#@䙫?=i:�e��S��V���z<�/�`�#
��$�e>&���[Q'A/'J�����Y����k� -�����c�Z?��`���~��$�C�в���>�h��S�a�!��Ǿ�>��74,)i�	H��_��.Mt�J�wj�������9���P?����4k��i��uL�2�+�tid7��.�M�c Ѿ+O�%��S
o[?��g��R�~?��y4T"��;�6�+)�V>G��|Xb�i�����*a \|X��<q2�ŁV�n�_�	�>m[&�r���QBh�-Ya����Z��s�?��5��򲺣
7b�&Q\����zp��@�;��_ŵ&8��M����m�7�[���1��t�)��O�_�ɔ�L���!F,j���H���dD����=\5���H}u}OB�w�b?nWᯀ��T�z7m&1���'�;�\���,�#Bd�h�5�k�
7]BtU�2,ر%*p�|�2b�DK�e0�DU$f,�X�$ū���:�����q#����liD1S2:!����N*�A5�/|4�X�К�\�)^C�������pOF��)��s�_���3
P��R��ĉZ+�,l!��B p��?��
m��Oؾ�V�g�n�yk�%̅�FgvxK���DP��(Q�QٷMHQ�_�u�+�b"G!]�4��~���A?+CC|�+M��?]�C ���!Ņ�Q=�-qNH��d]�s�}��l+���
�J��w�O�+<�Y[>L�Hd?y!@)l3
tΤ�F�\��iN����u��h�9��F;���Ώ�gr>����h�X�@�QO�WG155טBX�ئ`g!kDI��ДA�'d=�.\RDlu�Q���=+��5���x�Bt ˹
�m�r���e/?�P�^��a�܄�+5>a,�)1.<��B��Q�7��6����K��
�h���QD�O���x��*`����:��D��VS��'^~��R8M���# ܻ�zFj�Y��gs�Q�w?�x�Y��0��yE$�]d������Ge��U�%ZrZ$�`��1�P�1}�!��G �&g��VWW{SBJ}�wy��mEY��1s�!�HgS0Ӓ��&���Uc�*6銐G>��\1sǴ
|y�٣�"���,�:�.��J�wji�Ip�F���G!<����ַ���t�@�c
M����g�k��(2��<3,./Φɗu��]���>>��1�{@9<^�]�����(TH�P�;e����`B�8�9j�:͑��U���xn�\�(�/�x��G�Z�E����47+3�[*@@J	kk�T.�� ����7G��oW!�r���(����_�H�G�1P\�:t�Yc�yNѰ�i��O�T��O���]�y��S�b�k��}�����o���ܱ���nf%����O�.�)VQ��.���t�T��ed��k�[�4�q/9G�uD9��:��ߓ	�	��
@4c��	F�Vyn�_�aㅽ�pl��a�;b��>�����h5ꋚm�o�#�߆��OA�����Y$��EL���^m+a�ͦn#Ɠc�ߵb2�!%^�n��XE��X!)�2)��a{��{l�-t�KZ�Ϭ�p�y};�1��aofk��f�g:KL�J�bQb���8^�����6qq�`� \^���/d�݂	#��Ѓ_%�oD�ﾂYJ#v'h�Ƹ����1'�
Y�b�I�S��}�	e��/���Tu�G��l��ŖJ���c.ۡ[~�5��c��iv�m�+�W�"cb|"�~/��0�f�a����Y���|G�v7]���A��u{Z�Zcn�0 ����Z;�l5�y��G�Ŷ�^�O�33�� �aE	�>��U�Z\�m>g��GX+L==����Vm�b����
�ϒ�)a�I�p�+��!�<
YB�Б�裟��"��K�%M�8$K�o�G�j,�_<�&���{A4 �2J��߼`z���������\�5oJ�KԬ=[dC�)��Ƿ����0�
>��8.M7@Q��Cc��{��m��᜖>����������zᶌ,i��j���=��NJ��6�L��l���G��@##������O�^��d��mNɀd��.,-�7,�xj���h�Q���jkk�Zm�@4dɁd���_����0#�	��������}0ȉQC�����H��4�������v-*��_�w��u���H�_�q�^��� ��~b��{ů��I�^E0N���+iT|A�$��=»͞�W�������-�з�'a�c]�|�Tym�iͽ�ӂ�����"<v�ō�W_gn{<<�ǈ�^���ެ���cY���o�K��f+R�pC�sӭ�X�+^H�H�R�R��LNvH(�}c�Z:,�w;��ȉ`\z-;�s;8Z��h���"����{{P[p��;��o�]�n�W��}��qP�<�o���Gq��s����3Jv~`1��#OW��Z�&�|b��˕�L�͘����_E&oƞ����*�Ƥ�^���@IJ�2$a�h�R�=ˊ� q+PR&��6��t����	R�u'�+#����C����$�����w���K���s�@�oG��_kw;[*�D¥�xg�_�|�>���`��o?_����@��������᭮mIZ�j5��5��MDlg��p0����'l��������F�tmh�3V|��8y�;�g��^?TVR�ۋ�ӆ��
��n�f�)���G�C�˄Z��E�'���;%���$	� �`������+��*"2��K5���U�D/{�Y���8��uѼ�5�XƬ*u���7��45+Y��=c��� i���\ԙӷ��6il��}B�`B[$�6I��2}?��j���Z
�zK��[P�@W�������(��M��R����3]�!�GV�l[T6#��n�z�bB)���
���cF�_?JQ�J�����8O��Gխ({"R���#d�N�{3ǜ�8y��:۠��D�g�Qp+%&wݥ�(�������M��dƶY� f�3�~ŕCћTD��}EۖD+{BU�-�F����ϰF�jZ�S��O�&9q,��O����Ҁ������a��6U[�����*��vF����� �{�'.	\�)Uh�xN��<����4&�I�
Jhj�\@4T񔸘8�6�J��p��F�P?I�i8zH��
@��%g��V��=�~5�\M_W�V���E+e;��D�p�IKN �YN�>����e�~���Ǣ�ŖF�	�_��"hWM���2���L������Y��1{���3��1�'��z߳b/�=e���
��^}v�V�������"F���Ĉ�^��� �?�)DSD�dr�ôl�@c�*V,��*[�U@I�=�n�O�j
,$-o��_f�'#6�O��K1Ӌ�Vm+���i��Ә#���rPZsm��ɍ|��TK�(w0��zÈ1����V�h�~Ý$��>���&����+��d������#KD_nc������і��g����@����U���Ȯ��o�y��0Q�Ρ;�0��|tb�����9<�"����EMvzo�&V���޾>�b+��1I��{˯�E����T�]D������_#�#-����-N
�Z&h/I)ɭQQ�D!��m]{8��43�����"w���{�\�En�>�9��?Z��l=��cx5��eBoW�]	-d����$!�0C=�(z���!�,�H|�nfg%8<�
��]�N�n�^�8HǓ�r�A�v=4֠X�,�M@���?M�AX�W���/ypT��ܚ�2��
-U��|K�^�� ���$<�@.ѕW#�1F�}��<�:w㌉��ږ�������^"�!tBU�N��>��ə䟺_a�E�h�L�]�����������A̯ѩ��j	�ک��$%e~F!��:2�H�>\�\�X,��K��w\���=��v��"#S�袂g9vۮU���O?%��~�B��?=~���0LZ�`d�塔�P��J4�&/�)��<K�Ψ�t�?��"��n�lJq����˙P�⥂���C�zB�ӕk�x��ESk�D�
3�is�*�I<�b5ɲ� )��4,@W=�Y�1 [��9��Q�#O���njnn ���K�`a����QX���Ĵ��'���u�n�P������X��25��O��&<Wc�q!��4�*D͍@�cV�t�������o���pu�n� \/�e� ��D�9f�:$�c�I�`��ch��#��}4g�7c���cT�tt����$��i��Gx���/
��(z�$ǣ�z�0L�ǚE�ڎ����Z�C��AK#��8c���Q�si����M'~���1�KcB���=&��`�H����#��(��<<�	Z��h([�!q(��Bq
r~�
��f��~*����m�����.qj����V�$���=XT�cQC�f,HZ<5J�%���f��-g]��Gnp��s�̕�9�'�	_���U�\����97&��Լ�E�x@ɴY .|����l�+�D�S�G�[���rx_����\�]`~j��!n�[�^�n��`n�JӘ�G`�J�o�U�tY.&ࠀ�����}.q�s�A�� ���ZD��0��C:��[u׃�ee��]+��x4ʸ�,5���&
�b���Eum���(Z6��T;Ǖ����3Y�����d�䏫�Hڌn�5[0b8`"���Q�C�#�w���c^�Ba�}o,K���Nu�l �'��㴈k��f��ծ�J.'�	�ÂC*+]�j�l��t��ڬb�*�����#uT��K�������C"�E���(s*�lh�2���ǀ��C�m��0&��ۂ
5����������L`��~�n�`.�v����,�RJ�{�n:�ZP�����\�HɈ̘�-H����[Z�:�w`t�֒TH)�\ԣ�۪�S�h�z±$�Rq�DӺ��`p���dhik*;#R*���<�~h6 ��X�~'���vFC��=-��MwEp�o�;�&����4oE�,k�h�ǈԡ��d��������L�*�e4�^#�����3�?�ѹV�pü���;8���pj�y܍@�B�F,�f��ߐT���u��
�+^�6i�̞ݺPS_A�B|)�s�0�����y��Ϊ��P��8�qń�����+:0��8Y�K�K�
�
�Kڕ�Lc�ݭO��-Twf..\A��٭r nb�άdu(T�0������\n5~U����-����j��;�w,y�zK����3�g�>\����^�qL��x���_�n�~KPx�$u9x�� �kަ���`������%nHx	��:���Qe��ݢz\\��Ǖ_P��!������]�R��;f\�8짯i��ج23�Ԅm��n�Ib�t��޶�7��k|-Gy�o�rh�a����m��X��'��ȁ[�.wv�]Ԅ[��M��.k�0�@�%2�FhcAqTi����?�=������Ap���8��&��#񪚒P��N�^�.�k=c���6M��x؁U����W�[N'YWp�ǳ�AA���Sr���E�h�(����н%͚9UF
�Y���4��b��b������Iwn��ٻ��p����������S���v-
��kO'�s�l�Ў��ik��v�'��� 3����@������a�	�WV��YRFͬ7��۽��5�X��o��N��g̥���Y��zm����!O��tއֶ��i0���g�Y2���}ꣃ��pσw�#4Q$tp�XX<�Ã����*W�eD'�2|����F`��T�7dN��#)`�E�ڼ��_Lk�^T�V��P<�cN�TCV+у�$�Ձ�N;VQV�W׳��e���'�����beO�Kס#�����#:��mZ�����|W��Pu|����{�f�ә�N�X��wB�T��5�}~���������f���7����2�����Z9�Z�k͍�	pzh��k����V| xE8`��,#�NA
����e�l�q7`U� N�Ih���{)/���#�����FC�o9�C�\�|�P�	���VH�4\�u��uk!:�u%���h9p.�&�-#	�{�#) D��s��-2͂ōae��[���q�6�(��1st�@��?�Gς�j����������d����4�C�˜�o����!!�s�A�7Z���NƲ϶�)T��f<z�qr~�#���s�Zv9.�ZtT�PTm��"i�\����Z�ѻBN�ݨ5�!-�g�Hш"��h����R�9]�e�=��%��#�6������_ ?��I����8l�ɜqڕ:�M+0UUm���Y,�}~\�hc����_Q|����x/;lu瞡#H� ���R,ml��`�V0=�`՞f���:\ŝ�mٜ�̪�BOp`�F�Zg���#>I�`����>ئ���C�`C�u�&IT#�w�*���ʀ�0vu���i���I}L
�Vu�ld7_��H�� ��!T6^ܒ?����Rt(���r��v�*H��ef|Å�0��������Y��)$0��s�u����֐!���:����Vڋޚm"�mf���i����0�\�±A��t����q���}.|%ɺx܌��,}m ��u�+Nq�1h�	s���<n�h!��)�j�?_�>�`ya��2a;�Y,�tJ��b4J�`nF��b�JK�ߍ�bO���BXO�f��Ό�t���ץ��:�Ma��#�Ĉ�[���4��	��&��݋?k��эΛF� !����:�Omz�o��,�3{��)�tx5̀������&a]fI�s�U�@|��+-4�(zV4��"t�h!H��ɲ���t����6����p�����>�cW�eVj�9{��%�ѵlįbA��d )����i��9&Kb՘�m�Ab���j"w77�0P6����[Qb��(������7ݳzP�Y���Q}������Bv���i5n߬�����H�E
�f�J�,>vv����oE�~1��yy}n����1�_[�j�^��Ȩ�2��W�_y%0pJīK�ݢ��P��t&�H�cA����=}]�c`K�o���� !_Wd�d*B�؊��ǵ��J�3M�-�Kt�va�n��(\�'H�-�c��.6t��ߟV�Ϯ����6��W��լ-��ԓW_lfcgm�"H��q]����s�����3ɾ}Gb)�b<쀓iAQS�	B�e��/a �Q�ܮ�l�E�vb�Q����xe�T��*P�Ō��N{P*h��� Rb
���P'�M�h�U�*�d������$M����a���E�MO+da�V��d!ȱj�/�r1�ij ak;��/�/V{�h���B�C�ry�);O�(rv]����S�(ɵ�j�ڭ{Ch��'DS]#�3��1I	~�$d�)���{0���<,麞NJ�M��y��V��i̖��{,�sa�'�9���xh>�����A�!sȒ��2H�Fz��s���������z̓uo�@�jf�h#��ĝJ����[WIxh�T�������@pA��� ��QrcHjw�m�����U#b�̋�*��['iQ����d�"0^�%>�<p��f��^�wxYM����s���>����%�����}S�G�Pô$��c�OT!|ߟ徛>_~a���5�u>:��O���3`�z�AI�bK�%���iͮa�HHa����Tj��P���9�&�H(xw<iR7�G,tyf���c����vZ=QYY�'�6ud�*�����M��>�%��.Q%�#|�\�|m}x�2�����+9b�����	s-�2�	�eW~o|6�R88�@�%��^�ޅ&��٠~D^��D���۾�m/�yCJLI3� E��֫�qu�f<�#�/O|fʻG�O��7r�Kw�.)�}�<���HC�(Tcn�xg?���5���K���&Þ�z���L��;Q����$׸Ń�Z�J�X�\+k�ٙ#�D�Ĝ�u�R01h�´KFH�������%�^?��?!y����_1UH��$���d
�B;�i�������8P
���~[�YY�[����9���>�B]BB*��{\���`կ[��Һ�=�Y$���kή�H�pg�I����c��ӄek5`�N�r3�-��?��������j���n���(��b�-?*�F���nC�W�Q������1m�p�N���d1�!Y	ǚ��]H�t�s��X���pk/I�|�jV�Z���*�?^f]����T;!�O��+Ⱦ�@#�mJd�t�_���y�}�f]�G�?�����O1�M/�G
mxHg�S{��iH��YȪ�� uCū��AغN6T����h-f3փi\��������^�aI��m���'@+��DvX���yN�]K�_=�����G˽N�bHL8B������ȣO5D��p'��_utZ��=l�L���1�al��YS��x���2���w��=j�X�����SsӀ\���xl�/�q����#��ww\���rX�$NX���u�
BK>���]ac�;ʿq�j;��*���C���(]=q��>KeU��Xi��i�q�[r�u&����e������`x�}��Ir�S+�;�MWj�lD�T#d%s!)�=�U꿓[�;�$��9�W�_��Z���VF&J�3e���*�����gPլ]նf��.�"���la��AV�s�,��MI)�E�\�H�AR6l!�P���,?����d�^_�_���lP�b=����c��n�eG�$ѡlJ���7�!;�-�~�d���+EtE�0�ъkG�����P�(T��*�F�/�u��ZsǱx*�7��J��v�z:�|�'xl6�gba,�`���Gϓ�~�׼�=t!F�0��ᘷr�Ud2�� ������d��S����ma8Tt�(��������6�y�_H)3����HC��$���ݨ�m�|�F+����zW��[�	["�0a�B������<*;9��'��9�t�D�IE| �m��%�i|�L|�~䝦clå�M+�x0��o�g��#S�{O���n�ʠ.o��'PH�i�<��Z�`���N ��8뿝��ə�P2��2z�_�ܦ����T��{\�N���]�+2�ѵ����Vhs�ς����G��ɬ=Tܴ4����H��iu;q9l��& �����$�N]�����(�E$��"r'V�|:���^�VI�;0����bj����S�5kՌw&�Y��}<'I�H���*�?nvHDӠ O���UUE���r�y�ά%Ӓ&'�'�� �ɷo��8����b<�Vh��;c���Q@��Ĉ�� ��ϥ�T\�PB���`dϯ$$�n9�0�%Wh�
'�	Z����a�i	E.
-2�9�$O�!���e�=����P��6�<�IԌg�bt8V���]��Oɜ�b�g���f�B36��tZ�s�(��!,H$AU
�x��f�)��h��v�@���.��{gz:P.9J��J��[n
@I��82!�H��s����q>��ys�Ie=�F��|���#��\�G��exM�c�j1$�>��M� ��)8��B���` ��b1�c��#z)1������"ow��]�vQ*��x*���:QB�M�#*d�*���bvO���rZ�A���@k���Tg�;��,�l���"'.s�6U t�	�X�� �(�	,�%YP/� 
*H�E���8��*����a��}a�8�<՘q��� �R��2O�߸Y�����?�.�z�	C>tj���ЉG98���H�D���Ô���TVA1����[$��Fs0�#�-fM��T�*+�=��� @���.���=�V� �yaˈ�4 T�q!���+A*�,��cǗ�
a( \#�ۂ/�s�d�7��@��p��}I9�B��xh�ƍ�~�&���#��ȃ|y�E�a2����1C�n��倓�'N�1���a(|n��t^I��!.i)l؅ɝ���Z(��g��+��b��Y����������Q���]�������4J�Nrn��"�'9G�M�y������������ �C�A�,Ģ�dB�����g԰����3��Mܚ�HPCK]uݵ�t��?�MO��dF $qJ$ŉ9�?��=��y���vz��gI��tf-e�Dy�f�t��{I�7Q�0�ra5mCw
!-"%��]y��<��YZ�y����{ ���P��0$�u���~���G�B�ALs	?��
@��/�T��b&�ܗJs��o����G�	Z�~�\����O|�{\��x��<�S(E�Pz1� �1����ͺ����曯s��ϩ(���N�s�n���"�F�ǩ�Y�9�#+m�������@=}�@uvv���C^��ED��S��ZZ�b]t���OF�}x�)�6��<#o���K��8�n�� �	Ӝ���O�铧hf�����Ό�B�*��.���7q�^���!����s�M�%�����`"_Ժl)��vsafOO'��jJ���U�����%d3��F� ��	$G�@�X*�0K֢3 ��2���fo��T�@G]o� 8�w�������s�I��l��Y~xi8��︑���a�#c�|���
<0�
�����{f���3z��'ibl�;* ��4B�����V�YM�S(��brY6�ug�h�$i�rp*�yL%����_}�z�{�q ]���H�59��t�}�S^��ha��pC�*��YG���y�	)��0ؘ��a1�9l�&����j�{���*	T17�ھ�bJ.�BF��eB7�f�����H:x�0>|��zqH�J-v(�w~$������˩�������cv���<,?�r����j�Zr�\���x4[��x�,&��,�
Q��������0e�V�V�x�9������t8J�9ǘ��+λI��i��B++D"lS��Lv�����S���s ��s��b?�XGIv�2�E[�ii�l��CNY�����8z\�HY/K��ɺn[����+�閛n�rW=��3<_�9� ��M�ޢ��	�J�i͊iى�j����)���H��Xa��nx�U��D;��Cy�����4�F<��l�� %p���2ir�z�b�sڭ7yʟ�d����U�=����BdB��R?qekBXk�r�(Y����4U^榛n���j׿uw�
���y.�*8���d����m7�B5Օ������Mg�{Q�Qs�c��!�ȣ�u�Z"��uj�(��F��k�u��Q�t�g�I����2P��ڵ�c�U���P����ˡ�gQs��X��s����d7�B������۽�]C�L��CH2a(CH���-�b�\r�4$�� �L!D�(p���N���E�A�T�e�8iIc]{��42<H��z��f�z磊PǀRh�S�9]���9�|�@!u!|@Q�Y���<t�)"sd��xV�?:7t�CS���S�@d�3+R ����u��S��kГN�V߬�by���5c�@I��xV/.-���M�b�O���pNƷ�\8�p�ҖV6*P����n��X��Q��$y�՗id�_��\-���`�d!D,���Mb%>�q���A͞��Ĺ�7]=���FG�9e���i7��`����C�Q�(�Α@I�
����X�y2�����ìLF8j�a��F@ퟙ	6s�K*}	���s`� ������ΉL,�R�TIbz������O౦C�8%�@�f�4?��R�
�(
b��ۯ���ߠ�B�shgg����Դ�]��n�.{�&蛯���sp*q6 ����D����eS7 ��Fst�1�Z-�!���.�:;;}=C�����M2�'g�r�#)����b@I܁�qsH# E�1VMGna�Y5.�&���h���,r3"g�ֆ%�|ͺ�x�2�DHvZ
3fN���Qoo?uvw�|x���O�Sl����kt�gg��ϓ�椻v�f�O-�Y�qJ1�=�q�38wŊV��*��n��BN�����a_�@۾�@�7̉C8��C��;�H������K�8���D\�ؓ�JZ�\��Ř��6�Qd�%w���γ���&QC�f��Pr&�7x͵;�a��9	��rB��5�]�>��?C�O��#��㙰��1J����7ߢ�Ǐ���:��E	��Ew��Mi��±�B�t��qL��E���CM�!r��~�Z��`��n6jC����*�s�l�1P����@=,>C��Z *g��A-�����@f�E�$��\�z��Gk�K� K�23\�3�Q
j���8�A����뮿����t{=��/�ф�,NIQ��5ki���TSSG㓓t��Q�w�~�O��}Qt#Z���3�
��
7�s���P���#��AX��L�|��׹���j�$��9y���j�H�ɠ�-�Y�Ի�/}P��:	��,�
V���-�.�����,$It��ݠ��Ǔb�$,7� #2Q���F����Iͥх(5�Oe����ʫh�ڵ����c.�\lc���Z������a��9s�)1z���#�܆ÔQY��p�����]��(F��sl\#׀dY��ˇ���ޣm�D1���81w�y;����TL
9��G�<�K��$G����C���*	��͋��b�$�}*DTϱ����������/�`�
D�% F`�����laDN�"���X\�す,�︩e)݈��%|� �D�ڌ_�ʣ3�\�r�_�b�Q�,f���|��2��CP6�'*/��[4#�
�� ���vx���̕S����k����Y�MMO2��[��*}^.��(sa�����j�//������Ý �bu1��{�fs��!� <��c���p$БcGEѽ�DK������ʝ.6,�Y�Q�9�4�E"(i6�H�DQ�=2����u6r�����(<������`2dg^I�2[e�ë�y�ā#��@�hSU�8͑U(Y��z���K�H�DR��&!��������e�-l���D|�J����[�a��NMsv�����K�����R8�ؘ8(.+N��\_�җ8Ŏ��}������ۯ���Edr.⟁��� ��B��8�����yr�ʩyi+��5pY�5�AY�c ��K$ENT���Rpf���(4� bBK2��G�w�w?���YGa(>;�8c��f���H(��P8BVBY.�5�V���Mv�a�n6?��]|����]]�]0&�Q"� �K�5*�E��ָP���*�\~�_d"�~����Xy�w7�jr����k���;���t��;J�S㬯�<_��������Z�RdЛ�P���g�qA��}�`k�e��`�&�l4���P(�c��j�뭢]�?@!�BB]_T4�m6�z�N�3=Z[�q�!��� �]]�(���:��t�V�u��o\2G!�������ؘ��#I���SX��8��g>��������|��_fpp�ց��08ص|����;����x�u>�7��ʱ`1��I�s|Nt!�s|�h)E�M�ZH>�)ǾΣ�.�&3�Gp�W̯	@�rU�ݻ�T�gl�>�3Y-�e��Ƃ�o���W�!�Q��-p�4�����Z�ԍW8\;��l��$��yG_�> �C�x���16��*����9Z�HE�b� �Ų�r���?�b������"��`8�۷�˃E��𵠴���~��_y� sB?<ӕO����a��N�nD���)�rg:��)������q���@����H!a�Ru�t��܄E�s�ԷX,N{����-[7�Q��0�ĹX�]o�x��|��*o�]�v��K�P}�pqnŅ�:���������D��D�	E�d4��Z˖�2ѐ����lǮ���E'���^G����Gޣ��,G��k�Ő)��@F�7j9{kЊ��}�X�N�8ΟũrF:�ƭ������q�$Q�Rs>�SYI��q'���u��G��K���F��n-�s(�#��
�韜 �FK��U#uU�W;��.��������} 
�P��K
}P ��譅8+w{N��bF(;9v��jjl$���ā�������R�RU�4<e|�&�]q���רU�rD�AXёH���u�ѝw��;���a� �s�ё��;������9R*��}��W8��b�Jί�'��\}�@a���h�`�L,�f�KZn��,�1P}����G�Dh���h�u!�;SS�~���6����U��KK��t @�d�0�'x��+��/����5��	
 �m@9��H��l壃P�@p�%��*}>�ۭ\sq��1.#�UG#��{vR[�����451Ʈ8�,̓�VVs�zU�H�|�0��O��7.Y�4OfŹ#b����*q�-֊5��124��˚o��Z�.���������@D��T|�L<Y(5>ט(�(�G���
iuit@�����HKpS���Q��AT
��a�CX�M0��A�B$�q�n��	}�bL�ٴy+�56ҡC�xr����T��|[6m�t�������m��5������k��̖��`ꨦ���g'1���Ç��ɓ'ٴ�d����V�-"�HyX=�m�&���"˜�onn���j���@��s��Ύ�&�)7�:�8'��=��-3�g�bw�O2E߫^�J��H��aA��4��.��Ur�����C���b������*<����1�_���lq4mc}3mٺ�CB��y�[k[7o���!z��YG�x"(�X��Z5-mYA7�~+����ګt��^Ӎ���-��](@�8J�9è�u4ܩIOJ8�M�u��ʬ��e@�m>O6�,��%�狷�>	��â+$�51����֪�
�~N��.w�%ǉ?q�$��������Do��&�w�=6�JԸ��{>����u�6PM]�h��F���ǹ�W_z�����$PkVo��v\K3� x����ssZ��<{���(�Yւ����{��J��<�܊�.p�{/l�\����-YRdQ�EJO�����%�������'�lى=r�(E�b[n咔�-܎��m�� nI�����w/�%&�3��`�ny����)�yw	[a:��)P����U����6�H������E�Ό]��Qn��(mk�P�����) 	�#kg;�'�ڀӥ�j�^����&CwŌ�P�\˥"(��-Dc\b���Gd�����]�.#�CAn�������=+�8�x�er��۬��ɇ|
rsx�n�W���%{<*o��M�>��a�-���݁�
�4^@�nx�:9]����WRR�;RY���|��7뫋��8=53m��Y댚�7#��a|?a�-�ײ.m��ښ�g{kD��7������(�9g���^mޡԃ���	Q#0��@%��;gHQƎ^M�ux�z�JOw��ݷ��y��_���{_�cf�7It�H9t���%�W&9�� mhj�k��`��kZy��#�������졆��+��o�ʮodd���������L�K���G�����U�L�֪V(X�y-����=iQаQ-	l9��ɼE�����+�ȥ̤�����fQ�cJA^.�������f��N�)UYUK�T�;�7��L���
52�z1�S��ZB�"2*����fݨ��{�ڗsgC@���
OF�(2�8�Hb"�R��jU
�^<��LKI[�e%���/z=�^(r"�y+�4S^V�<e)	"��P�}bt_h���-���0�ߑR$��t8����_l#�e�����0��h�2�=R�A���T\�6�]l���F����l��#��<o\���4n/��eFwj=����q���_����{�8��Q��LL�C~��C��8�J��*;C �Cr���ʺ�!���O��lhc-�ҷu���r�&Ϣ�<3a�1�ʕ��]�n,S1�s�e ����sޯ���LeAA��5������9m��#?;�O�[S��=;�l=kJ'�E]����3ȖچtXN	�ʽ@���r�b0�YZ	6��:Z���I @��������zRڐ�Q.��e��"�[Y� 0�wXQ�X,�>�8I u������YO�����ç#����( "ct1mQ��e �>���	�Z������$�0��NM[�(Z�E#�S��}��hDC`U��	���2�|$�q�T|]}�re岛�ka�a�@1ǳt]֖���5�aQ9�Z��ϗ����5>֏���6��?395U�3
@��,�̪�ES)X������ү�c?��.��z��z��l<��,k��e��k�d7��27&0(�̐��I ��� �k6���ðo�vٱ{�Ė�T��II}\-�Md
�Or�fqa�J�k�e�_��3j�V��բ���K�������5��O����D�H����H�ٖvw�}S�� y��4���@�g2`�bH��x.K
n��������xYCܶs��E��ypG�{��a�%=/e:��{:�d���I�������e���χ�O��a�>h�ځ�-�*�H �6�y;�e-�ֺ�v 2�
���5ClK�~MW�������c b��"0a��zL2��6��vxezn�y�����G�������4�����g*'�H��}F}YY�!7����~������E����ȩ`$�
��ZH�Qk���V��-�ެ�L���n=����z@�%�-���S ś�������V�y���7K���%;�@�=�4�u�Bl��4TD Zx~�4����c��@�u?�Un��:�� �/kۚ�v�ñ��*�=�{F)P�p������d���,%L�(J�ыi��ݥe�]�Q晦���[��#>��fF�iK�E�L�
\��E�ݿ_[:(��N5^�n4 ����t\)Sk���A��D�r����鷪SY������p���Z�p��b]+]o3D|�+�@���/�K%3�0�:�M=��e��>��A��5�P��<#�',��0}^Q���w@ZZ���X�)E�s���@���\�̡nvÔ=�;���������49F�t@�R��/FOH����&
������V������o�������vNe�O;P�(�&LB�*	V�*PЦeu,�[�c1)*-�=����f�!h� �T�'��AF�MV@(�cd� >BX�Ǚ��"�    IDAT����8��umd�d(jKv����[K��~�
��Le�^��̏>	P
���������\X���2��Ok��҃��"�F��B�U��t����r^��D��-�#Ci62(�Wg�	���3JV�9��EAұ�(�_nki�g�����U,
��7GO���V�>X)�@��ir��V%2]��<k����QW�B䏼�$�Y��c0��4�����'��W��1e��i�5��TZ|�J����ih����E�f�YR��sq��^Z����FR�2�I����[[~wC�9���߾��ԢX�C⻰(+V����\���E!�_+�M�EI	�o�E_����eZ@����jdh�$L4�с:d��JPh�[�#f��oZ@?���Ҋ
ٽ�Q��o���E�>P��y�K_\��K=T���G\�D�S咢������_8��R��&\�ԮߺU5<4t2uL!<�Yf���|�V�͢쁃�?�ͨ����p8S��A\�J� U"�.%�iA1�WT�q�"`39����'� *���pX-:J������H0�}�x�L������đ����+/����2�,b��1[%	�Hs &�R�1��J]m-�}}���Uy])���-m-�r����n޼Yyex�D8�����F-
@��j}��x�;T���h)�&14�����:@A���E�yL��������/@�l##A���"J��5~�>w}`}+��Y���J<�г�m@�VTq8���'�+	*�0��f��l	��"ifW,Uf���L(�pe�RRZX���t�~k=�x�����ъ�#� ���(�Ei�/(��
.�Fq
��钐��_����0�d.Y�?!Z�pp��A|�X�o�ii,A׵^6��q���[o���,'x��P��zL��F`�!�Sʫk�~<��H�c�2;?��܊��"��w����{T����2��	�9aT�O����m-�z�@]>
�{4�Xˢ�e?�4D��?$2|3?�֎��������{��\kk�#�� ����׿�v8&���H� ��j��O>-M����+�J&0`�4��t
@
@��ZzY�'a�HU]�<��Ӓ��O��/d��eT�P�q�
���a`?/,{bb����*��O�������!�����oܾy<mZ��3J-G���T�	iڊ�A���Ӌ��^N�3M#<�cz�g�����WV�W��U.��W_�����9iii�C����Ŀ��oS�;˃�� ��9ga�nCi����Y�|�nXH$9)�-��8����^`Pq�gU;� Y��A"o�]������Z7�:ohh�?x��ہ`��a@����(�nM�sHݟ~O'ӡ{Z����cX`�����
N*�k�K_��x��28�9Z��(H���c�����wI�.1FQٚ���3
[�qv�OR?����@	vWa Գ"='-�sr��e���}�%����A��H�ih0_��K
��^_k�mȢ ����ǂ����3
�F}
������&��ڬ�&({�4��C�t�Ǌ�x�;�Qijh�5��󶴵���EJ����z�c}�d�N������_s��|�E���V�@;���EA�������b����JR�.��W*'O��C/}��=�pf���{7���Il�R˾�¿�����j��c
�9�nP�����3J[jQv7��c�������'
� �a��������o�Ɨ�M/_����C����#~y��WY�C���!�޿{O�c���$
�
�	��Zڻ8m�ٮe|�uL:J����~�-��G��`Q����);PYnY��sSSӟm������{w߆EMbq����@a��(3˻*^�d�$;3I������\x�#3�nF����$&��%Y��O��Q�fcmї��2'�1�7e	�C��_X,u�524p���8��ʖ��\y��7���+J_\DJ����p�kvq�	36`0��b}��-�������() (������u�b�~��;��bC@���B
Su(�jx��D���3J-j���@���ޖ���;��%�0d̚=R�h��R�D$�A%7K�J��.(\��hm���"�4�"��!JC�/;/[�f&)y*47��k��5�4�@�4�/���M�~�9j (��T��V8}�$W�a$�珤'���MAX�(\�,�,V���fG}��T@����GP���}L��ي��]��2�)騅i���K����nnk���#0AJ2xv�Ch�VЭ�͝b��çf�4��\^Y� C��c/���$ ]������u
S����L��ŕf+^ON.}�0��L�0�[@ee����3j���C 
���U��@űl�,T��~�����n(D}�H�@M��f=� L@��ث�d��鹳�;���Q޹HQ���̿��,Aq6ڔ� ��u�t���������(591*j(�X�,���c��K@����9�8�ͅ�_Wo�<tX��IYBg[\��?~�3U�{�L���p"���ں:���r����/wԯ/]��b=5<W���-E?R��r�ݢ�g����ϥ��3\J:�]tX��U$2%��n1i�]8?;˺�G�.G��0ZyV��;/W�p*kʝn�� �z�$��$�|Q�ЪE�rs%�J(8�
8����"ٴe+wPE&�%73]x~ z����Ӏg�y�7��� &7��� ��H�U��_YWJ�c��s�x$�U�GH-������e��gZ��<{�`����%Ώ��"ini�,)������q����-lvz��$�P𐚀�Ƈ�+��1��,x�&>v���M@�fZ`q\�ͼ6��_7�ԙi��
�|�R\�=��e���d��F��N�;]��[o��:���?q���M���G�>�%sU~ߗ;��7*��o�=55��DҮO��̣֣4ۭ�nQ
ȋ�n.� $�U5���*y����߹yK��Sye*2IIj�,�P-��)�Z���h�Emݾ��Gu���G���b��4 ����9y���s�4�C�p��h��;��lZ�YLZ
Y�(��>�ԓ|۰( ��PH�	�35[Q��rWCͺ:H�(e�GG�M�L�R�p��+�c7h��je"�k&��0*\�2*
��R���9ҳ|X�ZZ*�uĮ,����!u=p�*�x�&\`;��O�D/&1�*�U\I^\���=���"/��� ����ClÃ��!P��M ��UU���%��l���I*����ky��I	C����q\��v�(��H�T��~���n�u���&''�"�S�Ɉ��M��[�H��7�LY'�����zIf�����2.r!���f ����G��T�k��5B��o�)C�|M�E�
5�v �C�S(hc x��ɚb�&�C����|�+_���R.]��!�"�� ����/]�ze˶�܏A���ɜ%E����c\_  m�����RL&�JE��FB2���3>]�/�\Gm�+�
\���[�"S�}��im�f�Z�LR�,;�'���=�[4��P���Vtf�

	R^aU�0*�_�+6���d3�P� �`�����;���L���	B�(���`-%i�Gw:�r[���g���Ξ��\')���D�쯨���wK�-�K�77?+�,@�3'[�|�����K�~�ި������ȣ��UHɤ产�J}/��խ���c��q���k��f�� �Z�Y
�@���n�Z`�[��V��LZ[�9����P���9dJ���99<�!�;35%c��� �F�Ά��zQ+��{=�Q�����3��SP}Fm�hy�_�]�J����ܼ}W��T���������W� 狍E��x���{���ef2�cO����/C�äP�2a�"�َHE��3�g7�G��Gn_{+�l!S���	7b�(d����<�
�s���@z��g�	1r6��P�.Q��{��0�>��)�+ԒE������	��F1 ���"]]=�/,B�1K����p�%Pv�ɑؒY҂a���Eʹ�?Q�]��Ko�f�[4�ofv�EY�({��	�h6�4�SO=�J��;w�J}>Ȋ<n�#RQ^�bgMͻ�K��+��F� ������В��hkk��c�	B0&@Б�)xJ����K���"k�ިѠM�Ca���*/�Pv��%{����\*���.(xi��m�t3���|t�28RC0��aSs�lٱ[ZZ�djn��8�S�,(7ai����z�j#�=�OH��4��`pT2��d���׺6�����n^�~,<9��(5����W(�������2��5�U���Zd��ZL�k�A�޵"���Z,I��� ݞU2:�SCs�*2"D�8ySЅ͛A�x|%��P9WY�d���d��G���S���xF��!�B�2?/GF������q~a��Î;(	k��Ch�{]�H��Ӹ��q�����g�(��(X���w��e��vW���Z���}P:A`�d�T�\`�`��b'��C�nBY��(1�},k���dҌ�X[�p������9Īv�{����f{ejf�d9�ܞ�}��-�?v��y$����0*�9^������������`u�z��ȴ�(�Ë�3��Bb�Q�6G&wB�B����^�ex٦�g����A��}
�@��i��l\�U�������<�a;!��(�b���%�A�>��u�2@u^\NHCs����'	T|�֘Z62A�����#�@�ڸ�HX��R�m�g��n>Jŗ��-P^Rp����܆Ψ����C�oá�Ȫq��+Pp} S��Ŵwy��=oJ��,��4/k�Eyqfֈ���,��kk_�R(��-�(�b ͍&B��|ߴ*�[�͕᠗X�4�P�!Pb�R��-m�u��mh��3g=0�jmE��כ��"�m��c֓��l\)�c�V��T��6Խ{�JFF����(\<]��@iԧ	�=,�[�Z�O#3uc�|�n���왂���ʏ�<�pb(Z���u�˻3˾��B������<������
G?�Nތ����8���/�e+	�k��ݲm�^�������-�0{d˲,��48�N����c��H+P�9�@���Hku��Y��9iQx�@+2��z	�Z�z@�LA ���bi�.��y�sv  ��pT.�:�����	uCT��:�)���d�@��L0�A^���Ys��	�{_ff�������6|g�fٶk/��0{[�5��Z;Q�e-Z$�Y&QG�$�^�Sr�\�ʲ�#-UUl(�Qw��M[�d��(XJHƊ��Y�zn�5���֒~ pQ����;����r	��-�dg��r���;8�N�tv�����(��u�h�#�3U�l���NҾ��>h ���Sg^�Y_�w����E,�(� �1P44q�Bg7�;��!ms�A��I�F�+�\��������&��%$���
rP���TfNeoq��,e�\!��J�w�'�ɇ��%�Y0Z�c�n��w�.�zM�	��fg�sG����n�wﾜ}�=�I�YnN+(�F�g-qk�f���o�-�H��y�1T�S)�ۺC6o�%��<���K�on��g-E�X�iz�(�$�t}^���������*+�!�P��7ߚ��k}v�L]�tQ����4�S+�y��$x]� ˲ઐH�̚j����H��	����-)N�׌�@���/|�7���I^}�u�L�M�*<�v���jy^�SxR4.?�(���gNK`|�{<8�Z�w��<ota��Ǡ��>J���
m�� �sz]�k4�T���"�~����o`t���@ }Fiԧ��p�M�|�~�z�R��)��/���y��/ 855�(����PS^X0�s؎6�m���E���P���xd%��C�����;6F��ё[FY�e�S���%&5+���E2Lߦ9�曔���&#���`�CJ6�DAv;E���*PL�S���Cp��)e���N2侳���lϧs}�������cぉ�L (]A���P̝�i{ۭ0Y]�=4W�V`��4�uʑ�/е�Ѫ[Dq��4Gށ�C3��P  ׮\���W%?/��&$�r�_�>ڶ}���ԚV�̼LN�>���3��b������'����~A"��_P ���{����)��� S�:8���Ԓ��w��A�����QB^�0����l8���(�=8�v0��a���B����8�(F|��^]�gMX
��Yj_���7��Zۺ��_���:uF�9{V���[JC��q��\XX`��G�em���{�u�KV�����PO���E���0���O#Jp����|}��$����ߗ嘑H�ېX��lߵW����B H���Q�9�H��d�7�u��S��~E�셮�� ;�:�~��3
@�:�6(��)P(f�z,1�t��E�"Q�*�
/Hkk��#ϑ����J J�F�*  �p�b���g?�Yٳg�D�f�?}�/d)����EX���� n��\NS��ԑ+�P� f\k��z!F�+����P��S�f��@���Ԧ-�I�P)��-M%X)�Y�R�7�j�Z3,'h!�`�y^�;\U�{n�����D������px��Ҫ,�P�(�r{��T$JW>�ժ����"\%�Cb%іm[�f`p��,����h���Zq�3�>EJ��Ę��_�'�3�HV��h���y��
y�JZ#�Ѫ���"o���YbSh��C̵掔�4�͑�{v˦�ۨ���������bg�WNC�y.S�uqފ󻜍JHa~��|�X�� *��I��<(W��p�T'�~N\ �8 �RUU�u��41`�� b�䊯���jf� `���o��ی�*�"TLȹ��b�Zj��=* y��A�[[S�ј��9^�+�o�޹��w��C�+�"sSLtA���	Ւ�����xܜ�� ���e��� +R^����,�2~@�Ba����*�N�4KU�Q�m?������\�p��:���5�ո9X/�~]ÿ��.C�K^��b��c-��� ������W0G�f��m��� �%�,�X��#Pyd�>y���αC�������͓m{���h��G E��07�� ��Flw-
�l��x-خ�<
Բ��|����"���Zkj���5T�<1t�� P�Q�C��h����'
��E$����R)*)�PZ�3-������Q�6�s���_Q)AU�����yuu� U��>4eA�F�?>v�y��/z�����@.���d� �o��c�>5;�H���1:Ùd��C 
����O���0݈-�Kia1��,	W���o��`�{3��=0pb"�2Q�"�n�<�G�&Ʌ�-�R���ř�;gZ��[ �լ9_���0RC�\ϷV{�B�Fq8����
���?���wt�e4|s�b)���hre���y��m�8+_8��|���\�]�̥Ɛ���K8L����ճYf�Q�r�)�f��n�Q0V��o������Iݶu�4�4Iqa�'��\��<O�_Rvt�Q�8;LԷ`*����Q����^�����	e�k]��cX��`���Y\���E���@T���fq�+���H��u����{���30��e���L��1���bp���=�|�{.��G�z�sz����!P�k8��.6`�#�+��K�6Er�k���7n�և݉�]\w���<YY^��,+�x��V(Tugp��xp��X�F}���ϛ�:f�(��t�F�ݑ4c����=�C�U����\�_���\�O���踳%k���ŝ@m�^ *X����'���S�͠�0��N�cXȜO<�T�VqI��x����?��\�t��EXJ+��8�
v�? }[vHpr�c�J	�fm�Hd�a��)G�(УmߺE�+��(_Q�xu��Hcy���Qw�ܩ�u�Ι�P��Ttބ�
\�����	����Lf�~��$)�8    IDATš�`L�� �msT�n`aSԻ���;
�TXI
%��o�}Z ������ `ൠ
���,_�¯��91�����O~�CĪ�[��C���WJ�6�m����|���`�D���r�T��dRx�N�X<~ks��l�/��ؐ����l"��,?�T^�ᆀ�w�^��3��d�bN�M7�2��%��n����Z��In��L%�+j��G8;444�7cH���P]M�}T�Q���A~�Y)USF9�0M;��K�!��h>v� �n��pp޳����::�����{��O~"�FG�;H~���S�/������-��#�-{��I������
N�,l=�Y���ae��y�g�.)+.2��,�(�<�V�A���~��͡3�P���V��@i�g'�ث�{�<��оOĩ�7~��\�p��;�6��ˮ�;�_YA(�%���ϝ;'C��@h��(�p�I�Rτ��f�ۘ<��oȥ?d�z,}/�Ě:T.j؏��ϞyG�߽��S�W���Rv��/=}���R=���"��z�da~�����d�歴X�X@�����V���$S67�1^YV���;� j`t�@0�`�2Q�2y�YA�Us͡�۫�.]B�	��0:N����.������9yJ�|����?(G���7n���Qz�x���Y�����S�ddhP���t_aQ\�lf9��%���s�H
B;��2�ʬMlx�ȥp�aJ7A���|d�*�������ahj�HZ�и�I1:�˩o��� ;��v�`2�t7*)��#̷|�E�\�k����R�F�Q#cc�����N�uv�pX�*P�����M���"kщ���X�T[O�|��_�S�NqSeE7�����o}��w9�q�.������^�������I88A�=�	�Qpi။Fp�뀸1'א:�iE�ADMN�T�Q�Zт���� ^+,j��Ǥ�{�"�t}+�1������ܴ���?�_w�&iln���M�� �be"pO|B
�s$?������XQ���wl�����P�g,�0���^���keB�%X�(ܥ}�wɑ_$m
+�:�k��ϯ��
S|�B�`���Ȃ���/șǸ�"�����{��5���X)�(�#A��~�A61I���p����9�EU˞�KGO����\���TAA�,��ɅȽ;wd�N#��$\�e{I#�{�4��IU�_��}�J_�g+J��P0q;p�yx`�P8\�ʶZ$ʹ(����������-.-KmS�|�o�,9ٹ�*ʥ��G~���������&\���XL��oв�(���~��|@q�	�C��u�V6����͛�=@p�t���//�d�7�` Q(jx�q����*+e��sS���,�U��y�߸��}}-�4��Xu�f�8�-h�����$~�:[���|G��uW�2�\Żw���	�C����o��0Ns�FE����빅�N'�V�Z�u��an�O}�qijj�G0��2m#7G�՟���	bfuu#6tb�X�z��9�ĩT�9�.��5�Tt;H\�zc�r�樄C!VP���:����?� ^+'>����چٽ�i��$�I�ڞ%wnޤ��D(��5��঑
��ȩ�7����)+)���w;���~�6��u�֭����S�ɩr>u���Cr�m�Z�a���H�%�N	;� ���Kk{��Ta"zz�L_�u� ]kS�<s�9vTѱ���9��?�����at�K�r,�͓O?-=�����D��9	r	�	�\�t��#]^s>��@����ܹ5��Z�BLj��o�ili%k@�����r��-ijm�;w�}b%����@����3�A`|\�+1�nn��ly���r�%_j��H���ᓑ��RXSz�ׂ��PTiV�����A��5��̥�DHY�&�����zGy����E9��g�<��!~}��y�1(��rA[��;�^.+���|��+W�1�N���Y�x�q����]��ҕ�W�0lh2���[������ ����iÎ=����E�IS�:}�ܹ}�����'I�FΉ�_���{�|�d|�.�0��	i�*��j}���z�%_jtt��x���E��Y�>p���,�����ڴ���f/#��
���NV�$��*ܑ��(�͊|��b_	���dDV��e1�B;@���deK{G���o|��̉���p��#ee<�0��y��E�x�"��aN�^��~�ZFpY� ZTt�:�<��4�u�x $���ٳ<׶�������qZ���	�.g��b<��<3H��hhSK����R5���0�� *<9�S�؏�Y,+(=��%#��^��l�����\�1���p\L
�2ca�B,��[ha S2:�;+�5om됯|�k<���:���������]�7�Hum=���E����[�������������{�il�_~p^N�9M�
EKLj���B��U��QV�(rC�aXa6*��J_�P{Ká��5x������d��\��
�b����Y[��*�ԯ4�t8L7j�:Ȇ����F@���Am���ጢބK�kk��|Ub++,�|���Z���*Gb��VX�SO?�@�
��?��?��H���ˉ���l��g���������{?�%	��	_RV����a0%f��r�QT��ըP+��T�u�6>Y��m��m�:��.�[��D@d�3�^-רO�I-I�R"@����(�o�5�G���F6>�t�0<>����2�?����#���cǎIt���w���n߱��sQn�ELG��O��
YlE��?��J�=�0 ��_�gq�<r��!VM�Zp�rr���K�RzL����D
C干8?#���C]����G����S3��
�[�e��� ����EeZ�^���jYhw#�@�;� g���2qE�A�0&�(�2�@n�k#ΫP�����ԉ�.���^cЀ��
z|�A
FD[�:��b?��閟��U������N'w˶�R[�(�Ȕ�>��y�E�TX>@`ڂ=���\���
^�Kǰ>�͞��������ΖC����6tF��>8�����В�~�����=���~>eZ����%fg���i�#7_�	B�>β��A>H�r�
�^M%4�j	�#�M���!9\SL@S�,��z%%2=��a����a��x�Ɠ�&x|��Tc	�G�H[[o�Ĝ��� w����z�ݍ������B�Q�Q���m(L_��oi�!�FL�N[]��wg�q�߰��
.\���ץ �粶�"�s��e}��s�5g�Q���g3��ԩ78<Z���Q��z��Uâ�5n��ɐ��]omkz���"�a��q��=�˴({�k���YT&P� �U��oD���j26��;�z��G�]�pik$�� 0�3q%��ʚzV�Z����B� aQ���5�M�u .�p8H P%W75����6��|����~}�xdj� �ή�g�6���Mz�2AZ���)���?��<<�R�@�-,}g��;ݸfk����3����]����p<��%*U�uһu��44K����A:�0o�@i�o,ɸ`�$��
�ZTEI����'jkk#������oG����@��iW7Ӓ>)P��j�⾖E=�� ӿ����E^(�樿��H����k�X�����w뎝�m�>�����D�L^�ֵFTY���0�X���� 9Z�&��y�3����ÞƚCuuu������ ő[0����(�?���~�vwg?sp��_k�`) z׃�oR�x5��5iU�������{dˎ]RX\&���K�}���;P�� ��Y\���QF
�ƥ�����}���xjC@]�qc��@����t�Z���iH���|qi��n\��A�k�<
�
�j[E�@��*�{�$��p�(Q{U.,��9$�n7��[w�ޭ�%��'�&&���H.�:i��Z-�U+�E_ 
`*Y@}о��p�Ϸ�^�d�x�����oMNN�jԧg����^�P+[�"?{��߳4a���
�=3ߋ+�e+;P���Ԋ�Q!��\F���x��l�I�iM}�wH^��,$j�fg�ԉ�����Ʀ��IL"�U��|�	�IMy���-Ow��s���/?:04����lF4�}��2a�J$VV��L�ʼ��ї��x�z�<��V�s�4��h%@k��$�z ��Z�hf�l[۬�aV5Y��<��<��(�Ba ��'Q�[n��0��N��@$�@q�ōҳ&�xl3�aH������줔�������Ɓ�t����૑�lUm��8=��,�J�Q偮�U�P+�_3�Z/�=�6����C�K�4- P��G�*����8s���&�CY'��C�L�e�r�����+Yy�M�P�� �SL�R��]o�)E�:am,��:����lOy���,�����,<5����ڲ(��Tf��\�Uژ����J�����@፻�%����v��?2U�zt��Ja7;Ba[��T���K���I4J����ĕ�%P l�`,�<y�&�wg�he/�Ō��@	����̶���*++�]���3�W.�������\�Z�C�X�&�j=v[�z���[�������E۵��fhړ�{f�v�UeX�I�(�5+P�T,��ֽ��nr�~�	�a�#���E�����p�y�%��5��犥2OE3j�E�G����u����^wY�C�:w�Ҷ�7����g�\�r%���B}sF�^p�E٭G/����H�>C���+���AK�<ܹ����j���BkrLL�cJ���F�Z�8e,
@=��$]�LͲH�V��y�J�Qu9)P���f�a�'q^a.+K��ߗ�Jߙ=�z6nQ�._�q�ک���
V���n�L���)P�d�<���{kY����5���aoz���y��UC��)MY]�~F�D�����HDײ(LÃ�	���/JK{�R�/,��m�P�$g�.-�܇�FC����V|�b�k��*0q_���ۿ����KC�j�_8��nʴ(r&��6��-J�Rקo>���s.���̝�g��)PjQ�~k�J[�>9 a��VA`�&i�I���~�>�3j��3��
��� X�|���p�+8�x^�X�[@-�4U�C�fg�b��/�p��iS7�n@)`�rK(0.��eg��v?�a�w��5ߵ��7���N�Y��T1`|P�hJ]�'���P����!km�����Ɏ];�4�� ���6
܂�f	�Vr���ek�(�K�+d��K����9��l��|���WT$�SS���������҂��6��TTPH�r��ĸ4�՞���r���i�=�=����������������eS�����x\l(`j�d/������y��qm��o����BR��_{ԧ�� +������ ��B��r��	NU�t�ɇ��;�ns��P�2�5�K
@E���qF�7�0\W�MD{)*,��B�v�*��8"j목l����"��m������dD���^אָ}���m�=�
?<�Ω�]�|�ggg�`M����C��0�L��氃�@�f}��7��c�P�\k�o�<
9��.@tu?��_��Ǐ�����jK|�_� ����彳�����S��I(1�� \zQv������IM}��0�a��aQ�� /_���<~BbKfΪ���cC��^&��$�-���N:d���RS��Oԕ+W��?�'�H�U�p혪�FzvK�,�>V[� ����0�JT�wW����І#�[X@������ӟ�L��8N�BK����}�n�֋��S�a�&�Hz���ʕ��-C<��g_8*�-\>���
Ɔ��Hx" ?�����v2������y�N����HwW��.��)���~sU��ܰ�Í-��x��޾}�+�#tc,�:zԪ3wcf���y�r�Š��V��`o��o4�H[�͢��=|�PL5�	�8���K����t1U�� @�]\4=C �+F��T*L��ׇ�C�t� �pz�����V�_%�|	rG�6	�L'O��C�?F����H=�f&)�����3����U���ǚR���T@�ͽ��>;<2��'&&�`U�O[�*��	�=�S�Ҳ��Mj�T�{{��� �s0�+qa�P�T����������s���B�r���_���p� ���h�Y�`�0"+�;$_�:7���*��B��F!�**̗٩iy����O6),.d�{��IY�EyF�5��p7��e�ꪫ�Ş-��?��jT�uN<�z���ҥ����¡�B�����Y[��v����<H�j\h��tX�[5%��P+�`B]�!�F׷��	E����",Go(�aP�G��ò`Qh�An ;5���ܥk��~-��(�8=r��	Tt�,����$�b4*�f�؛oq��(��~����I��BCm=\n���^c]�o���>�>�o�����o����;�~ofzj��| S���VE�֬�i�i]	*��Q����u�,�8�U�s�ǀٶ0��m�v�~�]�Bs/�J�
�h�����^\THkBB#�큵���:!U:�rgɑϼ �-i���܁���̬?��LOF�}��&��6غ(q!�(��D4�0=��P��������zx�c�>��ɓ�ᛟ��_Dv�\.f��w�Cֳ({�OUk�� >"j�Eŝ�dK�wH�W���۫��r�A"%�-J|E�p����ok ��H�3S�4h��<����Y=�^8����[@a���#G�����),N��!ˋ	���w��bt^z�,Dv���^�v� �Yh"لTW������>�y�C�8�OdQ����/�Ö�Wn��Rl�ɂ��\\�H(L^6\� S<M'�ܭaH ��m4W�m�)����]�!jLj`���J�H{Z��)Ћ1�c���
�7yy�ᗒ��<.?с6<'vq`G#�A*P��>�ꩃt�ׯz�3�M��E\�Tlnyo ��a3����<� Φ.S��ϱ�Ji9��y��������@O�Ci�v��+�?��w��r����w9���E)Ƅ���:�a�@,H��J��!�/���vKO�&�z(�@n`��(=�G���<r�T��>k'�i�ItaY˳�Kpt�v������D0XÀ��\�혶��8��x/ǩ��+)�]��S�;Ρ9S$΂vl*��`�2��wt�K��&�f)LpB|%%`�N�+��j�o��n��q�ҧ
����7r����נޙJ%i0�k�<�е=�c�L\�[�O�r�1�E%<r�B`N����Y��@�	yݔ5��Z�(�x]��fo��k��<�5n�+�6aC)��px���Cf��c:Th-A����^���-yy�
J1|�X��(�����kWHU�JE�rP]R_S{����O��k�|wW�C�ak�+[��A^y������E"�����y�yE8����C�8#���=+.5�r������3�/���r%t ԝ[79��ݿP4�gmo0?�U*3��q� ����� &
�ǉQ���	���3�<<��Ό��<� (xlݾs��Xv�ձ�Ȥ��!�ò/F�^�E*��'�[�������*V��-�� ����]�_�����mrj汢¢���B_vvv�I^��������p�y��U\�p �䙘�ƹ�0wK_-g	���B��t9..�[�-(���"4�!���-�7o6�a�K1��EDVTR�h�W\�H��~�`B��x�x] �o�f)*)������S�[W(���Ay�ź����//��3��=���q ~*��|�����i����ڕHĻ�W[n~���v�Tg���dH�S�g�y9bc�����a���ZB����i�Ғb9s��U��A�-��3�4�5��"�}��\�g��k_{���;�OтՍ�U�|k׮=����a�PdR�>��Pr}n�w�����_z��W�jCc݉�;v<���q m(������|�
����������cK+�T��p8
�Ng6[�n�d��H)��$b  �IDAThn2�+	\N�4D���XX��!��C���~eC�*A1:��S"���C*��C2��.Z[ss#����Q,�-	�q--m<���R��8$>U��w����ryyٛU����[[�﫫[�������T�Z�	���ogMLL����
}х�X,֜H&�R�?+++�������э��/�����\	��v\>C�o���Ӑ���DXr��Rg����X��H��M���J�j���������A^T��Ņ�x<>���	�r�������T�/o�����)}@�����@e>1δs���ދD|���u�h�=+?wwnN~���N��e�D"_RN���t���{���\�"ٛB%�	Ij�$�_R�t1G�K ���_F+0x ���c�A#ѥ��幙ٕh4K�R�n�{���x";'g��� ��Wp����BNI�xuNs���w<���i���ۿr��z��JN(�L�-���V/,,6/,D�cK�x<^�_)L�$��T������qa�֙r&qW2�p�ەr�=�DBQx.�����^��$S�x<���W �rNV����ʲ��X��=�YY�hvV�LQqa���?\����g����<hfr�7}�� ���;������zV�a��Ғ7���H"�]L$�R���T*�r���d2�t�xa�qg
����7��$�w�r~�;���/Ap�Jd����"�k��PM��_����@��^�?�H����8�    IEND�B`�PK   F�X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   ﴣXSW'� �� /   images/aa6b1763-b16b-40d4-b079-865cc7d3b61a.pngl�UPLԭ�kpwwwwgp��������%�NpIp9�wq���sջzWWwW={�ԊQW�GC&B���B*�hBA��AAAK#���c�ZL�_�)/U?C�
�
(#��m|ѫ�h��A�6#��/IӃ���U�B�V�ENDL�PHRI��IJ
�p A�Z���d}4��z=I���xű*���s)�	�B3���~�|�y��4~��a����~�+A��k���Zׯ��Q;S�3SDb����!����E�8x����L��L:�EI��Wn��88�������X
����$�0���$H��X���~��P�K\�l�x�wKK#�MY��V���kr���%F�h"�:>9Y�+���%��
���^}ڌ0p�����h����oJX�г�[o5S
Q
ߌG�c����E��ũ����g��b�l�8��Z�=&"�i�������?�vN�<9B�?������`�7Q��;��(M�������`cC�`�b�9̱��%����t��H�V�*z;`�FHT�Ί�}�!�0�kvާc>�Oc����6'�+:�t���V_��}��|@Nw�EXsoU�ڳ���z�~[�zO�[�h��"��^~u�fEZ�L��y��?�����~d��R�Q\c2�ԡw?��]l�?%����S~Oj"B��mX�k�23�J�| kRȈ�VFj�ń^�f^���ΐy��DѨF��֖�	5�N�|�z�!��
�����Ì������5��C[���R��ي���8�ee��P�U�IvN�+~���Qk��S���?��_��>o��s��׶���
X�w	}�立�%�;CӾ��$�L�WlF�@���R�������/�5t���)�fh�P����E咢����m"�@"��3!Q��N���׳	S��$�}�M��V�ÎX�2򘭮��R���9�F�r,��Iś�"Í�>�cj���/_l8C� ��Ř�%��}S�����W��r�M��bD}?K�Ӗ�o��g~G�u"I��xI�E)��º9�8�=ڭ�<_��d��1�����M;z/����
r�����%��*������*(�_FՊ�_��_�n�&Y�-C/3ۤI�񼈬���(�a�E���\��8Ce��˜̦#D��{M� �m!	�䓇F�,�B �036��
�7���qzA�RBW��>Z�ڃ�O_u�_X�����?����|�a�)�	E;[� �+�p��~e���o�1�KLcs �Zu(��]f"Ƅ������4� �Y��{�B~c��Ｍ�Z�1Յ�1 �F�\�4������t����"�I*�a��A�>��YC����;��`�����~b�0A4|���&{�n����,�Z��R�7�K��;pzS���7y�d|�z��8/��?�j��[Pffc���������{Vc���n֢�2N#��Q;T��I�f�&\
C���X��̮/�
�GS��g�hA��'Y=�Gk���k�5�3	���~�X��k2��-��qL�V��ĮbܲN�T�BZ=����no�w5.���B"K��?�*��N���R�ᬐ栎�t�Pg�x̱_ڛ�V��4�������H9l"���BI�p��Q;��:��iy��6X �k���d֒���%�� �F�(��=hM�|T&*wk��=�L�JÝ[�M{ۤ~��D��ŉ&�*k�,ai��k�a,�Wa�H�8���.ˣ��y�Or�M[r��h}wuE����xk�#I�r9#B��oF�"�Y(����k�f��(�_�����,�v(�3�k��a�nQ*�nB^�'Z�f����=vZhx���2S��n!D���y:%�^�^�xcm�KN��Î�!%��rU�m�-���R���/'S�2~Y�2�� ���wR��6��;�N�←���%�����4&P�����K���Ld�,$�C�I)d���a5B����P� U�H<��c��Mu�[�QQH�w��,��;���ڹ1�{��}%���&�����Xe8�'�F�=��x^+E4����D�I���RZ�R����'����(����'YC"R`�MB{�-:�~#�ے?�Q����]�"�"�\��n��{�?���\�.�3�`©�]���6� ���YB#8�����C㦐�z�m��n���7��0a��}(��K[��k�d剓'Tm��鞇���W`���<7�?o[3�%���D+[�G�3N��C�������D�6�;ڱh%�������Kĉ���T���|��CA��~Q6��f^"(�x�F&y��)�����O;�w�7d1X�=�{���,=g��".G����j͠љ�'�$�ފ�X���p�̌[5Ҕ�)�E�'�E�S�uʵ�����I����98�ja+���zw���jޕK3�t|�̝����	��������f�$���W��w	�ۣY�����	�jj��5�ⵢ�h�3h���e�&,l�ҔЈG�~k�����K�u$�p� �9�P*����pGd�Z3��&���d*�EL��RY���Wg��a߫�^���
R���y~�%O�̆�gS�7�l䶸�:�Y�c���a��b�*E3��hlr҉$�+ؗ�r�n�sT?��+i�1�+�Y��XΒ;YBR�Aa�h��H�g��mC1)������M�&����C���a���R�@|�g9_��9��j�k��A}~�3jh𮐥�+c�J�WV�wNM8r�}ɺ�&^&�0W���Z�b-���"�����8mu��U�s]£�6��	o���/��c�V��"�IJvB�~
F��w�S0�吻W|1���V��vt���,�nh�+{
�<4x6��Lq��X�#�\cf	D~��%����`�JI�M�6���@Bk�04�{������Q�����#���a�}�zh��e�L�7���E�S��mv�`��@���.���Y	�M8�*wW�aNp]�9R1a�s�}��p<���glpa�]�<��lz\y��)hX$����!0c3�翽�s���8Ni;�4Q�C�x���6�-�|����NC���n�Iڀ�a��/?�N�'��bRTd\Ԭ��b� {1rw�����̣�4��0����7�~k��T.�_��R�� *��.�������!���$s�o,N)�;��9��!e��E;FN��t��	��%�M�N�����=>���Y����#��'B8�r ��$eR�&�\��dvH��}�"pSUq�{H�G��6�cNʰ̹*��>s�3��A����E}�/��B������_���Hn.+KvaS��n��=3�`#/s���B0����UM���-� ��\4e�SxU9�c���fbd+�ۓ�� ;��ØN/6��3}d��v.���Bd�p�ތ�Φ����#��	�f9���{���6OEk\��u!�%�~�W��xCg���?�@� �����6��|'���[�.���B&��[�Wł�=[B�FQo���zX�hkS�$>'�3u>�fSMs�Z!I�l{h����F])��%�9j8������]/��9�|���RgD&�X���6��Z�񏝄ó�^M���Z�m��=�9�)7m�pd)�T�|{�������a���j0�D���D�؂���w� 3�c0<��;���Q�V��yK���;�nq�0�^����Ժ������T[[_Z��N�yd[�xJ�5�F�u����w�7?�4A�A��m����Y��~u@8ujAK^j��
I���곖z��:��h�O���Yl��3J/���$7��`�AG*�2�	���)3*܆�uf��6��rU����rt3$Rs�)�:�"�"[)�\�m����w	u �VIks}������2��cL_�y�����ׇa�G�Rq_]0�����Xة:��a���@�t��]L�f�hCZy(t�(��R{��s�����u-ղ�1fτ�ϸŹ��ݯ���Q�t1>uѕ4��<LO�`�.$��j9��<�� nlF�cN� ��f����Uab �|щ�K��1{��G��5��W+����Ρ�@Ld�0�b�I9}��A�4��_��r���Zzo��+n��@�k�\�yb����$�e�1�022��S߳��iZ\�j���Z3���;�4���2��̓ab�M��J�ߔK�0�G��=��+�<�(S�f��d�������fA�&~�u��Q����B�}v��U��\U��a����'�R�=�ٱ��Vv���~����H���Is�0y���{�Ϣ��ҧ4��Y� t����A�!��S44)l��5+0~�G�Y��%rM����5oQJ��=b/{�ȃ��K�Z�1�V�Kܙ�QP)BV\��,��A�$iU� *�>$g��FX�H:K�"�Z��W5�I��7���J:�J<�ׂL g�Dm�>@R�� �κ�d&�
cH}ʴ�>��p���S�gڂX�
���)q�5ɘ{���V�
;^?z�p�dȍ+�B%�f��[\��"I��r��U��~~���pZ��𡃣�̈́7Ʈ�s�.�m~B��e�`a��D%ʡ�t)x���@����&`e\_i��b�h��%y�&�\t�W!���i޿w��XɱM�[�,�:*~���ԠJ��]`,ݱ����w���	�LmUΘ��~3�k�vΕ:���@���f���Ƌ��9� I���m(j�%e|&%�&���N6��x\:L��b�
ِ�%��j���Ά"�ڒ�U<Jf��/�U�q������{�=�r�J+�Fs�dڍ��7�O����4��U4�(4��!uvZ�1��cf�?���˾�v!�=��|P�]�"�삿z��|�9���N3i�Dh�S��~qz�h����m����1����\�i_lo_h��6Dih�i}��h���9/)�=il��n7���%^��A��y�� 2Bo&�y�L/�To\+\;/ƃ�6r�� ��%%�I�gQ�6���V��/=�]�_k�	�S3�m�.��@����`�}|�|�
��N#��ɏ�8�t��a�B&y�"I=4�"A��H�{�?�Aa��yy���!ww��3���M6�Z�_������M"=�/�����σ�JK`��Q����m;|���pCoZV�:���5,��=��oH�2T#�T���yߝ�j�y�Y�K���nej1�߰Ca�Whb�INN��G��Ԣ�g�䙋b�O�N�7m�')`����,��f3&K�M��*g2��4�5�)rfa�S�I �?f(e��xF�
w�B��p���H�Z�TV�	%�#��8f���.���.��2c�i�dĴq)���A���v�Β
f.-@�n�VVTgs9�0F�$����NC�,�i�i�z}j	�FJ)L����=u�A�D�HP܀XW�+���~�E�,�8������Z��"j�l�mb��mÈ6��8iBB���P*�(Ɛ9[׃� Xf�����/֛3��(F6��"�P��u�z�F:m�I��#-��G�t�8>-�@���tYm����*W��W�s
;Ά"V$�R�/��Qߚ���B�.����Bqb���[�Ё��A�<�{�7"'ec��^S��e�'�-�ӂ��>�|�}�����Y�k����CHi��4t\|����98�\�A{`�V��I�_��u�ftR���a�~�YH�VfVB���U�o���StLc��p�!)hz���l�L��&����'|M���ÔcsRRPaUB㰒�ȏI�-�|�?)�_c��#��c��s(��=/B��o�J%���ߓ]���Un尺�M�8��F��u�:�y��l
�ˉ�������BϤhEݻ�&�~˂��H�n���.�b��y�|��u�\͵���|%�1Ie	s-�û��3	\�]ji�3����lYmCj��Y"�Nܐ�������05�2[z���d2����������ud��	��M"x\��A���ߕ�DH+fIU���hd9a���K(n�f�1��i��gS�(X�Ť�0�np����Z5�8&�
<�`}4���~S���fI=����qe9H�Gev�6�Z�r"����t�"{���?oЍ�2gf��v���nP�6Z��t�ۏNg�`s��:\��l�L����wC�C*�`���F��	�f�t�T�H�Lu��jn3�zn�Ʒ�����`�4X��g������D� D��3`�;BPtyotezNmɅ��&I��_2��54�"���7���[�\F=����b�E�V�\�-�(E��I1����6��(7�1V/c�v��pCh���vR�qES�d��3=8R!�;1����Y��,��M{�E�Č�M.

�����yM�Ie�>NN"����q�C�v
5��0�����㮏���W�Pe3��|�;�?����9+��Q��Pʄ�*T?n~Ǩ�����d�Q�)��*���D��GZ�.��5hSZ��n���&@*e�[��x>��׉HɌ��FK���J��AJl-�R�����Q�-j�bI���6�<�0dP�B�mς#�*���O=��������e����y,C���s��e� �L�^V��&��pH��-�pad�   7��� ��iDc���rT�����z�A���@@�-���$�>�����iE��k�{ѿ���'P;�r6�	pK�.��n��oD|�� :�`�Q���Y�J~K���8TھAl1)t�#�ly6QK�C�y"��T�&aH�9�Ѳ��b�	-�;0���k�e��&ymlA���Ie�Q�owQ�?`ې`�2Y���]���ar+Dy��;��\c9�Fi28��ڌz|����^�@:�Y����4��iM��(�9�m�"@�7� ����@%t�G�9���U7lff�(N�M�IWI/��Cnn��	�cqn�&nX4x{{�M�6�S�Bb���S�5�&�DO*��he���x�AB~~&��M�K�:�Ai9{�h��LP+r2�]��*��e�����F?~�<��ӎS��-�噕e��9L>����O��e��K�t��5�7O-Ql��L㌔k=}��7[�F
_��\�[����6D2?Y<'�t+{7�`�YP���'�H������v��d'���h�M-��=�L�_�/�ύ�U&m�2���Tg2�LZ`��U��@%�p���Ґ] ��uOpN~��v�R�aVxp��a�W�!���}�"�B�W��LR�.��A'�Mf������id(����.�K�»��i��$i�U��h�ha�M:�qI(R�����Va�w�6>�[
��7��7��l��"��B�'�.���a@B���D�ǣS����jR��أ���a�_D�BH���(�Tj�\W1 �2��u�h��Tz�Bжb<���
S�r#�!h�7)�8�c�on2��b=�x_AV>���4�m�Qg�fhɠy�Nu:˫4�V��ڑ/�;��6�T�6�V�~Þ`�����$7�l`~�ռ�n��g��۠���M�y�}x�|�0Վx'g��I@���W�[n���D���$�� E�X��D����"������N�Jx�쁫��������Iv(?��v��ϣ����ɘ����1<�JDI�h���=�n�(�伡/��m�~Ԟ�4ȮID�bSB�jK3�ھ;�ܮ#�����v�rbG�)؄��t��hcM����jklp����~��ݰ�Q�T���No)���J�V$�~Hm�08��Ԥ�q�BT����Υ��R���c^��h��MoqEC����KBm�䐛7�� ��u3���H���W�H�Y߭�������=&>�(r>n��?v¼v�|_֜ͽ��c�H�a�*p-�"DA<�d��:}G���2��!�\@��^��ˡR7U��̟m�Qe��m�1�)C�@5,@`}#�Ph�f��y���-z^�Dj	���q��Z'�H1���s	�S!��ON*�bBw���?| �t�
+CV��y��̊�P��pK�)��,$�a9�øh����_3(���$�JbH��r�CxoL������4d�Z|���#��X5#M��F7�t�Q�m��!S��ā�q��,�KD����Y���	��8� Ed�S:eY��P�Ӎ�8h(�'�x� �����꼶�S��
|җ��%�<��:Br�3[}IG�U,�k�&Q_���h��y]��hY���U�g3�!3^�H������ֿ��ac�<LR�0|rp�#R�e�����9��N��\�����������ߏ��gr��n�3�E�i}�|�C5j~��ְۏ!704A��]���k�����?oS
+�/�	�	T֣��A�;�$}����������Jǹ����v�(Kڛ"n��5.�[�.���������F�,'@=R�;#�qFK�#E�>�}�� .�KmM�ЏZ�����}��_H����O.3���u3-�曏��:l\~������zm���V�7l8\p���V�xO(A��S`s("��k�+��B�%��D*�%x4�i��rbw��4'�sE������|��`��?>�C�5��������1�.��u�&�`�.�<�▶Ɉ#��@)�P��4�~8$��r��6J�ڗ�QЏ�.'_�i�t�`��z�jkb����B�'�F�b��$,��3��ŪuhA�%��X^����d>��_��fh0����-��O�<&`�����t���|�H2�(���0i�]�k_?-ġ��ü;\�WW�5N�J����I<rm�+}j]{]\�g�P�yF��̷i��2�����)r�˜1���Q(�O�+��씜2�ճY'�2�7�1�E���֬��\[���t��5���.�,ߔ=����-�Q��x-~��q�wr����c�h�λ��7Q��DƧ\_���!8�'ã�@�R�U�Z(���m��Ơ�ȖL�,��1'"�N���x�V%[�_��,�tӝt{,4�hH�'Վ�4�*M�%���K�*ur���X��#���+3E��)��bJW��#0�������W����/�]����z�����?Q�xUU��ʎ��7���ߌ�+�H�k�W���������0���e�!K*!��j{��J�Ҭ��|�,�a�hl�uξN���� �-�F�:d�T ���KD u�V^x��>S����ޯ��f�IHef:jn�OG#��=�*���?�Z�ɺ��^�����#��^�i�cÕ���-/�������F�ՠP��e���2f�ޯ���USB�,.=�)��w��g��ٷ^+�D�3v��~ٺ�!|r�*V��WJ�0��g��w�h3��w�E*�� ���vK��������B�Yz�:�~wP�G֬�u Z;Z\��*�c�"���Ee[Z�?�c;@����;=��������z�JP�j�~g̥��F�X�rj���`�A�f�lw�/���?�/")G=Sw��d�3�~5+p0�0���Ք�,n��g 3��{y�P�9�����b�NS��Im��X���Na-��=d�̽/��z� �3=Q"�,�L9';ֿ�$�񵷖%�>X�o�Ӡ����p�Z�����Ș��j�a��C�M�~�0 M��t���'�i�^�ZnZы���Rk��L�:�|�ȱ?]x^��A�@����9	U��'���"�	��0����%և�d�9����r�F.z�.��@��i��gZ�bg���p�����:�Q�����׃�"h���Fɖ��f��&�(���� Wm���U\�O�+ug�219�����n��F}8�j��m����{�3�E�Px{��!"39f,��������g̺פ2����o�J�F�*sLgI402��g987��z������ì���W�OP��>16?9��w"��Sa%�F���ߋ��/?��]�;�ϯ�"Z�]��1#sN�⌕�ݪ�P:�]�2\���6g\6�7І}�W3V��!}4-W������/��nN�׼��
�(O��'��1q��>WlN`x�7��K�����9}��@^*E��͹#��R6]�e4�\~�{bedӭ�ҙ�pC�N��B�0�i��O%��������-�_W��#49k��q�
%IDL����=���낱�ɔ��<�o��	�%��4�����Ϫ���J�#4涢�-{�U	��v��q�L9V]H�N��#���#
v��;Еe�س�1�1����KKU�D��h΃y�q�=���}�uq��8��O�T����x����&�n�W��
�*�Mā�dDl�k���v��\{։��ґC&>Ю��<.�&".:�u	M�Ӿݾ����=�� /��Ho�m2�#"a�a �=��G���I8c��}��������Un��N�p1���qv*2B24�Mү庺�;=�V4g��\��Iڛ?�h�L&#�M���\^&P:X��p}���1�~a9��t���br3(m*Ďb��I?q=��j ��zt��h�����ސ/_��q�l�����`p~���e<Lw��$0����5��-�)�-O�"�Y�}ԀN`���΄-Er'v�KK@0�U��B�k���ଧ��Ч��%$
����^iyv���c�RD�j�)�%jTY��
�(�Y�U�V�^���LaUQ���b�K�JSbg┸BK�/��������9�ǩ��ڠZ*��>J�=�O ��m/���F�]W��j�|���>A�����y���9��w���<_�x�-ص�v�ߝ"������	e1��-��H�ee�3��i�rhJ�������	U*V�����_Kh/YLvz��7��ѷ>9ҝ�C#�0د��h/�ݞ���TRaW5��C�������n�o�aJ'��n�m� {,�<e������;n�Y�{&���P�}�#&����0T�r����щeǃ������������������7���XrZ�Q*������1⎿�9�/8�fP��2W����5��M:�����(b#mK-��y蜶'��(�b}O��7�X2�@x��w� x?�W���V��H(�����b*�1����_�8d��p��/\l�/\����5r�h-�Z�@��q��o���K��%�}qB�*�����8b�Dz�������/#)�[������C�|k.�<�Oݹ��(\
�\�M�&�!K)�gn;R�p�K��K�DMf�l�!d)�m�	H��4��1l~�9�QP�R]�g�̜��!�0�+:�ޯ�5$�ew�`��t�_A0uT"�EI�����>���Bt�z��^/��K~�[y�ӟ���Ale	�`T���&!� ����"�юJ逃�ݫ�M�2�,cBí���9�E���yjo�����R�>� k�*��z�5E^�H1p:��}�);Ax��>�K�J��	�Y���U�	V?��B;�2.���M����-K�h\_Mp�Nz�e�s�v^�X�%#��:$6V��\K���Z5�k�LM�w<-�	����=�x�f>�Zh��N����K�v\�k��È�p)�Z�2�a��^��%2ӝ�͏'�똊`�+��jl�x=��]����U��Qj�J���/q�+�{9;#Y'}q��'M�����GR=)�]��V�^x��LЂ��B��-)��BgV9Ʀã�]d��OM�_�/������(���p���Wl4z��U�7����B��b�?.�rois�i�7˯���%��}��}M3��˦��::vÕX_U�bV){W�mr@�F���h��l�M��T,"/8d/g�r�Л������ 
� @��>*K�?J��=�ʍ.��ƌRM��}�"��R�����B�{�j�ɰ�m��O.��))a]F��Xʉ+�Z"�wX̖T�:'#�8�9J���U_�=U:�}�n��w_�2��*�L�U%Z�0&:��V}��j3�>�Լ:�8|����F���f��.���s��5���P0����
܄�/p���q�eEgs�y�|���z��p�AO�s�g��5�9���H�)��_͵C>G���f���:nS����a����w
'�<,Xye!z΂��T�'e��ws�И?�B�C�,��镾hKO�u�X���E� �S����H'UJi9wl��	�S�Td� ��"g�5h��_�hp�~��tD��c�
C\�I?�Ѐ'3���Ri�c�w����71�7;��#�����pǒl
&\����w�4�'���ጵ*�M�G��	%('#�5��A�W�R�y�z�YV��x�u�fЖ9�kR��b{�[�l��04���a��{܃�����v�_a�u1"�3�5��%L�k�["D�iR��3��&�0ʕ��&��?�U��̑���&��4\��R����O��4uqX��#�>�k�ʿ"
��-���M
�w(ξ�w��1�.�$��{a�����j94݋��q��,�~����k����Q��5�~�b�y ��� ���|��1q��%�8f���{ܴz��򮦇�K&���LR�
�w^�h��!m>��t�'�� ��r::;��+�S �^�c��kD�i�����`Y�+���;���������P��+Tz��Lr���&�99)��}i)|*����,�㗒02���T�<���$���;���[�9 �MC���e�T����`3�7�d��wc{�b���6�<�w�d�Ϲ?��[G��9�n�� ��7�;b施�^�LBrP#=b��vCW���Lƨ��ݯz�O�#�1ID+67sG+IL�EƂǧ�g���6��z8⌓),#�0�Э��ᜃ^�lꍇB��fs���#-�	gS��,TZ9{l!�_uW-Pm�(��%h�\|����Qm�]mӓ�i*fԻFB�(.!c�W�ЈWT��蝦*� (GI�[�����x�~�\���Ъ��*��bFh:@]Vƣ⋵�;7�
�-��W�<�*�Y-g�au>�ʏu�K���p00�p/�m��?�O$�\����dh�����a#�9�W��'k���� h��Z���,Sây��}Jgy�7#6>������Z�T�S���Z�x�a����NC�-����!ܒM7sB(
x.�dQKŞ�o��TJ��+�������y��~���`-����Y�&�䯜�u�s`Q,�QA)^#҉�"�8Y\�)̡�H\q�� �נn?�ᲈ�!��p!0579��7	IQƯ�������;��.�T'�c�n����wDx��n*u<�+	��z�QƳ[�
�.����X��̰�0q��&���RO�������VX�(�y�����}u}�S�k�~��=f0i>[�^���J��ǦL�=;^�V��#YlH�� +����)p���2q�n�+�ys�I��~>-A�X`�'��nwȞK�%O�����E�oH�U�k/�#�&:�Ɋ��J�C�K��i�د@�5��B���_a���X�%���0y�|V�"�#��H���� oU�/|�A�x����^F����g�k&p��T��N<����������d���1^���!�v��1�dO�7���3J\�v%:��}����MO��XT���t��qe='g�.��/�<�Y�r�Pg@������?�M������Wo"r��Vb�������M'������!4���]S���iv��d���I��h3�^n\��k������1SX�%_g��G!��2D�nް7���Y���J�K���կ��D�'$�cS����x^��;�� �%���&à����c����wO��:�oƾpa)�	�x����͆Q���|�y��"&��iv6�ε`"Z{�*�^�kď:��ϔ�Z>�L���T�e.�.5�&��������V�`:����1rچ��p7u���A����{:���k%�U%7 [�u*-�q�@�R������˟4|�kO��ڦ�2f�<���ޜ._��@DfZ�&A���U�O*�p��ʌ�J���,b7dO�oU	���\,����4
mJI�r�/���p�����l�z�`���L�vϓs"=�^��O�0yb,F;�D5A� (��-�T�'���(����K����6x0"(b��}���'w}��j�l��6�Nn��:�����s�\mEM��	�ˇ�6	s_��]��}����c�樟�ޖlfD��o$�ji��l_琊~�9�VtJ�6?�:����L'��b�a�P��l�#i�Bo��g�YP4����Մɸʻ���!�(�����`���Ҩ7�gS.�Q\zK�p�'����W��r�9���O�?�G�x���	��b	������nݶ���C6x1u�Ѡ��j:�y�i%+���jp��f�/,��'>���_���C���I.4�@�Γ�K�MN��� Ռ�Md��O��	�$����iX�[
t�۸�O{��>ܜ���U��TGL���A7���^\}�i����Z���fS.��7��ê~>�������T�5J�����0q�k�CBܿ��뎞0��x�Į����I��v��NB����4X�r9r.ƙ����~WJ�^���j ��"��QZ����>��?�:>����8�58���@�;�iQ�-�X�L6�������1Tq���
��ﳮ��b�eU4��	Њ���׉�bۭ��oK*�d-�����xŊ�-+с��2��3��<[������E�8Bwa�f��IIs��c���I/�O��K\����K_�w��w�8�ݽ���]K�s��(%���E:��E�rR�{�f���wNzd�7��T�o�@;�����>��]bx~�%�] %�Q9,��9������d��47��3ds}�r�廙��J4V#yn�"B>�al}��v7ǐ�m�><~���F�|��"�G�)Ֆ9�T��������z��O��Ũ����a����j��_l��m��3�A��)~Ba#/g�B���M���IRۚ�Z	כd=��/�6�k��/ޓ��p[��we�< #A��&5k�E��- ���H�!�|�����@>�܎����5�f�Y��ܕw nάh�%�N$�f0r�*��0����eJ�6ɠ�/���h{��P\�h�=ml���O��}r8�nU��*g��
ϕ6���<��!�����Q�I�:��cM|�\��J�VIQ�S�������W�U�%&
:��8���B>h����F�"�\��	A[�}�=^&��:+O�K���N�fC:N����o@�"��a���=+(,+�9����=�[p��t�m����߱�¯և����e�f�O�������<nFmS'���j(�x��xSSԀ�������~%����y�������~Qj�O����h��$���(�g)��Mu��+��ЎT�m����_(��et9�wg�e�"��R��!���MGTG�xՄ�t[�D�_}�I۩�/_��͹�s���g{j��A���]��6�'^���o(u��.wډ��wB���9��Q�
F��ſ�c�Z5� ��9UHb	A|�bQ�x��75��.2��Jr����YR��ƌt�C�	���s6]1'G��d���NCs��m�ń���~}���dK��n&hV��4ų;��Ϣ7L�(��[�x}�v}F`/��rӮ����H~N��k^U{�>�֖R,�l�"���3�N>��`��6��B��?����@I�����6m�c��xk�l����,5��C7.�z�!���l���~�$gM�׾��@I�j��*�H"�Qv��ĵ�p����o�:�k����dL��={5�͸7���)��>��d�N���N;4P��>N�[���W�>�c�����������I����)��-Q��HsF�7��Ng+lk/�1���i��&�7l�Ì ҭ(r�c�Ut�D�/f�ޞDI9��#5����)��-���#�%�㬒	�|ԄT�ہ�~�+&�x����Z��P���v�0}+	����A<��\5����\�~�!�?^*��>�m�a��BAě�dW߈��+�p.\(�	0NK1��I.��P�A�_�
#�ع�/O��7�^��vc��*@տX����@��S9)�e�z���Tvr�%^D*��f�w�]���%�gv���	w��o�vI��AU�'F
�*�o`��>I�Ӊ%��7q�Y屵�!����>z`���^[��o�'��X�Xt"+��Ʌk[/ב��io�%IkT�aX +>���O��W�#� �0l�fQ�Q!-���t����wI��mkdG��V&�u�����������3$��X�40n��3鶔4�fR�ڎ�4�d�ˍgC��p�=��O<��?���=Rt<�L��Q�dk�S�U�w�����{I.�J*6���Om�ဥޜԱl�<���?�S�Hn^�\T!75"U"潢ikB�>�E���Y��p]r�t�ݶ�;3X�5nP�I��[�Ɩ�XU�~�ʯ�{�#r��������_�S�N��q|�+���G��9��p�ko��n7�1�WWq����|���Hj�9�}�F6�$,���+��w��W_���g�\`
k�\+�!�7ׄH`!3m�L
�;�Ht�4i[����˵�m��Ł�{��/|����H�{��=����r�������D)H򾴏�V��dʷ�[�a���e\{�%�����<x7ny����ǀx8qW��=��o�[lI�����#�0�����\^���>�͗�G�k���G�?�(p�	`�Ķ�Q��^���lO��	+�}8��;��B>�k�W����d5����=��?x7�?��+��e|�����{���.]��'0������9�������������?r�Ҳl�Mě�I�&�l���m����I�[��M$(J����%��K��S�1z�{�Qu>�h���C����c��Q�/{���{���?�iR�?�����}�������gϵW~���kH�Z
t�5�f�?��ggD%�����ɍRY7��O�v�i{#�V�V2��5,��i]J�7H����z�]���M�D����4�N��#���< �/�^o�9��^~��_G��F!sطo?f�s���Ȥ=_&�Rn1�`ms��@������wF4����@�\E}�-��W�n��SWH&�}q��b/�k�VG[�f���F����Y��1�z�|�k��?�G��Y����AF�c�l��X��Mf�����lF6n����c_m��d�,I0�eط0+����w����ť�?+�s�dX�Le�vThɑ��ɏl7�>6���>{�����8MpckC۰V��L������oL��	h#0��%���o�Qoob)6莆�8�&.��<gN��]GN�+���m�WW��n� ����voN�'O�~	q�G��e|����{��<�[���.�ޔ^�����boڹ��Sl�/{�d�}��}޻���r�4=ӓs���H�"!�jI�]ym���Uyw��u�J��������"A�9g� a&�����������C�PEWᡦ8�_���{�7��@�Ŗ��g��v�*A�W;�L�2w�#F�9��'��U�ĂU��8.u|�w��R�=������l�łۋo�nnx�;t_DbJm��:�<���"a��,ıę�ȤL��
Zu�
})_�
�d0DT8%ҟ|���&w�,�j��[h(Z�~f�����nm�^P�ٓRK���*N���"�� w��;wѢ�pj� K���������~jbq���RJ�X9�5kVum��u��t%T���CF�{��O?$�n�y��P+�5��n�_��	f]���n��y,*����s���0"_����@ 3P�)��\��(P�����Au[�J8I�Bιe�0^�\^��'�ԙ��6*$�-��">�M�RK�n��c��S'cC��L뼔�y+ʁf@��(�$zL��BJ�t&����7�P5;S�E:�Y@�sF|�}
	�.�Y<�Co���'�3J�Ly�b�� 8[��Z-�:]Yv�E�gm����Ȗ;$���;���ù]p��0��Y%Bg{HIl�霜�?a�s�#M��܋Ţ3-~{�Asd�7���X8}�h�L��T��T���ڈa���IVޫ �_VXA��YY�5�~8�h�N��T��d���Eϡk8������&����#�{�F�C�ћ�~�}t�N;���&G�(pt��\�\���Qͦɥ�ɧX���F�����_����v3=��+/��������z�˾��5k�=R��(X:��pLAA��>#S*(`�YK�-4ٸi����ʽ�Q�G�\#5?���!,�����hò0�*��Uj�P����"�5����ǌ�q���U�f�����y�o�6�o�F�;~���
i|�&eW�������z`!G���x�U�<kn����k`�:�����)-L�d�I)��6�~� Z����5�6A���⺗ҳ[j���H�E�F�X�r�z6M#�"��a�n�׬�i��f��Y�.���ho�N���i��>4@l�Z<��f���5-m��Qb����/9ǦVS ��u-���!��HŁЅO��p�o�0t���7�!�i=�C�a�D����?�x�����)������w���������仏�>~���W.t�|t���)�ZK��j�'][í�y�e��U]�S%�`�����^�I�a22��X*�Z&!�&c6�q��$�eɆP���6(��x��%�s`-�Gٽ�L,���E��exz�ᑫz��Z��e˖��ק!���e������`�|�+W���,�~� V/'�1�
,���~F�� Q� ��Z��z5YR���v�T�H�^��U~��ˢ�	P'	������-�{v1۪padH�Wo(I4%O`��e���b�3��$�bU���Z�\!K&��X��ӕd��ex�Y�N~���^a����d���@�8��)� �%7��I��� %o�����������8Ӌ�L��.#���|M�\J8u��5^����1��drz�ٹiB����2)���'>`��)_"Ь�����l��w�U����z
����T^�M9+L���廿Eh��E�g��(��DbQ��S�.Y�J7�3=����ԪUR��L��W�*e,<7�����k/(�%(]zѽH�R�Q�Pg-���2nn�P�L$N��7q�����X(Ix��Mפb���ϣ�~}�.4i�;S�$i��g���?�M<�#�a��2z�8co��=6JĮb�eZ)8�,�Wr��X75M��ﺩ5*m�J��_��＇v4�|�L����Db�g����چ����6N���V��
痦�!.���UQ��O�9}�O����8�F]&��,큖��.�P��L�@��&c	m���;��[!�$U,�p�x�A�d��Y]��*�Լ�/#.M�8.U������3K>�s�J��=Ϲןŗ��Gl'+%,9Ӫ�%������D�#>@Sm�Ťf�1�����7���l�)����)�R�K�՝:�u,kY&�J�b�#����U�Z#!�m��������k��R��^M@����YFL'lO��l��F�|8¾��:��[I� �Ų�V0��F)XCf�W��E:`]�������:�#6�rI�f�Lb�Js�{?���a�f��bg\�\ʩ�h ��PT��I�y����c���Vrdd2) )ݚ6��?4)���&c�]{=;�z��T������>���iC�u7����Yv�֋���m��M�M*�"���l�R~�r>��Ը�V�>����w�����<,���ҋ<��c�LN�^���ǟR�$�ωv�+�υ�.bQ��Պ��u*�wŞ�r��ٹc���os��w�˯aY��Y/_��]<UP���S��DO�S�}��h�0�5�G8s��W^�9q�S(�.ګW�-�`���#06A��d>|&ED�_�O��Q�7��^�Wh�����/����{d7=��^���O Ow'�R�Kmi��	Ôf�[����iJ�<�p�hD��̤���	�=�h�D����9 9(���jU��$�$��-��%�fY��t5q�3E�;$��b�j'%]�L�F'HM޿�
����*�8��&Xwcͦ�����ۯQ�z+�3	mހ��5��05�_L~���������Rd~	
~Q>�������cUG��Y�ʅ���>VP�:�J��ta�.�����pr%����	"ڝta�g��qW�x��u�0��F��պ�	�R������.N+6T��z�׃IB[�9x {�N�3,H��ҷr������8�D\��ʚ��)�:[8ކv�b�rS���:2�ǧ>&�O�n�*�n�Ⱥ�(�z���`��w�*�閍_�R��V�-I`�R��B��bC���GPu[LK�c�Z���?b�Cߤ��jWY��Ѫ�Y�!�x�����\��g����wl�T`�)U�\�ctj�j�Ķ�kX�Ӎ�8�ȱ7���˴��5*��0ε���T�>� S[Ƕ�%��"R.ﲵ��A�<�03�)>��-�.6n�B"٭�,�8Xt&?��Mw�P��.nM*���07��Ą�pK� m��<dΞ����ӎ�f�D�QQ+J��6��L=:SXᏛm�LR-�������_eՍ7Q�F��,R����D����/���t[�
}ZL9�>�f�
��,�r���@w�����ۯs��h�aeRةVǢvɚT������!I�NA���I�&��;����t�=̴\Jm�
,P�|o$�����o]�Q����{#�fM�H�R ��:��e�nz,���3��2����'zW�V���#,�j�tߥ�u���-5��<k6q�����71Q����T)�I�������$��H�T�����fQ:�"�^��Z����2]� ˂&�+�|���,|�!�j�`U��B󓦄� ,�"y���X˭9��b���7���~V�#[��!��G]܌�M��"[ ����sTP�5�Td��s֯�dm�5���N���k�Iz�,����/<N��I���Ew���(R�4d?�c����%�:��Pt�����]�v�v�2RRP�^�,��y|2�!�t�Uꬄ/�d���&_2ݐdV9?$�6n����EN<�(��E��'bWHb�z׋N�Y�
��ԩ�8�I	j�J�~����z����OI������^�v�lNt�����u���_-�W������s�B+�^{����3t�m��*�8�T��Œ��K��|2Ѷ�*հ�xqj����3)���TX�A�v�Z�AS((���zz��H���c'�t�8��4�V���#l��A����T���&a���u�F]�^�2�b���H�RLN\�v��w�[�qrs�^?�&?|�o�x�R���*X�e[hU�g�ӿ�d=�4�Ѧ�N�Ket]��~B� �R���4�F�Cv������|3xB�j2�\�<������E�kNG_�DЩ�V�V'\�Rd��7�'��1���r}7�
v�@��)R��J�g�	d�ɽm��,����P������1��y�ӵ�՛h���y�2U9����T��6�GNr��jT������N�	X�f����>% �Rkb��2�#)���x��%�N�~M�.�^$HT����I��L>M�T��&h ��-���X��P(��Cܴ4�ɥ�j[S��� x�j����g(~�.�AB����w��;t++J	㑠���_���s����O��m��;?�fc�ҟ�F.v�~�	��I�
j�$�Y���\��f �<�*]ǊM}�w�}e����Ӱ''���j���	vr|�e����P�����?�_P��i�`m�Bi�&�&��Y��0�6n`����ti.�t�pD�*�R��K�l���t,3i�_��9��_�cͺ�|�#t5sT^}��^�3:J�\��)p$(���%^�[�Wˤ�U�tZe����Od�nn��oڴ��z��![���V��?��]m��j���!��
�:vw"B�W���I�R������}��}ҧOr�g�~�]�s즎�%`IG���}g�6v�r�]9�",����~����{�"�]=ݬ\��dW�>W��{E"�r.��
���������	(�p��
]ׯ`]2�=5��{�0��1 {Ky\"��n�$k��}�J��8�J��tQjy),�����oS��s
�K�\e�	�Y��K�yB�XҶhf��^-�:I�{K�2��>Y����/dR�̕�^c��c�G���f��V��X�J�_(-��(�qB�p�\Ӧ�H�������7���P*�aH�C��o��{1"ڒ���H�K���}ȝ (EuB6�ܬ2�I�J-*(�������o���O�"�a7K�X�:>��'}��֚.���t��{���?���a"��X��
H�͋�g��Ȳ: Q���u8��(T|/ W�r����'gg��jtw'�hONp��k\}���4�j�E�q>2p/�[lD��Z�ר���,Y��_{��7�E5e6[�+	� e���]D���U}�hbrgkF�#�� ��ځ�Y��(I؟嬧���{a�K�=��[�`΍��\��.��Ȩ�s]��	u��2�{��`�]���M�}��,k��f޷��CiǾ,n�1&~�*��w�@n+����*T��	�鶼�f�t�%�?���iTI�RG�-Ů6d"'�O�/��!�m;�q������L7~��$��|:Av�^5��5,^�z�
pq����hr751�U�]�פ^�$�%{����!>x������F��Q�l9a��F� Q_P�w[��f Ch���N
��i`�|�)w�g�	�K�YpE?�]����4��*]"u���9�A���Yw�x7��p9ID�`�V�BU,��h�@����O�83��4{`�}����G���S���O|��X^���~V�\C:�a|zL�b�6m��?@4׻J@��3�8��k��o���l�D���������������an��n�� ���7v媂���O0��	�!��$�Bւ:�5�X�6q��b��a�*�vEi���+X{띎[�; ���ʟ�K���p��妵y}��n�H���$#o�z��t��Fb�n�+7���%A��n'R,m����!�� (,�F����4×Α�,�y�z6o�H ֮}�"4C�������JV)W���$BNT�޳�nIko
L]�
�*�B���8�t�������I${1���9�2�ב�.��hh
��G'�my�Z�'�(�<E�÷��."�+�Ža���[���r�u���߹\_҇������m���[?�vm��٣���OOR��,�n�ql���ҥk@�f6JU��w��;z�N �3ѩl'S�s�q����#j䯗�PsT�,=��-�X*�7�T�1���w2��t��T����;ٷw/��=j��-Z�ޖSXɨU�c�'?���ϱ��ixl����\�2��s��9��s�2��K����h6M����Ҟ���{�i�P��6U�am�ȶ<�6����8���9�N�hؘ�Q��D H� 9��"��ƪ۱+�"G���蔱��n�4���Sdri�)��[շ�-+��K�2��1�?�4�����`��Q�N�]'�K�S���M�m�q�=��Av�� 36\���NtO_}�˜b��G�����J'P �MmՌx��*�[�����\�X)3�r[W�
.=�����KBHp�((���IMx�
L[�Fæ�2�l���

&\�v4H�o8�L.C'G��X}J=����9�N��S�8]�z����"�B�H<Do,@�Q u���)���.�l	����:�h	)�u%CoG["ְ5�f�2��v��y�+H��"���/�J	��C(���*ؕ$aG���p>K�.�Ii���,fR
nK���\k�u�tA��	���dOL�.kh�t�E����:k���b�*S�I;�ǚ��گ>@�!�6�&}����!��N���"    IDAT�1��N�|X���Ry��Ld_7jZ�N�LSk5����	0�T.���OBmh���~9�vӔ=k�G��O���-��:5��D�A`�.n�֯�u��ۏR���/�)���4E�4e�#ZY��9�Ps��]�D	 w�,�����2��S��/�'$ު0��k\z�Q��g�T��㐢��(�����J��^93@r�5|�[4z�R&@L,����� ��H~I���I�j�e�iX��%@�P,���`�t���,c������H��j��:�N������+�`ف�F����:��_�e�k6S�b&���	�H�@H=��A��׾l'�{ɬg	�`W�25;���{�z�K�K:��'��K��IOw���N�*W	�lb�ET�-�.���嶘ɦ)�*

ĥ��ᖟ�Q'���!�cƣ�I"+�S5l�"��F��v���~V�q7�#�A�ʒ��G �ӎp�M�T���Q-O�@��cz��l�9���{�Ӓ������s��������;�[��[o����w����{oRk׸��[���ۺ�e���ra�g�|J),����b�N32x���K&���w���߇+�\mP��Ů7�
��!2�O)ubp���孜�M�Z�vy��W_��Q�"u����5l��i�
g�'N3�ʫ�.���Y$�nQ���w����G��r�"'�~.~J�l�{`���c��H#���l��6E"��Rݢkl�h6UX�����?��Ks��>6o���{�.���@�[�nd�*�B2�2e�J��Yg�ْ�^�pT�YN��2q[ްL�Uf&����9=�˱����k���4C[��4-�֭6�i{��m��y
�>UPP������`n�D�������<!Zf�?�s��Ol!^_҇~!>���㞫�]�����`�Jl��O)���c[�"ct�[ɜ�I:�NM�4?0��tyI��lT'��D]�u�4!X�*�v˹�U�&�<��jf�|0��v3�5k�)t')|l߷�+W�����؞6u;�n.	�q ���V����k�Mjq���1Ʀ��]\ ]ȱ�&���7q��K����t��$� �}2� ������D�&I�Y�$޸�k��0�����Rx�XF�t������`u&.22P�%'U�iwC~��ӹ�y�g��C6,_Ɗ���3'��G�g��'��eBҡS��p���t��5��8��.�Ȏl��Dvd8[��Mϲ>�ɯh,����<T�w��1ѡK�v�s�>�z�|6���f��}�:V�|d��ɟ���~F\
cq��?�ܜ����
���]�:�X����7��+�0Vo��J�q�U��D�bW�pA�6���#
� Y�:�r�t?[��J�٩yK�Qw"̪�Ecb���D��oa�@��T*�_w)��j�)�"?	�Eg��"�q���:�݇H{���. �Oh����K#���p
^�pt�|�RVU���YXXP:O_"No�O��YF{����D�UPNv�%�|M�+�O�����$�$��%�o��շ�C����9Z��^�bkh���_@��d�ɜF�~'%��/ _��;\.3>6���	�	�#Ӏ�>|䯙=��r�^�K��:�P�sF~�keu�I5�|a�d���ØkwPp[��ߙ?
U(`��Dhڰ��X�$��3�h-]�:����Ќ�ɹ�N$ɶ7��ۢr�g�!�'�&\�a��&I�N��-Dq�B�q��xȻ=��I{��?~�g5��r�`XA�]/	���N0W�T�+������ϡ��!bJ � �+�����+!X)3������Fpq�D=��Q���_�ф�Z�蚐�Ir_�0Q�Ɖ�?��{Ľj���^�vZ�b◯7�Ґ���9��.�;ט t�P+M����]�gѕH�����Eξ�,_~���q�DH�Z5��&���;J��a��y�~jm��R��ݠ,�1�,��(�mm!��d��p4��N�)���f�@��T�E�Ah�V�|�~\�b��x6L�b�3Z�fպ6>�"�|�lz�rn�Rn���`�=�۵�jݱ�t{��>}���O�wN�>�������{���y��Wx��%�7�� ���oiV��O>eM�J�����I�n���ؘ��5+�9����;s�#����.M_1�(fsL����!�(X\�$@Mt?�9���dIV�҇�M��&��g�~�U���%�a/���Yv��z�
��b��cxO����8�i;|����|���\z�y��E�ۤ��b�v��-J�3Iڦ��Nb��,g�Л�ؖF���IS��]���SL�\a`Y���'�h�"W���^��"���N�QM���K]�Ē{E�"T�hRtIru]����u2[d�L��1;3��m;���W�����lM�Xr(��m�w��)�.��@�N}h���s?�ͩ�X���c�⇮�w�&*�����"�m��/A�Ϸ����'`�?o�ν���K�����ܩ�dgp���Z�֤]�4R��WB9��h��\�'pu:
E7$_�Å֩� p�(�n}g��$����p�5qRBy\!��|�R��ýe;�5���Gi�St�ٲs;�{��|�C>rW�5$�:K�V)V5^����+��Y�033���$��3�,̳a�
���Ś�����}�ޅE�')�(�������i7dR������Gl�^��� ��-����]1���������<�AԢT%U�ZK�@DU�
��dE©�V��S)�星]�Bg�@/kzÔ�.����g�w1g2�d�,���t]�3n�RlC��%d�>z]ϖ�~	Ϧ]\ZL)5d��
�HH؛#�r�fuH�T�j���P/��0�.���R��WF�:9A�Rae��/�9:�٧~���W�/.jJh��H��;�l��.�]9g�I]:Kk����m�8r�r	$c��}2-CCz�tK|�%P���ܱ��<'��*\���9&g�(�k�t�ذ,���a�ǹ��0>��&6��^,���n�d��5��]�<n
���ν�����6�c�eҰ�c��P�L7�X�_�����I�.�]V-=c������2??����Ǥ�+NW<@u�O<�������J4�c*�N� 7�����cT���{9�ǿi+��D������.�%�=�%Z�! ԡ6�%n� X �S��x�н�,��&v�M/��4��+����53�'?y��O?�=���Q�"�h	ؒ��L���#|]�2����g����X��Lۃ�	(5LD��` Ї�)��3v���79{�����u�q�sڨ7��w��D���/^��W��ď:�"�b����)���I�ة:�/-.�./�X����z���z�a�z���K�z<�+k�3�Y*�,������\'�@(dB��da1M����=t.�g>�Ϳ�?qM\&^�h�>��!�M9]p��� ��>�����q��H��l:����EHփظ9'�g�Q�0_x)ӬG;����fr|�R���]q6���^���q�'��^&�,l�1\m��j�Or���|�j{|�0_̫��*g��4V*�[t����~	�t�A��l�v�f�L�Zׄ���o�D�mwc�;�M^�D\�&��KC1+�$h���Y&+�4�@��6n�ʦ{�I�7���)(�����N��r57^�ʷ8�֛<���y����o~���)>���l�FO?O>�$����1r�,��d���~t�O?��k�;���6��6��F��)�
ģ���	q7�i��n,z?�/����6��+�N�c�WtR�3JT���aٝ���-��έ̽�
�sn�p�uR^����D�r�
\\c��(�&O���"{��^���3څ�
�H�?��#q�� �"�֥R��Yd|�
�R�-[�Ov9N�������*LC�W�T�o�ν!I孲j%�P�����Az5*2-��gi(��q����W._���#GF�z֊^�%M�Nd��l4
��W�Q
(����2��Μ�u�$L�'�r�ް���k��YJ���=��q���$��r��{�Ȉ����S���0=�?{���,v�����]�έ:6�T�5j�c]|�e�*莓�Cr��~�o1��\=ǫ۩"�e)�;B/��R�N<���GHy��z9��y3��m�]m|�8;v�`m_/I鬅���� v�~�ӹԗ��;�'�Uǔb��ԄÉ�	Ʀ��L$#lްB�S�wޡ���tML-�p�e����s٤[MR�E����a�`l��6������5+�&b����|~=���Ҧ�g�b
���W� ���Wn�p�k�Y&ǘ���rӿ��-�Շ�ē�p�ŗ0�ӄ�B���)����VKD�=�r-�����kob�mw�Z���l_(̊+�F�Τ �%�NI�W��R����NV��ڙ��Taxd�!��$�a��ܤ����������!���0�.��i�є	�2�?��Y4��Xk�����In;@JrxQ�.WK.��ΣS����<��ӵ���

�P(�}f>�bp��&N/�K��'F��a��g8�ܓ�/]$P� /F粑�eH��Xf��ꏟ�E���=Ȯ��'�q�B1Q�L��Q��8K
k�h���@ʑ/`��t2�T���q��ɞ8�=��M=���0�W�@ގ6Aׂ<[Y#
`�M*��~=G�#�q/V�J�fh��K�zo<�m�g��Z

TV�y��`7qa~z'���I�/䘙Y��2H&�t��57����?=Acf�Q�+fm)����g%ù\��-����8ʞ{��{�&rm�z�"4��:d,�nv���q�Z:m����g942�WB���R�-�B'+S�MW(H�߀�i.=�Cο�4�R��[��+4�eu>Q���ܫ-ȋ�p���C׳���q�oԂ�k�Uj���QI*�8Fj��Y�K�`I0/G������(ps�s�/�5�uY2I��"�$��_Ls�����p!:�{�����!��%�"�����t�?̦[�RP��ũ�ͩ�I�Lb�Ȕ3A������[@�Xy:f�l'v��S3-�C�Iq8�����m�>�(��ě�lH��W	��l�
����\��B��B�D�hQ�f�L�$��X�Ӭ���
	�%��C��`�P�l��Hh��6�X�����z;�#7@� ��ťЭ��I��j���cWJT�.+�C)��}�z�z6�܋mU� \w�����{�u�]�x�����{||�S~���3:>̝w|��A.r��9�?t��������7<����s��7r�ݷs��)����Z������o}w���m�O�ri�B&G"'	;39�ex��T���� �	V�I W�v����q͍�w��Zx�=���e��䅟�e���i���H#O�� e��9D�_�=ׂ���L����_�o��6�ع��u

�~\�-�Қ�gK�K���P���'N����e���j�*Έ]�=x$���)�S>K�,B�t��5�Z���.�K����"�a�-�uu�j�Ҵ�`)5�����L����n��}NJ�Gh�2����wGK'	�b�+/��`��\�x�4�+p��и�i�YEd�!|Go��iV��{��˜��z���$���{��������mMMf�\&uiR��^��:B9��[�h�0"�`��<��}f�BU��6$���.�4����ʐ|}A�Bk�?S� Z��7�ł���K��kh�_ǩb�K�4�V�{�N���'u@����QF�.)X:�0�z���z9(�.*��̬
&�eb0�n��b��3�N�}��3g�f�X��?H�����b�I�Q�d�4}&%���ƪ��S	$1b}�ݲ�P4���c��t�E �#ʎ� }	7R@�܂�z~��'��J�����#��Z6�=Q6��!��s��qꩧax�`U����;V��|�ա�O��o�k��Y�����7݁�a�un��wu��tZ �aE�KݿN��� �)'���ΰ<}�-Z�#c��̱�/�Tg��u�+)�_y�3�?�15E/�����2�p@���m��n~�z,��n;�o������ �x_8�ˮa-�N���q]��
������@�N��-��^��6���4	�3̼�'��1��!��&��rE���iaF��y��"�uS
G��s��w?@|�>�� �`���qՕ���9��b)(��<P���\������-6�l���r�"�.��KbO�1��3�{�1��<V���M#[��`I"{�e�~�Z,�{�*V_s��̈́6��UX�s(�?���Tb�*�B@��O��`�B\
4Y�zb4k�KLO�S�]�"A��6�����&�SYL��5��Z�-#:Y�����$��w-� ���N
��v�o�������
je
����K��g���N�c���vy���a~1E�(^cha��� �����k/,�����TKSJm��y$�����M
B��J�<x�mw=�/W���ZMJ���'
�F�
u������G��3�3:�	
 �G��mr�N��_�9��s�J9��їI���Cn���%0��������;ql��Q�����!��$G�ˡIc�
*��+��Y�03>A>���Tl���0�Z�������?�9|�D�L@�A�C�T	�!"�
�^yM�I��"]*ѐ$qѓBi�(qW��}	O�V��b�L�R����0
E��E�1����)�������91��/��iժj�Q-����T�ijż���6�c�=x�1<��}\8{F�CO?���nn��+�������'������ٓ�q�W��޻�p��/_�Λoe��M

^;�+ׯ��o?�������GＭv�������m�FD�T)[�ʥau-�E�:)0}&n�p@��M��Oã���"�+R=w���_ǘ���S`Ѭ�f/�v@= �]d��穟��X���F�Ё=���K��F'�l|���^f���x[��V�߾���ոz�	&���h����7u�-yE"�;K rSsO�v�H���Q)+mR�b]��:�>�AS���q��p�"�-�0?���e���H&z1�����P �Qɍ1d�h0z�"�Ԃf	�Z��cK.7��5�u4����)b ��F\Jg6seJ�P;{c���A�,o���2"{8z+v��Z�E�����.�r�������|?Ϸaϟ�z�է����Ĕ5����Ocd���m,)�%-"-ӃG���.�Ւڥ�+!-T`�l����)M�%�\���Cj)��#ɲm[������7���n�`�E����X{v�J�jT��ځٵg'k��-� ��Cr8����3�t��H�δ�-ANn	�qS\H151�����#�M�q��\�i��"�c����+�f�;,� ����&%>���v-�7�I%�=���{��������M[G�C^�ɨ
��Ҏ�>)���ҩ���t�j_�j�/��&�|��I&'f�U!��aM�.#������R�4K�.�]C��N���4!��������j�ٶ��Li<^�j�����(�V���y.M:��/t���
)��m5FFǙZXd!["`�\��D+�ȱ�9����>k{0%��\Q.��R�ɔI�!m���U���&��r���Z!|�nu���g p@A']��{h)�[m�v9Šfj,�� /����XJ�����W3L���>�cjÃ�+�vݘ.S�ǚ!�!�|5Q�ɂ�PЕر�=�<@b�~2� M���n�*�;wܜj(�;K��K�@�n��բJ�B�M9WTmL�T �r I{�*�O?řgŪ,��-�9qq���t�װ�~jF�nk�܀�l3���
Ѕ�!{]��B�.��O�KA�t7�9 I��L
dd/����w�����,ն���;��4��z���a��x�(�����4��v�'2tQr�)#�v��_�Ǆ6�!��P�������
(�[�**���5:�sim8T��6TP�b.�V�$�H�tL�#���0x�U�(���#��bm(!�^@

DA2�q�{����{	o��lۯ&2��l�
�&zN�� U'4R'�1kY�I�q���i��􊱒�    IDAT���'y�o������D���9����-k�kQ���kc,�&�{';�W5E��<�
"Q5x�m��O���U����P�� E���%P@�ɫ��rB=�K&��|��\~�5� 3@̿=��B�]GfUJa�ױ��4ļ��z$z��t�N�R����Ǥ�4Ċ�^!j$��L��t�JC�z��,h�g(S��n��a���:tt��}�L��ըש�k:��D�r)K��Vk�V��Z���ٺk/n3��&m�K�����ܳOG�>��~��p����G�g��en��.��+�`ph������t�v����sγi�����+ü��S�]&���7�o����Z����WH/��5L��LR�@�c�!�Nq�@J/�����P��Sƞz���Y����}�ƺ��Ç��<�"���x�e����mkX}�/�:�t�TF�	�o<�E�u��vlµa޾B�e`�iY>5�&�4d�/G��R����D-==I>�H&��oE?��
���KP�?L��J�Q&�lY�L�f�����]N,څ�Q�8�9���$nM^���\<w���9�[���8�����|'m;j�O�Δ^&�V�F��(�p_<�k�2�f���J������D�>��+��_ϲ�%(�yV�_~���XX�N��?�̌������GgY���Qަ���>t�
P|���m�.<]qڐNL�Z�T�)_�c|!��8��z#�5ҥ�˨��t��zK�ģ�t#E��x�A�~+Wal�NiY/�&#����bϾݬ]9@$�+E�9)�-�&m��ɗ�V �o����
!�M1�fz|�ɩi�F�9{�4}��}x����'��O�O�����-kd<.Rv�t�J�^�,�ސ�t�H\��(FbF�����ĺ�D�~b��&�a�u��!y�'v^���ZI�U�t��F@�Й!�*^���ke|�'��2��E��u����8�@,�4{����Բ�EQē��ۉn�CJ�ׯ�@>��a��{Tct�=9��^Rh.��-"V����I�V������|�[�wo�{�μ���1M�4[>��k�NJ�����vTE�mz�G�xVo`���ҳ�%#��@2<�M$�
�^�`i��ũ�$�s�����h{U���c��L{��������+���r�>/�ݎ��\Db_[r�XlݥnT��{�x��%P��S�L�zb	\�ܛN�Z>k-�E�ٹt4IU���['k�X�-J�"�s���
��w�h�q��'8�����i^�m����ND���%AV2i�y�����nd��k�Vm�ս��Ct%�!�1�M�9 @͑���λC��)�-���)ɣ�~mlC�KC��K�y��9��CO�d���Nr�GȜ�s!�4��-���R:+�zPm��M/�-
��]����~C���֤9 �`�p8�y*��cg�~��D���]@�<r�J��n��|j^ݳd���>z���K|��~�u|�4Q�nі�f9����'�F�����(��[Y�mD7���-�����$�Ѩ���G��D4� َ�D@�@��`Zl[�`]Le��鉆���̞<�[��K�C�IT+D�|�o)�A<�.{�G�բn�i&����g�}�v��7A�$� �pT))Nh�3ǒg&���[����9}H���&�#���L��`"F�r����ѓ?e�g�N��l9�@��B/i,�H��X�L��m�X���Vhy=��P��b��iO�B�]�(��L��l��PK"Q�L[�
�Z�@����;��^�;�R��R6����1����,�nұ�P�\1C�Z��e�+׭bӮ=�O�ۯ�+��.����y����;|������SgO�G����q��^��[����A�x�	�?|��t3/��2��s�:p�t6ų�<�Ջ�I�̲v�
����k����x��J����(�E5
��8Eib��Քf#�!Sq^�EH�>���?��?�:x���H^&Gv���_ƽ�0��p�*�ϿL���%ܞ��7����;0����0�e��q��x�rv��8�=;�lٌo�>Z�_�0RH洸��wv�$%�#k<�e���&FX�b9�׭��S����>InW���Dk��,�+�s�j9��#Xf۶h)�צ�����"�2�����(�i�i�6�ɤii��ߗo���sI�Ы]����y�5j��h^��w���e��5�NkE/�=���r���&�2�����K��/K��'�� 2y���);:�{��Y���JE��G}��]B����5LG@��M$��E@A�Q���R�dԉA
"�'W��Ֆ�v��A�V|bg)cv�x�Qn�uL'�\��.~)��,�j�r{v�۲�)�͉�ì޶�����z�jb�(A�bJ��pl�^m1cI�%���;�x��"������윂����s|��xJem\����I�{���<�t��A���&�j���)���h��œ�7ҿ�B�[�`K��7��X,L$�tE�M-Y��u�L2�����^n���l�)e�\=7D>_���)�X�<L�0Ʌ����7(_M�4>�㤷*EZ��W�U�3��x�n�Ɇ�n#�}�uIy���� �ɤvHt*$.'G��(p�Âj�ȭ_�P.��k�X�Xn�k�����Co>���/P�r�1D .��|����c��*)�^�z8�g�ZV���Go&g[X�n,X��HX�N��/�N��t�>�g+�șȟI������H��b�g1�㫤z�1ξ�4�+���b�'׍3�Vz����x�����i��%�n�ҝ�w��(��` C��=�.�.P��_<PPoP�Y�g5=9����i�^f�'8�������ݰ1[rٙ�R�?[-4���fB�o�[����HV�
̾���e�`x镔R��uD�2�q"˴,D�S�:��L���Ԩ5�TS%j�&�R�v�B�׀�!>}�՚Ԛ������tO.w���p˹�nS�M�kbn��u��t����TW@CńB�C��YXu`Wǋ�3�ж��U�![�z��Լ:�ȺI�}$��ӟp��'���}���VS�O��~I/�r��M���ݠ�c�]�ʣדؼ�{%��2�V��$��;]�r�n;@`� �a�9�^�d���ѱ�+�l���v�2���UrL�x��~�=�+D�e�r֊�B#�)8��:i�5�q�A%䥽f9{�{��n�]N*��4	�B�>d��$\N7�r�Uξt�u�� O�u#S�&�ZUE�r�x>�!?>Y'�Wx�{��ŷ�&��H�Y#H[�D�dy8A\����
�S��F���1Le���kx�U(��ăQ,o��d�m1o{ț^캍�X�r���voTM��y'�`F����bgP*+(P�c�B�T�X�P(�TO��-�]�b�*��܍�Q�!��bpp�?��?��S=�u�����?������r��)n��V��[����Ǐg϶��w�3��*qp��{�8/=��м8�y]<������m廋w�Pcrd��ܢj�HH�vx]���#H��
��/{o$�}�y~��:����@�q�$���EɲeZ^��솽���u��>��>l���ڱ����N�/ɲK2�$A �h\}wu�]�w����Y�sHt��`�� ���������Α^�]x�Na�M�����Ɨ��~0+��;X}�m�'?Cѭ�P����#z�1��~�T{�|�1V��3�nEy�.��v"3��bz}-%��Z������-05n2B��]=}�/�C�9x�ч061'
���kX�r���!�D�X��n��d�j!�Ǆ	����S���f�d��Z��-;wc`xT䖜���an����'�Ѳ(/D����k�H��@x���+Ȅ���&P<p?����+G�Y�������A�о�~-�B|��ќ��r��٫��Yoa��Ux�1�(#�M����Ce�N�I. ʌS7��9��w�i7�m5Әt2�Y��w�AH�i ۀ���`��ij*Ob�n��?]�D�F�L�a:m����8�̾��w�B�\���9�q��ݘ\��BE;��H-"��I�)���/��8�9��FEC}��������XZ]�g���q1f�ؚ��(ǣ���D�K��2�[	�� �A-7�OR�U��Mn��}cp�n��F����Q@�\�]��BS �I�^�E"`0W�Z�(bc@�c�
���[hw\��������6��m����3~ g��L���AN��4���C�|��-5�0��b��`����
�z�'�P.P*�)�d����4�aA�í��r���X�:E�c�A���s<t���Cv�-�ą׿��O�֪��Z�Iō'��ϔ`0UBf���9d6n���a��_B5�`���I�H�Yq��Y�I���Y2�W����"�E���޽�"�YM�d%����� ��{��<̮+�a$Ի��Uc��>NDZЄcr��|Q�k���%bs�C�WQ*��R���r��:��w��ܛ���P��Z����C$ɲ1��!�}���'����!�6aq�NR� H���hN��G�tu�����u�u ��<�m@f��<�N
l��Xy8-��y�&)6��!�A�*�{E��G���xzkn�n׃84|��/���;ķo��u`�Ě�D�>����7��	�8�[?�ÿ����/#Z�F��Rޣ����j��Ƽ~����b�
�>O�OQ���P�/�t�T�J�1�����9�>ο�#t�_E�݂�t .I�N� @�[�˳���Ʈ��{�Ø8���
뷡0�V~MRrtCCC�fr�ٸO��'�+�4������</�����BB�&*ԏ�������䏾�����H�dY��ϗ \'�X�D��@�V�W���o`�/ 3��M=GA��`�2 ��)G�fi�^�_������h�VC�+}��L�`��1����	�0�y�"�J��`k���xa %���ibh��zPĿ���!�ЅN�j�#�W���|(�Bٴ٩�h�6�g��>7��1��=�������>�sC��&Qi���HC@-厽N�V�N��F�2a<�sY��]K9���Wo����_�7^Á}��}��ַ�=|t�}|x�](���|�;0�$����'殽�$�a��]�.,���3X��Ã���?�g а� ^�|��-�����t�X�k�q�n���6""*9R�,����W���Q{�>�{�����C��y��|���ȵ�`)=@o���CG�{�E`b���}�9�G����U�Fn�6$���B�0��&I�R�WE
�[��0� ���_��[_�Go��ٛװqbGz@<���J�jQs�K���@N��Mk1imL-L�8�FT�	�z~O޳���D�c�(���*��/az�N��PM1�{��T$�\H>����1bF;@rs����'ixY.i@+*0�nB��C��G�gJ�)�#7�/��*�?����)�O�V�`����M~�������/���[�Щ�(�4ڤ�V�9����Ac��Ӡ�H�T�fO%1|xS]9e/"�H S�0\(a�P�0�A��kk�u�������`vT�MЈG����}*GDwbgWfT:| ���*��sE������H�����^��j_�,ɛ$���/`iiIR5o-,�^]�����f1ʗĵd�(��;F/o��8��d.��cjcJC�L����=��uMd3y�oތb���I����b��'��>+\
��E��SVX|��1�T4�u��/��8pVm�"�{�6���x���?�q��jJ[U�V��e�q��Z��Yt-����|
�x
5Ò��48��#c*T�P*�^�M��l
�Yx)�:�o}�4���vK��A��F�R�u����'p���3�`���,�/�xl6Hq(Eu�`��r�7-��0�����t���� �P���-f��QS���ʾ�6���y�����)�B�/�
ꏘڑ�
���@Oz�,@uǿ��h^�,��H�`�R���c��{���Zгt���1�k?v<�<Fwߏo�|I�M|���>T@�r)�X�������4"����\�Z�����"�9`@�c���q����v�2�VS��������H?�"������t�i�p�d7m��g�
{�X릐�Et�Dd�� L]�4c�x�±a[���iYȿN�X�K�^����N��EbK>�Pt�;�>>��_�G�u�3E<��#��s�4	M&�'ua��b�]��^����
[va��#T2B�<F���ЀԧLYF�����{����IMs%L�B����1��P|k	���q�'?�ʉO`�W�v�JI_ ���g��	(d����5�PBfj+�~���mDnh\���G�(U#o�}*q%�X�4)S���H�!��s����=�$s��-3Q]�3p�G��§c�����4W��A!V��5b�t�IP3c��yL?���ۨlُzW��9*v&���	O�}����!�bieӣ˙�1|J/�+r���i�!,��?�s�{��P��1'�=Yn�\��MY��J(H�ZOM�_�T��`Rr"�_�2�́�H�|d�<�b���0t�0F^�:P�@|c	3?�W���Ľ�����O"�{?�&&��qOJ�Ii�i��m��Ө�mw�4���l�Va�-��0��>�l��������p���Б�;��Ml�4�V{��9|���[��ů��-۷�v�����.�̙��(����"m�..���3X\��G>�/�h/	r�iu1w�.��U���Eds����(����mUE��U(n����7߅{�4�.���޶il|�k���� 0���GQ;���*
:���l#�=��cO�ܾ���}��?z���(�ڄ�����
s|#��0�|� R#d)��w�$x֐X1�)ԩ�ǰ�x'ưw�6d����x��I��$@%ANK��GM q�4,S�h�h��u�Pa�A�&�d��La�&h`�Q�bvn�z�w�]�͈����4��+9(|!���QE�X�mx��w�3���CM(ƖIi�p�!�P����1r��R*վ(毛�/�7�+�����ï�������Z��!�m�N,M���R4�W�\''|a�}�e�F�YHq�����$�ϝ��mE�`��A�ɳ&g�;�QVU���*�f�C��3�z�2�u�ݷ��i�!Tq���X_)` �����)H���b�
%��3��ڛ/�!�Ч��S��F��g���"x7/úy������^���đ��ӳ�*�����J�8����J���>p�[w`-L`�o�����X��%)��۴*e�M3�*��̚y�}
��#|����եa��.^GVu1Y0�ܼ�����K���>� �BU��r23�PN�����dD�����o/�=����pw��X���QY�ږ���Q��L���H�L?W�����:"?�HNԂ�E�X�ΡbŘ(]���Ջa�<����(�ɓ�b����r&zJy*UP��>ly�EX7��V�+��6Kh5;��(��*�DL&�`�"�����+PV"�`�:�Ȇ���w�l-!�0���s'1�λ�nނ^k��)Mp,V����0X��ve
5���±��m܊m�?�]O>�j�!Η��
��%ȱL�:����Ѡ&�C&�w����s
��� �P�TXN+9id��xA�ٸ�k￁k��w{v׃xĐ�>����yzʥW5�t;�����#C���J���L�\N��j_#�k����)R���z�X8sÄb&��(�»�q�g?č�ހIӮ�@ᤏ89VR�'<`(c�y��h�*ڹF�������G��JۗkĆE�䘼keD�Μb	�<�͎�(��*�1\jř0N�B�A�uP�"�c���+o���N��I!A	r���{ )SR����A|���&��{�@\�4�L����XEֶa�m�&��x�&�#���C,��	z����g,5�3�<��Lzm�_�!���:��9d=Y[!Cs    IDAT�X�s����x\�F*�L�fڱ�i�h�Y�K�W6=�$<��F/��N�����ڰ�%�L�欰)H�=
�(�4��@���X��W0P)���V�B���m����O}�l��r��r\1ǽY���] �de��&詉<kk��z�R�&��$Cq+-rLz)��y�aL�)�������4#��9�xp;&�|
���eQY���l;���}��w�Ú�jͅU��,�s�`MlݱG}V����u7�����?�{o����cؿw�9DaA��իװ�TǦ�[%M��!��wgg���$��ԆM�y̍d���겄���3x��vU	/�~���*�l^���a
剩�̣1,�(D�Hw�n���)���]=���GD����=�����R��G탣��Udu*&�1�ԗ�=��n��a��h��~���]�9x���P�'`d+P�Bݑ�)+�4y��y��˔ʃi���}K��l[���u(0 (��1��$�W��O��u\W�6���G��)!��H������$D��=/�j�%���}%%��&���}`�=8o�(`�#�ǌ�}� �*Ȭ�^�����\=;X��K�mـ��A�+�W��e��?W���_a	������g]�x����SSo����y�������l&��n� ��N'���bh�E0q[l
�S�g�5��o�3_(i�I��7�r������{!��(�&rd?ך�W�`5[ؖ�Q��ĢX�38�hj#܉�C�Z���`߶�(�(�
B�`�CqӀ�tRy?ȥ~��M��t:�/W�:�P���0�8���0;.Z?��=X7.bh��BǇ�Pv$��&M�z�ja�w�3��6��8��ۇ;��%q���;�&����I��sP�?�7g�ǦQ�_�<����b�ut�,3cظ}�*n޾�� ��x�$Z�Σ;s� ����x&�)��m��֐K�b�ǥ�v�!F86.�#/�f�`�0:<&)����R�R��<e�K���G�'h4k�5\���O��kKwQ�T�f>���|��wQ�'��
Ck�)I����{�ׁ��9�u����i���#O �a��0L�� ��m&W�5�7QR��ʧ̾>����+����PTI
�~������ �����^C��$ssȴCH��|iK1,)Np#	���6�����G���~��ښ	�<+[��43V0�ϋL+�"�&?#��_����r���{� �{=��k0�e������?���+"�)3K���)��(>�&�)|Sr ~O�I:�� �?�%��՗al܁��G�ɝ�r��L��|v-S�V�,^SgA�y�E���]�IS�3:�W���.��l���ώ�����3�S7�'P�h꧅�L��i�t��n��l�1fʺ	�<pO��(mٍŖ�����$� c�������`X�%�w����fUH�n��L��#� yxH���5fO~
�l߇ʠ5�=y�Q�v�\Ky�ܪ��M-����=��ϼ{�6Ĺ2r�ĉ"8D��z�ɻ����r߃���%ͻ9D/pd��i�a�"���KI�|�$>��@��y�1ǁAN�ܓ@6���6��܆1LŖ�N��p�uSE2���|����ӻQ�"t���ٺ�2�VQ>��c��ob�`S�a�`�V��(�358�u�L�Wõ���'�WPPB���@w�T�N�������P����y�4nW�%�z���8J)f�4x2�x~�0X&1�ԣ8��o��m�ѳ8�����(�/a��C(�ۏp��zŁXVAϕ��=���X]X���yTgo�o/b` ���C�=�X�vG�HΝ�����o��f��L��a逢٬����IƆeɐ��I<�V>�m�OH��Q�����o�&~�W���[���_���ZC��|��O���a�9I�
�H�T�"J�ΜE�տ�r�

^������Ϣ��a�h��2j�����(��0�.�2�vc���re��n�o���9����۱��G�L�28	�$-��5��)��2$�00-}~BȖ�^[ÕK%��Κ�ZZJҒ��)� �Y|��\�(�[�e�}�.8�,Նf��<\6��։�5`fl�A,�!��B���v#�/�airv��S~fAS���W�HS���Y_�]�ܘE��ch]<�����
an���#G�)���$�#-7�O������uS�E�&~���pu��w���{o���\�|q��s��kY�uئ�z0ןb�D�����7R��j�%����: N3���\�I��'�h@�E�yÐC?n�����u��l�(��@f�ep��:c�X�u��:ضw�� �G�g0���L>Q����!�q�X����/�gu�
���deN	�#Sc#(�!�g?G�׀sg0���\˅�r���G�X�L��=k����<;�<��<�M�ahj+��(Ƨ�cx�$������U�rvF�Ѣ���0D�L�@��%mt�t�D����.�D�vt�[���}enj�)���S}9��'�>��qB�ʿ�t��3B�(��x�����NԜP�"4N�i�Nʓ�/�`gӰ�{�����Dk���ɋ�@\�6T�gt�0�֮����O�z��FE`�r)7�aaF��=�4�8}�(�a};�hx���?�5�~�9(�atz*�FF��D6B]u&ì���5<�6^�sh�9j��0@1�t�ewo"��`xu,_:�ӯ���[PWk�t��X,�(E�5��Bld��"�Ε��j��q�^x;�-HT�$~�e�j�GD�*����ў'���9s�65����(|n��&���mdIm'^�.�}�by7BΏAl�uaX��R�r:N @��*�Kc��0�oă��-lz�K���X�b	"������2��?�¥h�/Ij��@�-D�2�������`�:��I�V��-\z�U\x�i夎x� �m�*��%���I�"HB�b��+p�E�Sx�����_�"�ڡ����<,-��LV�K3g	�&�u�!M�	&��n�i��K�m!�50�7���'?ŉ����W��j�q�ɦK=逄H�$r��&�K6��C�g�X�U�����/cx�(cX�	�JҊ)�-�W��
�A�܂*����SU6I�S�����L��6U��fp�՟�ƇoC�UQQd��2���	�2)X�[�EX&�Ϩ���KG���=����繗�Pm�P�3L_� ��Ϙ����$�3z�G�te���������P����R��r�����8�ӿ�{��]E%������&����ec�.�L�U߯�Ǝ�P�${e1t��u�*!3�T�W�'�8.J�
9��Q<���)�-���>��_�={�������1���Xca�+ö�0U�/�Y����l�o��ʝ��/�B9���=;q��%D���.><z�����x�����)�'�x^�A���6����k�j��R�3����O/Q�c��~�ۯ�w~���:� Ԛ�^�\9�s�*C���y��+�	ѽ�-l�	� 8w�w�Dr��l�:z�֖)L��e`�> 1�3W1����/]ƈ4^M��U�=��^|`�j�sq����D�di>�ߏ�'� ��J���Q�R#�L�D���6�t/�x`uu�+U��L䆷Z]�����.©-B�b<�䣘ذ�a�:���]��3%�n@~x-�í�Y kcp��J����`Z("�̙�Q��H��޻��X�{�3�Ŏ<�yf#�f���,�|�օ��:Uĺ}z�����
T�'f)����#K����G��)�/�l_��4{����O���{����/]��n�Rc(�b��/�v(�H�r�ˍ�kn~��V��6|�3��B����ty�n����!/�d�M���n4뺨�.Jqr��
H���ۄv�����9Loل�۷`�p��K9!⏇(��O�B�H��Y�V�b�-���h6�y�6{�nDEP;~k���SgP\�"�E+�k��*�,��6ږ����:���?g��ih):�7m���P��
�2������	����#�f!�ծe��{R� mb{bH��������V�f`�>�+wp��Oq��	X��n �v�K����4E�Q5�"����&�#��[�#��Ïb��/��NW0oc�lf��֓@��`q�-���������m�Be�2rf����ZY���a��Y�~���\?��$�ˍ�8��%5�*����H����g�
�|�l�|G^�M��y+�V�(I��ŉ)��	*�YVV���>���	��&�pi醘Ɩn�"g0t�Em�"�}�����"rN��,>�Q�V55����IE'r��p�I�D���Q?��a<��� ���	�`O�i��!�>�j��L�5�K���5i��i!�~�Б�d�0��X�t��軨]���� �E0\���n�b~��b��[З	��XhƥjZӏ?���};v�k��ashf�Y2��6M�ːT��������Gؒ� 1�{��B�%��뗱p�s�|�:7g`;Nj�fPC�8і��uJ#>�)��!��5Rg��0DP*�G�؞]x�[_���=h#�Z��zy���,�^1Ԝ)FZ����dB-},�W�(�g�
���K��`��ii�g??wyQP�Y��Ġ;L?5�p-��ܤq9�!6��R��5t�0�k?&>���}�q z��zg�R��)a��{��:�&Q�Ӕ�i)=��gz���E�R�.����pί��E��A���_'��Q��M*E}b	�M@�k�s�,Qȶ��8F�RAy�^��+�<p����JC6tY� %0��
r/I�+7~��*��%ȨYX�	�T�ă������p�4���{�,�	�\d"&I0�{0� ��(Al�ů�J�F���Œ�B#���&����U����u�4�=r���������E�ݟ�?X�tn�A��N�͗q�k/b-�`d
(�+";�g�a�^��V���7f0w�*��=95�=��ZL��6>��8��/��ӧ.@SMd���]���z��gR�ҧ��4$l!
�u�-�4Yr_p�*�"��Y���P.��=4-���d�cR�W���J�C0�9��O /N	���g�����Y��}ʭ�к-���L��0��%�?�����Cn�&aPǼWGf����𓀒E4��3?}���Z!6>������e�]��	B��  
Eɍ��.Q�I(�N��jƦ�^0�D�6깰����=�9n�=��[X?6�W~�1�u�N�7�©-������0�lߍ��P��g��Gyz<��d[�x�\^�`|����!�S&����V�� �tBXh��6=�0:�[s�;�����9�P� �����@;p@�.��3�d�����/~M��V�Z���~�7����̝-�6��w��A1h�K��4��9H�S�[��}��y(9%�:���!����Q(RްL�H4Ml�&!y��j��,�FEC�ɖ�;�@o��{�2ɗ��G=WF8>�%/�Q�a��}ؿ{;*����MNQ�K0$�8=c!CV�D���@�f���Wp��U�M���#j����X��kH�]F��F�x��QttT�����a1�Ј�"�[E��� �R�4�~I��v� ?P���		)���k�T��>���t`�*��4k�h��)��4��Q�{z��@&�������}�2�.2|��{��Ed��ҋ�I��Sp���,�!?�	/�����\����Mo݁V��r�����ܴ�eE���(?e"�jX\P�EJ��|.�^/��j�K(����ʱ�������u{=���."�#�B/"m�/������W��� ���7b�����C62�&�bv� zT)X�H�"�bs`����f+��L�=��zu�UL�K�,������͏߇�� �Հ�ŰӅ�#�8M�.�0B")I�"�a�Lﵟ����m+&����=�k�6���>W�rJ �ɝ�n����5�ih��.��dU�=̟;�s．��g���i �B����P���7~B�	R�������AbX`��X9��������_E�ݨ�z]��g��Wi���ס�AU$���M�Y`'$~i�Z weg�}3�?E��-�E�=Z��=IҦ@�q�[JJ�U��3$T�T*l�@	-K�W�a���W��ʶ���jh6���Ɇ+_�	�F�%:R�ҭ���M3C�z�T��PQ�深p�ν�*�N}�VC�l��b-*�U&ٜjz�X�e;#�Fܚ�q����6��.*�va�s_���G���ǰ%I���>&���sB����񾒦����`27>����-�8q���3?�݆ỂL�u����+�Zh�ʹc��'�}�sd���8	`��Q����ai��%���!v�-�^�M�����'�A��):2��8�q9;Fجc��i���Cܹpfہ�p`�h�s*�Ct7@6��CV����(���B���Fb�Z	�~k�/X�M�s�C�F�����tp/��o~��DE4�]�_����So���:�����|�H�Q�vQ�BQ����#r�E�mܹ~3W.�z���%�Jؽo7*�Ò	@����������h�	%�3B����ad�g�&�ܸu����i@(����B�hՊM	1���q`�ndmʴ)�k5�rEL�߀u<�7l�]�L�)��H������q�~v
+ￏx�6�^n�D��>l�+���L����~�XׯaX�ꮠK�-1������IX��ҫoHS`k&oA�����) [�Y�wp�p��F2D�����RY*����PJF�!B	nI��(k������q���q��yl���<-x�Z��Fu̖�]�05���X�7$�1�� �;X�gJ��F�߷P�gH���ؽ'�K�9�
">Ӯ�㊀��^ܙG��c��;�BgUrL��!���z� !�T�5���}�������|Q��_��h����G/��?��O�:���E0�͆J�#q��`�����s,"�X�4�i����ȃB��2�M'E���?�NOms2�
=��KvE3�a���%�u��,�!����#1�c��y��p�%t��Ŷ�[�q�$6��nd�z��&G���X�����+趍V�biu���5W11Xƾ��@�zo����?�qs�jf/I�0|�f3�Y��*V5U#F#te0s�0`IZ�5���bx�6I�e��re�R%-"}ʚ��DN�<&H��%7>�L[�����"��
�z�ٛ��x���A�7�s#�>i)��M�@?8$�T��i!�g����%��0F<�O?���8j���2��q�t��4͌��>+��j�XC�>��hc~����e937o����
V/���w_C��e�*�
���rr˕9�e,�h�l����><�?�S#���K�
��i;�<�,v=��h��'���+��&�Dԑͭ���=�R��k���cjp ��[���[���c�6���}���c��i!p�Ӹ)�������Ȓ�$*%)�,�#�����������ȌM��p���Q�0���־f����f�W�#/nh()�E]��\���_ŵ�>��k�b��)q"���;`��/5�V����M�,<�-�p��C\��a
;�x;�y�T�j*�Q���DGF�HY̰@Nl����ߤ���j�"�)���](�n�:��G?���k���l�}?7$+\���bA���1�78�l��N!�m4�݌���(v<�~�e�Û�p5t|JZ")�(34y���4b��SpUy㞇�����qk7/��'�6Ν�E��U/�曃n�����ܲhpd��朔#^�T�A�1�eCEhi�p� �=�<M�͚�������%݂n��o�̃�2eT�AEln�Zw���,/��;oa��)tg�Ă���̉I��U+��jD���
�F��W�TK66 �M����b�tw    IDAT�FƱn��|�	L���2\I�ӥXKb��H�A2�����ů!��ʉOp���z�6�Ny�d� �$�����P<g���m�u��Xb�����=y����Jc����Xq��$��?f�@�����ڱ�� @��O���W ���M|��w�:�؅����ˏ��W�����C�����d@#���,`q�.n�̈π[���c�AM�s�^kc~n��%ք�ĭ0�W�
�A�s�A�Jќ�L2i7I$���k�B�$�k����#�ۑ�
\�-�C�ە̡u���ތu015-2"��ĭ3���VJ��\�r�����4��ρW�B?�{��ul
�gq�?A|�2���k0�La�_���V�z8�����1�~Mcꑽ�wmEX*��t�ں�:�K��f@�l�����#��0ͭ����X4㳖���@kq7O����a��U�9l�C���I ZAQQ�0���.�KX���F��駠n�	�Jo��~O��!(eM}l���dtOB���@���44�Snj��K`vޱX:~��
��mb��;�� G'ɾ�[�?�V*wI%����uS�_}	�X?������~�����ǎ4�]����C�R����B��OP`쐥`J�)�%5�ޓ�́� ]�I@yv8��RY	u�4cQ�Ír>P�� e��gp[@����8�۲	#e�Er�֮\�;� �56�phwUC��cE���nC�Zرk�|�	��O"NL1e����8i-db�b��x|Y�XZ���KgQ4c�߸��C��ױ��Q8gfP�yȵ|�s�P͘�&ִ���Q���̍c�+e,�vN�����3���s�C/�037�Z�+�� �ƧdE��P!��k�.��I�ʨ0Mj���u��:�u����ڳ��a��"��L�?�rg5��)E�)�<dIZ�A�ů�T�=G����0�b�|�ey�iOO���h12�A�,3��\&_s�L-�ۓ$%X�zwn�B�ހ�;ظa��La��:58G?��Ӱu�(;�):�O�Jd9�&�u�%��z�A�i�j_#�0Fl��x犈J��������66>p���u1���EjZYd�9a��1H��馣�nam�*f�Nsa��}��P�B�}��������]�ݮ�qB�"��Z6ȩo&��ӌ��F�i�ŭG�1�g2��
��8����g��+�8!:~�N�G�8Mf}�Y!��e�-��*C�4J>B!X%��3�p�؇��чH�u�~6ю͏�I�+C�d�p���ϖ�?7'�Г����ʡC*O����)�}�K���C�H�a�%�w<�%�pv�0)���]��J�dH.��
��n��g�q��O.� �(jb)���Ag1JCpr�zA$-�E��#k�(�X|&p؈R���	�|���Uz�+�O�JE�n�^O�W^ߐ�D�d���CvP��[ǵ3�����D���q;5�Pz�H�� ����>"u�|H(I�xA�Ȕ?Ro��ڦ�`S��b���a���y�ID T��tU�P�3 �����r �o
��u�+�x�$��8��kHH)sz�)��	Is���"�d��XL��d��7��rP���~q�C��H5��`?F=V0}��x䥗1�kԡa ���2�1�N��XP�T3�J�xv�.�Wq��q|�ΛX�=��b��;R$��fa�P:�Cw]�c83 �e�,�мE��J4��'�^�mIZ+"t\�c_rC=�\�F�mb�	��Sx��~��= .ý8���������d�������/H��	q&	�γ��ׯ����0�!	{�UัP��k�vI_<�vO|�p#������<�V&ͳY&�PQ�ƞן�;�ꄃ�Di�'tQo�!=�n�y"bM9?9q��R�13	�F��,��!����M��|�m��<����~�}$�y �_�md�����ǧ��_� ��gP;�:�a�{w��7~c�|�#Xv����G�|�ux�9�m��vcp�6$��j]i��F�s}�c*O��t?M�z/���V�`ddTB�(id#[[Z�ҵkX�6���2�@��wI��i ������Ů�aU�0�g;�|�(;� 側��b��]�uH����}��`�X(R]�PA�g��j�5`�
�����@Y^�f��D�}ې=���zD��w�\���f�|Q*�_7_�o��9w����k���W_��+ot�|���rS@Y�Cq� m�/55��So�=�˽-ٽ4Xa�r�LW�'/�Q� �FJi�� 2�9�O���$�H��r��:��e�>:/`��q`i	*�:�ؓ�(�lX�z�v�aaӶ�p��lݲS���e����O�y�ǻ��jcՅ�Ȇ=�B�Ҍ˗����X9qV�C�ס4Sd�Eԩ�C ��1��5���]�C�Q��S2bY�Ii�ݾ�}�%<���h;��.�ҵ;0�"���Bq`XQ<Rbz�����d��F�ؼ~Y]G��M\?u?9���
��*�FG&�e[�ߋ@���0��0���*�Tߛ�S�c���dJ� �6'��
Tʜ����'���C�CH4� �H�ݕ�N>k����$n�D�,�WW� ��Sc�:\F�]���}�diF�������&�,�t��{q�������.A�J�+�$
���|�۷a��O`��!;�~�n/��r]H="{R����S&�Q /�N����Bu�d��;3���?D���H�h4�>@m��<)o�g�D)`�h�����')s�RON�"�a���z
��[9�D(�uBt=++m	e�s���P=l\?� qą3?���?��g'���l���ʤ`��#h����O�.�e��e���gz]x�΢�~	U)P+��5=���)��3�MM��@:jG�!Y�J tDXW� osr�@�t7.����gp��ed��^Ӌa���.��&�+����JD@"�ս�jq�P�ؗ&������E nȠ;@)bl�n�z����C��uC����'d�mI�g�6Jy�ӄ�VEk�&n_���}���]�n#�r�qw<�=ph��
&JM�")��JK7�Ds��i�T����J�P������`྽��S�~��q0��m�JA�<��\SE]W�?�U�^���K�p��y(�.�=��;i`]�jn}�j��ds�L3����d�L��fD��A.'2OzF@ɭ3�I�Y!�K7���`㡽�>���qT�����Xy,�<d�c �Ta�[]ĭ3'�x�7�`u�*��C�:l/D^�@u"9�
�!�%]C�ȡ���g�(��'���������n�����4�*�������"�����ھE���/�#���7��_�n��c���G�Aـ9����$�\N~�!Co�"g�:���\0�`J3'4<�_��bes��&a�rEB!C�1�z��;��R ���7�ߔ�1����~l26���#h10��xLH#�#�H�*��D�^�����q�!5.�}����BdU%UGE���j֨KC�н�{����"�{'h�������b�臨�l���).�M�x��oc�7�1P�3���������܆]T����8����ݮ���Im�3�_$��|_��d�h��n�ҀL�	�b�bA�yn���A6V�ub�B�D���j	r
P�U����ϊ4aM�Q�o;&س�@
�7�
%%��q�x/�ǧ��O���1Ri*�q
T��h@V��j[�����X<��d3
z#9��E��C���#�ލ���ˣ3����#~��R.�㇬ͽ7�����{����}�Ҭ�j'����ATԚ�����>�������/	I�#?��<*}�_����'����f2�������w؁;4�q�UŶ��8�w'���vjh�?���g`,�	f3��q4�YDc��&Ǡ��	�/�mdrC(�`t�:JE����Ea�^�'�ד�nC�v#���-�]+�/��h]��d�;Ƞ��t/FL��П q��~#3Bh%�1:�p}4�k�@`��QNQ,`x�f	1�s�ao،�̯6jY��eB�Z�"���H���r�e���������]�A��K��	���ۓIR<���wF9W�^&q��PK���q-5��J�.�?�Fb�Q�����Ķ�`|�6I��5���繧#�9�|5�kBwW:�5p�kP�F��J�l��ε����Ak���B��CӤI�W��:�'?V�KT�T���h����3�C�~�,SC����0��0��>l�u2�Ι vʘ�_�S�N�=9�-4juawW*i�ݹx��ݾ�x��x���V��bvA=�U���K��FM�5��Z��n�ŷx�Q��UA7	�e30�FP�ވ�]�0��>nڊ��G/��*�d��	�����b����M,_����ѾyXZE��0�*��/W�$���齦��1_�iS@x?���9~�F�Ϲ�����{݀W� �n=F�ۅ�����Q�f��sA&w6+�A��"w���|ͥ;X�}��E)V3���`�F�5����7�&��U��8��k_��F��G,2������H�i�xd�0FGP޴Û6!?<���:G'��V(C!��gX���Ǐ�⻯�[Z@��wm9�y;#Ms��^�k&�_���I��%��=�yY�2P�dY(f,�4�*:���c���0F�g��z7n,�Fcbr�F���D��`qa�Z���F��@�Zȑ%EP�e0�{����R(K���O<�y<�hT���k��)ic��O����0���@���T�z�<{�@��F6Mab�l9x��r�cP�"d\?~��/�p�4�n[2�$ߥ�y6����(�=�z8����5(>q�)�&�H��c!C]��F����Gd�%�4���F��F��^VEa�}x���-�~	�c����x�{?@����a����{�q�i�O��U�L�{z�	zR��iV3����D�]�]ܿ��؋����S��Ό���HQ���aO��Ѷ�|eeVf^<�r/����Dhv�P�I�MUf~������!C"=a�F?������Y�c����4�W��p9'�r	Mדs�	�65
�R�!�9���D�|�%�yl
X��Fh��Qc�j�S$n�(�j0�Sy�d	�MW�4�$	,�1p�A#Fh��?���Bɦ�hxO����#�"M���J����K6��~�/��l��������y��#��7=$b�]_ņ{�,C0���_��GE��iD�"2l�S���|�l˒F�{N���$P�&���}4��]xBE�| �-�E�J!g�Х��
u�nC�z[o����а���~�(D���yH�[���b��s;,	j��&��
�|ϓ3�:�}�A
����^�h��hI��1}���M���!8wyR���}Xx�H^��T^�xEK�~T(����"��6�}y=x��+p��7�=�����o��s�l���)H�f�qC��Qtǉ�2�[-��ǝtc���&��`�KM� ,C�ye|=����Pſ
�	��B�S���hcZX2D��"L�S��Q��5dC�T�����)�@/�˖@���T=f&���H�H�u�jh��fK�U��
�4�b��V���C�pv�L���`H\zr�H��� ���(��CX,��Y+�tKHXmI�#A	f��n�Z�		m��Ѷh�4�-[���7"K����\�>��6�:Z^i;+D�������p���g�0�l7���:��a�	�i�l���	7U�/�?}I�&�KeA�	'�1�B�|K�����^�#�7�o�2�,��� ���7�k�a9�|�t� �f�5�΢u�$��1�3S0*��G��kIC��")��MK(O,��P� ��lX���u�4_\d���,�u����W`źMHz����({9��)�f��\q���c՚��v,�>?
��YTO�CT,���G�6f�%q�a�G�Q"+D�"A6|i�ؘIc,��)s"�d�w� ����|�B�J���B��aiz��^�Ī[Ѭ�p�62Y=�����kϢ2v�l=0Q�u�u��ul�q�y�b��<����=�U`5-�L����@7bk��&����7�P�}A�����vR�O�7_��ۮC�E��m�9(���Wva�+�C�N!���[Q,&�6ȑ+�T��_�*I���Ĕ'������fG {>��])��5���X�Ҽ(���[��`�.Y���mǂ͛�� 2)�p:>�W|�_V����V�Hs��e��Aẹ�P�x�H�d�,&8L�es�j��xԲD�V
Y�Aְ�_(�N$�[���n>�r�P����pjt��@��O���l�Y0�TY��ƞ6�Y3�S�1͂<�4��X������dZhC��HI�E�"��E�O������ﳓ�@�}�d]��p�zd��{,ݺ	[o��+�"��$�&ŉw��k�?��c'�5A�r�!��(h!�$��Z6�)"ゥ��v�ဩ���*C���ъ�Ҥ(��B�y�p�!�q��0�(�\TZU43�[�c�}߂��z4�&&��ñ���u~�㘚G`Hw�`R~���,
�~�����iLN�#��ȤH�Ѭu���4..LN�Ɖ�x16���jJ�:~�0�Z	Y��C���6�-�b��&��B����D��!�7$Z��f�F�h0�.Rq��:*�9��)V�ٜ�tPs��:����)Lp��h��$mG2i�f�)��7o�f���l�������;nC�� 4݁{�$^�78�D�V	�7�&�p�z�f��x�7�Z�a��������xsgN"�����4�Ź*f�sҰ�a"��dڅ���N:V�T��F9�"OQ@�5ȥ�+d���S{��B�h��L�ֵM$��;h �����D����BL����x)�y� ҋ`H�G�^G"͍jM�|M�XPE.4����p'n��4�\?��9=���,�g� �{�˦�	͘߅�+�B[>����+�N�(�=�M�?���÷��\���[�ӟ�����wE����Z)��a�U�	��S�9n���f v����ur�JؖL��'qi�=�
G��'�S`�>��'l�
t*��尸��l��4�hz
��A��W��˦�|���B�y�0z�P3xPef�h&HV\y
+I��C��KCW�/���4g�8�Ǝ�BB���ׇ�7"�p!��' �{���P,b��è|~�����aJ���h�"Lm̸-��N4�1���#'�rP��2�E���6^*�@���܌js��쓏pl�'�(,�X4�8uf~���,�W��b�%!^ؔ�J�'�|�tD�E�21��1�w���v(x�xd�ZYh�6�\�"�4�|^<�=?@�ZG��b��-�x�r�&N����(ڇ��,�-t���l���<"�f*�r�g��M��*�&�Kl���&�-�G���^i�.��OY��]bS������[�Pk4�w��	5S����waɲ��L$'ǐu�H�]D�2��)�f��J3P$��іգ�N���1�X�k���P�l��Ta��s
�fc�|�� U�B�\�\�;w~���бt��,�����o��֑m9:��t�_���Su���u�l��9�a��%}Xx�1eV
lu��������H���\��J���pa��Fb�UW����D����M-D8u/?���9�C�]8R� �U�[����OR$��wf�]��bv6���`1P���S���Q�M��r�Y2Qe._���w���mW 7�'B~�J0V��O<��G>�A��O�{��n��z"���nK�MR�H���{̼�i�a ��)�FW2'�9�TNh��4��6Z��L$����R�x��D�G��i*-�NZ��,�t	2,�����vF��Ĳ�	ym	�p�\����|���@���I��-�w&�J^3�����д��W����<ñnX    IDAT6��4lݔ��V��D�@j0����ż��o$P-�qj�a�9��XGX��(֦5��-]��(�I:}��ܥE��!RQZ?vSS�mæp�W�&�81��#+Бz^�$��-�dZ�'M���m�6���[�V_�@���iWZ�*f&�0S�&��|Nʑ�!��V�t^��r�,)9�D��heɇ��M�4L�Ф�H))����xhNO��=��!�=Y�I;˚ v��D�ۺ�������µ��12]�AI��%I��sHS�T�9 "��de�WRp�*s(�����9�t�rذdsrv&��{�����tw���H��%m":|o��a�z�-�Yh�,�ZaWkv܄�_�:r�7z�����O��-΢�M�n�fu���0>5))C2�zR\�R���_3�z�.�YD�L�L뢽��SHe��g�ڏ�Cubf��{��y��9���$��� ��]�a�4��eː]���pE7�B�T��rM�
[��Q��?���:�I���L��-3��I;	�hg���^E:6`��H邘X��\Z�� |N�e~���?���"W������Ϳ�?~��϶��'Y��T���2]��MC��	q#d��L�)�숍��[�)Z�x�b��mv�l���dJ؝_+:ir����O�pI{,�h"��a�53��K-���P*��n	w�|�vʀѕ�������yp����'�qh�Q�\yI�,9&Ҧ!��.ǆW���Ә��E�Ѝ�k6bh�2�� �q�$��������O�?��o���O`�^�I:�%�F�`��ު�M�KY�I�ù� �"+�yް�}����CwO�|gOǫ/����}�
������R���MNE�*Znb�#^C�*��HQ��(J=b�bJ���.���N[��.�$�!0IH:��A礑���:�g�0==#.�7l�u7߂U+W�9;���1yp?�����61  p"�D�}M�)Sv�7� �B���K!tm�xЅ�J���f��
O����t�	���@����B+H^w>���,��S��%��,�=L'1�Ԁy�#�)VÖ�Z�F�ҥx+��#�8�'Ť ��;�� ����&��Ů�����n��s�͢�p���JI�ذ�6^���>O��D�O^{�OBب	%C��m�UAϢY5l�$�,.�Ua-yR<��b�,�iU%ͣ<kj�
-C��54�*��M{�Z�O�#�Hf�0�(�O�������!~9&S3�Ɖ�M2�W�a�A��&�)ֶ�҅�~���_r%��FG5���a���=�[vB�h��Xf�ZZ(N4E��t1V�_���.$�6\RK�q�835)͜N!�d,�\�k��?�x����H+�8"��b�(��ؼ��Dq�ȧrH's��z1G1g�D��t���NL���1�60Y3]*W�P/O�J76���vd+S�CNo#ᖥ���&i&4)�KH3L�s�E����"��;z�4�1[�Pt��3}Hu�ʬ�S�i)KG4M�"F餥Y��2�j���L��0ua�y$��P�T�>.=��LZK��E�&CC^w��Ɂ��mB"��&�4C���5hɊ+/(���1�e§��Ndv�j�n	6l�1�Ւ��Sv�����j�Fr�*��x3�f`�%������mF���Z���/�%�d�Ӳ�֤�Q�!��n%�0�b>��&�U��+?�{|�ƛ�%�,i;J�3,p�X]=�]���y�����(�$�&y�c1�$DI���}g���j��b��I2���k�$a���0�Tׂס�������O�ݰ�*L������a��;q�]��Y�03h74��09	:�{��x��ʨ4�2�L%HÖ�Z�9"$n���݄�dQ_`B��!Y�zf�@�G{���~��＆�x^�9���t���rO��C��Q��
���<�`#L^K��I�b3.��#>�Rj7xi�tH�;e��,v�b�$h!<$؄������y���⛔�g�L�ϵ?X���������C{_X�������}�5�ɼ��d�G4��r1��SM��,�Le�(ݯpѕ���,����J��CC�t��>�E\dX����Rhp��d��Q_��B`0l!���o�-RH�[$��-z.ڤ9�F�����F��%�Y��U+��!��+%��z���j�]-�5q��	�;uՆ�������X�H���P.NnK����"��#5���| ���C��71��K���ɘ��t
�PǬ��j�AKbwp~HP�\}}}X�|)�ѝ�#�N�N����{����S0BKDȥ��0� 74�-[6	z0y�8��Ieh��*AR�:.��ƫA�f��t�O�{&Qܸx�l�FK
t�%SY4�=y��e�N,�t+�T�
fJe�LQ-���߇�EK�`�<IJM���a��Q9|�ٳ��f�=�w!*�G���t �Ň<�0�M�HP9͉�ƌ��B��m*C�s%��A�+
ʈZ�6�n��V '�+�K?,33ӂf/X�l��'�15[A��Ƃ��!���p0�M#���5�P�H�)�0k��S���.]e�\����B����b�p���%T�p������������$�5�ļ�E�H�����$��FEC�I�I_���v�oRVZ�Y�/%�es�Ƌ/���c�!�;~0X���5z��L���U��Q�E�n�ũ, ѕC���dw^���+����\�*{)7DE �s��麧�o�dgL1�\;��O0���`l���I7m%J����;�7�[>_����1W8j��)`x�|葇���@!�!�S�&J���.${ze�Z+�b��y�UC��#�A��S�����g��<�������t���LnOȵ1�YD�,\#	3�-�����Y���G��.X�܊u�/\[C�c��"uQ�
 �E��H��W����F���5؇��T� �S�̝Bw�auB=�Fb!�� �F��"͉(z��b��c��7a�ڭ��$M�RY<�)]B�L���9���g�Q<7�Y_�'���0�m��+�V���f��'q��Q�V=�ѽd9�z����U������+�^��#W�A�4�LeI�&���|^�0�����o�ˀ\/�GGa�8�4�H�)���]�6|ֿ)մg�
tm��p)�.��]A�� �
_lR�����?KD��{);v^&�k˯g�+M,�..�Y\}����4�y����h+�EH8Z�� �qot���пl9.�i'��]-�*�YlƜ9��rh�d���me�3�ޟ�4��lGG$�����CG�����v,Rk��+���O���o����A��BƦ3VŠ����ن���M�L�����y�˕JԔ�YmB�_R��>d#��Y�w~';��|��W~3����g���ȓ8��ps��Ј�S	�/d��&�5FҀ�d12LY޸	�����:�?[\���R�]�;6�qx�4��F�yV��T�'�^n�a��f���bL��I�Ja�����?e��!����
�_���Ί������՗_��u=��)��鋮R�6�<�� -���#�� '��Ǯ�J�(� �%���-r�qf��Xb�G�q6 h֙���`�r���(�@����@�o�U�C����a-�~Zҹ�!ȇ��(ք��0��H��p��-��L
,N��6И��73�d����4�檰z����;���k@� �gO`�WQ;uF���\�N��|7�e�����^�I%�؏����ۯ�ć��F*7P�}�[�<W�I;�Icb*"Q���@O�Ƣ�A�fRH��l�u妇�bc%Tj!�mu'���#���q��m�8z�<�$&�C�36'�>K1Jn�����]"U�bP�9����S���K�:K�����@�L��
Pn��[�
���,��f�+/g3�-����C:�RD,�@�|_h`��������=��Md�P&����B���mmD2=,�d* ����\-���fBc!����mV�����B�Vװ�^�e6bx���Y���b�޽X�hۮߎ���p��=����� �z�ӧ����ϭ�IrLJK(��P����	|L���D
�xḘ(9"��B]H:����>�!:�T/�\�%+���j`���H5k���P���ⓒ��}��\ZH&��\��о��*�6}cTѢ��_�u�����4���;�Dr�����p=U����3�'26Rv
f��L�řR	�n��@#�E�aۀ�0)�x<��_��E���O�0���O�1�v�֗���c� C���mN�6�
(�8K�|�flٴ��8&��$m~�>jXp�{�^��%����fifJ�Ǝ�Cc�$���-���l
6���+/��|�AH��N
y�FҲ�nG�,�wy�&-\.4�3Ǐ��G�JE��� �l�kv�)�cZ�R��iy�VA�3�*8��OȰc��gx�g?AejW]}���V�4���U�{�wH�U���eXx���_���Y�:�!&?{���������'��WoRʖ��`A� 8§R�i"ߍP�*�+�H�К���]O��Ob��1�ۋ����w��0�����_�3O>���0.��&���F����;��%Ǝƚ�[���{еn+P�!8�)f�����1�*��2�X�dm�	D=��,Y��57 ����̾�33B�I��u�^D�1�5�e;B�x��7�X����p�΢:�Sj�&����5o�^��1 Eڙ/�9�`��4��REPS�L�7�ND:��������jc�8��G�8z� B�bJ�'t	.ď��¤���V_q	m��RRE�����@G:�V�����w)!<�$��ى���I=�|��*�.�"�M�,N^�T�WC@��0���c�p��}��C�hX"BM+c�9-t��eK���kѷv�d���rN�9h�~�"��/5;r8)�r��s�ΆA�,��	���t�	e��&�0�j��h%�ӳ����b �3�aUr2
���T]l��-��m�0l6����n6����`1/4jN�9��]59D��Y��a��B_�}�?1�ň�6�~~��d_�Ѧ{��լ��i'Boh�{V����m��(	��~�܇��.���7���������󻮦��N,��N��h>,���$=�M�W��V���PHL�?�-A�OJk6bsɔM~�e�"�ȶ%}ѧHM�U�2�ń��a�e�֧C��6Jh4KZ����"��6��` 6r,v#z3��x�SL�s���0��p�WA��VE�o!O~�
�8Ƣ��}�ׁt���μ�8�g�:�`�t��^�48���}���
����B���0�����,V��
�zS���^��eL��rS$�5Eo�Z)h�g�O9H�T+ZZ�}��/{��z�mk���a�[q������P=��?�$��"���)#悋�[8��c����`�ʍ-�Zp;�o3�-EI�Mx�&�fZ���M��l��&\v�-@WA2�f�����w�Ȏ��lH���L���8}������ko ը"���xx�X�F�!�"���!�S
�z/�T���k��з���Pf@��ܚX��r�ID�nl�i'.��$� E>��~��y�.Ŏ�r�PqPm�)ѳ���C�u�3(��+e�k�e�E�59�Z=��CE#�I!m��à� ��@�K���&}��T�[o��'/���͛���[�Z� ;��ｃ��y$� N[��\S� e�F�?�I@�-X��1
+��c��҆�Y��TSpq��u\��&V¢0P�A�*�1qT ��2�J'��y��d�wC�mb�����n�#7=�ГN�hU`jLVs�l�<��r��|Ң�P�V��S�����G�'��:��6;��nS� ��CYOa�����`/�Oc��_7����WlC��7#�'���Q�ƙ�q����k�0sd/�̠f3�ͽL�R��p��Dc4d�����bQ��t�ڰ	�-��֪�cto<����L���p�]wa�]�J��"$r���U�|ē �/��,��G���Gyfw�u/.����F?x����P�p鄆�WlǦ۾�Ԧ��2��z���fΝ@�ЅeWmå��z/�\��Y,6�Ш)h�[H��R)����� ��*M���4>�S�1�0�|9�o�!6�g�y�>�4�C����{��޻1s��?�G�|�K���~�O�ޠ
�}{p��g�ڿ}~yKC�5Qm5Q%�:�A��k�2̻�.`�j��ǹǞ�sa�[C��n��� �-�t�J��'����~	�d&B�[�JI���ǫ7�eF	�5)�YT���{-��s�"��nK�_��<3)&OdR�X��p�Zt��V��X�7]�^m��N�6MEQl��x��#Z@����\N>���!�����b���I�L�d:!H$��.)7��"Z��vcR+C�ؼ�Ҟ�1��T2�d*�j�7�`�l	ΣU��jЧH49ô�C�n�5���pu��yY�R���z*Q�m�g(��L"��Bq���v��m����1��� Y�0���|�Q#]��5�Xl�[�O�ќnb�������-#�0��hS �2�ñ�D�&���Fg��D��x�Uހ/��kó��� �L�+�����r�
�qMQ0��EG�CTs���'��������|�+�?���k~4����ߗ��M��˝�g��(��Ӈ�l��/���^ziM�R�l�#�j1Q`$������|\qWa]��'�A��*���_�`0tG&�t���K�m�o\9�H������	 =�٘h:C���Ѫ�w���Q����ɡ�q`��0Bɴ�l�G'���6G�U�?
�Et���=���1`~�*��q+���*��O=��=�c�@����s���\&�Ů,�n���}?���3���#���C"j�$u�m�Hg��pέ���4��.�1ǐ":���"C\I
��)�eT��6]'q���\dbʏ����o܃;���;��������6'�*�I�$I0U���+O)�x@�ȅ���z��#e�`5���t�tG8�%&��pFз|	��.���tZ��k��G�#,Ob��)|>:���K���˥Al?�]?�N��2r-O,�,�����f'�rI'#r�OX�N�}��<�Fr��ztx�-:��B=eߕ��+^�j���K�ĭ?�sd.�h`f{�x>ލEk�a�W�{�* j�������ud/Lbi:���'���y�c�n����l�12q��=��f:(�}ޜ<����8Sh�� 5���XS0?����~t_y�d��L��
��!�kHYi�F'�5��:
+�cцM(�pl���:��ʸ8R�"��Iis
H�XO�%j��:ȷ̿���A`��¶j8U'�C�0+Ӈ\�0ʁ���%H�!��J�V����'pf�>d�n�*rY�ÙU�:�!jR�gV��,�8���j;by<Kc����G'�ً�}�'
�Y����e�C̻�j�ÏD�G0u����������kE�-4
B?,�[�ѓx����ȫ�0����&p%t�Dʎ;��D��M�If���-�.B��l����0x�׀��r��s���c������1�t�ܼo���娝>��S�aN]@cvF\+��U[�x�����:�������qݝ��.6�yq^���Ay�0��Kn���.R[�������3��0q� 
V��q;6�w�k��:qG��ũOv����^���d�f�[�-�Ɖ#g��a6�gFQ��L�ߏ�{�c��%X|�UH_�Ž���C��"|��߇5��l����'o������?�!ҫV��o�,N=�4?���
�a����G���C�� i��n�X�8p{�ϑ|8'�\�m��Q��ێ�"2`�A��<`w0s$*����3�b>6�?�8�sj`|Vs�����Y����0��PN���J�ܣ�HG����k�	��zB_���i�2vL@T�J�3�Q�)[�C2�    IDATt٢?�JV��(�e&�&��
�V(���>�r���
�˰��,2�v;%ַ�ɋ��I	��xp=:rq���MH��yb�a�Ҽ)-�؍��q����*��J:��!H9�+{���;���ȍ��l|�L��c� @�^�d���d����44�H�	�\G��{��|&L�Uc��(��1����J9�ɠ�V����H��4Ut3�k�%��zc���uwc�λ�[~�]�Ϭ����?��W��Q$'m�Zb��/T>:P�1��俎T�@�i�0M�R��i���W�_+LN�|sϞO��ԩ3Y.$N���jj��#�}��.(<���D��J20s��K_���/�u<����Z�����9ِ5N�Sv�j�!(m6Jި���>��e�G�\�?7�Fqa��6N�\/z����U���4k�N��ށ�l���@��!���Z2n(�",�B�y������7�d�<�����X�T&���}}�U��,��������<`t
x�=|��o%}��NR(�i�L���c���hyneN�5������,�4,Y�}Ã(��!��c�w<z�;j�-���ʠ�$�32�V�@���Ň����|��B��J�F���TbQU��TZgr�9�]ğ�&G��&9����	Ҙ4�]y4#�̜�[ʛ��[X�r�~�.v=��<�+�߁?����N8������o~��	�<n��5c���q�@5"9]C�0��Md)9@cS��<`M�B�4�V����6�zK�߁��6�Dc������Q����+��M��;(��������̛�+�����+y�'Nbi��@�Fڦ�!I����|M�@��c�k�����OHXMĔ��j
Ho���$1�#q�h�5x�x��q�7���w��`���zI�2Ӥ%a2%6׋�V�����ko��+�
��|�=����Σ�\�(3 <i
�쩦\qe;4"�$���$$�O�
	SV�1���)!Q:w����*`��-X���E����~��ѩ�b;Z
����8���ϟB}j��\�(da���ub�"̡@Nrq����Ɂ+�C�IB�=��,� վ���mPX�[��#l�\Gu���Gb��q��),��䯽X̦�����aಫo ��eB��G���a�YA�ME�1UL��(@R��#=�L"�Ή-�亐�GT'�By�V�s?���
EA	g�p�W��������n����#���'��ٽ{���5���2SX��&\s�}�_���g��������މn��8��Kx�7� �x�6+^�|����Vп�v~Jd��&�Ξǎ;�����&2+F0}�(�~�8����uY�m�������nDS3�ҋ��+׋˷\��\70>��w?�ޗ_E�`V�܆�+.Ai�A���гh�}�{��!��^z�i���3�^�7�y�񾏍a�w�`j׫p&'a{��d��;&f�i�A����z��K�b��=��0���%YA�ً�"����pl�%s��twb�ڱ��X/t�Ɏ>K�sw5T��J�%:����Y"姦����5��;���8T�3��,6�����)��q ast�baʽ�t��NhJ"(���4�IȻ2Ie
�ŔF5�q���4,^S\o��P�e�R���+�c�`5d"`�m4I�s��J\ݣ_|��ʞ�1�K�N8���t
��5�������=���oB�m��p�R�� A[���M��$�A���O�0C�8�}���X:��aꘫ�f�si�;HS��w�rt��9�b��$3�����\�(5K8?{^o�v��Ċw�[m���ߗ��HA����S�w�K\e]P-��sv�G�l4MC�S�x�������;A�'�@����fah�a�hQ���7=K�4+�"K�"��ckY1���v��0�0
me��� �B�h��j����v��4WY;15�i���)�����XH��x�"}TE��ju��F	�R*~Z�^��e�RG��4D<&�kD�d((]m�Me38GA�h�4éI6�Ī���?�Z���9���	Z���X�qv�q���O�h�8M�	�|��o���7>���)?;��r�&,��%�(Bm��u۰�������:5+r�������O�.2L<�eR�^�������g�|����]�f�W���Q�sE�՛(1���j''��9��_������[�(�@K�+��ݎ8���T���H��P{�HhW=��O?��z�sg�J&D�I��m����U��řEd�u�>���ݔ��׺c�r_%�ζQ�kM��!�T����j�5X{�5��n�	G�z	�?�0>�� 6_~%~�?�5z{rx����c��>zY�K� pZEm�lF�$Jp�,mҘ�Z)�T	d�J����D�C;�@��1�60Sw��ù��q#�e7�Ď}K���O�����7�g�������+n��~�8��q=p �^���<��a|��#���$u�g����с)��H&���|���
�"L�mR<���B:z�s&b5e�JT��o��7�?�s̻y'�,���C�c�F�b�o��l�31�F]+.���WN�Ǟ�@8}^���N��'���P�>��$P��x��zs�{��1�	b�Fh4����ĂeX��v��v3��a�����\��*wYm�\��"fΏ�t�>{��O�@����ESc(��MD���(c�(�[i����A�`��E���m�]�zп�Jl����Y����p���7~�[A}����Zq_���&^�������!GG2-����k��9�s���D))��{�#ΡF�N��>��O���?ᡇ���0Bex>V�y7�ˮ2�x0շr�~���'O`����?�6��,���ϰ�՗�-��-���.`��w㦯��W�A��Y<��?a��Y����b��7 3!N=�">|������G��#��{?Ƃ��"M�}�b�;��]��l�l�ηѿx>�N~��| {_���N�B=԰��m����b�4Zm<�����{��`��^U:tG��@��G.]�e۳/��z.��_�:���B5<}�(��'��߃E+V�K��P�;vO=���?�L���|7��.h������B��Af�<t�YBU7ڟ����o?zf7���&4�-� �k�h�m���p�sN�Y0*���E����T��O�幻�������'����̊��܋������#ğ��?�����6]�Fw�Z�Jc#�}�%��gi:l�&_���b�+k_P�>�*L��]$M��H���uf|QJ!�,�/�ʚ�pQ�������ų����*?[9��AG�������
OU��/�w��-D_�@C���`�'u�@"�|�$w�X��0�!=���f�C�[bkvA��?��cj��J2�<��Q�l:/h��<�G>�*.T��������.������\{�٦ RO՗�k8�b�U��T>O澄�$�.,F�'�(-��Z-���⩕�����뾦��&�t��O�q7��(69F��Fv�XGM35-�ÀF&,�����C��!��ŻnGZ�Hc%���jZ��-ti	D�F�;m��Nhz;���͌J���zEF�,�L.C�ع�����\�ڡ�{�5��i%>��6g��?٠4�l$�i8N�b�~����)h4����C>��y�!���:��N�`j���9Tk���G�� �8I����i���S}�K���~��Õ�l�����;gN�w?���3��b��Kp�7���;�f*��]��^�>ȕ����w�����i̼����@ґM����@-1���K.���}�;�})�g�@i�o���?�l7�C��ہ�O�A�w�ܳ�ݟ 59�)����=�(8U*c����J	m�Y���_�m؄{��� �������|\D��bj��M
܂J���'�<��v�B{vZx�kE�'W�SE�ѱ��A�ΤF�1�E�j��I(a�%�a���ڢ�a��I�������k��m(,_��o�9������������/��H;�{�|�����M�%� R��~�}��T�(�tF���$�m%��n��pl���#��r��l�701��8��0��kp���#"�{���{gƕ���^�����ʯ�	=�ƙݟ��'�`˖K0op�{��}
�cG�z豀�BRl`���dH�{=�BՉ�!�x��&�2���nK1�I�����w��>0�BG�$�_q�~��Xp��@��co��������n��o�	X�R���NMap�btvA�?�8N=�03�6�8Z��"�8G�EO�N#�s[u��q�mȜN��ͽ���"M�YI�a���ˮ�e�|�+�
�*�5~���+p4��8��C�R���/p�W��j � M�	��X4�i
$�[�US@��jf��M�������RH�Fa C�\���X�y�s���o���D���K��ޯ �6�=;�O�z>�sn�?��_��FyNϾ��x�Wh�8..i���	+�b"e'ЕȢ`���]$i�<,�&L>M��UD#K����!u�U@o�
	�7��9|��[���'����U,Y�
o��x�чE��r�d��G��C�^�ś.Efp �sx�_�����~�ش�&�\x�m���bn�3�z��Kpş�Ko�@^9�Ԫ�N��o{e�Í�݇5�7#=�W�^�1�^��K��{d	���c�W�u�g�x���pnl7ܱ�׬�n:�5TF�$0+������ v�ދ��!\~�u"���P+��hU�~e��4�^ cb/����=��T
�6m�5��\7����Ҋ����p�0�?����������o�`���D�y��qk
�4�k%P��_*�;M�Z,bK܎�s\}(���l
H��Ţ�g�*2U����^�Ǯ~_򌖵(h',j�@��|���r�*�.E�U6!��JwC*�B�P��Z��Ha��}I���(
�U󭬬�H=��C����_d��%�|�8��H� �����|	�F��Ns���������e���*�=� ��K-�*|=-���{�ؚ�hR[�`Q7":bur����x�K����)�@Qw�Iͦ���I�P�ND�U��?�{��r��s�i4�����V�~�_ikn���D��D�ړ��F.��y�1Mm�C3ԣ�惆�R�=?���$�iF�N-�(2�02��D�ZV4��E� ��6mG�+�bvd#�
�XZ�q��G_�X�3W8W!32�H�Dw�1���ŷ�b�O�7�j�|R-�t-�Y��5�oq|��._���BΆb�?���R�e�������&̦&�!).���}ѹ+���8��o
��0�N��*Nc鏬���<8G��u�MA�C�-���%��#d+��0O�ɵR�S'L<6���"J5:}p�u`��O�0��d�z���C�םM��~\�u��Eo6���$>x�5���V�+v܄���/��:��$��Ih������l��J�3����/���(�RY��hm�̠�|%�������@b�
��Y�ƙ_��?}Y=�Ko��ۯ-`��yӯ�v�0�cc(�m_���.E*ݐj����9�Uk���ѡ%Өx�U�,ƥ�]/!?8� H3�2������Zэ(�v#=o�� �����{O?������/b+a�Ǔߋ�2_�y��CLǈ}��솓��Փj�K�Q��!��[��ߎ���ѿ|	�Ъ�f���Sx��7p`�!\u����@����<��~��'N#M6�A�����U��˟� .n�:9�!Х���	A��!�I���YZ!0Ws1��_o"�q���Fa�ZL�=�~��~�W&6ڂn|�G���_�Yl?�m�:t��^����1������'0s� r����&u�%�r�-"b�t�PS	�.�Լ6�j�jK�Ǩ�PAz*+�T�&tc��a����p����%���)��=���_`��!4K-|�O���w�̟'|�\A�n���N��'ƅ7_G�R���⸡�B�r�r��{_@�����->���M��/jmU�-1�j��k;�ö���UwX�J���g�q���=�)�3cp���at�ڀ����Y�F� >}�Q{�e$'/ K��ޔ�%h{�JAz!�xBס1�E�b�"��s�=�.��4��<�$̞A�lڊ�4X����x��gQ:z��,z/߀M��	,X��}����Gpl�A����W��[6	g_}o��p�A?�'��'�)'��;+{~6P	��ژ.��Lq~�<\��`p��@� Z� n��|!�jؿ� N���+�`�Ux������H:�;�Ckף���AK�`�gO�~�3g����܎+w��IT>܃�~�8wd7`61r�&����0r�-l�1{�<��	���Μ�UW^�5���=zO��q�p������ہ%�e@�w����$N����m]��E��q�)l�U�����<�s�c���a��e0�3
|᡻~C��tu\y��L��.�<�F�b�����+g�ib�(U/o�Leqv�G�¹]�����c���s�� >����Vϲ�r��E��ƙ=�x���<a�P%IM���D�
�������F�w�	;K�8�3.��_\L��4�g+��rڔϲW+�Ť�R��dU��sVܼ:��ؑ+��O�{߿n�!~��z�
���yͿ�P��	�)�����)ῼ���/P��/�/>D_"$?Fx�����hH,�Y|sf��|�l
��Ցe��N���%�M����*�ҬPW�n�_/�z���bcЁ=�&
�p(J�1B�ҕ�A�;�!]�h�2�n�t��R����Ć�w�X��_YSE�VYh�˃v�<�A,k�^��iIN�)t'� 4��[���oS��%�'L'B�X�P��j��0
4���f�K�+5��".v�rO;��Y���a�8)툅:]��Ū"�S�q��"��ʞ ~�jÑ��vS�$��K�	���a=��R�+5�|�t᪳���hJ�o6�O7,�ڀ�(��\jו�v��'B!i��U	�L��"e�a*��i�i�u�4�$�р/���RW�Dyv�8?:��cS8Ǧ��"�x�� )�7X�����#%�b!"E)6�N.�v�l2�e�b��,��5���o��G����p�M7��w��K����pf��(}~�j�tB|ҍt5���]��K�5�G�ȯ��(z|�ۆ�[���0�`�U�1�c�l�
�P�B�Upa��8��]X��UW_��-�Ѫ_��=o���+�Gjb]4N�1�Ð�����Mq �Ф[��&�R���`���B4ǆM�m%Y�H_A������:t�{ѷvV^�v.�Wo<�8��ϠW�pB��١��"P5^�<��I�L2bKY9�b�&��v� �9��V�r3�R��5��g���m�Yq��%T�3Ѝ ���� �ċ��39Xa�֩�8�³�����E��05��&8�!HìB�q�l�����9t[��-Ϙ�,:Q�D�mc"��TF8���_`h�	��:�9����eFp��;0�v1����k�bf|�v�DϺ�{������S��@�G*
��.+�����
��L����MYP a
4 	Ѓ�l6M�ͶS���Y�Yi�;3�1���4+��h�c��Z�نd��٠w 	 A(x[�eV�{����@)�a"�ЊP+����ʼ����|��L�`�8�h��������Skc��F��§��&��*�F�ౄ�� �u�:���Wq��~�������=��^yM�����p���e��I�nh�^<�C���_�9r�&L^��P z��k�8P%,���4K-�Jy�4G�G�����U�⳿��c���A�XQ�    IDAT8�쏰t��/|�v}6�;���:d6�ĮǞ��w`��Q|�ӟ����(Gt��1F(�M�8%aO�^�5�MA
��5�^'�}0����C�!�e�}�i��w�=;��_}�|��F����q�=w�2��z�|�{8��!��o��������}��[o`��z�Ǳ�6dҥ�zț6�sE���f2�D7(�Q���uj�7�l#��/c_�:������"���w�-@������ĔL����?�?�1�rx�����T��Q%T�p�����_��<�[��m�?
B���:�w~�m,^�]�p�cc��4J؆����o������7m�[�0���Օ5(�&>x�|�?@o,�sO>����QZ���ɣ��6:�;]8V�,�=�f�N�G�~L���B����)g�R�����cs���`1�fE�ڛ6�>9�c����jlݷG�~fFxK5���zkT��Ѐj�ϝ^؏�_�f��"ss8-*��c5��j�=��iJ9�I�/�
�KI���)2,��J�N�jr?��)W�⵫=^[�t�O��\��Y6Ȅ/�#��O'�<�W�L�e?��/3D8�Uw��2���)1޿�h�ZE��J^g�n@�.(ꌐ$�CW��)S�[�ێb4�+M� �Rs%4���'�ԇ���J�&Vy+�1WU��k��k�1�P����?nH&�]�u&k1�i
ŉ�o:���׏4�Ѯ�KS�R����4Mr���K^�
x�L6D@����<�T�p��DF�G*�Ir �i�E��4�yK��=�<�������?M��Zmbg��~����zݱ8��q��(�9�]I�KNqZЦE���S�+�k�^��+Ƒ_��9��M� �,���]}��O��k���՘ިi��iʵ%]��E�F��2T�f�U�8�p�[+c,�<+E~b��4қ��*2��r�I��B�@H���F��\���5H�|��O"���t3�m��B���=J�Jey���"�eQ$���7�wD(�u��Hn�aI��A�h,-bfj
��L���,.O.�V��*���ɩ�3��%2�)H2���5�0����� �ux���ظvY3��������Ŀ�?�w�d���o�ċ����#(.-�/k�)f�zz^����-�Cut89����h}xβ�������Ï��ч�������s�G���.��<X�#� z8s���0��Kh����,�
5S|.:l^+9�YMC�2BLu�X�̵(`�L-�G.�F�����m`�r1`�:�
�h;yL�>n�F��ͯ#�(>~u?��yL~�!J~�܌}�ge�JC�R�� 1�2,����ƪy /�'�����h���V�O��?E������ �A��8�7�u�ny(��9I��^�������?�)���(6�(��gLY9
'J��X�S

u���a>A�=�ӂ��d�<�2Yq%bz,�7ظ��]#���Ǵ���nS��]?�=�>�c��t"�+#c��ő_������٨���=������{p�ݷQ�pef*Й" 2lPt�f%'�����4��)�y=?D��Cc��F��POٕr�B�?���Bd�|���N7���ԗ`o��N���O��������B�y]�:����j��|�e���aח�{����i�RnVP7r�y��^��O�t�"U�*J�I�M�Ǎ�\ƣ���}�	��.N�⏟Gpa3��m���b,��Q�9�;����)DK�x�{������&�7N)�:�Sg�Д(�@�z�k�+��ĵ�Y�L%#�) .���u����������\������-0�������k��O����=����?��a��ο�����N�c"Km������pč���f�a�[�|���v˾�ܪ����C��������^ƕ�p�{��Ɲ�o݂���9L���U����#��Ʈm�P]�	�*vmA��넶w��W����g�'��7����(¥�|���3����W���'p��mh-�NO��g�l�Is<r� 5Mmq���ￃ�����4vl؈M��#�n-��:��x#�#k��������L^A{qz.gp �� ��~0H%������=�(ڧ�`�����t�1��l��^B�Zņ�u�[��sgN �����m[1|��@����	���%�?@��1��.0bf��n��Wa�Bӑǈ��M(��:)(Z]M@ʵ_�^=�ٌ��������4�&���%t��I(
W���X��B<�&J�|u:!wv�YpriIb�j
Tj}�ԕ4R`���/��{ bf8��$�^�|�+�+MAbjA�k��w��(�i�P�����M��~�jt��	ic ��C�k �В�@��sM�V	���4�nĽBi��vs?ؼx]Ğ��d�ԛ�vҡ:����k��]X����TU��[tS��G�]�Fr|�����u�ݾ�'c�}�O�Q4q�ns��n�����֝�fc��Ip͖SʙK��O!��'�͵���N/)�Ӣ����Xgm��z>��[Vzki"h�%(|B�Q#|�8�հ@���i3���5��y���/�4�;��PE�g�+'��4���]��k�t���O�����a˧ g�B��ԁe�HU�Ej�L&'���[.[�f@|v���ԐD5+a�l�s�4(�����Q��"���q�Ҵ4�,`��"�m�z�bQ�.��5)�qE$�E�BR��D�����yU�X�z���0c�������;������/ȏ����o�����GGQ�^@�k#F+�g�1�d���O�'R|�cGq����яa�[T���5��Y�͟����y�)��h����P z���^�~��g��� ��CާPV�	��s"��,\��t�łK��57��r�\_	�>�4Vo؄3g/��Fܸ�b��u��"mX�
:�<��Pڽ�~��֍`��ћo����#�z���Bɉ��H��'�P��Ѕ��������<;cIa��t�F7@;WDߞ�q�|�]�Ѻxo=�C,��6��ˈ�n���������_'�p��E�;�N<���M���RT��2�6��s ���)��H��T�����a9CG_&��\A��T����X��%,!Ĳm����ѵع�>l�u��b�#>����a������8s�C�زw��1��Qt�&D�L�G����h ��*�"�vF)��N.+�h������ZW���'	��^�G^W�A�����b�֍��~����p�b�р�DQ�b�:f�ǅO>�@���ըn�,z�ŷ�A냣�ff�T��K�K�k�S(�&@6'���ޥ�Hi�Y�0�K�ڤ�whp	�d���}�k��'��5h�����_���.Fki��r���wބ�~���n����$������b��g6�>ĩd��7	�UFfj�{-��kZ9�(�D9g`�TA�]A&SAh1g;|�>���:9�\�81�2�
 {��������0��:���W����b�>|��G8��~��CZ�YY�F��"kȘlʕ�$�6{�v�nu���ߓ��8_�О�p��"'����<^|�gزe=�y�1���׮Q�a���˿�k\x� �ټ��;�#޹���w���#������F��o����{{
q����]|�gp�.�|����v?�$��v�;}���w�t���ly�v8#k�.�A1N� ?����'�`���=C+0x�M��Oa�7�)V��yc�^�����0w�\9sQ>��;�cí��j�V�N.�HN��g0s��]�Eexh1ࢍ��q覅�1��͞�_�j˗���_�g�%�P�`í7c�C���;���#s�<*t]��jIh2R0&�����:?�� �u�t��ï8��eH�{郒I��X�F1�CT���q-�E:ɀ������BQ���N7��I����RH(	�B�i"��؋0)�J$�*E=���U%-PL�dZ �z&�h!�n����B�c���n��xC��w)���V)�z��q��u>�����i���{V�W�ٵ����i��8�q?q��35Z����˔��e%�}Me��
����E�z�@�.�V�Lrm\��H�!�q��(9��1�w8��$[hm�லT�`��<�8DK1�jȤ��������q4���;��?}���me:�p��sU��hy��d��8pr���=���Ե������Em���Q��1~��\����)�KO$/2Zvug�A�-�L��{���PED7�'QX��X��l�ɤ@R`�&��L��F��Oe��Ђ5H������)w�_96��JU�H��t��r�	Q���rMH�S�9E����z6�G&��`��R�C[H�QAf<^�qJ�l�|k�`�7��Vc	���tq
g/N���y��7���a��-�*�$�CMz,H���V�"ѐV��4��ʥ��c�H?�nE����_~�'Ρ]�`�M����Ϳ��[��W���7����_B|��W�.��
ʻ���/=��{w z��o���~4��h�l�^�A_��;��|�`ۘr�� BW�`J�@� 9R�\��$�6>��W_E��QZ=�Xz1' rF�}.�(��Kθ��a���x���br����?�k���^4gp�8��X�p�@�g���n܄���X����z�o :|��}��>BD�=��+!�H�$I��4������uB�2�����h)�ND�J%#��,f�0�o�֯���и2�����+��v��Y��7�$.:��!�nf���s�|� ��PZ��@�g"?�m�
�2(]��-�l���zh�����9�AD�'���d*�A�2E��s�Ȱpʊ�c9��Gh��1<�u;oDGs�膨-4��P���<�\���b��Mx��ϢY_�?�)��Y�{.�F;�a��+kb��
}�J�rN&��cR�	K� �,4���e,t�h�>.���
P��X�u{>چ�V9���ߎ�}���G�P�������@m��N��ԉq)~Fq��02:ZW&_Z���a~����IH���@$�3�Ŵȥ�S)��L�C�i��y2�WM��ŵÀK�J7=�9���灭[�<̿q���p�ƒ�!S��X{�=��K�G��3����|��~U^�� A�B�����}��Z�_�#�kL��D�ɂ�k�aM1�ѾA�u������0J}�֭��p�pׁNӟá_����GP�a���x��~�����C���~�}t�ǘ�K"j���{,���l6B����h7<4=�0@�v�L�f�T(c��[p��{�W����3���g��4��������@n�F��P��8s	����p���*豔G`���&ܾ�>��SG��[��/��v�����>�8�F��*�����f&��O=�}_�"�ƀs�x���3�b��1����X��&����'\8yo��W�t�����j�nύx�_��;����v�A�����K�1��aL]8�vl��f��.FV�=!��m��<�_���o؉�w�FuU?����;�㯾,����nCa�v��@mf��q��X�p���ЪA�m@�����D�}�ҋ�ϝE��;O�x�59�pjӬ8�1�E+n8��SE��U�ЍE>���c��WAE''י�9��R?���G�;,��J��3q&�_O�t�de���5r�I>,f�I�9*,/�)V��I��꽉ui¯[i��0)~�I�^W %k�4���K�&@���*�4&��Y���EC.��	(O�9�HZi0�א�l��f%�Y�z�j�<�)�Q�$
�|�@��WҘM�	���y�h�9��4E�y�}��L^ A3&'u�k���{�I��Pp���85r=��8v��'�w�VǙ��\Kl
]���5,:�oz��?)���@���#�k������=�m+R<m���F���v�)����?}1��*��t�<q�> E0�u�&�iM�l�S�D�
�TW��n�A�u�����U��7^�ޮ"��R���$&��d"�N2���X+Q�_KK�f��7R���sCL>��ß�Z�H�?��leR!��Jg ��IC�f���r��Pb��c��̦��Rm
n\W%�
�5$�C�����.]����py�m�	#S@�X	
^�$@�3`QGJT��sSO���8Z50�͛F�{�z�L�\</BㅓW�vzشc7��G�>����Ν���o�v�$�܆Iu��ܚ��n]��=c@�	\:��/���]t��C�2IW��v,��`�Z����Pk�`��PZ�k�m���a�����O_���:����&�Q��0{�l�}�ي��&B�Äg��2\.5�8Wo�o�o����ǟ?�`q3�N�̻q��P;;�-�w�GB�Mc�6��:pe�7�g�*�%�G�,�4]�I��D�B�ĝB:�$3"Aa��HS�UMA�{�`���oX�ѧ�@�ۤZl�������{�=sYM߲������u
뇑��+Qt� ��z��II�&����o�b�>���E��/���z.��^M�h�=��/S��#�6���jp
Ed�̝��X�c�}C�E�A�efOt]X�� ��v����n��[n�����8�X|dl��T:n��XcqAD�4P�9��
"n�0�b��Ag�Zlb�u1ըc��D�ׂNq���k��G�єP�F#�q#�x�i���.aq�L��"4&���0o~�r%��je�j���"�1�xg#��a3�D+�g���t��x�G2%�(�b�"��P,$�(�J'�t�.6g�MtB_�@��ۇ�|w���������_��c�Y_Fi�&lz�q�|3���h��:>��3��C���+v������0���#Nɚ���M�J�${rZ���SM�U��T�ִ`Y�l��0x�]��j<��������k�����F� �oނ[}Ccסު���C8��/�>���1@�,ϱ.�f�"P����E���-_����I�܉��=�
��;>��?�+�|/~���6�v�6���ob��t���Qk���X��A�݀�5aes�\�jU��su|��G026�lX�a㮋�s�05�	�ӗ17N9�=܏��h>�g��ۘ8�1��zh/�x�iX[ocd2ڵ%�\�wa	��W_F}y������]���y���@�����j5x����j�֌�<"�\�:\:r?��_b��1�}�AnY,60��8��g�_)c�#�p�yހ��<,ږp�%��)����~:���+���9���!��ȦNT���ڂ�dSe1(��h�
{LD�
bO�~�ǿЈV��)�=A��iY(J��f���4��X� -?S~�&�d���bk��O܊x$׾�~*��W�s�(Χ����K�J���p��1E�DD�(����A�/J��c
/-K��0j&U��/��-�	�ҕ�����SE���T]���_�:W�&�a��_���N
RJuZ�I'LR�����XI�����M1_��L'��Ñ�"�N
j�MTfC�����jB+�G*���D%l~��w�_�mx�i_̉oKM�x���!��EԳʷ���M}�O��B�Ngqm�u�m�m~-��<-��Z�eY�� H3���j�tmq.ɸIÐ�,FyPS$]]W'iWy-j��<�0��Z1qZ]���C"}�t�>���"+ϙv�)�/�H$�.iK�.XH�E'�z�W�J�$A;q�����@͈e"ȥ+L��U�'�7���.C�(=��u���ȗ�@�b=�|N	\���QXd�j;&2�%��r1�b�%�ad!�af��j��ᓅT�\B�~O���:&'�qer�3�XZv�u�)![�ig��Z�M*f��CBs�ϋ$�%$K��X7���܂����w�p�$>>p˗f�w#�\��?�Y<��/ap}�M��$z3�/OG�l�Eg�ٝ0w	�7_�ٟ���9��ڈ�fHNa�f���.�0k�`X���oö�n��wނ�F&����%�&.��;o�;~���+��    IDATI�K-ܘ1_$�-�^�	KS�xW.��,�|Ka��X�E��3��=� ��}6ݶ���d�ټ<�#������رcn��6E�����)��`��Dӓ0;]��4�<�Ȃ�#ꛎZ7��&�_�ɽ#cT�Q/:4N�� �P�?f�i�k�~ &@ٿ?� �|�I���pf����z� ���7l�ح�1t�V o�E`��Ç���#���С�q�,$REU
at#v�'��Ž鹘�40�P\,Q#c��k(���L��[e^�.h[ȗ��وi.�Z8>��� �"-2Gנ�z���]���F1�qF�� �Sx���3�x�m�����DӸq�9�.M1y�Q��dɦ����B����<�Z�tc	�e��'E��}�dL�!l�;w�o|�w���x���̙cX��^���Bw�7�bC��a��A)�E�QOD}�O1�^�IE���$KM�(fs� �#�Is"�pb���D�H�c�0��uQ���:��}7v<� ��
?��[���;095'Y7���[6�|y�>���=�!0=����jȗ2h�K":N�����Ce-({�2K���-y>�鷾?����
���؏��0�o��c+�m�ˢ���('�ӓ��8����͎M���J	�f�Kp�gϡq�#�<2�b��Ye'd�d࣋.z54�.zm�#��%��$�qR0�u���琹c��i�����f/��S����|�y���$et�VQ�@{Y9y��H�H�>q��d��T"$���޵��8w��?���Mٲӯ��g��Ѹ|a�bd�:<��/c������9U���.-��@�0Å�b�%����,2�{�_�(�g�"t%s�;�X�]�y�����5�øa��m�|�o���/���r��{���U��*U���l`XQqH�ᇠ�0�����_ 31�|����	HC=���IVGj��K���j��ғ
_ө�\r��5iV�����2I��$��!����IFo�tӭ���(0䴋�vE�����V��T�����jvD�`�	�B��$��kP�|��Ɋ��8�f��5ͤ��������I9dJ�2CL�D0A����+�apq^qPJ������SMUb)*0�����L�$m�����S��h�=�g*���a�9�|���|�0�e�_$�Y�$�w��Ns\h�.�;U˦�0��H5<6�(�ǰ9��/��*��SL2i��J��I��!���w�m�� ��P�g�����ch
�V�-Կ�j-���io��(��]��:pI����Q$�"�+K\sX
�#�9ꠦE|:�IrrX٩]����,� ���;E���s����[
紸gq�ғ��;J��[�4��l���[aźi������D����1	�&J��Z4�2q?�I֋y��)guFZL�oh�u]Y���.>�b=�4��=Q�h�H4C�?c>��Zj��ktiE���6������� �>�s�{-�3��r!/��<
��H����Z}��54�m�2�ZPr�}��.��j�:��X\n���a�"XD&W���)�aW�C�Ї����rC��ؘI�~��Cøi��:��L_>��3g�-6wcdsU�۶��s7n�w'��o�&#�ū�Ґ�	̟���C�z�u��?��s!J-�x�����Z1[@+SF�8�VΖ��~[n���#@�u�.}�!�ϜD<5��b��:�ZY�<w6 ��䒌)2K���c��0��a�aڸ�8��\-#^=�Mw���!�|#��
��K��-���pܝ��쉣X:�����yd�ẛ���Q�h*�Q,���� �N��}���I�$|��Ƕ�����tO��
M,YYx�6`����r�h��`����`��i	��"�iM8\���у�:��983��5X>7�c�Y�H������0�,2N�cKSU�:�h�1�YF��Q��;��9<�1@w-�se�7`��L��|?�F�p0gf0�s�6]��M#�����f��/ɵ�+�ј���?{K�/���pz�r����ǉ�2I0�VȦ(;6
�rYǁ�gG�LA��8Ģ����"��5�����<=Rg��CC�-��?�C�W�z?�֟c���昍�`P��$�ɦ�ƪre'F���aeDWBms7Zq�9N)6��Z&T^#�1���>b��3��e�4�r$2h��g� �(Z\�	o�k�l���P�tхI̞���|�w`�c���n�zN9�o�}zV�.���Ѿ�̼�iD)}H��d��R���'͕�M��j#}(8UDN	�B��Px�!`'m�������RL3���*�6)���t��r��0��;�\.�f���Bѭ�t7�ЈZ���dJy�����FF����<��U�pｨn�$�}��)|��X��+�Ea�v�s?6�����i���P�HԮ�u;��0��4���0f��Y�����%�rSW.��я066���6�܁��ҏ"i�lY쪃�=����1��`�h��m
�V7Ʉa>L��,��s��pV�������B/T�6|]L����~�����K8��[8���+�qþ=ظy#�V��B��8���m���N�L���E�ٌ4�%Z2��	��]�f-����#��[XB^�6�T����F^gHW���s|�-g���J+��+���'���k�ϒk��>��i5i�r/�L��ѻaf��r�W�jN)�6�1P;�'�U�;J�%@b�*��F7)#���b��Ӟ�6���hJE��BTsyh>��1�i ���_�2�&׵��R�s�B��^q�!]�b~N���PT��)���s�ص&����*�J=8mR�W�rJ#�w�
^	I@XE/�H?�j���~s��K��2z~��rc�F�+j���H�|)�������AL�H�FjLN�(�ⴛ�U�KK1��<�#X_��I6��,�N}�L�@�]=¹�)i
��'c?�ǿ�����p�_�uy������EQ0dFδ,y��; u��\^�Rh�^}D�T�:/h36u�1�����/��\��cǱ�C��z�gUE<�K5�4�@�u?ִ ֢P#�-е؋c�܊��P�?�j���O���8b���A��3z��u�4DU�ߌ,����ql���xV�eZAi!�|�q��z�zhFǽ(
u�,0M3� �L34|?�l;r�P�Y�(>��8 �s1^(���8���3���Jŋ���/��z�;R�'�=�~Q�ܭ'O�s�ռ�O>�A�!�I@u&3���f��vǃ�R���NPd�����C��qCx>�<���3/���Q�����s	$�C��\H�
dZ�,I7�U��9Ћ3XZ�AcaqÅ�C<�W���q�m7c�M�Q]���h�T�w{�Q��f�?B{����q]˂Mj��&z���l,�94K��mߍ��oB��Mȍ���/,DO����a��8�SS(�G�sQ�7�o�P��<���y��Q.6+>І���tr�4���\�a��1�n�t��xh7?�(�ʗ�7���#n~Q���c�`��0��~��Z(u�ť�H�FOG&���ΰ⋜���.Z�j"HKF��C�E�o�#����9���.Ԧ87pЊԌ"s%h[����F���8�7 mr�rq�О����`��8�W0�X@�����2�4TS��)��h͆C�ͱ%[��Hh@�,�>ڑ�0���V@�R�bG�������FǠ�nF�v��j�oߊ�PY�<�y��4Z�ϡ=9���.L�Dki�. Ӌ`t\��P�D'#�'j�R�Ҝ�3kR���A�.��8j�HC8��1߬cni�+�!�cc92�����<���K����1����A:.�ɺ�\��
.��bDX�_B�`KQ@����Ƕэ",,7��h��i�#ׂX �e*bryO�xl�[��
TLG"j*��9��ߖ�;��
�*��נd���l���4PwC�t�U�V��mY�:�f�~�/`������U6�
L`VEQ�Pk���.�Ȅy!�{LGG�5łL
��2�LK��p�zL�sXI��6�.��l
��C�w�'���4�f��"�2��S�;�UG�A�@�"�����A=Xƒ�� ��(6�86h�n�Gje��L_?<��^���^GШñ)�w0�n-��Cadv��L��b�,��zm^�#S<�6ݖ+���Q�ٜW,7j��궚��jsh/70?��U�C.WP�2��C�j"���[1¢%���n��k�Ip!�ȋ4]���[�&:�s��jK3B�p���JEX�x����!��\�,�U��W��3g0�,��yTr��n�J���~q�))�E���d��ToH�S� ��>�\�#�=W&_F/�\x�3pjK�[]�	�8-�G��a�\���?��J��ತĕ/�{�J� ���� %6ڹ�$�S`��ą2�B��C��%4KA0�������O$� A�Ű#�=�_�(J���~8e�$��zL������B�h��C�ta�.�z,l1i)�b�]�ϐ5��m��ajqK�M)�M�@�筯�����q�z�� �:J�jx�D�S����yJ����W�#�n���ڕ*@k��E6��"�O�/���'�P@f��W��u�ֆ�%С��$�:�d�睔���%,	M�>�Z���X�Lњ��Iu|<����ą���|�ǲe��r��/!�w�cP�k�������
���[y��5+- ���3%��w{ސ��y��J��[�	��^��i��5����"���A�Fzl��n�pׂ86"����ec�`zZ�G���qlF�Eay˒�Y��(���M�b���H�!-C������+m,TJ;�b3�1.E1�g��c°y���n��^�H?���d����C�����}�y�?���+��9��ː�����4\x�!��.��H��Z-y�<��/
*��<�PЍL�K�t��mKmU��Þ�B�پt4Q�̀mb5�v����ӂ���瀕C5[��f�p?���(�*��j�RAP�)DU._� �wQ�X�w<��� ;�$������^����(�-۰���w��jZ<����rz��C��%���^G�M�{�$rK���n��M�"Z#~�U �.,�]��Up�,fs8�\�	js�����q��B~�u�!���?}������_Biy	���4��"t�߶����SR�{�p	�"��BGT�.@�4�IR�A@υ��J��:#�8��_�8��`lތ��߇�݋��ʡ�fȀ�^����8��̾�������j�� ���ْ�5�IZn�4 �і0���W�%u�.5�E�Ӂ�C9S^�L::
�<��~x�>l��p�^�N>L�%�����&/bq�C�^���\GmiZ29H3�S���?4cX�贒�������$y0C����B��>�ͼ�����ք��쑢��R�)�_����^��]���w�/}	k֭�w�,N��?�+O��9�b��U�T3�s&F�JYVƑsh8��s�����Z]lk{�D#���'HX�bG�]DI2�`4z��2|^�-d�H�3�l��C�9(��$��B�|#���;��e�������[0w�8>zq?�gN�vۈt���n�)M1Y�����&dO�^eB�&oX[.a�XA�, ���0�ߎ5O<�������p/^F\[��e
�[�������y��nە"*�u�6J���`��"�� ��ż��r�B;��,�:���L9��i��X(�u�/��d=t8���=d-��/K�OK1�\��L�ò� �s���ӟ3�d�l�&�Bs�m���Z�]�O�h��,���n�V[M�頍�������d�� �F��p�m�N�z6�Ș������2|4� M_�.�vC�WH�[]��(�o�r]薬])wQ�2�D�������ڵ����̜(D6��FW�u	�,C09O��7���!�0M_ѕ	x	�A�Ŋ+)��gT^RR�^�ht+��Z��>�*�PMS��Yf2pM���<�ܺȬZ-_F���>i2&��"�]�B�(�+���W]h�!z�/@]��O������2��=\�:BM��$�1.����y�SS0�-�b"�ie��)�)�j�&pe~m�XЭ[���jkQ1mۋqD����Z�F4	):q!�~�:7]M9V�hi& bj���*J"
`�:�H�"�8Y��&<R �mEq�N�)b�EM���o�w.�z�eH�U ��҇�+f����wM��C����q*F��B�ES����S��i�A��qh���-M��5��O`!oc஻~���/�q�'S
ȫ-��+�᫚z9oj�L5�O�O�?q������_���cG�ahQ.c��kR n���xCp�5L��C@��E��C�2%�͚�-�Y6�鴐PT�tT�Ffs�
TN�Ҧ��})l�@�4��4�:0h�u�-7��ҳ��Y�����`�-�T(��#:7��������t3��>��U4��+/�{~6<�c���(ݽ����`� �=x�y�����B�*�KJ�|�K�~�C���F��c	A��ӵB�B�6��E9.��*h�ʘ��v5��F1p���{`��w���pI��� F֭�c�|�
.�} ��s�����N]A%kʦ��3���
���h���B���E/�ϑ<UrY�P��dl��(��)i�m7FK�0�&a�Zl��v\�=�i'�WV���1e�Y8u
�_}�^z	�s��r��'����f��p�:J����Ih:\Q-AP#�D��a����J�]h_��>�Ձ��#Ȥ�/J���� ���]'/������ǎ`f�&>G0߄�P�(X�$:ә����6��z��WI�)�9��Li��Ѯt(SA�E���j�h���=�R����9�7ZX�|,{�L��[��׾��O>������|��ӷѺ0���U�RZ,)Ȯ�`ö��Tl,���=��_ ]��8I/gF�!3�h���t�F�����JeºĔI�t�~�G�9������ۍ��HXF�N��z� G&�2�2� ���}���/`ݝw ��`��Wp�W�t���;�I����.�TT�dT����y���0����)1\�����`�ZF�s+�?�8��̎�»�=���އY[�C��p	F�O=6M��9�/�1��a4��y����uР���DC�uѦr�K YL�%�9i�Lٌ-:�̣���4��j�k��.ێ�Em��k�zNs����{.5K,-q��
�9A�mK5E'+�C�^H}�,���ȉ8R�y�QYD�Zϣ �8� ����p�,��N��]�A8�v� ���v1�^��l�������H�%�x���pr@8X`�!��|�$j�0e3"+JM�fH/%цŭK���(��74M�����7�}u|��D����М*�ݦ@����j٬(,)�_}�(��h����T��R�ꆁZ�{���v��ۀb��'�BW뺈x&M��5�����&�Bo%(�bVk�Y���X�h1{%	�F-ߓmF*q1�5��<���3�u�(�P�'�@��o64z]�����9�@�Z���q1\,`��*�s}��Gd�����K�D�}SM��B�w��q���U�a�q���Uw�$�
��W����Ln� t{o�y�@uH�̤t��@���M����VE�6�Ƒ�)C\���3J���*V�j���q����bN8d��z�p�����i��]	����D8]��b>���?���_���7��U�?=�?�xh��y��c_�����Q Dw���h���J"�v&�:�%M�ܠ�Z4e��t�1�cÂ���)ʥ�=%iT�Vb��q��!�]���n�&�8n��hOf��^G�a�.�'8�迮9&tǐM�z�E�eb)tQ�c�}�q�N���Ǉp���=qL��򺃮_�;���|��	�q#BZ�1f�b� �w    IDAT��n6L8VQ	�X�O�0����a��_���$�ZKhQ/�����u�)�9Z(���CӴ�Ȕ�^��~�k(�u�nX)V�e��}����������z�v�}ذk��(�� >5�W��_���a�������g!H�hr'S1<�����^(��$�]�F�V� ���f�x�fl���Xj{h��v݀=�?���6Q�������=}�U��Z�2�r��s8��K8��0sr�*�,���� �Ŗ�&��V����2Y�gt�'���kfs�m�0�j�����P���z=F�R���"�Tp�o}��##@��6���Gc��e4'fq��QL�_@{b}^�*��D�"O�'&;8I<�O��l�	G��As�Az�CV�ї+#�Ɨ�"D�Z��L��fC��T������l7<�y<��߆NQ��4f������ȳ/�i�`����S���n�c_y��
��ѷ1���hg�_���q���Т��q7���`������%ˀE��%�H�(�6���#E���V7��C�Q��DR��;ײXݷ�L�rv�����B�F�p����Cel����^|����i���:5� ���([g,$"�Ԏ��B�<�}H�H6�u�A����!\*��ڴcO?	g����&^���IS����X���>C�D�Q����T(��D\,c���a������h�>B�I2=�Y%,�tC(~Î��d����u��B!z=���B����teI������˖��$�� �r�	�j!�D|����]Wi����|�<���X�����Ď���/Yz����!yЊީ8�>�J�%�i��A&cK�D�kcr~��ڎ��E�Fޯײ����LV��B��N�C�	iy���b-Ɇ�{�ձa���M�nK!f۠f��f��7�gS ΅����>ӥ����K:�㎸�\�0�x���Jy�P���)N:��|���N}K$ζ�F��;P~�`� K;��7�1�s��,����T{=��� \J�щ��*,����Г�F0�@)DŎ�4 ��@�E<���/a��1��M�&,�2W�G^�!�L4�.��b�Y��cQA���FCrb6��I��Y��^ �ƪIR"]^_�h%�S!1����NCl9�KA�7�ĕR5mJ������)SLN{��`��F���n���V#d~����~a]�ں*��|��P"VJ�%­�����K(��&I�l�	�H�B�]y�m��8�y>�r8{�x�����F���-�9�X,dп�g�?��j
��+�z¿w�w��s����X(���<��1�#Z~��#����T(����gQ�t�����I��pS�S����q:&�Qk���f&�Y��C�A�qo��`�� �%5��ϣ35��C�r��l��P���΂�F�ማ"�:�j�*%�t�����=@>N����Bn1����F�d����o �a�j�%qC��g�.�v�,s�a��~��?A������Џ���D�CY6rC��#Y�.,n�@�]��N�v	��Q�����ہ������c�x�}��ҫ�_��ǚm�q��w���at�u�&���>��/к2�"�Zd��4]�6�$6b"�ƞ4(b��  G��}�@��,�q`I����c��ރ���Ml�w?�jE�k���'����'�B��i�N�{/ʃUUULN���G^~�r%�F�Bϕם�l��J���l��4��m��Y(�NVl�A�����NOt-=�]�<d�I����z���{��*(�� �<(�i��E���,5q��9,���s�E{r���@ΆA����e*T��	EnܜX�]���qM(-E��P�	�y�-G
Č薌�C�ļ�b|v�zMx}���ob�7��4������~���%����Aup��AL,-a���M?���~�� >��wq�o����"��(�ɘ5s�X��Y,�[��[��݈a����׆�m�f@D����!�l�9�'�z<�ֻY	��a��{04�V���f�>d��dMD���9�F�v�Ξơ~g�<
~>�:�݄3MjS�Ӌ���%�K��?B�P�^�N ��r)V0X�CX*b��E{�jl}�sp�oƕ��a�w����I��mR��-�NH2r��k�0�WE��I�â^�t���{�k��ܡ�(
�wn�+�7��I�h6��h�NS��y����ʐnE'$����!�x'C{��$h*+f>���5ehc�^�\�ĂF��|/q�L��C�)ǫ��)p�ɂ$���TF�.)�\��֮�#���-MG7���4�h��lձ�k�m��A�!��4Ť�U3��f�s'Ī�Sdg&���+Rn;)%e��%�&
-#~��c��K@'3��b%�&� �)��B^U�f@�]T�/�A����
>z���,���:lȬl��I�)KIj/U����Yp�������ٷ�z=`fjYi�)�U���W���O�Z�H�x$�j�Ԛy��rR��Lw ��BeNu�$լ@���N��	L��h>����~�v�4�P�d\׼(F�mc����v]^�L`�Ҽ�V�����F�������<���o};"&� A��$�$Q��e�G�̮��;^�m���ښݚ�ڝ�����^I�,���(�b�(f�@"t��7�{���~�4Z�ݪ���J�%�PH�{o���{��}B<P���A351��Cj/���	��vW�?�+*��5�����s�5侥�F��� �zƅ����¸�Z��a�����d��.��@���/��2���Z������^��8�gݓ&$�4��*�ON���Li��� �8��3�~�%L�9��:���i�[_������?���|To�v^��]{��;��?*8�z�Pzn4=�/�JI�2�z$��M'eϵ"�$Mk>��T��Z�l�����(.�j 8����G��a��R����*�&g�9qa�#���U�q��W�~�����R����b!��g�ZD��:��/���{ǿ�u�o�s�� KQ��kP��V\��/ �C��e����Yi�+�R�î�)ƀ]H����W~��'G��n�|X�#"��r�y)ɹe�МH�M�n�c0[��ո����5���L6�`��a�-L:���N�!��+Xw��h�Ÿ�M�.���W���O�}�(�D�c�D+��ח��B��8�?K���,.Qp.�vD�
����QcH��I`�X}�U��O���]ס����{����_ｅn�)@Tw �o<�o�
�n��6�<��?���=�y�-1��4�<nr7��,�&�r*s����m>u,y1�:�dK0=��	7ta���/�^C��Q�A~l��8���~
�6��)�V h.��_�̻�q�w����o΢J7��昪I3��V��`)N雤TN�fy�344Lu''B�e��%:7l�H����]4�e\����?�Y�9�������;~�a���c�a��K1���_�� �U��Qݼ>�(^�_�-�ɓ�#��Z�"*Z8����K�.������\���"&�Eu�ו�@��tF��L��N*U�	�PC?�Q_��
�/َ��@����t̩T Dy>Y����d�?�o��a�x�qT���!5��A�഑Բ4��Y���u�ş],Jui�WYy�*WѨ�Dl8�(��z)��v'0��o�#=�C���|ȳSdZ� ��*�Q-�P��sTmG���TZ�u��Xp�X��1Nd<!Y��6i=�7�aQ���%���8��\+♯+?uz���	�R[��QJk�%��R+�>���R9��JͰ��`Q,���
�1�gV�K��Ʃ钗��:���t{
1e�ޗn/D|M��p_Z�v��^Dw����)����)���f��/�aQ�,A��R��@S��i���E�]�Ϛ���F�_G
�)�OE#���m�-T�E��21�kt�p>���,�U�,y*HJ}�i�ގ�r/%]+@�s���Vz��{O�i���ґ�n>ly�Y�R��-YL�b��Q����[�E�=���h���Hڬ��&w�#Xj��lp@J�ŉ���ʆ\��.�j@�ט�@u�ٺ�A��Xx�Y��{�����@Q��Ҩ�ƣ4th��4�:�*i:�
E4��"%�X�ȢU�u&��'M`���](01�i��`�$P?ٿgk>K6^�,�+�CA����kT��)��V8W� �Ԁk��X�辸&X;�6Cz��JH��>�܅��&q��!�2�L�j�Kh5�jZ���%�>f�$�4�D��EH��G��k�`,�c��a�3���i�D������{˄ƿ�%�G���k���{����e�J��eAD'@a��2JV�*����f\���.]|��x+�eݽl�򴤂'�|tJ�u�&�U�E!ra��b�F8w����7��ܢhh۸��Kq����W�`�VcW²,v���{2�;A"{|��D���~ޛo�8�IS��j�݈���`�>l�P�?���۲Q���*�,5�ZR�bh�Y���9N=�#��2�3-A)�6�*��a`�$�]夀ɉKF�qL5�q��ŝ�!)khzͱ�;.�3b�� *��(�V("x�����k?�1f���t�NN�8�H�;�H�%Hp�ҍd��r��aS����$k��y9n�761�Nc)�1q�U���6^�Ϝ���0wt��Y8DǺ}����Y-��~5v}l'�;���������|�Tx�r��M��yy�Q�H�hIj��� Zj���`�ہ��X�#�w\,tzh��5�Ub6��Bђ�X��22�\Ce�:��w�h#$��^ʴ|D)�ʫx�����}�jk0H��=��2I�ONϤKQƴ)X��s<���LԝJV��C��P+/n]�ea>q:`��a���-�ݏ�c��ғOb����?�D8�q������]s�A��?�'���[6���G�/�����~�5�*+8(T!E(�.��[D�ˌ,�{�owЏcI?V�Dx8�q�0Z9�ZBF��H��F�i��R���Cq�u�Z��E�X��$r�
�w� 
5�����?�>N���(u�#�� ��p:I[�P��rs�J��Ȳ
TS�h�N�`�61Q��^�Kasl7܌��7Ch�;�G��8��/Ł�k�$&�����W�j��\$Ye��B�zp,:��`���B�����ҍ��v��f��)��J��z�,�#-N�/Dp3��I��LRZ�22e�i��8kyV��Y����[�B�rl��!����T��=��K����J����-����W<]�L�'u���|���nK 6��>(V�K��B�ih�*.�Q5sB5!r*H>����DJ�9��S�峈璑 `�$�reS��i��2E�����"�,��*��I�T-�j�V���if��č��^�ާ-����NL�:��*T�P/U�C��e�aG\	1Zy��Fo��n6_�.!�8e1�5jڒ��-�tE�!ҿ��S�]�i�.����p������@��Ϡta���ב����sp��'M�	Хdy�;c�D�>]y}ו�YGԙ��㡰�Ѩ!�GGN�S!pzOٝf�q�Kiq=(�5�*�q6=�H��"���)8�b��/	Х�Q�v�f���6�;nDT����I���XN�&I��JB��g:��������2zt�@@�ׇ*�FoFA3Qb!p����1����������HFDs�b>砼k��/����[aI�QY��}���O�����c���[����CG�3y�俥������4}^��WL
�H=�B;-����&�(�p��d+TL'�D�<u3��%�LfZjB_���c�L�bL�߄��c��7�*F��B9(��Ǡ�!hR�c��y`����|��^Be�3���ˈ�݌�O}ÿ�I`�jeQ�^P4ڊ�݇��@nHv'�S|��~�#�~�1������C�J�?�z<�9���PO`1W��b7��?���;�~%��t�����^lzm��SЁ����c���Gp��`�y�,�D�vԥy���57��F����!JC��ܿ0N97FAjx�� kM7�Lhbb��x�_�.��f����o�;?c�Z��;�>�WM�b�;@���x��_���ހ��IcF�\&P�1!�[\����Uh�ɂڶ�v@ʁ�"�:�8yDv�(�lk	��6��C��'Y�⦀�Z,�Vo(�t�T��"7>{|�s�ä���l��ߋ��	����!�ɹ��q����kL�T��5N���kE��z(�@�\`�D)�Ʈ��S�b�d�ˡi�,��n��;� �^>x�m�������^F���ݟ�n���`���J���<�<��]������^4L�k%T�`Q4���S�i���@��ᆉ���c����p匨�iK\�T,�9�RH��5�`���b�%��M,������\��Á�? ���\	Ս®��9�}O?���=}�8�A[R_'����Et.n�2	ZFU��<[Y(,�'l�2j�Q�r̎�;�Bq���j,���{�x�O���bn�h��������h  �زfD��Q��<��Y��)��$�&�C�E"XJ�\/`��>X��g�+���Z��̳���S�Yѳ�dr�u��,؋��D�Y��"�e�40��L��󉦧U�[��9`�ǆ��39�)
��/��`����E�Gb���A��9E�yB-���Z�2yz��H9�r����2!�	�>�e���L"H��闥�섓΃&T�8q�K�+Ӯm�H(YJ�ʾ��*>âO��8��I�M2���"y�<oH[<�na��c@��m�B?�8�D����C)&�,ļ�=����oC�[TS�dR�Y��2�,uhŬ(�D���h4�I'l(�WZ�-"HuL�L�4�f��`"�!����� f����0����)��9��T�!�/��~��˲�x&��_�!]
}'���++����Z�ˎI)�xe��J�}eS �kz�� �O�����W6�j�s���Q�uP_�'�%y
YS �3x��)`Ð�'31�L�Vح�p"�l� $�B���(��)�>u�GOIS0���X����;�O�JҴ��k����?�ߕ��2�Rq�r�M��}���+��'�~������tc�\n���KMI��5��\����I=Yw�	���r�Y�@G�YT� c:&%�����<L߃�y(E:��wv����c�ĄCg�\	�5�P��|�#u�?i41'ڜxpm�ku��6`�5�����j�p���!�|�)��a1�Q���X���`�OI����~�N�`��0<k(6֠cձ@{B��nXL���S��{��Ca�	��4F�^�j&��!��Mt�"�k�8Q����X{�բP���zg�D,�1|���,�rEB��f�����K��`?��0��H�P�R��ʦ@�]J#�{*ӃTS �5�7�THžh1���հn��p��1ν�r ϑ��-�o2Ey$�H����Є8q�^xo<�4Z�O@���$�$��7�+1I/�]�'BN�EF���]@��c��A�(�hc.�\FH�v�ż��|�+n0�z��Z�	���ȳ@�*a�K0����0�@�p�.��q��~,�� ���=�|�ه�Ѿ ������K����Q|,MG�̲�e&��b#�!�<�ȇ.W��LYZk�`��!��r����7���G��������S��0ZG��
�2��	�����3�C{Q���#O޻�#u���B�,�@V���6�,�bW*M}�"LG"q%J�"���%
�*ҋ��(���k���"��MTke�[�Z�$ןֆ>;���%wݏ�s6n�o���'~�����-������t���VW(7�܀��Rǥˌ��� (�>djbIZ���W(�Lm�o��믇�~#`$w"�u����}�]�U�e-\>�|�@��W    IDATs�~�<v?�4�qp�d�E�Z�O[gl^�OX��B�*�Q��"G���5�>�̂a�p@���A�4DR�g�m�*�E���n���X�픊æ@r�����$�3� 4;�Ż_25MH������)�\�	�K]��)BSQE,�ӏ�� NY�����;� &@ٿ�%_nY8�"ɪJiB�~H�"j��4s����G��˯���[�ŒY��	O�E��.�����)�-��"\foI�N��U�F�y��L�h���(�D`��{]���TJT�H�}��am��a+������P��[o�\��.!���Ę��R&+M�
u%ƞ��+`"���:��f��	nUS@m�jT��K�6b�f@
K����{D��~c1�%��4�Y�����Y�3���0�{�8((�r�s	Ζ5��u���T�M�JE��VÜX���Wu�C�A���M�����B��͂���u�?v0��QB�6cl$M��}�)འ�_|J���u�BG�%e�zNFx�I��kyR����+e6���8��G���/0�)󬠕o��"No�x�w.��sZ�����z��p����������/�LOݨiڪ��	�Xd��>����1y����lT&�f�S�B1R�Ѵ1���D��	� S�H]БT^ǁ"~��+�c�Cn�C��(�@-2P��X`�_�៻nI���X�c��K����E�_t���~ݵ��K?yK��:���1�3g�s$ܱ1�}���x�AA��|쇘~�9�s�`�Ui(�U��1,XUt+ul��.\x�@o�/^��o��(�}XU�L
X��J�T�X2<�M��J����?���"D�~�e��{��F>�#��~�%��ޓ/���{��f�L�3==P��D�Y��E ��IA��l���2�
�R�D�:�0ѭ��n�՟�rL,�/���xZ�ts����p�G�C��ҥ�Á����Ж�0���2���>\RRH�1���L�R��$�aCǈU�j��i�\WDi�9$�����MbL/�����8p%�F����1���8v����I1p�M�N���1�\@��F�ߑC�H�x�KQF툺n��V���W8� V�,�8H�(m�&�T��4V����ǜ�	�`l�v4��ȕ����$���� m]�h�� ��a�!` �x�y�y�+h|�� �CI\�y�t�B�J�T8�� `��~X�o�7��x�#Φ ��O
{����㚍�.���h�@~�
Ӊ�m-�4�h?ŷf���uXu���z�=�ؼY�P�={0��39���,�KM���J�k���m�H��/Ѹ�f��i{�Ӓ�M�mb�TE�<�X�T����]��VX�mR|>v�nOU<�ٽ���b�ݖjj%*��������}��$rQ��#8�X	,�P�H�\�p��!+���+�Lu
6z��A_��mt�=)$�,�诅�J֔�;�m�r1t��9��L�d�ǥ�'t�&L�t�ؘAuRt.OR�e�îrj�Qr$5�{� ��C1+���y����ƀ��|�H"����<O5b2QS@�P��������^b;�h��[���z�D��_�AY���n�b�HX����s5Յb�e�Lс�?IU�F��	M���&�wi�@mH�i���'.�4vm����F��ƹ�֔\�cg,V+8���0~�=JS���g��C�ʮR�W�(�3��ل@�8���4\4F�P�i�\��=P(���>C�V _z���h��(�!Z�wc�'0س[��1���_Y��r���zHc��9�i�=�V�|�x�$��k�_��KŸ+MJ�r'k
��H���`2�N��[�ֳPϴ�l
\#Ƽ�]�o�#7����@�H�H�R��t̻�F-�hiDϢ�P6�l
�ִ���Ƌ��>+���S�/4*҇�+A�!D'��ȏ��[ob8袞�I�~��ts	s9�|c������5���J�����hR�_t�~{����.~����͞���^.�s�jEF\����y+7����D�T��r�/��䫫�YX.��)h��,]	�L��o�|���`���0;� �5�Xڨ�:Ƒ�� ��A_;��-�0m%�>��	��"r�"�����ጌb��mX�i�.8q3_{��z
��)A�b"�ã��N��̧�r?��7��gЧNI!%�����b��M����X{�E@����װ�[�A|�j�,fayR�lA3-ѵ�n�BtP�<N���]����Q:o�cGq��'1��3p���.�lG�t�ʓ�-�st��%��'H����E�HĆ�o,g�=EV���Ј%���W�(|O��HA+�D�b��]źnƦ{�&j���F��w��O�^o ���Ы�P*�k�����m����P(¯Nt� sKL�m	�J0F�J�D)ʲ.lL�yTa�`�� 90lS���[phX�=��H~J#��`�Q`�琖�׻T��)�D�ێ�#̷�$K�B;O��\͚"Z�t����s��b�怇~�t	"���1`���*�0R�"o���HJ��'�6jm�y7�NwPcI�&.��Z���c�>y=��Ės�~��7��/������~��CzD�Ve�\[L�(9)Llr��0��F����TSe)V��2�8G�,�ㅘ���Qf�F\��l���g�������h����+�c��m��BT/8��U����|�W_�3;������,�}r�=)\Y�q���'+�ƽ<�Q�4i�R!��F
5Fj��6`_�k�ظA&���I��gI6
9������U���cRT1Y�:�\iN=�2���7?�<X��L7g���1�̔�-��r}r�KbZ�m������,p]��)-�$P�np���Z�
`�8W-�Zo�)�<=�5(�b�*�X�Ҵbқ5BcJE�2i�LpU�xܳ9I����D���R�KF� uOb�5�
%�[y8)��yb���؉����e������I �_�=,z>I"́L	dsMvRa+�J��Wj����1�(����#y�c58}&??M��Nt��<T�:��@�"L;�6'X�7�*��ہ�������rpθ,8��O`՝�lE��"��M���m
�Ե�r峂�T>N���R�3���Ϯ�ؔ�� �eeZd��i
�q��6O��`F� e����K�Nj%�^j����ʳ�pMi,�*Kay$aw�߂b!���Y:\���*�dL����,G�53i��YvVwH���X�[�Z�9���������-� ��	���_�Z-g�!I�lN�?C:5���ɞ7��q:%qѪ�QS7Cr<(ؗ����A6�؂~r
~�#tw�+MA-���`���9�@e�5m��_*_~��oJ��QS�r'�?���?���������^C�X�J���1 {��a
iV�s�4ѐ�%E��"R6*��yl�C�b�0��IU�u������>ra�B���y�7�DC-1��)#�B��"F.�����d�(V��/K�N�������[9h<؎ǉ/?���/�0;���W���07߈͟�4p��}�Y�>��.Sm�2�У�Z�Ďm���{a]��=�������?�F?���n~�ds��U���s��%hY����\���C~�*i\N<��<�8
�`���D�̂�(gb@޺���[;�"0�J5�OԌ�^% gaC-C�%cfrdy�c��!�st*�k�N��WTzճɋt,%&��#Xs�͘��F`�zﾀS�>���_��\D�2"I�Z�������CKF�|��=t�lBuS����9t}_����^0uqp����i}�ʡ�Y�K�&�踡F�!�\� D;��&��,���9I'*���Z�I�����Ke�q0�i�F��h3���f��<�՟�Њ��<:���y���r@Q����W��C�0QB�.�X.A/�1c��c:��_���[�!I+�џ��~{vF��Ct�:k�|<�Ʊ_�����D���$V�8���0P1lvG��H��d�H�i�eaG�ԥ�K��/N'��t�(Xk�U��p+ο�:�w�6����Ͽ�{��G�P���\����m[�z��$�����1��kH�ڃa�58Qj/b�=���Q�b��g��ۑf��b6�T�k$��x0Q�H����3����54㢋��S k���x�٧p�7E;�j�
�p����3�br�⮳�p�]w�:�_|/|�at���r��vH/)a�J��	�*
�! � ����b��ƙvSPn��sCd ��#�ȥ�V�<fߩ-(��B��\s�_Ӧ@8�,�XĥS,���:ÉK�r�Yħ(,�^�(d�����ԋtB���6H	ޅ��H�B�!-���]�/bT3e�E	L#by�=R�.'��*
�_���B(C&f�}L��hy>|�L0 ���D2?��S�!���QUם�h8p����������#ݒ�j
��UQ����?p��|6�|=]�BL��U.���G����2��xz��9���9l��~��~'p��H�Cl'�0�\r(�P��rc�:�e(yV�fT!6+)8�:m�	��IQ���KS`�!�Q����IS��݃�׆�L*�1�d2������IՔ�{�Xe�p݆��Wq1��P�1�謝h$�-�ϖ�r���4k
�f�l��!�f��+hͼ�l�q��׍c�]wc�f����K|�'��%,=1iO���E�UR�'Q<s)�|l��|9�9����ls�ϯ�ԕM�0��3���`��}��=T�H�WqbnS���o��e�y�_��#���~^~��K����:y���\��ݔ�K5Z�8��S�,���ٔҦ ۼ�Xp�<��[�BHD^��wş9���8�\q q���5Cð�c4���w�g��TkX{�U8��������,*�sV]$p�*dHg�(���)t����a�8�s59�	���O� �y��y̿��?�*������;��a��p��W��;��>p�C�y��8��HOb���R��j&?�X�c�d����9�*�a�؊���`o\�:�W��[�A~~�J�+fI8�4
w�)٢tJD���xN9�d����M����/#r+<yZ���@1�l�L	/�4�j��ꦛ1~�-������9?�(���@?3��D���s@J'E�ⲋ�k��i�gZ*
����t)������e�+b�
B����ω��YV�ʨ����Ѯ���Dd�F`�BZr=�w��(3��y�3��w�Z/�JT�c:��<r\�sl�c���l�����A��k�����+��I��'����Fy��[���3Ut#fk��XS��82YrMSa���t��R�UF&�b~b�T��&[/�[.݌�Xy������?�������#N
�YX�z��eSG%��̒SD>�W���Z�O3pfz
Ӌ"|夀�$��|���l��8�`P��_�'�v�'e����E<��qb��-�oí�߅�K�W� �c����:�_y��G���p�&��(D�G��\ϕ����C/
'�:\��\��>��1b��W��(��7�hV�o�������_�2���
�G�V��_�<F��c8����믣�bj�Z������o��g��w��{��xm��F�<ƇG�)�3�G�:	=�	|Hm���<斈�*�?����H�	�I��i�rzaPs~��v�-����0u�L�z�e�WtN>g��gÞX�ۤۥ��C��.�{>�~0��;�U�~ �	�wi%L�-j��u�K-ʤLD0��R��q
��Ҙ>Cs%�)�?�	Ӥ6&Rz�F+1�ia�G����2��)�u�?��y	���FWt#L[�CI!�}�A�Ra�v0lrߪ�#ͤJ���c1K��(p�i���`�������XB,~����US&�9��yh�ںwdc7݄���\���"H,I�Vf�s+'8��g�+�$r/���Z+,�	6��X�3�"mC@�6̈́�f��GE���=�~�'����զ&ME��L�O��P1����_Qg�J�P"��ˬ����
eI�DYrtR-[��Ȧ �����we#�l�׵ �~>�sVa�wb�O�7-I��M�J��F��P���V�<C5�[f� �������i�*NU��x�N��?<ϸOr!A���}�bډ3�|�9t����ߒ��ZB
�O,�a���];���S����5���>�Q���o����G~��C>t��b[�Ҍ�G�V�J!]���u����:����򐐇<��	��z-a��x�%h)7��[�u`�4�R�F�8!c%|��*[�Rx5�5k��9�|TV����.Gex����G�[�C�4���F�����?ġ<��i��j@���>�\��{P��&�4�3}L:��G��gU��F׎ax�j`�ۇ��~��_��w"?�F�o����2���YS ԟ(D�0p��C����k`���!��|g�y��6_y�˘��W���dS�)�r4�$�G /�Պ�%����)�%!n�+�`r"��P)���F�B+6�����b�����!~��8�ď�{��s�%9\syr��e`�7��U���Dq@i3hB/�� >�cL��h�Z��~���G���'�g'�7��Q3,�9U��"��ѩ�>���~c����#r�P�g&փte��b�1&GZ'�TDlYX�CL/-a���Bg������Y0��{�Q��eW�5� �օ�f��X;4��#L�������'Ob����5��g���*l��R\|��Y��l����%�g��}�UG'����v�j�SAkQ:¤�gZ
�Hѳ�2��.Űa��41=3���ytIH"�H��ω��âf`b�|���+�_�I������~��������[$�`��i��̡1�
��	�{����~c�XE(�������r�&�K��ľ�^*�X�^�	q�r�i$�FX]�c�8�~b�Yh ���~���N��.���1���8�V������.4����⣏a���bf�Y���?�'ش}����y���F=��L<��LꨕʲG�Q����4C�����n�X
\VFW�$A��t����*uXG0SQHφ�Sq"M�Kx�T.3�|r2&֚��P�NO�x���<�ٞ-��i�!���:M8NB_�}�Bz����*��ی�=I;�:������Ȥ����?��fam��a�AѶ�cF�c��%�!��(�fs�l���z=��ƩV��K�Kq�I��av~��N�G� 8fA�etU�e�I��O�m�pzj5�+�e�9l&M���q�>_҇Z�Z��)�/����T�M@��%!PҾ��@װ��X,0q�MXw�]�e;�bM(,!����(��%�E�G���æ@�r�L�Y����q�GM^2D�{�ω-\/A����h���I�?�*�)�Z�p:C��qYE��N�*3Ynl��/ ����Q���)��q\iJ�����P��k���,0��Uj�_/�r��
�`_����]���n����ι0**<.��3�T�r<<idbƳ+Q��T����'I�І��D�x�ʕ�9�}_B�ci
8)Ț���w0�P�Ci
�Z M���]����3��cW����Я�$�蝎�{u�c�>�Ї��trr�vWƿ������a��G��eݾ<��[B�#>@i�7S�I�Q��A���Y�y1JP!��0Q������4TY��r�9��`���5��Qܸ7|�>l��"��&�x�q�:�W���o�������q��g᜙A��D@I�Fuۥ����W^��*��1�j׌�<���_��^@��a�[(vi�ƂPĔ-+7�z���,�?<I�%"�s�\|v���s� {�ǩg������u�)��8    IDAT�5�g�J�$J���)p��O���gz �nVu�ɢ�9�gme��D	eppX�PfL͖���
W]���� p�*�x	���	��?�3݂Z0I�2hY�+C"����f���a�[���䐫Ԡ�r�&�~,�`�Ϣؕ ���/*{8��P7I00l8b�A:�P�i(�cꪦ�yX�8v�O<p�BZy�UMC�ȣl�$K�"dA֘�]�!��E:�:h{�������B=y���i�x�b��f�*�9��^�)�6��4��6"ڑ��w;�����''��c�9�b��J��|�6l�jP/��ӹ���i`�zG�w�������i�p�{�@}�đv�����::-V1��1f{J���&&��u(�$��|cScQ�����O<�+�������f���?���Q޺����Å�
�'��퟿�S���K���������A��W�:�0�DV������5��i��fCƂK�"���pz�a�u%��(������!���ЋM��J��^��l
֭w��_�:f�*�ɕ�n�j\p�v��r��O?�S|�]L�:����?Ķn�̇��ҷ����~�R�������|'��u�N80�<C=����"�[K"�'e����axD)�)`�C��<&�@k0��%E������`��a�W�}�,�\��,���.ub1Ƽ�/�-s���G��}��|� 	�D-�$[ ]g
y��b��4l�c�ƀ�BvI�#h���.�vO2:��+�P/�P)0�<�"s���S>o9��V^����ñ�i�?�f��B�T������4��I��J�C�(�m��HC/��X�t2�`�>�fc��q���|eRhu8R�`A�#8Z���F춱�8���T��Oc8S���!5�=�>:|��b`ڴиv'�}�v8�w"a��SA�	��,XE�%�_��C(��u�J��V���{��� ֤4Fg�^�U:��"j�a�.:{?��O�Exh?Ɛ�H3����<j�R�׬R�&<-�3��W�%�E�B3͹H��u�hX�Գ��
4RZD��K'�������I�]IOR�0����	�yݱ*Fv^�������,#��r�Q*�gm�Y��������j
F���s��1��f��[�f ��Z�6�J���MA�`���c�q챧��`7F��4"4fS����Fm��o^�����莻�S*Տ4�)w��s���g�}��:���NN����"n�D�L��fb���M��>�Do)Ҕ�/fT"xb�I�2��W�gt~`�c�t��]����f���(%g�b���CC:4�eXpqmm�BP,#�ȕ��n���hN�«��{^~[֟����[��3��k����o��l#�g��[��%joF岭�|;0T�v�f���Ak�E��~�������`�-�Љ�s8�
-2�D�wn��fO3��gi�6Z��գ�p�N��%�������j�����%�Tf�R,��tfw�\]���LW#2t��CqC=j1X�9J8,>��X1kGB"�3C]_���	}r�+Uh�oĆ���A��7p���Q=>��BW,��X(;Tr�wpw���&I��r<�x3ЋB�b�I�F'�ѢC���Z��R@F�SF�a"� 
Kk��F�aPe0��%pj@/o]G'	0������$�(���3����3yxM�&�5�7�`�K�,[�w:�̵�r�P�@d���Lgq_����*��Y�n���v<XE�ih��x�*7�w�����ȣU�B۸��qԇ�PEmxis�@������ۃ����g� �y`���^@���j1zI������S�V���8��,L���`0��6Ź�LGδ���"dR���~�5�z����OX�85�����L�9��7^���� �m?��{�>�0N>��n�w�wdzr�ￍ�O<���T;��,B��nXC�ו�\Z��B}���f#}6�l�v�`m����0�a����\�q��[��{��z�8�ȓXg8X;:�5��A�����۽G~��0��������J��O�*&�zc^_2 Ƈ��sʒ���"R�.���p����.���\�X�f�F�{.��佋:
�r弍�늈��UA�Iz.C�H�{!,�(�_1/�%����Hk�-���ꆖ��BP�2E������C�O�bC)i'�Eē�maydWl��3��ԃC�/$���ߏ�7đ+4�t[�*7b9)�1�B�^G��K.N6�v��	'}v=�8�0�#S�X
�je o˔�A�z���Wǔ����aj��s��`�0�qq��A���4n�0:=$�K�D�4��GF��YPh>���1��W��]��O˴�(b�q��-�2I�'�,L�/J4x�����_�r;��C��]��� t�`Ѝ� ��� u� ���� k�k\�� �XQVb���F��ԅ���l��e��RMm�^��M緞v^zчP�~��a:�q�y�x�A{fSeiR^}�{�,�;�r!���pM��8�-��lRB+T5}e�%s�t��r�ſ��%M�p�Ns�7��h�:�E�^�����"2h�\�fZ2����2IM�Y�lE�44��&̆`�σ�������^��fY�Tn5�a�,kp�}��M����I���3���D�CɊ>�����F�L�w����}�������������_\�������;O�����3h�rP�	Pq��Ȇ�+D)K�\D`�6
"�I��O)Aϓ06�a���F��#��h�9�t�0B�룪EX��1�(��8#'��n��hx.�v��Х�#��\��?�W�xo=�<6���{n��囁ǰ����n��(	4���ˡ�ihU
HV� �ˎ���#�G(�8u��)�M��0:��jb�^,#Z��`��1spBB]�j��6��6��pK9�kƠ���i��E�,_���!�i��T�}�)��2/X�<�$�,>�O�`N+�^(��PYD$�i
�TM��p�q�Oq x�%�8&±!ԯ���Ø?u����\B�t�P��9a��P�8�&��M�!=�+A́�P��b����MtCĘl
fz-���,"�Y�	W�|V1m;%LXeK����i�B�b_л�z�.�!b
��\0Xl��aC��2�����]F�RM��s�1�Y@����������\�b��|�ȽΚᥲ��M�[XU�c�4$�q�+�\	������c 36��1Ӵ �-�i��F�w7���9��R%��)�C�F!�G;����KQ��!�` ?��`�M�K�t0��`�V�L�TE�1������\7N
�>D$�H5T�A+6����q�g?\t1���O�o�{v��q\s���Ǌ���x��+,N/�����g�,�J{��-����IS�ub6���XD�URp����u����L��y&��x�!u��Je�k�Ph\��i��j�ζm��x��?�;��{���.W04�@T+	M�v�GN��䠏��7|��am�9�W��e����hkG�Q�VK�A�ani ���j.HI
��JY�(�n��'�|��z>������Q14�H�I0H�3�L6����+H�%��p�E����s�w{҈�0i4B1"��	�NG�N�%���6t�;UjU
9Ž�<�T�y��2�Ԩ�j	k+�I`��0�j��v�h9��a�pP4���>��/4a�sFCm`hx�rN>'ሱ�Eǫ�����a)[a��RDn�.I�������ul�E�*9h���(��t&�1�w1�'X5̅�R��8��S�;}C�<&��e�kU�j5����0gf�=�B{	q{q슑��7%���X�oR7,)d�J�Ԣ.b,.���W�t����Z��tN��gR��Lj%KaI����&�����r�L�2ʐL�S�*��Q�@=�+S��h�����C��W�|x ϕ�� ��f���H�N�Tj㚕Ԧ	h��ˌ�Բ9�"P������]�԰!�]
��2X���/2��M2M�Y�:ѵ��+@w����ad�5�Wo@X�él�,u'M9D��O�Z��t�~�� �~_Z6~xn���h�\���	1*���~���}�:��R�������z�爏�x(Z!\�hE]�l.JS0�s�7.�����G���J�_�`S��+/�����'OO���XZ�J@j�RT�gT��>tiS�%(f��?�[%�P�:IW	#i
8f+rC&���c����Q�fY��	"Q�{�k!F�i��	
7M�Y��ZCk�0&�oÕ�8rt4��Y=��v��}o���_�c�<���2T6��������7���]����xD&L��L~�BP������Z@�V�͇M�d�����I��o.�pP!�-%�����.d� ?W@�4ұ��y-	��E:4�ci�l�(�{����`�D:��g����&��P�I�`m�֢�Q���*D��!ʢM�R҄�,+�����D��e����v�C^FԤ:�9(�ϥ{R�Lt�Il��<�"��`�
0��#�������l���>�0)����hS7���*Eô\��Q����_>�s�ϑ_�q���R�c�;{q���U�����RE��X�=%
~�y��X,�c��(�Y��9�Q�����S*9؆p��E���L#vQ�����[6�\��/A�;��ՆX���.&����_�����`��&�=�f�(�*Dj�Mf��T�D�G
V$��n���|$f�e&Q5�)�0f�a9h��X����)M)\̈.�&\�Ǚ�I�t������E���z}����l��roZD=�}�<����c���/��;���������`�uq��8*�%D��q`Q��v��&��b���[~?��M�F�?��)b4_A�X���0o9Xn`�����c�P�^|�y��w�:1��cݚ�ȍ�`�8r���>�����>�	\��Qڰ8u���~�!l0u�+e��ȟwJ�]����|��t��~�#6M�Yp�kȕ*cG�ž�{0�up��u�41!S���i,>�|k6B�Ɲ�B����ۂ�s�C�1����\A�����8���9�l[��瞋���p��?�7�xǎC1_���(F&�Q��1<:��a36�*zr->*.[��a�^�JR��(�އ��wQ��@�-�Įi�S���;Q�d;P"f��@�w�%aR��yF�#p��&�Ь��K����k��p͈�`�	'����f1��Y=:
Ь�������q#n�+A��f�/���W�{W�3�~���fa�%"a�΄å>��vx{7ܗ_F����>��� v*HO�XD�4L��?�im�>f�U�q
�\ox��8�BI�u>O�_���SG2A�l��)`��)ID��Ww�tZ"D}�abjB�0�(�!-$ФCspg�������>�����S(��B܇Ҁ�_��_�k��8�,�S��G�$LiP�K��m��55P VF��N�@���JAp&>Vl倘�1I8Z�w�����4|4&�M�a�!���?��	1����86��p
��+��*M=���IF:l��Fs~Ǐ���ؙ�T��Ѩ�X�H �ShH~��1:Z��u�8�>�$��b��dG�t�x�SKMi
*;w~�O|�_����G��_kU���7����7<�ܓ{��[���137�^�c1"IJJ��%�U�"5�NU�+����V	HU$;QEA��x��*n��bHrrI�B�L�P��zJ\��30L#�3v`U�m������Q\�F�}}�S�<��̙Y�C#E�jt_G~��"��F}�4Ւ�s���,�h�Z�a��t��b8�KH��<�'��e�)�s���8��f ә*4Hɍ��IGظB#'��$g�vbD^G�A\R�:9�D�-���$�
",)BC<ɦ���y[�A2 &�Wj,����pAt�G���\�J3��#�a����`R��������>��/��Ϲ�vn��I�4Y$	+$P���\�rպvk6�N�n����o�^۫8�%Y�,$�D�:���=���/�>��;��?���454�ts������}��	��X�r]¶X��r�ֲ2B.�#����#�@�#�^�ZyV��L��h5*�e;B]��Z�X��}t�P%���S
^9F'*O��0��ˎ�Y����D$��_�q�:���w�·gPZ�� ��e�'��Z�,�������)��8�ZEk��E�`��b5�Gw�a%�Xt���О���i���BU6tҍ߇�sj7�x��@cZ�k�3K�`����gh��2���Q�h�Zk�n��:�4���?~�n��h� �Ʈ�4Xm�P�0HȢP���b�v�n�*b����[�e#�^&��*�A腆��a�~�Ÿ�÷a��&&D��ņ�T?�'�!y�T&'��G���B��1���_��o�fS^��d��TS��4����	:��h:V�MyΙx��Ia���??g�>��Eɴ�r����߁����^tia�^zU�B�4Q�{�ˉ^����V�e`��bv��Xx�q���@��˘�X̹��nG����^vP�j�e8�����+���b�C�6���<3Y���m_z�3�e�A]&��&������n ��T��u����u;h�m2�%�����ߊ�Zt7��)"�ئ���.� W�w�������I�5:삫<K�0|��X~�1xk�FJx�+����-.= ��.d�_�Ќ89��q�*�5	/�C�l��J�i��[)̥8�3�5�#�-6�!�rY�~+O=���#��-��]�|��ց�:�!W&-\(mF�:ne�..�6�	�'�A��G���O1����H�Q��Kx�9��M�����N�4��pQ�s܋.D����$P��Bk���LL Q�s�$P!���1RT��0@D7��P�-|%@P����+�0�Ia�DA��F����0����)>��c�Q�P4T~���$M�5Ȥ>?�qB��1T7��+򩇀5� S��غ���~,,y�7����"6����ଥ�8A>�$�gl���(쏛��R��d��{�劫� ��.�r=X^�S����`$�mHS�QX�S1��m!���Ml6���w�z�6e�ғ���
��ԇnz2��M,dG1&4��8t��H����,@�����%�v붅ҕ�q��w�oo7�������g�s����G�vss�o|M� �8�[;�h#hw>ʔ&a�$8FM�,ߏ��݆(����dQ��������~�}�#�T���>��h8.
��Rl��l����C�A�7�P�+�V��ژ�=���&w��RZc�`��~����(�ç�vC��JA�h8R�BW���b���=S��i��M_m~~G/�eB��j����\�DV+B2%J3��o�V�2��B��(�T�yƁx۳��grϘ�����>���s���P9?)�85K EFN�S�r$H-��L�m*���`3Hk�ؤ1�}�=����A���ŸP��F�Ό�ǩ�j|h���~#�f8�$���l��s�	��>K�F����������P�M�M,�']������,�dSCr84D0$���
�O�_8�A_��O}�@��Q�
�;%����ȼP�������2�zm�I"B�0��%�%�Κ��&l>C�ʂO=��@��Qw�p�0%��A�����?��{r��)��S�ϛk�WV��Y����taݣ'0<���F1�b��gN�tQ��d�樇@�я�2M�Y�J����4z�,E����HF"�f�"�)���X�F�޲�_�\�.̳�/X��k-���������.��
|�7?c~O=�'��-��{	~�S�����Z�E�XV2Ȓ�    IDATd)�u9Ͻ`��h y]�\��@}L.�d�0E�[�5\}���TC�k/v�zt6~��!l��JQ�b�#:ZG@�(�:2ׄ59!�+�x�k_��_�.C�	l�2�������������T*2\v�����'6l�v�>@ ��p?�=L7������m��g�o�8w���{�9 &@ٿ�⚋����Q��,sQQ̓�(�#,6�O䂍4q~��e�<����E�S���q�y+O=oe%R�HO*��o���\�N�6��:���ͧZS�O#��0�����@g@�_Q^d�Z:�xK�%���t��"��5i����ɏq�gQ��~ŀY+a��W���2�6	�K(`8�D�N�C%W��Y��%��n�s�O�����`���7�&������9.q�QM�a��`�Hњ��=3��ŗ��w��J�)�[�
O4Q�Da�MPGqjZO�z$4,#��� �(Uj�����@��f[s�A��.�� �g��~�(ʃ�P��! p��=C�߹�_ %_P6)�USp64���3�ޒz�&2y��jrH�$Ն���?	�ub� ���:R�e�e<���ۙ�;��K��j�5b:{ӈ���ب�����z��\�����H�)��U�cy*���.�| ��JКv�k�6�m�64&jB��8���n��j�ӈ�h;B	��=$�O��!x�	/+�12'����V��_���_�_�n|[h�_�.�o��~�������>��x�|��"���eY��"���nHRA���R.	l�Qs ��
u���8�F29�8�h7i�m	�Q 3Q�3�#6���R:B% j��Jb�"\?w'v]w �w�O���#���/^��Ch�ֱ������7�t������ 6V�z��8����.�ctl�0���ۚ*�eNѮ. 9v��rX�X�ێ�\J�
�Ug���#��G��WHKn3���2%�(�_qF�zS@46�VTq��!�se�l����(�RP� AD�@D��L�0���F�<�<U�|9Vƺ�Z���,b�@ЭDL���cԟDJ(p��H�q)-0�P�{�>�+HYh�]v�)P\��6��"C�XLH ��~E�"���� 6]l�:�R�j�Z!Rh)S5�q�Px��beǃO*��	U��[F�:$�r"�9����C��i�*tL�>f�LT�z�p9q,�ѝgacC�Cz�)L��ni;J���񔴝a_�(R�DZ'�Tw
h8%Iwb��XG�%��.�`�oEq�N8����M`˞sU �� �`��q��>���/`z��$��"�&�67���e��nɄC���bM>K�)J#V�-,t���"q1�<'S�gƖ�#��d1ܩ)\|�ո��kP�s���3�8���x���q��r.f�m��?q�L����8���(t�@��C��B�|�r��¦+��\�]�n��m�t;�N'%!Uv�t3��)4��b�4�b�ދ�����\�I6GpAWN�ht���"��P��H�t�8|�x�o��=�ML��z�;���[�L��H�.����=�H:63���7&���yr�c��Z8����^��Ϣ���ǉ�gß���@���Z�%�\{�H�l�Y�M��Z��]@}�����` ~�h�0X>�^k	aB�&��#u�[D�)���HC��6�1ZX��K�`�WP�( �S=���]�8g�r���yw�2݅o���c�5<�"����wM-Kt�ڈ���93� 	� =���5T�"�*Ҁ�ӡ��.-���<�~����Ջ8o{��&1�}
�s�5�l��H֌�?D�v0U��t\lF�d��Zo=�|x�m@'^8��?©{��v�t�"h�Rxq*'p���Ꜽ�)�#a�C��#�24�_�W\%��2	�*�Z�azfF
�A4�_(�� �g�3A�^�'kH(��fs�VSh-�N����,��-E2�!�'�;�a�BW�;�
��=��)�=�w���� Wq!���/��d�l����sG!��e�"m)�#��đ'� ����i~����[����@��֒$<�v~sB�E;���{3�C�O2�2Y�F��<�F��w݁+o���<N��!�M%I�dq4*(���Ʉ7ӕ����5]��.a}e�w��Ν�U6M�bmcC�i��OM!�
���PFdJ�(	��M,>�(����Z؁����Cs�\���,A�+�v�?��v��#K�*E���C�*W��9VWW�w�����g>�ǃ~��.��X�X�@�,�[��Es�ⳝ;�)�Y�r)̻|U4��@�*]�n���$������!���u�4E5�(�wP�CT���2'��P��b���8�����q�$���pm�� �\�������:5�l8D���3�x	K/��z��$�z!,w�hpR�d"���b�g�b;�OL�`娈��)C~��yS�ƫ9�"��<]T�b�l��`ᮒ[e*m��2s� �VD�o6d�_��j��7ݥFU	]�2R�$�,�J�hd�$=���W4	bS ('L���*FG�8�S�H�w!rn�DαI1QA]��;�̱���rD��M:?��L:�0Y����v��	��-����Fh�BC�8@@>�\�VJ���6Q��<_¹���"Ŋ`	�Ĝ
�8��(Fs0D;L��ɛJ#��ed��<i
8����.I�L�*�y66��4�b���H�[�l���D���t�uI���c�+���`z�9,�M��d$6]�<\��چ����;w���P ��T���2���3�?���Ӣ�S�^3��m����`H\��`$�rLRvj�yE�ܢ���G]�nb����� �@<���(�^"��.Ԟ�"�94vl���=�v��^Fwa��&�nOi[J�:��G���݅�&�7��IbXQ�6Q,xB�Mf�H �\R�FX�IB�A�1}(������ЂF��M��=b�������X=��!��<�l;��VH��!���3h��عg��9_���g������1�9���P��]��07/T���>���e���î�1�VKqзn�D�7��� ������
6����{��]���#�Y+��e�9�=��'Ĝ�(�뀁M�bҡ�۰��P�w!4�""�̩���?�^y�!�>��t�lEA>���[Ė�m��2}�E��D���puC�К^D�*�=���t��	�k62:t%�uNe���������LOa�K���P��
.֏���=��t?�d��iP,"s�tP�J��N`��,��&�4"� ��|�%9�%W� .�a�����6�E��t����d����ѭ0�z�1)����&z�m��x�G>��=�#x}	���o|;�6�(���=T�XQe��󷲠�PX�%��>�h!���}��v���3a�p���|%nvK>t[QGiz�@5EEd�*M/�/����,6�D�0�E��	M�q���R���u1֩�2�$�4��!=v1'G��:� �j�Θ�@�)i/2����m��`�Cۜ�ʽF��|�\ &I$��Y�M��q-��ײ3�U(�A�77�P`$iS����ip�c��5=��б��84�`�7pͧ��9�\��XF/�r0LW���Ij�)�NϢP(	����v�������/a}}�e�K.A�>���U,-�����9�� �&jSS�uqc���z4�zp���6֞x�W^@5�d1��@���� E��k�q�G?�?n����_R	��~ٷ���)���>�����o������_��vt�(��"9_O�d4�����>�
 ��}�[�!���d���ا�M����;��|���.�L!�?�!*I�*'ڣ� �n��^V\�� F0��~�T��W�؞,R,0���fv�#ŢWZ���i E���KҨZ��Z�w\����rC;����Hz��'�D����W|K�����G�\��T���$:�[�h
�.�D4���V�oR����t�F#�v���q]U�1r]h7j�#�7Sl�6�`���X6�I66\�6�G/?&q�;�FH�N�;��y�,�r�H�u��|-L%(��a��Tf���~*��.�P���)�Q��~�������y^�Q�-(�oy(�>�2���v�Z�5��&:��a�nB��� U	�Y�+i����J~����)�Ymu�)`�:��ΓB����&���Ǯ���+)��]�(�vUS`��B�h��쵰N&K�I�Zg�ר�;w�45���,&��-[�OMa <�3�x�	T�Q�x��n��Q�Q�a��	�6��9�I��7U���E��y%���ia����Ω�!�	����V�,�Y����&��y�VV��� Q�Z�<G���~���0E�2��T�a+"��KX�5Qq<TEӑ{�M`�he�n}	#��"Ռb4,�5TmC����#9�x��ƾ�����/����eT&���́�?�����=��+K���kq�mw�49<�7�s7��B�66�0{�Ͱ�;0�k0���ŷ���-�DqԅM�	�m�ad
e�Eŷ�(�"��k��MtW�����j���v�+ٲ�e�"�����-��O�:R�(��00-�w�u����b끫�M̨������w�8^���x��{�r�5���o���Bb��5��fJ>�jET��t76d�ܽ�qZ[_ob���VDc�4+�ѕ�5:�#
�#��M���Ͱ=7����^\}�]��<�A%�r?���q��~��e� �ǟ 4\HR	*l0żTF�>!԰�:��^:����Fxe�~�,�m=O���&�]�v�9��s\�dr/bz�k��y�ށ�~��1s5��<�T��~�W��%��T�<���j�I��� �:�r��ahh��v4�5Q�����=7�ݲ�]��(�%��#��B��b��A��M\��&�_B��E�\O��67�15�@�L��!��C���f�l�����ϛ=5`F�� k��Y]B��3���Jؗk�P{e�%y���!��)5A��������lf�07��H�,�"(k;���d���LD��6K%��'����'�9�E����D���UT+�4��b��kz��ګXs-��۟ƖK.Ɛ44�,_t�`�^$����w�^�P�t�(F����N;"�m۷b���H���`yy��HY�JSmcv�إ�X�r��)>�#��.��.ʛ=4�|�.������M	\;��*���5W���?L�|�¯Je�vS�r%~	�����}�׿�������U��2��}_��m�yS ^ɹo���0�/�a&q\|��\sQ�h��%��&zL�$��C��SGݲ1����V1�0���Q���C�ť]�E1�Q
;����2� w��J�-�f�b7�����ؼ�>;�HU2(����}l9��jƗK8�yC��\���O��"��C��y�Bؔ .� CW�\LE
��6�<Ii,d� :���k+G�LJ�ޡր��J��?s!���j��˩ ]�r��H'b�����*�Z>a�-�8l�5�X[�I�ϜE�Rds�3�OOW%5�!U��e��D@��|��f��-q,��� K��jI �0��>�E&]6$��P�u�a��^�A1��:�D�+ʘL������@P7�a3ٳ�.�T���R	n.�3��X�lc��u4+KүB����EВ ��+a��4cp"H`߄�b�-Kp)�mZ�6װΉH�kI�E�@�@p��:�SӨ6&0=9��k�s�6Bcs��H��(�)�:�0�m����C9GS�2eP��X"}��F�N$0+A����\C���4�"��&U��"��'j�9R�1���3;C�G�H5o�Nm��������xD��<{.�Z��A�B)��V�/��zՂ��m�m!�~.����{�;y������/f���έx��?�����0��{��� ��&����G����س8�������C���z���k���:��;������?Cp�L�	��*n#j^"iJ��dQ�d���#^�V�k+B�(�f$�wie�^�J�D�QE���$)V��n�i̲D����}�߂k��&.�z��$�$�OC���>�'���x�q�A��$������f��*��\�ΙIL\l��`yuE���y� u[]P�V��13?��*�c�)O`3�v�QS�c ��j{���� .��`j�y��~�/`kYC�QfL_�`��n�dZ���غ�\]?{�$�ū8N�4]� \`7�m���������][��!�m��d�,9.����F7�m�.�����y�]i>���ꏟ�+_�"v�CLC8�܋VÀ��L��h�� C�
L^��Ic�#��p�x�v�|f�:�uhXj���1# M��{��tC%0������A�P@�I�"D!�w5L�k� ~=ĉ�Gq��L��bvn<�S�͂FG�0j��^:��ƚ4�ד@܇d_'uU�䱸X�u��;�J"�g�ȹ�r�`'��hVx%T�2�k��"_���iE2�Y2J��))ցryR��L��1�"l�3T�<������x���=�-����}�$�/�*޻�[mZ�?�O�y�e�J� �N�����:q�A{���y睇��U4�M��=�;w�߾6��-����}�w���Pi��|�)�_~A����"����f����e�|�����G����/���zɷ��������C��3���~����3/|2MQ���B�\A�B�<*����h����M�1~�J�S#Du橄�Yd+�zJ�bNE��7
����(SCմ0�Y�P��o�g\�p?�0a��\C$�I+op,�N��}�������BfCR\���PR�W* L�%��y�
���x
��I�x1R���9������,/���� Ň�wS�,�r� uD����"9����H�xR �My���l�(��P�P�O�Y�#��N3��	δ�����+߇vn�!%7"Z��uՔ�H��O���� ?�/Y��$e��!Ln@���?��W"0njD����*g��ɭ�u%���"�$��
�,�tI���i���d�� �B�&H�8��*5�皉����n���p�S~Q�o�l:I���$�rb0ԕ�`2�C��<T>|r�E\�HѼ�ic���A!ȹ��LK:�pr3��m��*2|�X,�(A-��"�P�mYH-+řnk�!Z��йx?�v�7uI_��%8�I�m��	��F_	VK!×���w�:T%R�M[\��q"S�=�G!��t���ScMK�.��u����Җ����iЄ���Ք%+�Y�/%�S��jz� A?�U���@�f�ρ��=ʢ���4%���ԗu���Ǚ������ڠ�7��Z�`�t�m��z�C��8���n݉}�T��G��C���>��ޏ��b������x�@��3��?}�!,=�j5��?���������}7��?�E�U6���� �h�<�o��_`���1��������S'�a똫��ii�	چ�A����5iR���a�>V���4Q��:T�iB	�SqD
"��:Z���w|W}�0v�@���\ˆ�'x��G��>�����%�o�rC����dt���B[�e��Pw-q]YY_K`�D{��Q"(6s�����V�A���mK锐������L���K.Á�����}P9�2��N�g߽��s��b�E�d΂�p�A ;�d�p���Cy�V�h��/��W��Ѐ�u���܊��9y�B�����rQB{�����߱�|��S7 p��JK?y/~�s���U���7��޸)l��R����q��аi�84�b�e[���K.�ba�GW�y�M��2l��P���2��	؆�p
���H���0qzzZ�}H���imlȤ`j��Љ�an��UC����&6���"�g�A|�5��\��Hlm�PM���V    IDATg$�:U��c;.�\�Ơ��f\��{�X�,;%�|e��:`�ʞ�k%�倻�j
���L���sw<�d�����ԁ���odiXM�[�]�������*�������<r�q\�JY��1�m0�cyq	�^�a_�ջw�B�X��������z�����ܼ�;5-Eg4�dc��A��Eq���O�B|�5���l���{a��8���;?��������*U��M��ʕ�����w>��S��w�_W'P,VP�K��*��a`�\�#B��D�#��� ����A�\t�9��KS��E��X
�4��������UtS��9�
I�����(A�0Q"5�����28�r&BAa���O�D�h����E�f�F��K�Q+�}��7��>���7�7�i$��-�T��h��<��:/g��\�ł(��"��������8H���2���@9���X��X�
ү������3�� EC��:m�x.�2`A')��ޤkP;�"8��Y$��,�۔%�4P�/U�D�N[�8�kH"�$J-�H�r!V��`E�1E���h=W��4Cć<y��k���B7A��:X�%i��3�tO�)O���^,��n�~�b{mǕi��\-�mbs`���@�`I0�,ou:{8����E9��>�;lL��T�e�%4Ҩ�P��-�CH���2b���i�Ǆ[�o�p�)����eb�$b��~�#�Pqu�J��u٬L��F�af����jC�,�j�aLiS�F7L�&MA  �C�5�2|�PQS`�X�q��C��'���|��`sN�R8-$U���i�AǛ5�A��e�����*.;�H���m�`Jo��D)�<�S���bE���
�-�P����U�[��5�>�l�f�)�z���g���Øv��;�q�W`�dt�v��x��Ǳ����?c���������'�0w�Mp��^`�6yfN��i����O=���g�*L2�S���MB4<U�A��$S�"��5t���0\���p�z�����^�!FR<������I����c���v�F_�1ep[��/��c��~�!L�	���&��,5c��:����X����U�g\�X秘�E?y��ɤ�w=tZM,l6q�;��1޴ى)l:�:��ο���	������+���&^��^|����`�%����T�^t����i�Z����0�}�Щ.��c'�:%uy��:.۾f	������%�������Ms��9������$n���q���&��~���Sx�o���u�%C�Y(�
*+Q�/SH�����cB�D������`�毽
�w^�5�CMx�e��2H�e��e�p�1'�d�',:�%{g�Ι�i��G��x��3��P������Ԕ�����4o
�V M�9�";u�Ϟ�v�j�N:�Ѫ��߻�t��NzT�J[�А�U�h	�R��)����y����D���8��	��I�2y���G���	�|頶��4�ɠ��q�n�Ł�?�ݗ]���(�a���Գd��L����M�{�����3�~�jY9�GrM�����L�`�kcjr��GH���B�"[m�>���O�����`�=��%�m,�{X55���{��u�����o��?>���_�����v�ةO�#����ɉ�L��,�P��t�Q�l���Xy(M�(���	��S�LQڜ��Q-Qqh��/E2T��T��hh*`"� w����k6*|}6�'#7��>���4m薃���e�(�K������21��e�pu�qKV^5-:��<��Ӂ1eh,�7�����g^���6�@X9��.�oOKŷ�KE���)tE����s0�6���CK4n�l
(�M<(��2
�A��� }Rr+Y��0��c_���+S����%��,����b}J��8�h@�)e�i��H4'��v����4��Q����5)"��Q"g^W��)���ZY���R��`K<��D����9��+J`k&J��B�����K�f�m������u��>�d0uqW�P�-)�����[6CÙ~O(6����i���w5�xi��s�'��I�.&�(̈́�a�.�Gܜl�,Nͨ�NH�A�@���"�/�>��
*��O Q�`�l�gJ�ި�o�<��� �l�KS(W0��0U���I��i���r���L���&Z����0�U�BWc��AL�د<�� �AR���B�?h.@ޮ䗐�[ӽ���UD�Ti����1�)h�E8�+�DC�tl��0����RI&Y������,����(�ۏ��"~��o�ջ�ƶ����*f��az�^Y�6^=�7�Ɖ���k��M��v���h}�����@t�\��������W^�������c�x��Ɔ���Ei�]�MO"Ԩ���e�C��-t���3�h1б4\���}.E�]p��rc�q0��T�V�Gױ�?�w��o@����QD�"Shk��o���g��=w���P�M��B��ۂ6H%����/���	Ķ�a8Bw`�7���vh�L����A�Ϝ���L+2��!t�`B(	ͼ'7��8�|������a<����~�s���"q��BF���d8�05=���9'�2�Z�t��lT=W�Qg���u����0����SZ��e��idg��J�	�R�������4{���^���P_[�D܃�R;C�D5B���h��� ^�r<«�&ҝ[��]נ~��h���	�X�o�!}\��T��/j�i��R�O���ae����V����W��fSA/��fkn�����P=��$�Q�I0�؄t:$�!��T���]�ss��3S�5=zS%�\�RtH��=]�{b�@�"5Tߠ�Q5j�ﯜ�(���̄#R0�3�LP���9;!���N�*z�w�Ħe�p��#,ګ����|�e��iBM���"'�|/
��� �EҚLz��L�5�/�P�z�I�6���-lB��'S3p�e:�*�)���)���#������"&�6
���!�u����4P������y�ν�7O��ԱoO
~U�Ŀ�����b�?~�s����/��v�m`zjND�$�+�%N�敫�*���]R�s��|S���p��ǲ� �ϰ���!<�'��:"?:���c�K��)��T�I /ę����K�P��_hp�NaV}~cne������T6w�N�fYw 4�?@�rX[��@d1^U�f�(9c'���6��[k�S��[� gu�b>I�d�#����)+oҚd���9�s<�1B_2����M��8����<�&Ζ񥉘���r+Q�Ӄ6N�[�D����8��(X-���9n+G�����Q"Z�p#�yD�h�Ƶ��Y�a�&0$�y!���Db`�/`�PD��`�S%6���u��2)��z��I��D�n�!�oD�dR�B[�����mX�M�(��	��)���db
E��qCNc���4F�V�t�Ib����n�b٨�><R��%:p�� �� �\�5S=G���q?C���4tX��q�G#�T�����5�H�#3-�G#�i5ю��%"=iP�)�@Zuz���e×IB�$%ρ�����nI���k�4�,ӵ
j��!��JZ�J�ӛmt��Z�������c΍�Mt�(�S�@�e��$�k����+_�$�V�t��TR+�q�m���'^Lr�-&�f���b�P���Ԕ>���F�w��'R��&�Y�.P�mh�����ο�(��&x���q�_�9v<�W�(�.
�	e���q�����>�I��s@���}�C���`v��k�^q5���U�c�����g����Ӥ���@4;�$�����I<T�Q,�fyr:l�MC�f��G!��<�w� -
Q[D�ҜE\#�f��}]�^�k����}�-q��؀�D�3'��g��|��8d�R�RA�i���H��0�]�T���BU��=6'�L���g�q�֝X^���2�.ڞ$j�� F����/:��ݭ���܆��ߩ�� +/��_�s��η0���zDY킬�:3]�#hA-0Y��1Q��T�FUrH7�X'ڭV��nwЋ"����!�m��:l���ތ0L�]�����?x��0j���%�{G��UL�����u �rj&�L�j�ݱ�&�b��=,%!^h.#۱;o�3W\��_DgD"��
��l��h��n�]��Ĕ�l�Ǽu�Ü���n����1��愢���:�b�5�&)ե)�z	�VN�G�����cGP�iѪ��\/�<��Wr�.ϳ7Ƣ_1����dH#AM�[��h��b��
i�-mN���<�5y�@D��MN%�SR��Gh�`�F�X��^�l��-���_�yW\�:�)"�,8nQ���j�{)[ոr��y�q�܁{�4#��@A>�8��i
��И�B�ؐ���d��<R��s����Q���_�9���^
�bahg8�jb�2P8pŷ/��G�h�������o��?=w����ݟ���>v34��嚲�b��؍FVzVS��&"Ċ,���!�-�a2��*	�"6,z�-��,xa�kҹ"%9�50=��,�V��s�U�z&����:����0FQ'/�E��b�����/��-@uR�HHl�KE$[6hN��c���t�`��?y�W_���q��#�h1bȖh'bY�%�⪷�<U��7LyU�Vr[S>m;PY�����E�1�� w.�y���+^��1��cA4�36n9w�/�ꊋQi�3��5#b칈KED%���4]ƻ{D�M���k�#.Q(n4D��C:���=��tK�,�|�BI�,Yd����ݪmɔ�(#���]@�꣜�3T3�Nψ��s-�ǊÍ�0/���c}8g�f���)�crh���"o��_�)�]�i�r� Cq��$�w':(�L��	]�t���וi9�ԮL*�-V��>#�� ��)�lE��n�l�l2�qǴ���e�M����^n�����يS.\^N��@4��&;C���qs"̓nY�ʏQ�(��0�l��B�*0c�g����I�1t�\�T�,:q��(Z,�29�^�rK0��-���i�Ɖ��i5��t^#N=(T&-ȱ��2�o�P��D�h�J
������QOhJ�A%��2��kޫD�&?k�x^�L��85y�'�}�7FCi
8I����c��1S,����d̲�`p���̕7JB�k�?�ǿ�mT��+5XQ��ڔ4���M^:��,�%�܄�?�Ax�3���h=��� hm"�O�~�u��v'�w/��X}� ��ܗp���P.�
��)��"�]��&�V��R�½�djw8]L�/Ka�f�/��tȢ7��Ѓ:��P)Z�������n�Ϳ�;�޹CNQ�<����3x�K_�3����ux����,��9�传��H$]��ʾ�J�����=M�(�9��;-,5�щG�^ǉ�/���G�~�5�;�K���.{�m��;��9�_��a<��_��+ϣ��@-�:ۙJ<1�0�e��fK�(y�h-��"��#�����A�n��v���*��!���N�^xǞ{��t7E`��}�����^hU$?{'���x [�>*f �L����$v�Աq��2R�E;K�vL���D�^Ŗ����C۴1�L�N.����3ZH��Ч�B�$j�gF���@�sf^��E� �sZ��\_G��>1�Bٗ,�.i�a��&0zm��O z�$�De4@E���E�9�&�mA�e�9�'�,3s�v��>���f�E����	���X!��@��Г�C˃�:mP��z'�S� �j���4� ^|�u ���0"A�qpl���+�͟�.��z���g����\�'�����kj
%����F*E4x�0S`�*@�ߒc�T*('`9�re$��&�K���8���a��GqA�E��cdE�!Nt�8�iY��k�~�]�W�n��ۖ�o��3��o|��?�7���_?q�b�G�R�m�yR1��YH�P��>�Y�?�z�s?aA�ń���Z
1%��b& ���J��bR#������m8p�.l+8h�>���a��i$��p�+��j�$����z+&o�	����U8�z*l��x7�"����fk~}������paPD)�BE�+��*��Ӏ�fHc�O������͗y��%���0d�{����c�c;�#C�*�I�����^2�uI��I���TS�X�bֱC�m���TĨ��L�̨�Sݶ��Y��@�S��������fʫ������&\9@@�J�L��Í���Q<PV�Un�OH���@)�0k{�ޘ����a8�òti"9�e& ű+���o7�!�z��&�H}6FfIz2�$n��PЛ��(��C���c��Y�-Մ��gJ��M��T��y���G�*V�>D�+0�,�6q���2A�e�&c�W�I�֥��s��Qw8@���gZ?N������D�8��u���#�"	|�D`!Ku	��i�jѢp�Ӄa��
ӱ5�f`�T�D�Ϣ	�:��d��栋f�-y��c���d�&TC�
<�Z\� �0�I�&BW��,_�Ê�à;�dd1FQ������D�+����C��F��`���(�&L��&Os��k��KTt3n�~.��ФQaS���eHb#�E��t�l�}��`�4��pޭwb�k�����Xx�Xa�:��2J�e��o����a{@�����?���}���>��ԯ~*�����>�^��ob�����:�����}A���t���ik�頤�puS
p�4�ґ���P-פ������g�����67�v� =�<���=��m��-����/�́�U�R���֗��7�����et�P����k���[ދ�;.Q��^$�/��-IrQ�FH�2da�(�O�J!K�f���"n�ʣ�\�K?}�?�0F˧QB&M|R��E��~\��� �fE3p��G���#�=�S�Z����n\s�](�w��ә,h9<���fG�[���S=���[*\�L�W�`�-�f�~�x�K_��შ7
p'�w������� ���,��0���1��>L����}��A�"r��G��:��]�6ph�Ew���w]�-W]+�#�0�_���D��-�"��d©k�p��Α���_�z����[D�⷟"�"4��Q��QkTaq�JtX��B�"\[���������2
�>J�8�3-���L�4<���ż�(��Mq��вQ$t#~5�i�̦^�cʩ����)�C�y�ș�'8���k��Sf\�T���Ι�<�S�p9�-4��M�ob�n��O��o�^�"�ÛIѻ:��n��K��Sl�8	
b%�Sk��I��J�G��0M��noS��J�߯�Tj���z�2f����7p�;�����8�H0MG��q�:-���~�u_:�O���w��W��^�m��?�|�W���������?��/��Ƒ+Y����x���Ȅ295��r!��a����y���~��nh2iȝgh)��HuA{�"�H,�xY�=�i\�u�h����3�N�ވZ�,`�R��+���\~�ZM���P@qfU�1�4����b�/W�����ƃ�c�����/�.P��Il	�&�"%�b��8B=���'ȩ@�p��Z�J�#��]%�M�'o�5����<l^��s�u('n���)Z�Xl�\���3���VS<\��D�)U����aXtp���B��⠏{rki'��:�a&׈��؋f)<����|^F�K��7#[�/A�RI8AP�Ű�pF��l��G�~�Jj`�T��j#o
t�iJE�B�N���u���a��)4��i�N��INujB�i��6ӱa0�T��&    IDAT�Y�D"d��L��ʰ�&�~E�q6q���֠��l��h(���n��1S��+���Hn���:�@Ysh�j���+��ZR(dy3����l0@BKb�;>j�*J�����}l�V��5�;�V˾6Lh��7��^���$o�S=�PwES� ��4Q*�u���LK\�3)���O���AN[�Q�7`SwB�-�3�B -@ҿ��^]C7
�'O��9�L/h)��� ��"%/k�P�%@�h�I�%l`H
s������L6b
��}YIc�@��1�0Q��������`�e^I,4��b��#�0��a�w1�����p�j�e&�9N]������������bQ��?p^��7p.��X�lن�k�����J�z��q<�����_e-���y���ӟ¶�n�:�I�T,�SiF?B4�K3�t��NWM6���\,X���^��Cx��_��߀���q�x���>�.G�b�Fq��ケ����%��_D{mӻ���݊+o�����E)�DRmU3��Q@-�*zC�#�
��V���_���}�SǱ�苓��s�M��~��*Ǿ��3��g?��}5?By��K�����O�<����(�0�Rɬ�8Y\��Q�N�aW�$���<w��M�[�oݍo����3�����2ܪ�����w����n����|�54xk� Sq���GMם���C�S�e��F��i:���׺��LԱ������1,���x%y�ŉ�|^�������Y�

~R-�ܜV$2��P�4ۛ�\�ZE�i�Y�j&��F��k�0N���g��J1C�B��e��>�e6���B�ƍ��-z*��,����$�Q<��<�X�E�.�����-æX~��(�D���q������-���j�����6NVf�N���	��G��AG�h�n���p���&����m���>DV���i�̶�}�Ps}�T�4G*�����e]5	�!��M���'��1^�a�O�Y(.�V���w�C��g1k�(�̺����#�kh������ʍ������m���o7�*W�_�s|��_���������~϶-i
�ڮs�+OӖ"S(5�v���.d�����{� 9�3M��,����n�{  �� ��E#7#�����n\����F������P�HIK�����;� ��h�a�wuy�U����e503�����1?�" ����2�|��<�dA.�� ����.� �8��!;���cn&�;ϥ$�P�EA��F��#X�b��h2��|�'P�ahY%�!��U"�f���ĠQ�1v�t��6f6��_~�[$R��칏˴ ~�(no݀��'ṝc4��SǮ�3]4I�R���?������ǀ큼D�`���
G�v2��;�"�Y�re���*�P�,�|T���.b����˄����60�Q:9z֥;�SQ��B>�A��C[&!𡞼!&;�b��,]'˅T�D_4	��?��N�`�	����y/y�qǩn��dJ�^@�G�)/�N�$���IC�%I�u��Bce�HM�����X��D1��\��`�{2	t�z�*d�i��k��q�X�����N�NYӀ���W;I�tQ�$�Eu���ը*�bk� ��@Go;R�4b�84~���=���*������3u�u�+փ8U�<n�&R���(=��&�&�&���S�qz"�,j$M�O�M��e����Xҙ(ҹ�H��,O��� �0ɴ��'Bn:�jbL����+jj���3���s�S0�.�p��b�>Ib����0b$�м^��򳓽]��������s�k:�SY�Mg3�n��,�	"yGF�|�T�+T��;Hʩ���	�K�&�121�	��񾑩!_���C+�fQ��0�Fu ��ۏ��@�2ћˢ#�~9!�D
CNQ�agx]H����A�%��@��f�sDG�^���J��2p�-8fMuϩ�� �|�"w�
Vk����|�9Its�n�ຍ��ӟbp$ �W@����k��X�r�ʰ�R�S��,t�S��E�!�%�'�X,���	��|}{;�ڴ;~�w�f�teBV�<
^y���#���E	a�Aܺ��?��?� }]�P�4Ӟ^��Ϯ�����i,�R�	�dSfTh�Ŋ4$~VrRT�Ԝ{x��q���o������u��G��mUVaȌG��w� ���@����g�����6#���W¸'�a�믣r�$���A��F
�[���J��q�N����� ZX�c	|�u6��{�����p,4Lh�?�*'�
��k�nۏ�[�����ߓ���@�����E����ñ�oR�� ��q���� �,���+V�Y;�i6�<p���씆��wHVc/�.B�TS�$����]q֒"��s�p��A�1�������	y`s:�y7��2'H_�����a�jE��-10�&EU54o�g��3Q�^.ӈcxJU,��1�z��#���d͙�+'bE6X�(�c��JlT��,<���Q��KyԄ����'""ӚQI�R��!F/�w31�Lv"r`��c��V�I��l��hE�&��2���~GN6�n�.����\5[�����FU�0�H����-�)��?T.�/�M^t'�<axS��]�����,*5�5�P������Kwv_���+��?'<���"��(�q���e]���pj�O~�ӟ�={n���qa#e[I/vR�) ǁD��M�GI�a��r	�E
R�E�	�4���'���B��G(W�D�dS��R��IcP�Q��P�k��2�A6�D6�������k��7�A>/�~?z�n��U3g�.����G�L_�݉��8����xᥗ��;yw��G���ṕE���e�� deR��Ҁ���w,���n�Н"	�@x,8�,
h宫NA�4�|�������kR��ü��v(�	Z%3j�3H9B�J���\*6��@b+�-3���#�F����l�2Y�3���"��M����r�#�	eظ>���`2�G�떎jA���j��j����"�r+��t��f�+k�T��,C8P��p��*t�d�B=�]���TV P^=�GN�H�=�'�dM����۫
M��Q^V��bnF�a�`�u�t�C&C1_�Qw�¤	���0�pX%�D���M\�����������Ȱ�1|��1%���������k�r����rd�9D���m�'\���IY���w���-�,B$#��ʺz��<	�͏H��N�\g&��/�ꥳ���&몪~0���Guc2E�,

Y8hR��#�#�Ԅ��!��1M�'I�;+|v����)�\��c{w���[�TTb���0m��7�X9�b�������s���Lބ��
c���!����#�?~�.�]��;��C�$D�=�Ԃѳ�j�X��� ���>�?rm�O�m���T!����N}�NY
����� L�@U~r
�ᠬn_>��LF�ϋ��M-U�(�Н�/�<��r���z�$,�\����A��5���5�B����ǽ[W�H]U73_��u��oX����Ck]�.Y��S�����py�n|��=CiT����~C�2Z�٢C��,`Ճ�l�yX�@�g���[q�HX�@�=~�����ņ�8���(7�89_uM���sh^��k�a��u�-DOǩ��W�7"�Ehp&.{�W�Bńi@�E����(\�C{�:��A�A2te��R�]�'��w���u�JQ��K2��1h�t����f�D��D��7����qh�Z�Ix*���R,~�ۨ7I�\�m�D�������� z�w-��'����Q�����X�����0jH%��*�U��w�E͌� "�ٛ�ؾ��l�dv�`R"/��*�^7��ѧ@$C)p@ތ�-E��hz+"h�?��Y�PS:@���nu��K+��2q����ƜC�M��ې]���J�a�)O)�Ү�.��.������j
���9�z%5��Ľ}��}�u5�T�,_e��2X��r��t�NyI"�'�Í|*���N�vv�q�-��`�� �X7�F@.C�R��S��P��N�}n���\�D��/�\)�9����E*�ӼhOTA����E���!2�Z����3����|˞Ճy/���-�HT�X`�sd�;�0�J�N���ڲ����#¬)]�!WN�>���`B(R&�y����39��](��(:�r����ߜð�rn���.��Q���/p�Q]���fM�T�<��п���,
�;.�����Q�T�2S�S9���������!@��J���I-5�w#ۆ<t]�t��/��\�F����z��r���v:�e�����vW^�vc��#���h�#Η7�ܬ�΍� a�zǂ'V�Rg�
��aW%1���EKFw��e���&\�/��Tܦ�Z�(��,
RY�RX;���UQ�M�$1(P�*����g�a�/� InN�n7��������?cF�^��۶�=���!x�w�t����߳��O�ݖB�I�Ӡ�F-3#��9o��ɤ��@��h�RaO�K
L��d1E-lu���N
s���X,��"n�21P�h%b�(	6�m�U0n
�x���TC}�tj��ѡ��)��x��yp�EA*�'"����@ՅTA�VQ�	3gc�رp�Nf�YD��O�k_�C*�/į��Ll>FO�!�$P�]����7��őCH�Fe�sØ�`1�O��Hy�T/q�� L�Mbb�XT6�@e9
��f�ɲH�{�MF�s�W����΋��B��ј6s.��bF����c�,N=�K��!����aðb�*����b�]��FG���غ�Ct޿��PU׀y�����*�����F��9޷��_n�3�-��Y�᫪C��a.a�w�\���{�y����f-��񧞄o�8�Ϧ���^\9u'��GW�Yg��Fc��h59B)
&�	=�Ɲ�p��I$�v"��K�7��:�q�$ \�G#d��n]�G��;\<}�uX��jL]�J%�܀���;ځ=�|�'�Ȥ|FÈ�X��[������r9�_��w���-p�n1d�L,x�[��>[�}Xm3���ù5���-a�v �=�v#�B$䛜�P�4W�D�������A��Y݁�l�>�a��N �s[Q�*7��Ad�.D��*dq+�/�
��'�B?��-�1a�R4̘���V�;�N��S5�	��z����V�ظ���k�����x��Ri�9r�~�S��^A�L�n�p<��+���Y�dL�l5�nI��5f�<��FU��� :��b
WP�"��ؕ+8�n-No܀z�嬌�[�JL}�9�x����cʮl��{w�����c�B
��J�\���zU&C�������Y�xh7c̳�d�)�#(��O`xY tw������u0���`��|ɀM��`�w���Q���*|�1��>臿:��+�c�;o�j�d��T�gQ F�`)��8�T� C5�b�hOW(&�WKAE�iߴ�{��W0���4�����Ѳt5���Km���:6oFS1���F1���/�%ο�t075%�I�ǜf"f�Q0�M*���Z�,^�Ͽ��Q��pڠ�L�E�I'�r��q��sƖ���M+�^�>��`��&��/���V���#�Z� �<x�3]"�A��T�-��=�x[&O��i ���S 1�c|���UÏ	�@��`�����82�}�Oy#���jj��R�������<��~/-��#7�|�<�h����������;I��dhL�&��r��|�h���';�!��������^FUK�!e������웄�(P��-!VkҰ�'�Q�e�[��ep���\^xY��5(��a'���	��F�A�o��я>����b��FL�;�����rX�rr"���<U[�����;R���o��U�I0W��b����~,>�sx����v�d$8Z�:v���5�)�����բl�
��-Y�<�Ψ���5-[z�&db�Sz��/��4 ���Yp]z�t	q�-�Vԝ�f:M]s�ߜk2/+�#����;M�ri�ŉ��;��Y.�Pt�CC/��祉̔�j�6�-�,�\�,�a�S}|�`�P�L������hǜS���5Ӵ��C�ȌB����7(��4���
��_2��St�U2��Qq�2�L#OȍA�1�n��if7������9$R)1?����E��'�M��d��n�PY��뜣)K^���*��|F�L�XŤ�R	���/ӄ�����=�e��a�c��f�> ���u�̮�8u�(�*���[Ѓ>Ŀ:��[?C��/༗D��^���:����]&U�%U
E��Bi�P!A��%7Fδ� �vӒ)	Y"Cj>�`Y:UYJ%N��)~ ՞D��ցVE]_�1�R�]<X��@��@�4���̀O���\w�i���b��n=�75�Z�W�F��1�Q����ƭ�qh�6ٺ}��eS9a�}�u%�[����D.؇�Ktݽ'��)ë���P�=R	6�eq�mC�'�H"�T�-X[���j1���K8�{��+�x_�s_��/�G��ۜ�Ir{j��پ]w�J�5n"����#0j��ŴNaz�k�𓟿��7n"�-��~��z	SV�Pdua���&R��cǺ��p�$�LF���_�c/��ԉn�n'R׮���8{����H���4,}�T�CK_�03�I�q��.�߹N�,·���U/���)��ʚcw�@�W'qx�V�~�z�=���z�g/T�˥�r1#�0�����/�ù�_����W<�ǟ�PѠ¸�G��~�N�)�P��'��?����&�y��~�7�Îu"�)"��<m��:�N����I�[��	\ݴ�֭A��T�?O-'t4��!S%]�pM��]�)`Q��8�s"�9D��;��rir�B����2��|!�T4�q5ه��]�����Y���T�b�x<��%zl!b�n��g�������(���P3a2p�.�n݄��}�X��"hZ��˟jj #�[GO`�_�������ԏ��^{�Y��7���7 C 9[|c��+Gy6('�#ɷ��.�}	q���Ξ��5���̤�H�4n�if<��-�QQ���W�<��߃S��%Z�r	�*�0j�"Ly�T��gy-t����8�U�tB2u0I&�:#$`�s�38���	'�[7#�6j<��4�k�ыc�s/����m�˷��'[��߽��#�PMW<��o����c�b,%o�򎌝��M�够�H>��m)���[	��x�����M��7?A��%��ze�X�����y��v���	�]���nT�)��$�$��.��!�:��>Bu4S�co!�v#�k���A�B/�|�d@�"��#�Տhwҩ�p�~6�\�8�$�Ʉ@e4����r�x�4�I���q��u�ik�ι��x�3����[n��{,z���?��ݻ���,\�40f�j�IB�1�(!&��}
R》""�bp?�	�a ��H�� ϐ*z�ʰ��J�BI5l�R�~�h��8_@��s�LQ����X�t0ձ�^r���P�B�ǔ �T�J��É�G�~�fĊ	�]:�-�7q��}\�Lѐ��J� ��9J��O�J%�L6!h	�[)/򚸜^�{e�7�sT4��q�ߩ4Ya�H��V�'����Ņ�{�u��7�a�쩨;
fY)��X
��s]!8�|و�ֵBщB�X��x��4�p�Y��2p��e��l#���f�,D�Ĵ#Xf��0�t8�Яi���C���������|:�`
�n�i�ãi��4Ys	��ϒ����L��Mf���+ ����&�ղ,6?]:M?͢�4-�E�3wL|5��K%D�P
c����L8�R��3�*�*��� ��R�k�&�S3-K�4M$r��$�N�,���!V�hIj��e    IDAT�ݓg�]�51�QΥċ�a��|��d��ћT'�A�������-��������$�wÇ�y��N��W�E�Ȗ$���7u���X�IO�8�����4rH'����Q$Gu&e"���2�`BO���K$E'��B�lIn��a�{�c̎%�R��d"E�1�A$���DP�#�E���XM����|A��~4�����#S� ��TTH�9Crb���Bו��q���s-�`st?��A����lO!l��"����	��\NDJ�C4Qu{����4����c�.�+�x������s1	���4%P$8_����X	�� �ʖ�U�e�|��5@ W��o31)DmY9<�Xȑ"���F1�A��F{:���8b�W�BȚN��c�-�����ǞYP���S$�t��^�ڷ[>��ݸ%x�I3Ū7���Gg��(�0m��;,���(~�����n#À������c�W�Q^	Ӱ�3��7wK�����!��(UB�4&�����bۺ�ؽm3�z��	�a��x���)�ZQF2��(pj�z�l����l�M�bP������'~��^Y�q��sX��?ý�7�Jf��'W����<+@�V���s�2��S{�
�h˯z�u,z�5���IX'��(��������M(���'`Č�X���h�4E��ԆW�I����qh�F$c=�e�hl�g�x���U��I����cؽa=�\�(�z�f<��y̜�U>��%�(��%>y�������e��`9�x�e����
�����A�wⓟ���eb=>�L����C�ZF�ϕ�D���Цϰ{�Gp;r0�F͚��/��G�Ά��I���}�N����pt��`��A��'�7`����C:�gej@��z��ax�
�/���2�KZE�t�q���i�E敺��>�E�e�����T�b�x�|������6l�;w�=C��1x�������ٻ�G��]( ��b��P�r%0�Q*�{�Oa�_���_��^H��e��m�_��E;�n�;�LT%H��[��6N�	8����s�8]�#�kh?}�֬ō��0��-�#�-��_�s�4���^���f�?��?�)n�8=G���.ä�+�d��0|�2�u`'�#����������Y,TE�XK�D��-�ݽ�v��u_�?�υȨG0a�
�\�(�2ҭ]8�i>�뿂��CY}�p���:|��PgB�iA4r*������S�?Ӊ���C�
_k)N�Q�\G�l����27�cD}9,-���%�^�
� �IdN�ƕ�?@��-�S�E�4Qթ�[D���8ٲPp�H)�4}���F��ZTM��	O�@��)H&b��zb��s�N��96�mHP	��,A�	�p�[���}��e��x��z�XR��^b��S�
:�LnX`vw���eD;�z�`�4��zQsS�'�h�8ۍ'6��{�sbN�3N10�ȄKC����� ��^���|��(�"[$B��L&�"<R�+���
VJ�����O�jh*�l~M��	]��_C��h���p��E�.-���<�~?=,��РUG�<G�ip��,�y����;��
��^6��06?��-�ODL0z�^ٷE:�b�;���(�K {��h/�ʃTE�.G��D��������'�H�[w�y�*5��P��r��0�oz�Ӏ4�s�(碑�Ⲡ�5Ksj���;���6�������<]Y�p���&�����Z]]��BrJ.�\bZ��f��T�
���'�l���Y�4�xH"���UL�){�����`˄z�@f�U���@�-Y��%�����0�uB�m��˫�T�v�IV;&�:%yG��"��C"	�-��;�ǛB:ߥ��!u���/������3�s���M%<!R2�&�4�JM�%�qr�Rj@%���d�c(1�KD�R�Û��U >���NX�N��� Lɸ�?���J��e@���g���L����ۋD�F&�����e�eR����cM O)���!�$2��TY�K�Y\o�q�Ŕ��0���1k�8T�udz:p��E�w��H-`qru��fYm#�|
�]	o������UĳY4���@#��!����g�ܸ�/�~��S�ͻ�u�hv4^fZTA� ̃���2Ѥ�mpB\o����WT��9�������xc����ԩ��W�|��X��K�˄�
n�6��rQT���;�N�����4c����99�>���
yq;ُ�h/�3Yd�\~�An�IM�c��Ŝ�Ϡ~�d���ס!~�&�܎=�J�M�䈱���1o�r�|�DI�򰒽8{d?~������5��ʻ?�ϽOy��߹���w��-�`Q)��ˇS�+��C��5޵[֭C:����c�x���0v�t�x����X��l�ѽ{�y瞘ʄk�0oٓ��p���Qw6#�ů���5���ۭЋ:��&L���+�A˔)(𞶊0q\8�{7�GO�-d�)�u��>��~��&�DQ�*�z�kX������cЈ��t����U�-gb�{�nބ[�F6��, T])������y�����q�&N�߃_�@��>r�$"u��4�<�'P�<�_��|�Lm�Na�����\A�r`���0���0d�T8�eb�d��v	���^8��{�P1�	���S��WU#��B*�g�ıM��z�8<.��鋟��O�]Q#�^8�u>���;E���G�U���yx, s2d��5q���P��#@��
�Պ��׭T��$�͡��DC0�j_P�.]�:�s:۲idEd2� ֎���O=�(��ps�A|�{?��{1c�B�}�8�ꅤ�:�wv�+�E�B��y({n��h�D߹���?�Y��Y�o��o������T���A�\%�̽��/�1�>��F��72xT&x4��3s��t��i|�e3n�߇Aa�}^�X�3^~h�@Q� ��@߅�8�w?ř��ec�\��K�a���Q1a"rl9���Cp�!N���(��������-�Q�Ō-QM�\�z+��߇k�¸U��Dxd&<���.���H���n܉O���HFo#RW��+���7^��X��h��ZXD��Ԛ�(�C�l\.����P)c�ò!oQ�p��B>weL�޼K��{ϟCKuEd���^��U�� �A��S��_�G�N+�)q��K&g��7J (�!�`�'�K#��2\�d8����DU��ƣa�h��x��z�����/�p( ���q]���-��9��bA�&X
&`k�˰�Jp$�2^*�Rq)�U�!�]*��O����Lڅ�E)W��U�>������7�/�b�{�=ђ�K|u������)�TìԸ��&
D��Lf�w�&�<�i��܎y8j�cbğ+�ՌT�$
�̨DtNij)�y� ���W�E�JR/{ϗ��&3��H�T�y�4�dm�F�ܘ�ۇ���*�m�*E��A�D�p�BQ��<�L
�_����G�A6 E�E��Ť��#m<%�e3�<u>L��:u�@�9���p��*�E�P0���ZYS��������������N
,�r�u\&�����ώ�,����tAxQ�(	?���A��'D��X?x^�I���*�<[}�F� �#/M[��;+<I�T2�y�َ :xvK�7	gT��_g�����O'��etd������ �o��l�x�\(��(�~��:�ߏ?T7�fu���U�Yx�7�
�
�'�>����?gr����ѐ8lO�B#�`LV�`�����A(X�*���ʔ��M*��gǓ���}Q$1�R)�44v���t�H�dQ�ӟ@gw�i���+䧠���U�9a��Z��&S&͠`Z���aڸ4V�`ژ1�2���vItn]��\"3k!D�_�N��g�|Mf�Nu��%ܽz�.�C:��БS0b�48	%��+	�)�_�_n\�����wFI��4H�eM�e�����STQ3���CB���K�/	b
�X��'E9P��Lh\�R��87��s ���4�\|?���X(?� MN�Z7L��m��J;t��2Ԁ'N��>���>'n�w�-އ{T��.��'����G��@ٰ��=��-E㈱2�7�ܾv��n�����pL-�p%�yX���hh�@ȏL2���V|uh�������9����;X���UB*��[�h�#eȱ�楔�i�R9�\��i��u�:�:r�<(]�lQC����-���3��҄`ȏ\<�x�]�ݰ�>?�b�@8\������S0i�\�7B������#�g�z$�zE�&�/�b�P�_�4�/~޲
d3��k���p|�v�{:���E��UQ���b�(����]���8������K�DP_y���K�y�8C^$�1ܾx'v���o.�d'���N�!C0v�L���(���Sv��?��O����+�yX�m�I�cԌYp�W+,x6�B_.�8���!I��l�-���L�������r�}��a�G������@y5&/z����!C,������ůqj�vغ�)0�'L�c+�C��	W֋�p��+i;~�\
U4ף�b���Y)t�JkT����Q���k��R��]�� �][�Y4��hō����֑s����N'��L$2Y��IxC�n��O�@�S˅ ���U\��4��	L�;�̚��|���~`?<p�P?w>�ϭ��dB�w�
����8�y=�b
��1aœ��	8+Ò�LD
H޿<@1¢S��n�1!`�#Ttb�T=G26�oC.'ڿ9��[6��έ���rz'�h�?s_�a�Q�p�q!�H]��C?��ܾZ���J<2�q�<6uӦ���r��t�$�XSR7��z2��f�#㤗	�j��B�pg-���ݼ�o���彻�(����:�ki���0v���BU�� ��8�~���'��܄�̇)O>���z�q�T�48�ө�=� 'ɡ6d�@iMUE���[Y%�w��Z�p�Ě����/�vC��蜆Y���+��߃�j0ПE��)\���mE�Gc��I��Ҭ�n�0o�����-�����A��B���\��A����A�h2�{=q�m�Жf� ]�����P_�}D���v8	Ed_�L� �	��TM7��$�s�t�$�dE�S��`bY�O
ϟR	�i�%I��4�k<�K�i;�Z��/��U9���<,���<;W�� 	��^#�2�)5[����`�%F�!Qy�eS�")~&kK���'�:D7pz k� N?99��3��d��P�������=�\����N"*�5/H��JA�s*�{*��/3Q����'�n���)�g) 
�"��V�ȝ����Y劄�g���.pb�Y�>�r�
HUE����
���k[+�j�/�W����L~Q�������T��EӤ��M��a2i���(��)K#P^	u�UR��j��K&��`�-I�}Q$�h��'�����>�J��n�|��N������8k�A��vT�@Qfr��^J�g؍G����R@�3�(�Q�|O�(r\v� ϋb�-�U((�m�((A����6��4�+���C����'mj�ۛ��RJ3�pUUU(+������dKJ%�!��q�1d҄��k��4����Ggw��w��0��8�	R�+��JnKc9�W*����E옆�p&o��I��������깳���|�_t��
�j�p���?E㌱�꾇�'����W(�n��Au-�>��&��a�&��X����C�aݸ�@4�Hւ�vN8�]t���#F g�Ub	��(��� Ʊ4Q��j�(�w^�P�.1���]c	� �fDR��Q>��k;��,� �2���LMd}3���qIज�*1�ŝ*X��
�^��}>�\:RNm�^�)����y3�����
	Y�F<��IS���0e��"�K��y�
voZ�s'�HG7_�9r`�	�ַ���1PVBkg�U�ڿ�6�A&ڇd*��,}�E,�e4)>�-Ri&��ЇP؏L:�h�$���k)-���Q̠��U|qp?N=&�R"W��{1f�l�{bꛛ*A�'�����5��/��Vn������c��9����	G&řϏ`�����v#�	��/w�R�!�V� S�t*���{���	زw�^B(�ai�,~�e�\�5������q�̗8�wn�;7a|T*q�1d�X,y~5G���,$���7o���]8�����b�-�0k�"L��8�*����юk�����C�~E�L�T�`]��V<�@� ő!쯣'vl¾k��y*����U/a��/�b��}�t�λ�������	� ��p"��xf-[������.��{�&�ڽ�>��h�@!�.�������1Sg#@��QD����7{�!��f�<�	'�/�)�#bQ@�U��+EA�ۏgq*p8���ў�� �,~	GPH7�N�y��>�@W:���E�͔l^���xd�|~�Y�q(�tw��)¡�MpTU�>�_}����a�?_ր�.C��9�zhnfK�KWq꓏qp�g0rq����b��'����_H�66��Dq^�C�BR<��ϲ'�^�5��|��E�޾���@�^D���n�Y�����?f*
^��#�Ҝx��¡��'6~3�e�&N��?d�,h�
@�4C9��|�pF�_�)c�u*�Hr.�ʑ]�2��t^���G���C�:���� S#F/]��Ͽ"�7"�ڎ��mŎ�~�\���-�So}c�!��!�����zs'ܺ���y\�+urM�fZ
VE�	g����3���u[q�Ï�mkE]ă��EhX��f�|z�h�F���mX��h'��$|Z�'�N!b+�KB�
r�r�҅t�iͅ~�}!/ڬ,��$�^�����a8�q�S�Ǝ���cǢ��
�tV�Amwn���6����A���d%HeCDi�d|�(�Viqr��m%y�r
�f�|��8��[T�~@�B#<����ܶ�1��|J"�@�b`*�ubs|���'��!���<-*eҔk�i�k*9� >JE�-�k7j9%R{��t�����s�HTI~-����IY!r���$���Uϕ����i��q2�T
J�8)㢜��E��+ Q̯�q"`O�D���D��#>����W��#��
(]�"�vc��@��R�{i	���%�e�N(8t��U���/"��?W>f'ȿ���_ĻG���Lţ�Ԩ_u��"7��4��z0�zP�<�rK�7�qPw��t�Ո����8>R�|�P]��+%V��T��i1��M��j�� X:�J[�!Ҧ�@
L	(���=��]����}�G�?"���)�(��b�a�")ٚ˦��˞�����jAb��P�B4k�b���l7@e߭�m �p�HN�B+�����&\t�%N7�f}6�B�#/;�C�C�]=��ޅ�m���!_$��-j0��@�o�~hHDGK�Y9�l:#]%��@m �qÆbls=�4�3h�rU��H�dg�Q�Ԅ��C4>:�x�؃����h�o"G��F����To��-�h�ۏ�ӧ�uv�3D�a��p#�9� C�A�]S��s�ŔI!]y�l!36+x��M��"d1�v�IU��dj��˦�[�8��-<j�(b���x>�D��"n$2�N�����dvw"'k�4M)҉}u������$@G.��|]y,|��>�������~<��Sx�շ0v�L�n�M�;�`��u���o���ПȢ��J���?�72)�\!�\'N�߉O�+�u�G&m�3���9���c�L�`���'�R�����DR�&T�p���
�p�N\=��cߖM8�}�\<�E݇)���7߂������g�J`��Oq����m��{}	�8+_}�_ ((���`��7g����'ܸxTH�r������`�sp��X8�b�u�+���W8u� ���6���o�Nݷ�    IDAT�?�PY�s����7�o�'طu�����L�3.ŷ��]��� ��	�Kgqp�Vl��Cq�N��1L�?�z�L�:.:�$\��ikŎ������D���|z �'_z�_z�H��X�s�w���[>�~ʨ������Ʋ�^C�i�z�`�{���_���-Hvw�����X��+x��WP1|
Đs@�_�ٍ_���%R���׋�s��?�S )@ֿ����Fq�e���8��C\?y�lAJ
̅��4�z�Z�g�oT����D�;���u$�)�����6oʤ�����PU~�(t]N)
z�y)
ړ�b�< �5<a��y�B׀rBgN#�tֵ��0n�ڍ�B>j���(�1~#FI H|}�>� ��C6׏pc�<�	K��];�h�ǩ��r�nq����N.�%���qմ�	�g6+����;�����׊� ��j�<��?Dx�,�ްp�Jq]]��W����?@*z��r�N��Q���y�l���^�����~JLrO-��(�e�~��ع,uFU#���b2%E�����v�0��NԺ-�ۻ�1b�<�|�m Rͮ�O�������-p�Q8BN��?K_~5�Ǡ+�E<�E>�T�<"���t�gR�����iN+�Y��ؼ��rZ�_�IA���oځ����@E�	�c�i�D�x�]�N�MaWX_]����ݽ�F~3.�J&�n�~��K����eHw��n�����!c9���W�u�X)�X��0k�RT4õ���z��67c��qhll��v�~�}\�v7n\��0tH���tymu9�ȳMMjN$��ν�<`�p5��)A�?i�U��iC�����'�knW��\�T(���*�R�6�e6I�VB<�u�J��
��K�:�s%[�J>S��D�B�Թ�4������S8~?��H��϶�����l�[�(@r<�Za$W���sm��&<�N^9����,)8'�^�5f\�j��D��B�2�d1���r?�Mu�ja#M�Q�35k��� 9�Z�<��(aZ�D�_�<%$Q�����P��O4M��,�i]����Ls������B<�!;��(E����=(
LT��Ͳ�i�Ѷ�Y`�p��Xh�\A��t�>�)W-"�l4��1I��_`�re�-A�J�E>;+��RH�X-���7�mJ��* V��^*������leQ���8p���S:���`�*W�LZ���H��� !-�y.*�K�(D�e(��@(�E"Rh����|:%5�Y �c�u�E������v���{h�ӎ�h�"����[�I�t�X�yRаR��H������p�.X��-C0yh5�=�q��9���U�L��>�5C���W_��'�^_���O������z��B������#����9�0xd�{����ޱ��߹�
��Ώ@��!aW���Ș@�F�1D�q���˔I��8=ꆖ:��
9 �@A2��KQd�e�Q(J�@�%��2�b�I�A&���(�٢8Tk+��bjDS4��$��#LP�?فX�%�N��i����љO�=�VEA�DVw���ׄ��(���8�{�]I��NP2���v�a�������hokCo,_�V���_U�Z�L�4.܃���o��v�\Q�qv���g�S�<�dH���ɢ��S iԡG�����<�/��k�+��,Մ�H߿�]�a��u�����t�1k�x�wT/2�դ,��}�}[�����H������������f3`��N������g����{af`�3i���K�D���sw#��g>�g���H���t�����0o���ˤ��.�q{>�6��y�@ O��=�$��� er�j�
E|�s'>��/p�����k�1突���	Z�LR�*��({���ݾM��4�u�X���`ɋ�n��AB��-�[�;l��#��ᚚ�p����²�^���Db&�:�m�������Nqť�S����^{��!�p�%���7������t�}!�^f.^����_���Q(0�!?%E���8��oq��~�2)D\N�	94�g��E?�E��#>�tb�D�Ԑf��[R�h'\D��Q�i���Q����A��DW.��D��Ry����8\��G��y�|`�d��N�R�ϛ@[:ϜC�'=}͔u����6�U� *He�q�v���[� o$l����1y��0#��(���$�^U�!�?�~���By#�v�.Z
�h�	ݔ�ݱ_o]�:�@����?��G��� ��.��l�)������O?���=�� TS����0i�S<}R./������U�m�UR�l �A�<��^,������ĭ�����[���BcЍ|1�"�Q�ѷ��k�nŝ�q�����mp9��.�`أ31o�j;������Ņ�
�$�d��|*M䫉HoQ����Aq`�J�YD>����{pu��SQT��� �2{
V����L�<��7�ܵ=���6���W��'�6O�`�
6$�K̫L9��x�^�#tIap?���`L_��'�=�¹���1��U�p���v�n{�z;Dvt��1hhF-Pam��)��(=)
�a�!["t��?����v2.
9�ժ����N	�Q�}^T�
�^jw�}�Og��^��� �����Y����!&yJ�T����8WK�P%���~�����	�t��$���"�T��WX4K�W
��.�J�����PR�:����i\&S6�l>�k�S��Z�F�hr��Sa���jʤ�.��i�(k	wC~2�s�K҆��(���x��I���6%��D��'<+�;��1R|O�*b�wL`����Y�xe4����X��|��'\��mG]�N�V�C�8%�����WSe����b����s���+���C
������K�h0�D�(x�����K%��9���Ra�G��x�ҕ�+�����(��$L�ը
VMD�Ih
~$�[�u���L�l΀\X�>Ň
�����9��L����f��WV�
��+�����")i��r��gS	J�DU�ߝ�kv����┠��w�|�?��1��$|��X�X�M̀b˔��H%�J��t�n��0a�`���"y�ns��Q���s��.��~���}l&Ʈx�͒+P�߅�s��z��@.<� �MC1b�d���Hr��'q�	���a��L���6"_D�Ԑ���5�Oh0؅(q:J�S�0K���?����5��2��ؖ�:T�d�I�بӶ���O���"��ł`�����WM����c5�T'���.�[iX�������I]o�]��b�\�x��Ȧp7�@G��89���EГ/��$���a�o�i����븍��v`�G�ŭ�7���W���������R$\ع$��$����v�d�z�?c���c����x$x���$��{�{e#'��4��}[�b�{�8�s�|��"lk��c���X�ʫp���QHéqx�gرf-�߼)]��D��>�W�>y�$�A�y�,��o�#N��+K"�c�<��~�c�X�$
�)r�Ý�����_��/N ��#A������xl�r���k z�6v���7�2y!���j0gɓx������4���b�/�{7�#k�ѓN`��ex��������7y6���װu�G8�c��s�ֵ<�g���l�7��{V�8�y=v���B!���^�~�ۘ��*h�0L�������qd�F�9)`'������¢��!8h0���T���������JQ��Ì�K���5�����J1.�D��38��C�}u�t��9�c����T.0�p�d��G�OP8�G,
8�I�4m�P��:&�n�r���Qp�ѝ��n�q��X��z@y@�Њ�W��3���f����г܆��;]�8	��n�e��w�py|�*�>�ի��#aE�r�l�˿�#�iD�c�g1���ȇ�� +%4l$Pi�P�-�(<��R��Y�EAJ
.�D�GYz����[pv�:��9)
r�gS3}�]�,XD���"�b�T�=��iv��Who�(>ͳ�a��Ϣl�Xġ#�P�S6S�^�>��(wnI��`�`Y��C:�L�ȃ��#}�.؇s�6��y�!7�4�z�ȼ�����4����ا[pd�z8�^�".ԏ�iK��~�8�]�qtw���	ayL�(%)�g��s"�B7_��ڀ�fN`)2Y���ʉS�<sa3���ÕG���w���3 G9p�b;��m�Td���bpY98�_��J�O��"22#}fy�*y	drHI4�����͛���ݝ��77;��v�w���44���/I�#����T6��gDFD�}�ȔԼ�{w;��ͼ�Տ.$���E��|��S|.�)m2T)�@Q�C��J)�	!i�8�p���dP�i˄�Ҁ���P7�"�=:�:-�!�%��3;L;ď1��b�%���m�4e���w�e�4�c]j��U��2�/�Gi�5���Ae�^E�.ԫr�ϺC �lD]r �%��Kq���ɪ�NT2ͪl��WW�a��jyBϿ�h�J�g�"�������_<t�"�Gוc������ϸ^L�5�(E\���	�[��Ag�۲�2�������ypS�J�*j׈|���� ��J������b��=�.9���ߩ,8\??l��7�es3�]�_l)/)���q)���H�3-��9���Y��@U��5z�ϕX,���)��3�G'%SC?�es�,ˬ��垚G��|�s�O��z�v?7�gt7��\e�7�<��/���]���\���e�X��:��M���t�S�m�ߥ�/��@ۅ I�Oi���;r5o��F8�r�WZ�B��|�l�`/�����z�P�a�U7r"��@�
9:]���;�����8��Ǡ�s͒�.��m�mx�3���JJ�ʲ���Ŗ=Gjѧ{�W#5jYf�e�>gj�������u.5�V����MK��P*�\���x�.��,��ߛDw� �R�E	��ј�(_��jˁ�n���ܩJ*�����h"�D0��5j��3Hw&P�[*P�٨���AkU-��Q5y<�Ϝ����o�m��6���������(&�b�����ڎ�M�`�8-9uzCr<HR�TR���~�D��䀑8Dp�˔����q�Z~.d;�q�h��! �Y��r,1+{|zTD}>TGR��(��X�+F�oG��4�w�<*�}��o%;��0z��*������؄���b�Tjm5��xU��Φ�md��s#s��E��`�Vp"W��܏�w܍����(ņ�{Fn��1�:v�GG��Wܰ�~��+Q0s8�q��Qt9.�ڮ�,��[����_b���Dŋ =+4�g�y�Ѱ.���I&��X� ���E��Ob�gk��S�͡hy�c�S�h�-p�1���Ql��%�����:v�@I������;�b��xe2�����x�g�_m� �D�Y¸��q��3^��F��F����)ؼn�4y�a����\d3�@Е�B��>~�E�y�1���nƂ������&��~��܀מx��N odГĜ%��{��bI���"V4�}�>z�Ulx�$�z$0m���݃YW]5T�&��H�=�/V�����&�H����� �\q5��'Rb����lx�]�0i������;q�7 H���<wg�ػ~=��o�'��\A��p�5������G���,3{�<�S;�Di�*���H(����P;�`��J�$���FHB��rS`��8'�4����)@5͌4,�~8^zMC���c ]�P�>�è�&ٞf&VU#�"c��4[C.�G�/�/�F�Yt��Ȇk�5ћV#a����k��O~-9 :��Fu`���a֊�Q�jB�a���D�b��Ƨ$��p8X~W�S��03p���z�P���|��G�a��ʦ�^) �$�)�Pjiż[�Ą�V�[�,[��uQ�v���x�9��؇h}-F�]�KoZ�ȸ�Hs�`�Z@�)׆P((2"�|�I�4��!�ʬ\�9!�g����ۋ㛾��w_G��4�
��4��c0��%=}�cH�Ʀ��ÚמGȗ�/�A���/��Ps6�2rY�ta�<DTkрi.ښC5&�z�<�ѻ`n��M�d&�;�ί"s� �|�B@^�bČIX���4}�Ā�O"��'8ȭZ�_:�@l�~[�C�Uy��Reh�[@%�4���c��Bu&MB���0�|�� �?��D/�B�l^�8ͧ�mD;�.���,@�A����h�)1u�O�����
!ʭQ.��_���r)�.T.�M����],VdB^�^P��6I���ֽ���*����s�����y�!i9T~^$7��<�����+�.i�~߹�L��2R6 �H�B���y,�y}aSC<���Y{U��妠"����E�^`���J�#���f"�RIAb��8����!	Q�?��"Ŋ�<c�X0�7��o(	��2��.�u�[S��{e����7�)�`�`ӧ~]l���PS@\h��hk*58�2��jqP��h޸�(�R�r�5��/��5�� �=����&D��0�Ӣ��۶���L��sJ�ꈵ�u��uۣj�����W�w���������Jɣh%G"���'�`�_[����W5#	i��P�䂃}����7.���R�+��ro˾B-��ϑJ'�Ⱥ��d�C��_���E��]�J%۲��,�6O�.���Y~���x<��&�5�~��W�c�|����Tbb���S�ؚ(*ZJ���P�xr^�b�f�F����d[�yp�0�#I5b�q�!e�f.�!�I�q���bx��I�!	y�@._D:[@2M-%�oԞ���M��j���r��4F4u��`O�,ML�1�#��z`��,�6mr(@��Z@�u�0j�d*�>k.����-Ptaŀ��Yd{����u8�a-����=��`F�B�����y�(!Q4�b�P�P����n^��r�d��+b]+f<[��K4OB���"��=�i�Ő���Z�� �8�1�|��锤��LKp�lH/RŜ�T���`!'R��XJB?�l\J."�x7�XQf80У��ȣ3�A��Gʣ�@���N	��'*n��~���^��-t��tc�'����?�ǎã�௪â�7�{�/�]�c.�c<�i�~�8��C)�%)����_`�̙���τay4�g3���C61J�^�(�~Zc��ÞM���c�KZr*i@�T����y+�%�4���
d�ۯ��W^A���D���b�+q���a�8w����h���<�����۷�M�l
���c��+�h>A��'�<����q|��{R�4�������
��.�����B���<�5o��5o�	;��Uu���]�e�> R���U�lٌ7�r��L.���.��~�h9��x��i���X�������5���ӱ���q��WC�]]�a��ߋ��zo���=%driT55����l
Xlɺ@6�ןx��[�T_?Ä7�wލ�W�B����4A@�{p���?�5
=�������%���!�>R��Vi|p6��,�n�f���yTE�"�&��4/�f^�B��Ek8&MA�2!UEAS�pܦ ������)D-�FB��@G�a�3�D����N��>��5���ȱ��őql$R)���/�<fK��y�T4�D`@A*T��9�#,M� �žu���),�Εԏ�W^�9+o��8L��fYb"�9n�s$;Y����@Ӫ=hX)ds	rIi�I�Q� ��*誎��N���ly�yT�)D��K���ìU�c��U��#oR��AC��	l|�ql�M�>�HS�λ��X��E��Z����/d�������"��Y5�� �����a{���r9t�܁-�>��=;P���h ��`�T�u�\,X�m��1x��_���"��Ex#*���EMֳ    IDAT�5
�`�9qx͊ �����d��J.H�)o��8(=,C]2�4zOv���]�۵1'��*/Ld�6y����p�+:܉���p���O� �f�8Y)�$^�ɸEN��ph�$��q�@�d�E	)�_GB���Xz���ys1a��҈�Y�6}��P?|�du�^2=��߸s.B}c;,ŏ}^����!^+D`�fم���fW�/ŧ�&Yt����\��)�E���uiJ��וްq����6��T�92�da������J��2l��w�Mn��o��[1I��{.�|HS�c���UҶ\�?�E2=��3����e�M�4w�*qe���l��ey-��T���A��s�\%�#1�Ѭ�_�a�-e�)�&�ޡ����(����l
XÆ�[���D����~��D���u�r��Eܿ���:��d*K�|��V�����g��������YO�7o�0���}A���NV���_��wX3s<&o��:���_���8�j3����z�-��ƹ�#��q��^�q�W�;����m�c���t�_����%�y[��? �}8NX61�5�Q���(eȍ���* IF#����U�4��l�݌�xߑ��A��Ϩ㔆 �w��X���w��=i�q"�������o�>�-�0�bu�S(�d2�L�>��]���6Ǐ�%&�:y�g�L�2@x��EI�)f1/�Q6<���M�-O�\j��ۑ�8��틢���t�hT~�mfFp�MLu��~Hӹ,2��\^8��5�0"b�KB7r�2� �r��Q>d���5 �B6��D�%�b��è��૊^V������O����o �}���AQ�����>Ȅ�(�&H��Jb5�2�]�D��IIT*�&�e̪��<���eo&�k �~�b^�GSdC!J��T�K)��[�|gCP2L�I�w@T��C�J^Nb���ݔx����m�*f-7�tF��蔐�T�Mt�8]�b��0�W̘y9�0T����a٭������RL�}]ؾ�S�>pP����6\��f���ė fhNeȮ߱O?�[	�K�r�Jd1c�x���i��D���E����;�>|%����B2qg(��'ƍ���j~���Po?r��z�|�ݸ�;�H�cB�m[?X��_|�w��p� �\�7�u7��Mta��ێ4��op��>�~I:l�8|������w3(޲M:��G��?z�L�͑j���-&�]��9e�� �ۅ��{��&J���]��-Xt�J,��}���{DS���_����Q�!��5u��7����Ǥ)����1�ۉ�eb�3pϏ��̈́CO�#m�{z��/��g��Z2Q�M����<��E�@�+k�S���O⓷����NA��j���o��U7#�� � ��w&���7����o���AR$�E7���< T��v4W��ѳs�>�$�mY=7�U@��wu���_(!���j����������28�B��?xd+W������,0i?�O�Y�I2)�9��������#N�?SJ5�$ %���H�X6��k�� �!K�Z�U3�"|�
��M���h�_��_�f+�R�Y�܌K�_�R��@P��^����G�?'WDz()�Ȅ��@U�bBJ��L�Q$=b�W=�k��6A�g(��>|_<�$�Tjt>�<��f\��[�~�-�6�B�1����ő/���O=�C>E.q�P 3��3W�Dd���k���9}
��N#��@��0~�xDc1��p��$��љL�����	�h52%�L����6<��l݈:Ղϧb�SB`�0L�i%f^��H=2�O������7_EH��Tс��cpt ���!����g���M̶TMs�˭7�el�%����|*�u��eb+���ر�c��%�'�^O����Xz��}�*�z�0�f-?�jS=�i&l��j��I�=E�s�ؾp`FOC�R���?��t���ϝ�i�� �،W�~�D!��L����#�.�b��8\��Z̚���Vh~�bҹ��b59�$�_�_�Q��畆��_�qNݻ�p	WR�S+�UWtn
~�X�V�5箍n�Q�d�����J=s~c�J�*
�
X�����:� ����"�s�X�����Й�,��l�I���f��(����.+���d���"�蕤�pC�\v�+��������0TR����&ۗe?OY���5U��r^��}��1������σ���Q��#S�]��^[���T��w��|o��kb�.��m<<-c��_��k~����M�7��?��_�+p�Ķ��^�'���2v������&R&g���
�e��?ʇ�]�'Y��T��	�(JI��4�bp�'	����ޑ�\2�D!��H���Bs4%7����L���%-�c5�di�RC�"Q8���0b�eR�x���ƅ��� �ˠw�V���}���A��)xR4fѝ�dK`V�a��HۦL�TP�;��4XS�+Syو��8�vƷⶼ3���hy��W�nb$/ h�J6tJ~ŕ���E�g�70m1s����Ш�Bf?/HE�T@����Y6��K��{���Rpf��^�fg�i��f1�	�	)Ň�9˿�=,��.��]&�Y(�vb�������Gd5��������?�1"Qe�f��}�/<�8�8��Dǻq����/��f��y�f>���,Ñ8�x�'	ֹ���/��K���dؽy#~��~���=plj۰��{��v6Q���D�}��S�~�e���i\����+q�}��~�89�
zXN܇'�S޳v֔ ���.Ʒ�!.�{��}�3sȟ9���}���v��c���zS�/,���s8H��Ż/����6
��O�x3�Zv#n��~׷�7�ù�|��<�8��[)
��%�K�^�:B
P��*b��������{H%��-�1r�d����$CBa���NK��t�W_/<#�L��#�Ԅ��f]��W��Y�~�)|����p����qͪ57��T��,�o������S�2��c\q�R��Bij�I��r��ڳ�����܄�����U��g�r6�f���j����:��&x<��1�8�IaP|V
<�"j=%�D¨fnKI�/�Ͽ�9gri�XJ��Q����BLաs��㱠`�̢?������k�^4Ƃ���m�5�͜���U C�:N|����гo7J0���p�ʕ�}�M�5��2��*fp���vu��1�Oe�t�=--��~���ً\��%撄�1|�4�4�[0������ǡ�3́ǯ"0r,f��F/�v���{{U4m4�l؀��=�#֢��C���,Y.MA���P�QSI|�u��'��	&��c8��j.�c�Nt��f ZPkk+j���#�"�X8�e�>���ڌz�a"4��,���n��1��@O�__�ן�������a�сS�$��˯ļ����*yDFS��N	�E>s�"a��pbK�÷���|_�{�<�[�ٵê����h3�o�&]s+��������?�`�Ih�n:%0d����:��^k>���ȗ��W,"�7a����3y^�^��$b�̜�1��B�k������$�?�L�����(ym��4W^��f]�@�^�K��x<�d^='�$ĉ�����n���.~���YV.B�
[�W��2!/�p*�7g���Q�~��E��Jd�?��UD"�� �?άr5����9�罚�l�r�
Ѱ�-�ȗx]�u��6!�r0�L�0s���[ʯ[�[��S��『��e͚@U����šbA.*���r���t}��y_��A(/c.^��B��m�!ׅ9�
�\������i�|�܊�̞�g�ɦQ$�T��pq�&����DU�����7�q�P�@�l��VU��U��_�ɇ�u��zt�o���Û�������6l���(!Nd���8�+HR6N�y@�v^q���d�g����\�s��s3�n�Q���N9��I	ѓ��L�?5��<Ӄ0��X�nxٸ�V������.�>��� ċ%(�h�4MW�ưYSQ7v�`t�F����K TU�Q�����d�0�A��]ص�S�<$��!�Aʣ!����O0�7��"�5��D��DA� t�hh�+'R�ɡ�3��$O\�_��,����[��q��t�yR��y�E�,xK��_�y�lS�$�1�-���i�Ǖ���8E��B�I��Qbr�WC1�Gg&���4N���md<is$�*�����q�m�Ɗ�������R�=Ѝ-k���'���c'��a6��U�����/��D䶥�ܲ�<��<�����R�슫����h�T����d0�H
����PSB6��� ���U�hƭ�Z*�N`��/�O?�)z�t%/�5���ƛ��o�_���d�'v���
�nَ\*�R1��kq�}�c���݉�G��3��≇�{�n��'�ȃc'��{��i��ϴ����'����?�u�|����������	�-Zіr%s����{/?��x��[A$^���o�m�����e��m�8�u^~�ع���K.��߹c&M�n�3�����᝗�æ��G>=��Y@�����a�5�A�݉�e!�ݍ��x���I�<Q�Xu׷q��P�l�(��#�}���ͷ��>+�G���}�m�"���"��a�Ж-x���@��#��6�ì+��D72,Zdf�w�.|��8�}|�4�Ŝ4�n�WH2LQfs�/٨�jh�P�P���;�i�)����0!��|�!Z�nS����Q�����8�ϣ�fW��)j5�U�O������ʡ/�G� 1��>?Z�Q�uU���@�i��|��]�3;v���[�ھ���R��n��[oE�mLI���_n�\6cm-�p��`�5�E3�;pg�OASK���@H��	�wXS"6����S�C��aDhc�0z����:%=$�[�|B^��mú'~���+Ӄxc�/�so��'��*�:q'��A4	(���H�E�l�Μ��m8�A	Iu"?�ղ-�w'�88��F|���з{��l�@���YqF-��E�J�`;W����\����jh�U8��"�҆+/���WIhU�ñx�o|�yƕ��	�Y��"^�;7�*r}il|�}|����w`7���Q���тi�,��ew �)��ظ_��q(G��<-[�4�̺Wҹ%��T�:t�d�KȲ)0J��M�ul
H ��������~����!�l��D��!C�����M��+����`2ρ�5�p	,c�i��/|�dߗ)><?pP	K�Fh�;�r�[���S������]�lnlŜ���=�gȟ��W�|S�Q�0>��{�����9�x.�-U���ey���2�FdQ��Z�����8�N�@&��l�|>�zX��������� M�H�(M�ٺ�^����'�Ht�1�C�!&^�?}}�IY���v�%��j��Ԋx8"��F����|���yN��u�̰!��oR0?TQ<@�h9,�d�Ѯbz/�����B]�=�#��_��~�D��O5��'�ПJ�[���Ç��ݵ��-w��%W8�A,C��ڀ.E<?(�@[t��������Y0�<�ZLoe:.����(�l��4%����PJ��S����l#����j�1i�ht�5������8uJ!#�j' ��i���xƭ��)�c =�wb��>�>��GOJ�8z�,w�� W�ǎ`��`��-0�r%H����^/��%���tMGH���&�����i�p3��U]���g�<��J��P(�\@e�"'WR$'B���n�7D��FA
$��:nK�3��+�'9��<~���P�EWnŉ0�'2�i�"��5 :�N�28�N�t6+ȼ�c!M�:U~����+o��y�%��̓�=؃}�W�yG���y1�k�����0�UR�I����g���_�=�ޏT:��Y¼E������4k��rb����}��DJ����d���=(���a�%��!����z�&����������ے�<o��q���>~?M��y�'�^��� KA��c�8���=�b�uPc�2���٣�������B�U����q�}����ka���<��=�(��	SI����h��G�%�V����Ź:6�Oc�����Cf`@�ؾp�-�
w>� �Ǐ��cd;�o����cطcrF9�ĘKf���>�K/[ ͘4�E��GE�n�;H���X�jn���܋��n����=Y�62ݝ������#��a��\���K����EӨ�n�WF�>�,�{�E��>#J���_r=n}��L���/W�F6}�G~�K�=|\�P$�\4}
n��>L�;��b�T��ػ���4o]-5��C=/Ԝ�J�̠%"���5E��:��e�?�}E���3��Z�\� ڢ!����<��,-��B	�����iGu^õ �U/t��R���2�ڰ�����P�q�<%W���t����w�~���}����q��d�뭍c�%��;��bɂe���uo��
�[Z0c���6 ^���Q���EfĤ�5C1z�s�Dۨ	GsT�b>z�wH;�����)�x�XD�Մ�)B�`"�`��}�������7PLu#�P����o��0�Ka���Ҹutt���R9�s3j}�:X����B+������0��^��������[6�-���	�u&,���T?0�Ł�?���G��t8� ̀�� ���,���3��1<M��P�Ĩ�B�&�Ʌ1���!L�Ո$UTt9��W���o���#���u՘|ŕ�}۽��41���;����0�{+�d�h��4J��yU
P�"N���d�sLL�a:����)P�h<F̙'^��v```@� /s
D�����ZL�:	Sg\���aH�J8�?��)��FS =�4�)�������?W���,�|���M�bH.g4UL���9�yĨ[ԻyD��V��3�}	��q�I�MѕZY������r�Lnx�����{�[��pc�y�$6�_�ݻw����(7Ե<)��ϻT��<�5WFU��BT1��;���%:D���J_Ÿ�J���P��{ݚ��Ś�^*n���x��!�j�c�0�H,&���Z��Q��󨪮�E'����t�l���X6���I��z�����'�!��ءh���j~�����VM�/~���k����~�c˶{l@��C�F�榀HMI��H��
6/�n���Ws�]>J8���]�5\�P��T���!���a�[����bAA��v���a�x���^<��#�TqxP˦@�q�x�Xz-�W_�{6c��p���XYzȽ���D㨋0b�T�8���/��C��I��s<0�:�>�ɥ�9��uo�Bu(�(IM�_��>M#��"��1>�rve"s!Q��Vf�̓�2�O��`j˹�r�&�a��`Ć�I�4{�tfE�l�QÍ�O
&� M��k�m%!]c����܄Ȓ���'_�YG��͢�:�y�b�E(�����in}�A��E�+��@)ч�ｃg���/�{S�`��)�����3ϣ�K�}�L�|�鬉�	̸|>~�W�3�X�''Sq�PN>��w�	N{G��BUM&L�XN�*Gێ	{�,vn\�g~�:O�B"�)�%��w~�CL�s�g�Zd���1^}�9�޴�%dr����;���l�s�����G��~��k׊���V0����.V}��.C�[�b��w���Ƶk����J���+�mBnr5�C]�X�ʋx�����1Kp4?&J�� f.�o�!jd��j�z����8�{73�T�������n,�j	����m���>�������1���y    IDAT4�+�{Ѻ:\�-Xy�=��s}!E��n��³x���>I-��{�ո���øK����L9^�|�9�<p�|A��s]#��	�f��S���<�G�������>n4n��6,\r=���1�����/<��[7KB�Lxi2,�U.�H�a���Nc[�:��!�=.�>�i�MtR\�sS�+�U��5B�_�����#i@���|i�#m�� F�#��dS��rA��<� :@ſf3Hmf��h��Z��fw�c��OB���H&kH<�M�{
��}#�`S=�,[��܆Ј1R�:���~MM��0f��e;=����$��&�-I97���`6���C�?��۶���C���F+IHW�%Ӱ�G?�r1	_�T]&�~���'�٣�Ŏނ1xz<������D��)8�Ӊ���Iq4j�tt��_�f�b�^�Y&�IQ����GU��ٕ���Ԗ�x�~%��l
�joƂ���I�W �*� )x^��ð�z���X FPCW*��Q#p�q)�K��͛n����,��\X��	EFw'�^�'x�%WЃ��x����W����6��F�:��sfc���FM�h�聽m�?�:�ڌb�ހ�4�|��P��b�Hz3,�&��]�a�$82���{�0k&�\{-�H^x��<v����N�����[1|�(��0�-(:�l��sr��,�� +KlJn�wI6��܀2��
��Rt_�ȵB�@���h;�o%a�|��6�+V���iإ=������ƅ9QeD��2�?������M��ۄp+�cpp۷n�[o����g�R"���R}��Xq&��2��L��[&�
h���0�A��,!�eہЁx�����3�#�+�4�=*[8��i��h0� �vv�f �K}�-A$E{�4�4K�Ϣ~0�D4V��ӧc��q��8�H�T�	�l�r�����ly�A�J�/d�5��U��O�q��o�H��?c�O�n��gx�p0�h4�? zmN��������+���<7���.�ƬSr�v�ԋ��C�.�d((�s�g\�)8!�W6Uz -Uq��VC�&��<��,�*��-1�GM���9���0�G�����z��n؃&���d��R4�@S���Q�>�O���{��?��� _ґ�x��)�s��O���
�Q�JS�|�<��|�t�R\߅���ӟ�!7��_2�(# A�ruw�E��ގ[na��d��>�n�N�LN��[$��)��"|]�9 �bT�(�x9�s�3k�-���x���F�'o�3�G_�@_!�4),xC~Y��[�7�}�̺L�*�a�GᩇƁ}�%��ĝ�ѣ�����s�|7P��?����k��z��D��L�&Ϛ�;�3�͆Gs#�5Uñ�G�}�n�KFb>$��08�B{�(̘9[�&�X� '��΍_�?<���n�8�-a���R4O�5KH.����,�~�o��
��>Ջ��,���x�*,^~Z�d�s8u�0��)l�bb��KuP=�f�r��������)�8�>t/>�$�m� SGӑ6-,�y�������(پ���P����ɕ�M���&�[o��+.G8���Ǳm�:|����<z�ͭ��R(���.��W/A���n�m�聽�d��سar�$���UUc�«p�ʛQ��"��b���c����g�E.�v�u>f^� ׭��ǎ��$<M|�����w�)��K�瘩ӱh�
�0�@@X�*�жx�'q��qi�x�4�l��%��ʥ��k�s�b�8s`ֽ�
N�ف��G��{恰Q!�ӱ�g��4�@\u��Wф�!9̋ޢ�������/�����xU�&~6>|��r�o��<J������Uh�4��0�7�w�,�TR<F� "�ޣ�.�G(@��_��҈1�3�l�X@�"s�0v<�6���!�Z�E>4��[�9V<#D&}`7֮�UUUhkiG]}#������P�L�g��{]0��݃��Q�a`�6���_��뽈s��Z��2��#�f.��%�_��ч�}���3��"I�K��ī���{�Cd��8p���-8���F�l���6�%/�"�y�Ux�W�XE���4O{ �o��\m�гm+^}�!��s4�ș� �ކɋa�-��M"�K|}�W�/�[%��?�!�R_m�Ξ��c��׋���Ttv�3P&�˩X�ob�6�QpHEI�kUqv�Q���KX��0��1�1���"�14��k���m��S��b���2g�"���I�oނ߰P�U��#��P�EZpqW)0-Gr4r:��i��q	.[v���x������=F4غ+�����M�-5v�ZG�����D��I]��B�)�Wʬ�����_���oT1���\�=�d��1�#y��c)ډ�P5��^�rNӅMAl txJ��F���ω��[6�$�M���,r	<��S�����3X����������W��d�y��8�q�%������-�+9Rl:y�|�܌�9\��������y���MBu�
u5�J&�J���C,�#�"�:E�ͷj!R���E%�$	���Q�Tr�%d���^[Ӏ�v��ILr8%K7ߠ��	��C]�Z%D�n#U?����OF�[5���G�h޼?���/�N��c�ƪ��"�Ͳ̇����G�82�(�H�JÖi��(r�&�AN�����&w�^��LR��8	� �zV5��G�f�T����C�Ռ�W=R��b���1����E��˰#�g��t�:,�����~�M��.�8���bH:
�:�	�Ez���C�Â��k>�1�R	�Y���4�D�tב�`p�J2�5��R�*_s�D����k����� JR�)�E�Hc�����n(e:n�'�16����@�c�� ̐P$h���nS�5ЕΡ'�G�X��	�a|>t�1~�,\v�O���;��)�ݲo<�<��	K�4���݃	�'��!�#�Ƒm���K/����Ȓ©��2{,�c&�����YZ�$����cB;)S���@#G��es.GuM6�%���׼�>�}L%Ѷ�}.Y��_�XU�e3�ط�+�_�����P�D]c#�/Z���C��
9!d�y�֭]�][v �s7b�χqS����+�G��؆u�3���;oc��Jeʜ-�0��y�sՕh=^?�AJ�=s
;7|�����l,݋�1�0w�՘x�T���*�L���������:!2��f.\�i3桙�8��O�'�`ח�qr�N$�0, a̤)���Ũnh��i��$L���A|��{H��#�-��1yƥ�t��ok��� /��%�c��M8y�x���-��2w.�F�7�p>�ha��l�|�܃�p�k��ęӱp���	��1�F��v~�z}�����.�Ʌ_V�%�٭��mG>��~�45>��o�g�<��R ��V�1L4��cQ�C�3��M�����L=7ci
�~�
�Q��Dr�-��j0��bV�I��W6u���H �(�:�`
���r�r`�$i����`�Ob���,dlj��%�0g�*h4�r �1�i�����N� 7շ���	��8�0�����>&y�p,�y�FÈ�6��9>���ȝ<�@фY2P;y$�~�Ͽ%="y"<G�$�8���x���p|��k��z�R\s�w�2	O���;����T���	-������	R�'�H��n�
)نYż�
�� �PX�i'���~
gw�D5����6�\�����kb�8�n#6��N���SP�B-U��ŉD,�����aޕW#���4��BT�ya�I�I<*�R*,��(�$:�d	4Tp��c�������wa����.���8��0�͍X���P�1��c���'�ٴAHГ@�ǝ@tĠ�Js��`��C�,L�BҳCi������T�'O��e7 �:���&�o�����
SW`���VG��҈���u�BM}JJ�'"�11��~�-D�S��yO.�e�H�x�0kI
�2r�R�+���Dx6��@�\h�}U𙮬�Fd�n��6����T&����|w٪�P�ԕ�|o%�����.`7���%>H�� V����>��ܹ!��R��u3|�����Ŕ���h��M��9� ��g~���ϒ"p
� ��hm�P�u���(2ț���V���5q��բ!��_��yL�v��ֆ�)�hX+(���`0"Cbz��#j:���F�q}L)w�|?HxR_1���!T�s���D���O���)%���;Y�d���>_�X:�	D<q���!׈'�{��O�����.\[kh�;��,%�RP�.��)p��_�Ο�O�A>�А� sw�>!���bV�bz�B�j<�J�Mn��|�*�9;�"L�'�ES�,�z9��׃bȏ~�B��+W@V�
� �	b^����$�3�09y���8#z@Vz~��U&�.{�M��W,Ǥ�0ᘦ$%�l졩�|�B�
d�3��"�C5Ү��89�b��-Ǔ&�����&QE^KUj����U�
PS,"b�n��M����撅e²eSЕ�`�0`�>�����4'=h3���Èɓ��J�r%�����p��1����F��U7�}�("<�)(1���q|�ɧ�$����3�����mBf`C*	妍�3g184����ٳ������1k�|D��6a��lR��[?_��γ����"�Ҏ�\���& \�0>�zN�Ğ�۰�.d32�W�`��9�6g6�����sbP��M��s�6��W� �u`֕W����HH<&4�o��3|��.���I@޶qѴ)�r�eh9��y��������سmN�/t9N��F�´ٳ1j�Db�"A	s�<|T4�g�Er�O>k�bSf���Y����&Q4@���چ�_mE�N���D1l�8̽jj[�ɴ�.0RIu�ƆO֠�����	hw�TL�3m��Hc��W@)����j��%���E�vL�t&�ƏGU]�|>�\V*�3��`��w04�/R��*�h,,^"fQ�XK���8�q=���g��%��,)�5��?>8���&���@��=fA��D� �S&ה��#����M��!}(]��tV��D��X����D_��0�#����trț(�Z�h	�$� �P�y�󆑩�Èn .�,ԏ�#���Gqp�FI��Tc�u�1s�2��Ð�x��}�woC�1��ڂ�a#���ʡI"Ԕ;��#�_���@��k�!ʸ�������8��:Ċ<Z��kq��w�u�5@ ��s�a ��y�}w5>z��8�Kd*m�/Ŵk�Et�h��:�cݧ��AC�0��q4׶��DKh��OM�JP���Y���8zgϞ9jKC��A�H�������ECPC6���c�����?���'��7�ӗ_Ñ�;��3�0�@�!�����WL��&N�Ϝ?�Qd^�&�)6�B�a���3�;I��M�<z,g��}�]_|�R6���8��!��ě�e�9�Y�����H�ރ�HI;���~���:
⎆jMGMPG�ÜT�ty�Saȭ��°�)(��#�TEp�(\z��9�~[�X�Hԏ@D�Ԑ�y௉����m��`�k�Ѣ����((6�2��2�]ҝ�J}#t쏒�.���/p�i�Ԟ半L��3��(kg���P�#�r� 6'��5WBT	I��y+��6.�C<��>CDQ�')�J�*`p��S�Ű!�J�����e�E|�o?V��֬Y�\:sA#Cj�{ͥwJ�dw� \�浜�B�"o��I<���#w���TGJz1]��_��3��hh���Q�!^ۃ��8jjb��ECh���m �Y�Hu5U�]#���Kum�kf&^:���'k���FQ4]OӶ$�T�'{+����%A��Ԑ�
O1����p���������?�G}4��G���ݻ�_���k5 (�>�HD&��A��A�n����Z�W I�nroe�&�s�wr���b���=Wlv>p�<NSrY�pH#-��brl
L��PǦ���$�_$7�vѣ@+�����i�բjG/!^9��Hx���T��a�#����	��f����)/��8 ��wN*%�r�=)��$�>�p��_�Q�2���N+��,�q)��?��NM9A1��Ϗ1
*_bN�ܜ�j=��PL����/$�� ����W�����,�� U4ez��PSudm=�<�Ǝ��ys0��)B-�I�iÉ�N���ClY��]��D��d�JL�;Oh&ő�{~�G�����Ñ�'ŋ>f�,�v	F�/�(�p'?�p����Pl��y�u&D0f�$4oq9>o	v.�B>x�ܽ�=iXUmXp�b��4գRH�Cر~=6~�1N=?Ku5��`�lj�]�M��ؿk;V��:��E��D�q/���/E�hh�Ļ�R��������c��m0�y�*4���W\��Ӧ���z��(���ؼ~6���A7�u�HL�6�f�A��v��!�;�v�['2����dʤ�AL��R�\xFO���7N~�N���*���h�!?:&NƵ7݄�Qcŀ�l:{���.vm݊>����1&��kcܤ��̇�4~�S�عy#6�������Em[+&^r).�7��-��(�Ld�)����ۯ<��{w�۬`���㚛nB��IB/�5j����vb��a`�.�Y��L�%���\�� G�Z!6�^ZB�@���y�M�Hg`�d�m���XU�����VP
��Cӕ�"aY�9x���Q�	���;ӑJE�2dr(�覅�hm�Ո�C�i�V}�{�%Wy��>�v�+Wuέn�$��M0�0c{��zҝ{���s׌��9�x|���A �BI-uP��J;V���_m����ϻ��V/���U�v��}��O��k@v��ל+>��7��W���*ӓ�k�Gnvږ.FâE��(��F�}�.tϝ�%+W��g�xFĄ_�@PV�f� K��tl+��]8�i�<�1v�š�� 85��������k�u�
��\�Tg���)��"šM[�o�;=yU�}e�h�;F[3�M���}���ѽdR�f$�DI��'�X[r��wm�����������"<��;F9��o���#����hNU��,�5t.\�5W^��ˁ����wbǛ1rrP��t�����E�)�uF�==��9U�RQ�S�4WEe��RBFY����%�K���:(��ɇG����0y��9�mR�q:� �Yz���mv��;Q<|)�@�`�TD%���d��שs��e1��D١�ŇgF�7��hѮv�{�hX��m|��
Vf&�4�$L�͘=���k�ޤN�z4&��~f��t���Ws�Ľ�@����8�\k�?X�׺�Q�Z�i��-��a�+,���R�K�֧l2�Q�k4,ҥiV|�&��a��1I�.-@U�p�Բ	����GdO5�� _��DāpÆx�����W�;�����E����<��H�Z���3�]F��zj �L�"�3�u.�����Vtv��b�^�"��#WǞ�e���Ӥ��G:i!�ʠ�.#tR��Xu�-0,LVQ*L�X�F�\r&��J+�Ai��k`��LG>=n�L԰�t�៚�?��������'�����<�?�q�C���#��Y�j-rZ�4n�t��H�6�%MBn������_�+�ɳ�o^.b��
\��N�]�z���=(�Q)�b]i��Cڀ�!�0JE��
R�"d�[7P�G�⎅5��Ib!/l���}g�p@�<H���e`��# ���Q4c�6-L����ٮ8QU��)0&}��S9m�s Ԇ#+�c�^�x ��B�Pm)���8 WZ�x
p���4X� C������\G�35W���&Vb�CQ���MX&Әa��x�wK�U\�N    IDATvAu�bILG��j�S��1�F�����$e�������D��8���p�����@3Hq21=:��/���~Z�x(����/��/� ��Es<����xO?��l�"?;g�l���2,[���sT���Ӷ����6�Œ�؁�=5%��E+�A��`Zz��~��WO`�K����)���u��⫮���݈��nxz ARn����>�(�~�S:@�����J\s�-�1g��L3��/Lc����c���Cl���E����۾��˖I�O�C&=ٷ/>�$�z�e�ƑH��>k>�\r)ο��1k&"&��}�������c���^���,]��_=��.��B"f (������>�ûvK��;��:W�x3����DB,�RG?��}ooxUL�2�:�ϙ�+o���[# ��t:*���/�$�'$v͜�+o�2V�4�wI�-�t��1l{�M�������wa&�h����%K�/^��� �����S���<�˟a���Q�;Ȥ����vqZ�,t�D��0�� �<���� XK+ŭ	'j�}��e��Гɢ�M�@Y�0R���tN�B@�,�E%t�%��i�m+Q�Ҝ(9(�1\*���{�hܕH�1�D�9$�(
�@&��\�%ZQ�K�ڛ�H[�Z*�JV�T��V9����`����L�E�Ɉ�jsz�[��y0>�Ǿ�G�={&�8�3K�Ê��1v��JXc���9�i��[�==�S�a��qb�.�N���2`�"���QI�a5�#����^�
e _D��c�2��vl�.��J"�3���[ѹx1����X�	U�-N)#�B�S��W"B%�W���P�q���>�ޖ.D������o�F��h���ʆ�d�d�X���p�EL�w\�;�*�N��X?��9Kڰꂥhmo�BJ:�0��b���U��$�ո��"��\	���D�U�>�9��7���!s�[јm��p��A3s��Q�'&���P�DQ�T�0I�f�@�7��Q�5����L�U�ζ=&����nV1nV��4�k��֥���-�����+�e���L)z&����$<2CP�ɪI�iQ*�n�j������iǺBGW���\��zX�_��Z�p����x�d��CP�s,ͬ��V������5����0>AA���,�3u	�x�	
:�;M;-~��A��U�Y�xJ�j/�����ej�||��Gغu+�;���I�lVHa��@pZ' �S�PNMN;�(�QB��}Z�Psn
���Q��:�H�,�w������u�J���,�i/j%$b:2�8��9�{���YqD��є �WB�0�|~u����w�2��iK�5�2Q�i��Km��Q�V�Ne�~��V�sMk��|v��g�̏�{o���>�;vl�]ףm�t��-	x���H��ě/Ӳ��H8�����_�	�3XƓ�3�� r�^�AD��ϲ�s��}d�� ��x��N j�=���Ŀ�Br��Pd`ה���LEt��	�QL&�]�Cy�S/ו��k�E!AǍ��vc�z9.o|Y����^�M)�#����N���瓞æ	�T�J%�S�a(�t!��+K�9�]TI�~\�$؄�C>�G}�Bw:�.�Ds�G�WF}ՃY.@�*�B���� �v#�؈??�^Dl�Ɗ6��4�����
뮺
�Ӡ�0>�W�{��8�����ݍkn�
n�����Ӎ$���&�>ٵ���K�����p�9�k.��^u,]�\C���M�����o�H��G;��#}�kj�EW\�x}z4�� ?؏מ|��s?�~r
054���U7ތ[o�3{��4nv�`�W����ͯ�-�K���pn�ӻ0w��	�E�Tā=�����bë��Xp`�I,\�����a���i�C��F N;��?�4�y�1�9"���Xw����0g�Bx�n\qr\(O���'8v� ܲ/����/��?�z/��]��P��������g���f��R)�;kn��Xs�%����R)0t�(�|�!<��R�����m�<\{�mX{�eH74�=�VQ�O=��|'N��!'�~훸��k��9C]��䧱s�;x��G�Ꮿ
?���KW��[��,Z�Q3!n:�Ǐ��16<�
��hh�`��gㆯ}g]��Vx����x?^y�ly�)D�0*%D��`(���`@JzR:f�rh��B�+F�
NLb�./nU����\���$�k�$R8I�R,H
2�X��и3�D��@��=E>p0�8�x�r|Nq���Bs]�T��x
���Sv8����<4�a�D]U:�ţ��6c�eW`�%���i���r.[�;�m�4)�h��x��j�XQ��3Eqi�g�+�f#d|G�ߊ^}Z~J�}A�A�w0m�P�T�Ǔ�FM��'QޔL!mŤ�R�˘rlD�)�Y�W��x�C������$���<��h���-��7���T̉�L���05��hh`�@G^وM�<��C���S?�JV����ciZF4!�l�H��II�}jjG��bԶѻ �.Y�����B�JkU q"-�n��|�$U,��Hڋ���pp�~l}s+���lBS�Y3��|m��Q���]"2TY��&��*���#���t0Ivz:/�6������(D�iKC��K/�]�û�?��ϡRu`d�p�&�T\@�l�d��SK%���K�)�	$�	��K��8�.~��[6�T^y�|����Ы�T�܄�F�{�
���9(�J1��0���9e�iI�M�C��p�~F[�yZ�,l�O�����O@�B"���`�F�XZO2I@Usi��&
�C7@������R�P�����N©�4�j���@҆���%���b^����N̄E곯&ٺ�ܛtbG�r�x�VE��l�.lR��`H֫�^W�i�[�;�Q�ЅH4.�'�~5:��/"�V�R�9J��zΌ9�d�G�V�ϴ�����3-�?�'���c�o}��O�� �i��$k���)�V�#(7wTu���˿C�R����7�ܠ ��Cr�R$�.�x��Bk��'W���;5�\ �6��24σ�UQǴW u�H��F4$����XD�����GA��K���D�z�HU�]�P��	]C�֑Fy�B��1�E_�QJxy�IA��4�
�g��l�#e�Ӂ*5�:D�����+ѧ����,7��I
�.vy�|�'�rɐ��6����J��W�Q�=�����.��р�D4&���d�kŐ�Ȕ��P��?w5�D^���cǴ�a�$��=�r\�eZ}#����շ�"\p=���,#oz�����c�.�h���W��n��7���-�"��`��A�������q�o��$.��:��կc٪��%jR��P�����ƧF01<����KV��/]�X=��.� L���6���O8��(|MCˬ9��O���7ߌ��vT(@���عy~}�x�����I6����]�=�[�q�k�06�G|���q�"f��h�2���V�&���J�=1�w6����ܲ�a`ּ�����p�M7�{�\x� :���6��؅�����m�l�]�E���+��!Z��E<���`Et|���x��e�19>�h,&�����Rh	w|}6܉1�ƯzG���Սy����_���]�h��pZ�j@a
￹w��gعs'4���ŋq�w��u�_�XC�L��#9'w���=��O�V���Y=���+p��܅&^SS�����Sb��	����:ڱr�j\w�W�h�y��9٬t�
L����������N"��51�Wg��'4��Y��ↁ��a�M�a�u0U��@�0 �^����N5|"!��D���r��!�h�Y
rјpIߟ�(Fvp�N ��P`�9�B}.%�fŌ�hDqp|��-N�
�؅���,L���ގs��k�x%3��k�>ؾ���64t�	G�jP�(

�锢��uE�X�ǵsl���mێ]o��Hai:iU�o"}R(�ʯ �+2�%�"�̥3�6��Lw��E���msfAkmB����΅��"��Ď�Z��:"_Qx�&�)�Taz��#�T�@���6�yCľ��A�d�-I=��2�DX%(�����T�.t�*y������&�>o1f��TbbN7+l^)
��"��t `����(��DLDi2aWpp�~lym3FN1�%��dI��sp\t���֣ȸ.̂��\<�	P�C�8��e���EŮ��G���Ls�T�\P�Y�E���]��Uc��=���s���\NL1�D�l�=��57#]�(�-�[FԔ��{1��|�R؊�X��#t�ڦB�-�1�_�5��d���Y�kD\�(�:���E|
�]�BA
���{���{eH/
��a�_M�0P�긕}w:Bp# ��_�$P�E���x�p�$���ǓJ�N��!
v�yNx{��H��.��f]��Q�|C��!�:L��c�JjN�x�rQ9�RA
yfesi�r��{҉�<x���)KGkS1�G����k���T�X�s��1k��Y��u�}�hk�@�Q�<P���#����D�v"����x��?�mM��?��Mϧ�~왿߲�oG�X\�Y�M���?j���&��3�G��m�Y.���f��
��m�2��a
p���&�I���
$�4��L
rY�����!Q	e�/��5�Bq(�̂�\b7+��ɘ��p��a�ɒ��R(���9��.�	��<�ؖE�HqpR.��f���&�(
�b�(����jqϙ!���UK;��!h`w�7�L
؁���Wʮ��I_��%�ܴ[�cqC�Nǐ.�.��X��e���%0U�b�p��@A��+Ҡ�#���.��_���b��W�բ��(P�O������3���;(�\�vw���q�m��L�2φVq�����o}�\�C�N�{µ7߂;��]�<o�t��\��4�=�-�n��}0qj�DW}�&���B��8�
���ǡv��??��m��w4���;?�n��6$�3*!X67�܃'x�?��tf�.��z|�?���K�/MP)*��$~������p�p,3�������?a��+M%rc��D'p����^�(@u�9+q�-���k�A��n����Bt�8����_��^�o�(lǅW_�?��D��] �hG�*���O=�06���81 "��/�w|�O����I�"Hv��$^\���^�B�SH��||����L@6���|�%�p7�������$�/^�����c�eW ��tZ#��o����܇'��\��-����~��a���H&�0>�����>�?��3�q��5����a޹��'t���lz�q<������O���pS�Pd���d�����J$�a%�0u�iOD|��(S�]����aV6�@�iBgL[*���#�;A��:��>�(�7cHD5�+N6�\S;���8)h�� ����S�$U�h~'�'��]���f�B�|]�p�E��M����g
�J���ތ��=h��@<��
����4Uʋ��.�V�)��q����qr�N8'��M�!�:�#�'����*���U�
�m�\W�9��h�t#fq���[�s�x%���=�A2J�Ѫ8�0̋x5�Xf���.�112���!L��ġØ>ڏ����a��(� Z)2���oK�B���-���B��9H6fQ�وqwv���E���m����*A��˔-dE����	ŮZ�r�&�ө�{��+o��'f6hJf�愊M�|	=�4z8A�V�p����ᾢ��}��3��E��
�:�yp���V�t�����ܮE+;����/A��_�����ݍ/ @	F]츉 ��I��wf�"U� �$+�KNK7�tE@���һ�?���$[:�U�]��z�ɩ�#k�NZجc�/�y��)9C|+�A��(�([���jeQ��h?���z�>���k��� Ŀ/�Ϥ脏�k;,�C���W^C��/ҝ;���^;���{�Ӄp��2�NNO H�cS�6e�}�pR�ߑ:�'4j���G�=��Z��!Y��X�\�76!YW���4�ߏ�v�z5A�i��x�:.,�NՉ.�)��~NX	̚��l\��ί8*�@�:_���YѓI;���d��:r��iͅ�'�yi���?����s˖�~�Ն��d{�rã���8�8��z������$,S�u϶��O�Lqj^� �T�N�J-�����U���t$��\� �"Es@v�䖁���n�Ǩ��eA���k�#�D,�a���ec������$��8����dcb.;1!}��iY2���mMh̅������mͲ-��9��С�HHU
E5�U2n��v�$��������gw��V��h�Zb��!p��KhD).��G� :�=C��a�@��B���k�,:g��w����^4J�{j
���H@��?��B�Cg�������ƛDDMv�H,�¯zO��I:�' ��w}�ϰ|�*q��"�訖��m�V<��3�0F�(�:{�~]
K3˂��W���O�#�ܾ�y��m������u��� P��*�|| O>�+<|�E�ˮ���߾��g-�_q�CFP�OO��_?��{���aFpޚ��7�����B4͐1���xp��?�;߄��8묳q�J��������&z&�O����o��2�^��=X���p�_� ���`��}x�����/bd����B|�����W_-��ݙ�����#�݇��1:)>���_���J��T��L��8
���?��w6I�sּ���w���褓N+/oρ���۽W�c����MeƜ�����p�WoE��E΃_��<`O�����{��бh'��U�ʝ_ǲ��CO&��;�����\�_�s��� eZ��C�{�hÇ*ڢ:�)�6LdhD0Uqqh�&��Q�+h�(P��B��fВIP0��4�"L�A�Ew2��x#!\����H`�`ʭ��V��b
���Z4������$NLM����x^�J7Q<͡�L�O"�18Y�Q�ىs֭ż�"�ބD6+�e6�c��%��͒{�#.�O���'�����-��r��6Q,H6I<f��6�چҁ��)��&�q��}%j��K%�a�%������µ_@��	K�EٞP@g7��Ta��3��(LL�X���� �|����wj�����àX�!�T��<7tY!��@��7�`/0G"n"ޘBɰ�D0{iں[dR�{X4$�.#A���J�ҤM��2�&R�EA���������_ǩ��4��,��I��R����a&�bZ�P��Wd�n2'��/�&����S������}�?G�6�F��$� O�ԁ��@����Νxw��4�\F4N"�h6�@Aw�M-b�j�S�t�&�Қz_��@�đ��� ;�qE��\���YA�4ꦔF��'�a!v����|J�Q�`s�&*�@ B�p�}�.��j${)��5�A�m?s*qf����J4�}R��ܫd'T�Qj�}�5=�Y��ul20�=��4����s�F��.�����x��aV�����O�CN�	�Y'�qx]�B����'s�.�\,��Y�3Y��r����DqrZ��X[)�*9 ���i@`eJ�%�;{ҹn�OO6���9�9A��!��֬ȫ�t'���}S5�Ӈ>ۊ�?����/�pݞ��Y(�m�|�A���s+촚�f��C~�����1�H��I�!�z��ʄI��47��	��ٶxp3��9,&;��T�
����
�U��	�9$�@Y���@�[Y���B`�Q�a`�*>��+�Ё�n�K��&(BèS�T�$�[�1��:A� �)��) ��eʔ@�C���N���{$�Vg*�.Ȝ �B�}�L�� ��+\Ie$_�-\e~�A�	$�S@�CZ ��ZJ    IDAT��8&���`��&Zu�����r)<+�)MG����`����Qy\t8�ЅaR�*���\y�*rQ�(*�9)����׻���-�O���;�ÿ��_�V�DU+"j�S�c� ���(�~�Y�>�u7w}�;Xy�y@��H�,v��^��+x��Gqd�Xz�=�q�_�eW^%�CA�U�"���.~��~��>�/�x}=��p��u���@% ���K��?��>�)H�~ɵW�[�],X�H��~�39��| � J@��?�=zB,얯X�������B豸Jy�5��|�����}�`�{��5?cF/n��-����:w�Xs���x8q���?�l~�MS�t�c��������Kʆ��>��v�����Wl|�U��s\��Y�?���q��׫n:}MN�����#�ދ�ǏI�7g�B|��?��K/C,�Q������[��������m��مo�y���$�D�H�����>؆G��=��lc���9�����h�}���W�>�'}�'�ͤ�h�"|����/�DB���$%c�xy�3x��G1t�t�e�XU�ELE&'����6=�.3�6�H:x����!S����I��%'7ؗd�(�8��c�sP(`���g��
�zL��J��0�^�_E�e�=�BC<�D"��u�*ON�ojR��uR��\n�bX �I7���!Z߀E�Wc��5ȶ֋�XKđ�5���u�GaӮ���d�l�8OQ�#ԏb�<�vlx���i�`hH��@�Q\������z瓆��BJ`5�7p��V1k�X~�1w�D�)E���xan���T,-V��i�f��/ȴ���'�����qd���ǐ�5*@�Z���(���0В14^(���Na�\�Hqe�
-��un��Y����Rl;
�G);l�\Gĺ�ɾ!g��1�9!P֙\mZػu�y�=0��u&Z��L�5�k-T����P�BL�W:1]
PVp|�Ա1����X��0D��v��F�*�D �24��.��K�C��s�Ʀw����q͠�P,/��ȥ�=sZ����oB2S�L� �ȤS�
�P6|��Ah0�F�c�{�x���N%���G��q}faπMj3��x�x0�V�rȭ�2a]���>,2k�Au��q�+��3@�j2�P�3;�g�����	5���ˤ��@���1ytabp���LS��B�p����^,;�����p�E�+��ž�0�S�9<�50�X}��ي'�LP����%(pY�y8��=�$�t���q����Zb���)�۽}����n0�H,�X�&K�V��(Q=����Q+�Q�&dcsQ�U�1R�M)8=�"Q7����9��ϟӇ���!��׿�b����������|����3A��B�rk !��bj�t�(��N���aʘuzl%N
�Eh�+@��A�z���:_C����8���!Ŏ!�jq;v䖭	�8��Q�,LPT[��{8�@�C^,/���#��.a�\��N
(d38.$(�,�-�8�3|vJN/�,�����@��Q5{���@lHu(%������0	��g�+�ې|L�p����
��jR�ijH�ĝ<���)���\V�`N���"))-�\c���.���M�87����I5��s�Jx{����_`����(���w|㛸㮻�>�Њ@��gC�N��{Ƴ�>���1	�Z}����}�]u9��h|m%�������~��Fd"4�����5|��D��A](�+���_}?��?���c�YH���+��?��Y4Oܧ�L]�F������E�$i�yٵW��=,Z���i��=@ytw�}7�Y�,�N��?���/�
��
$(��&@J��6��~�A��`'Y:�oh�57\�[���-_�
q��ڃ��Ï������>ҹ,�/]�?�����U��BSZVU�����شq�X�����;�ĵ��*E 9Agq����7x��{024�^�3zp緿�����z��s�P��7���ߋ��w�T�[s��w��[nF�j2�6�mc�����#��wϾ �x��N&7w��M,g�Z����G04p
�������<5"�3g��׿u.��J$rY�s�ͩ�KO?���v=�N!�L@gg+P�=� ��!QS��X]��HF#��GQ�)�-�-�L��Ԍvv~�q�Ɠ�]��)3D�����ГɡΌ!V%�1@��e�Ї(���o���њJ�%�@<Fq��)_á����&"�%p� �Lq������y�]��_t���O`�\��� ����4��.�S�8vhJE3f҆s�<', *��?�{�x��~c��-�@�BMq#.���$��FP��&��\$*�å�sP�T���s��9�Y�б�,X�:8��B��c��m0�1,[�-�-���i�h�99��i�>���G�����PwQ�F�d�� ���t�+�aRidxNM�B	�c�b�ytd��.����Xt�B���u��`.'����&�x�-%_��hj�3�q3L�^v���W�B�HK��hK�I���R� ���U'ٞX_+�m��B��SRu.w.��2���
f�eע�3#���+��2���+6`�+�pa� �j<
d-�f̜�����7"�ʉ�.���B3;GQy�H�J�jՇF!���
�G���l�d�1���l�*�|R��%������B=�և4~ͽ�LPr�y����������	�D�LT�'��#�VF��t����VQz!��B��tR�8�?M��92����ӔҘk��|��Y"(6X�(�!YR�P�H}N Np���}�
�l XKf�:aސL1Ts���lv���U���#�̠��f)	#{o�l{�=|�s'&�Q�C,��:K���wš�$h���X�lڻ �i�Ñ#됚�D�b�۪�i�B���6ZE�M���ؚh���೮��<���|Ͼ��<�5<<���S(�����OG|�+��(rы�X�`��2�R�@$��ڝ7*m19�+��RT,)w��XЋ�0Y��P�P�1�X��l��4���(~�,�r�)kR��贏#�Wz����Q'�@ L����P��b�t�p˘*Pa(Y:$	�W!I1��XL@���� �W�*yح�&��|N/v5$���T�F��j�f�H�Z��\�(��!�c���2�p9��x��CGֈ���1�Бr�HUD=N@��4�5�(��4LBC�5�(ں�����BCC�x�5������)������6��2�]�v��-�M]C#���j\w��h�lF"�5�m��`7�������� �����u7݈�/�::[�%�vǏ�+x�=����b��މ/^u5n��f4v��Ν���8�{{���z<x� ����s��7��Φ+����llz���i�������y��sqӭ7�U+�H�$��.?��C=�-�l����R�,µ�^�+��"����}���x}��w���8T��s��ո�K�`��������m�ڶO<�8�~����Q�����o�_��B$�ض+n{w��s�¾��nSP;�[n�^z1:�{�C0<�wϬ������������]y� ���vA�$�k܀��؈��A8�+�����u`ɊejZF�d���>�dН;wKAf��3o�[{V�\�ű��11>���mݎ��!�-�͸��Kq�%�J1��	A����;�o�qz�Y)�i���1�I�v�J�8�tvb��h��P�p�q��lhQp�}�-n���^�y�����N��(�%e�T��yh�sR�F��DBp��
���TpJ�Q��Z�I���ֶ&���Nd�|5����0�UPpl�%���S5��t	,T},ZuV^t��l�ah�43.Y �ό.�F��05*ਾ�u���"Č�����������&;���#c��q��#)C\�XxI�P�*g�k���h�hŲ/@����^$;{Mf������?pcÈ�uttt ��C2A$E*�7��X)�HW�������8�g���$;�,��U.��{f�����%�}Ѷqld}#J(�+���c���Y4K�.C�D��9ϑk�BuN�� �E�W+��7#ֵ��m{���]�'���-L�O��;E�CG!��$�=j2W=I���!�~ǵ�Q7�޻�4�TN�DԹI`2�ҁ��8��dR��K/��?<#�ez�ӂ��B��-�h휁��Hd�a���	)[l")p |q��R�;�kiE�PH�L�m](i���&��=.J o"Ή��@5�P,��V��Z���[s
~	]�j!g��
�����)<g4CQ2�H�g�xCMcؐ$��󅠁�?S�6Ra�;�k�9
-���PmŘ�`H��t!�T��˿ädqt�V5�!��tK(�.ic��D\�����b�63Q�e�sϧK!58Mf2H$����<C�k���/���{?�L*Rbb��᠘/HУ�9hn���sWb����ջ�T<�M�/(>g�&�2����)�'�L���&��9(�P�և��s_���_����;z���p|N��`W<@U��*�p��\ x�Պ�ZE-&t*��vI�=mJ�W,�gA��\f�%��D��T>�d*���>�����(
�M*�9Tt�P�GjG���Q���>���)]��a��%)-Ky�9�#ol��p����XIb'�Ś될��y`�Żx=�/�x֬ڄ>��:-J �pn\a\�,Tʝ���xʒP�9*�s�͎���Ld(nԢ�Fch���k�xE�"4��TD�Z����{>�D�t�޽�&>۾X].Z�D8��
�1�Hܻk7���>�xJ$�x�YX~�J$3&��v�Éc'�w����c�-�'RUV�^��g-F]c�W����Ql߾�?:���)�s��Yy��B<�B�<^
�
ڷ��.&'��CK׍�Yݸ���1{�L�!#�۫����غy+�������9g�|�^����D2eq�/�ŉ�'�Ɔ7��~���s��5˖��ҥK�ʤk��'���㏱s�v����9��p�^���χ1��]��M�p��I�IF#u�n���7��'����xo˻<qR�_=M-X~��X�x�LsdS���}����7�{�.��#��HG���V#S�P��ajbR�Y�.&'�;����Ӄ����%�7����ٳG��+�rTGK{z{{��ۃLO��r���8p�8>9|v!/�j�TB(Z<f͌J
-_��/c���>��$SB/s�Cז�'n���zwd�X5.�q��Ƿo����ÞG�׹[@��Р=�:t$Rjm��4G�WP0�p�2L�E�i�#G�?A���o����
5�%�tQ�khO�ў� J��A!��q�@K
H3���`WD�1$�q����]}�Lw(��ʈ�����YD�<��4�-J���R+���g@�,קR�TV>���O��?���0�R��~D����D �L*1*C�H�d��r��~�y��
Z�1��vw�a�"�͚�)�%�����6��&� ρ�sV��sn����"��Q�Fyx[�x{�~ gbR@�N��2i���31��u�%fe�$���v#~#Z	h�йt&:���㔁�����=G�-�������N�Z��܂��xRcr|��ܲ���7�@c<%�NE���8ƀ@j��d!Dj!��і<	��O��mhe���i��@�Ɓ�0��=�o��.�������{�r^�C$-LZbMY���Ys��ցd�&袖�5����K��x�r�$��� c�LC�q�Y��� �O�X���IR��)��m�-�w<�C��+������񵊱E���v�O�LUcK�"�iX���!88�����!=���
jZ���L��i�BX5�g-��#��$ݚ�j�("t��(0yg���i�Bk��Tsh:�^\��5Z� 6.���6%A���u�^�ƑQY�s�z45��H�+���iIb~��c۶���	`Zt�" -��:��UX��q�=.��
̜w�f�É׀0ߡּ��aF�!�fG�PОj�|��g���C��?n���'�پ���P`*&>���|�O;�#�$*��Y���X�Ͱ�-NC%���������Kҙ!aB��A ���p)���CM\��)`P�Rj�!cT���È�*j��Gp�w����3E&JQ%z�G��J�$��Q�ᙠ�d�qL�����TT��j^�,��\���.~R܇B�Zg�7倞�G�5+M���0q����@�-�K���ИS��9N
rf�=�����F����������x�x�@�iZ��YsL��*�<d�rhkk����2�w]b�d�t?؍Rӂ&���"bTK1�ϩ�8]��Ĵ[�Ը��L]nkF}CNR}�,�t��SC#(���%ś���ף��CΉpf�ͷ��S���;)��4c2����bFO;�[T��l n��:1N�� ��܄��V�7��70>:�Ç?��Ȉ��5��գ��I�Դ���Y���0
,t8^N%�hnoiEs}��)
�9<q�_ ��H-�5[�Kcf�d�Ie��Q��bC:�?$�(n,ut�iiF]c�xU�\ܑ�S8z�N�f��[�Z���)�N2��IM��c||R��\ue�Y��bI���M Q(1:>��BA�J9I����K�@��TnY���N�����,����hhi��M���k{��Q���Q���vR��v�����#�FS:�u���_�u��ꏽ�6�����A�f�:%-:НI	(��n�%�lЭ�38���
��͌)MAT�
ٺ��A��$'�.mZ<4Ţ� }(��Q����a4��C��+�����F���h\G��COYh�hC��yȵ5c`z�N	��t�[�d]�x#"~J���j^h���*�2L�ҳ�������$���8�cF��*��y�8Jn�2��b��k6�L"p]� Ǣt$re=��k�l�Gz�l�_w!zW�-���w�b7\75Qխ�ҎT�ҩ$�1p� ��)h����S�;t���d�gsðb�̗��������P��*�a�O�`�\��_�h�� ��E3�8��� +���fQ�����u����W��T��-٢-��Eѿ� Nlځ�p�v�Bc����4�%��K6P(�����t�>i��(;j	��Z�`qߠل�\e|��j�	`[t�S�zw��������z�=�+��I��$l+�3�Y��ܹ�1w�B�ut���U��P���͉O5"�fNh9K<D�(��˕�R�S*�d�	l����ډ��P�-�!�����X��l,9�l4���n�\�t�np+�C���f���@�P�	E-�@���uh�f)?�v��;aXX�H$tYGy����Wt��~��A�����S���Z��?Z�� L��=#���TQS�Zh� ��)l���y|���a�uBh��R����	+����aYW���0�w��	��a߁�ؾs>�� ����|,t����:J��A	ɨ����=o�]�t�Y-��C���%)�x}���!(Уn&[���T�皂Ϻ(���??t����?�wom���#��|�Mc1��Q���E��k���L�˯6=`��uP*�[M:�p��`��W�@�A?:$��C�RA�n:��5i��JMh,��s<�ԫ�K��?5l�@!A����a�BP��N
L�-��XP�/6C�j1����(4� j�r
�QǠ8�fq樔�fIi�M��Iz�/(%���%�Y�D)�`�qD�1���Q��N�ȩg_L%�R�M
h�"����:Hj�3PvJp��Eǧ0�.l"	#��NG%����,�.'�A�eA��O�:���)�Q*r�e��@�"ګi5D�D�d��G���3B�    IDAT�ڤ�*bR3�����^`�ǒ�i�q5��Fe�������'�e[:�<�j!f��x"�T�YM(��O�U�ΦÔ�q�K�iE`ƢBM��|
E�e\\��I�T�;Z1J8���(���шp����K��5���)�?�q�5��d�d3Iq.�y��$��I㘙iӼ�8���d횷vm|���q�S��D�f ��99s�O�T,����µ����E��8�'�� ���7SS�cZ,j"7E��"���d��y\�jUX��x2��X��l�|�}��U���~���TN�$��"ɬ��ri1���k��w��z[Zpb����z�}}ЊS(�ax@{�L�Dh��i%�@`���?��%)�W_܇���n��J+-���e�,\^�.��1te�h�r�A<�D�룜N��cth��}HD+�dp+�8a%2i��S��w���^t�Y�\�X�F�S�P{��I�5'��xe�+F�Gap�?�Ƿn�>5��G6�I6߳��T�ݳ������މ�t�ى�OB�$�2$,0\�ʎ�S�<�����7݄�_�F��IW��0x�>���d���z)>	��h���+8�q#,ǖu����]IS�뜓�D��	�W��Ύ���p���a����&�cj|��)�
J��*0;3�X:ͳ�P�كn!��_o�Gq�c^���6](��I*�J�\k�'t�É7>�10�s:f�1�B5EvF/�s��:`p�;va��4�uYO�Ҕ�hD�B֜o��4�z������D�ve���UL�5Dښ��k�y�:l~�=���s�2�F�P��a�g��Յ�3砫�m�B[��I؞����2�Y�� c�>J�����T{v���oĞ]��&�2\�����-�+.�W^�%,:g-��^�����@z��w�L��=�֤�Y��y�hj5kϰ�r�õ�LPj��.��d����5�A�?�g��q��0��t́�'���ߔ�<��ƕ�P|j�
�NS�+L�ڣ�8�A7,i\��@a�.yC���4i�|��|-lq�ѱ���Fa:�r1/k4׵��t�����8x�(�9��S�p]��hU9k)�EEbfT��{�x��3[�t�,_y6�{ M�P�fK3�O���57�$_�F�~`Z�p2نhK������Ϻ*�������x�ޗ^z邡��l��<J<5�������#�3GfaϞ�q��V�
�2 �\����5q��g;ӉI�ȿgЈ��t=��j�H���tc@t�(������:W����v��0������	��`@��'b��b(����骇�k�.��(���/�R,.�Q#��3դ,P�E��7��.aM~g��`ތ*A��pQ.�B191�"�P�*�J�eH��Gz4�i����-KJn@{NT`"�D�@:C���-p���d�V�i����)�
?GĊ�H����dѸ*+6i��C;.�
��3#N5��.
�+䐲��n��X����&S�p��bLNI�)K�a��7�jCQ�6�S�VI�����*^n�!U�;˂��8m,���!#E�"�S\��X��C�W��f!��Q�]5����T�/�'~J׉���F���nja��C?�[ǮYP�t�P�|n�<w,�X�h�k�I_�b���?6_c��v�)�oRE�'�'B�)r��e E���465%��)nbr#+�-q�eǐ@�ɮ�+}
d�������Z����n�m^|Tv�T��)O�p�I�=*�o۳Qq����_{�j��{�Ŝ��ߴ	o<�ܣ�@/s���h1"h�%�O �G3r���/�c�.Iw<j��� �8:���ZI�"� #m+�0n�@C��6%����L�� �Y��m�.@v���vnǛ��-*��h̥%�4��K׺X*clrS�<�XvՅ���<4�Y�X��	M�Q*U[�GrJ�
�DX�zX�b��q<q��8��&��Q�Q�g�"4�R��e�=��8�3ѧ����s�����LD	$feڒ-gY����{���ǻ���k[�*P%J$E�)�)f H�� �1�`r�\�]�}��~U�!������9`��C�����>!�ŷl��;�"��ek��[�n�܏�^{	������v%��/���'�a�6���z�>�Y��(�x� FH���0���]C�F�+��q��Q��p����פAb����Ր��8�D��[��_Dl���`r
��p�WQ�;����
Y�TȄj-Ha��h�'�˶PTHR�aI���@�iM�.��E'GI���e�DP��r�����²Tښ`��ж}p�^ �
\���K��շ��s�Q���J��V�.��x�תy����T��"�����%T��	�s!��^���U�|�ׯ��?�C=�@9���
���pD�=�P����h�׉P,�Su���A�����+��m�1�D�16:�����o���A�II#��T�όafr �����p��bǮ���a�IM�/��hq���;(�]�J=�����y軇�ϥ�x��>�܅<����١�"��$7,7�b�v��j���.]8���4����0�?n�=A����z��y��|oY�����^wܦ(���@CnH�&L�E���e遨o�\��&Ӊc�V60<&{��յ0���L�>���!&xD����hQV�_��[���k%|7�*��P9)�Ʈ�L�c�O4�uK��_>
~�M�����s#ͯ����|��8v�xs�dK�L4����"�&�yB>go��������P O!�[Tq��@�+k��mx�����~�٪TeH� h.�%�8Y�#Eoa����*�(�{�o�T�q������x��U�}��,w(��j2��~VJ�6����@���F�3o*�-��Z�(n#�m�0F�A�#��(�[Z`(�s���(&FG�'�:�������!��J�0|A�:UT�	C�X�d(���f��k�]D�VF�aAt���Q���pm*�1ۏ2�u��1��0).?����rQ�\�	�+�6���<Ԧ�&GT5���IN�r��c��5�oT���`�6A��I�r,�aD�q-yl�S�V��� �%�C�2d*A2yղV�_���q<�2��e7�?�f��5͑���SY ��̓��)MH]p�U�")�>�z-�W�/q
�H�Z�k|��~i����È�8�C6�`���h��I\Jq�`��{C���< �wJQ���J�&o_�:��	���Ҥ6.���עR�%ZN�u���C����QE���79�����D��|m�<&���N�{+��C+Rn�*ȯ�ᷫ����`�m��_����%��c��Cx�'���!h�P�O
�A� $CA��Fݐ��I��eUۂ�Ѡ0/AK,��?(�B�LV�(1E�.6��*�9<���I���"i���sם��U���8�g���a��e��D#!�Bq�,Z�U���(؜�����붭h^�
�dj9a��r8u9�B�cD�i�  kl�����a^��J�(�%8��|4�}����fB��85T�^©7_��o���&�zM�sN=������G>�[�,"͝p��������f��2I�p�X玾��x1��J�a�5�||�4�vR3�؈5w��]_�#��K�L�������{��Q\�La��C.ĺZ1o�4.j�O��k�F5(����L�y�,�U�_�?�}Pa�nC��aҵǲ1}��|��1,�g:�ᅍ��g7p�> �\��˯��s/��\B�� ��h�JU��V�NӀ�W'�5�
���━��s" 9��K�
�z���b(�����:	-f <o�W�Cb��ҍ��v�2.�=���1������ׯCKk;鴄�qk+u�qk���僠ߺ��x��7���c�fJ��S��W�(d�15чJi
��/��{��]�>,�f�/�e�M��Q_�ףj8��P�\�����۞(X�?ݐ5��sP��Tg�4��Y�2|,���f�u*���j���x��a<���{�,���F��|��.���E��ה��gU*n^�#Q[�%WH��t��������ԓ�>2�!2�̕ZL +�l�s~��DP��B=�:[b!Sqh���ў��k�c��-^��c�� �AS,?9g�M��V,���p�~2�:��_�Ϧ��ݡ�[������˯l�e�D��M�����xY/AP���W�~s�f�m��g�1�iP�	��p�ee�W��ez1#fBl�H5�^���˲7�B�*
�>�EI��z�C��dDi�d(p�-5i�f��	�e(�j�d�@ �r(����t���c�PP��}��%�<��Ї������)��P��K	�ؘ��¢#ݜFss�𪛚�X8o�4��c�z٩)A��*��g��V���t�K�N�+�xR9�tC�@]�� �3�;�:y�NI��>G�t#��:��J��k��n�0"!�S�K$]P|݇�]���;d�Z�I������CP�������O��Fq�U�g�'�$g�bO�^9*y��4��Z]_�)BC��r�N��o2H�Y.-H���	W\~~&����(�g65bcK�N�}G^�<��.����v�.iJsK�]"��h}K�l���I"bI��N�NE*ћ���"�f��*#[�?�di��7:co["*�]1:/^o�e�0�0(�:
���KI|L�L��,�y�H;��}�"v�n�h*x���$�
r%����%~���6��yՐ�P.]��l�-��$I�18���+�}j����B�bQ����vۭ�ӿ�s������`��O�r�
��,J�q��|@kX�t�d0,��? ���Q��� 40?C����xI�a�Z�H��t�V�L�-�)l��Iɡ캁r���ػX��1y�^}���B�WF)��� �pSȡl8�c#V�}ZV�F,����M�_���;��3��ĨW�٨LL��=�+��C�XB�iH�Z�R�4�5���K_��=�m �a{ ��k����q�����L�"�p �` ���^F��v�z�S��৑h] _���NY��kd�P�ü��I1q�����FK"���a�@f(d�WP7tTS	��w/v�O����lӇ�ƅW^A|l�|cV}�);E��q�[��]��̈Pw�0���S���-Ui�@a���á��������=��?���(�;��u&��=���i �	\�@��C8��!42��z	I͑��r�A��H@�f���8�楎p��̉|�@��r2؀�u��*jA�5���|�k0[�H�^�5wߋ�{ 3�j!�C����N?�X�-��u��r�j�Y��F�#��]�1q7(�LB[�X��Z�����x���O#o���j�QȎbf���֬��{��Ʈ��H��\R/u�;�O��U[���F�Y�s(P4�����V���y>��{�?+�78(��g�	��Jy�#��Tn���������6FG�`tq�i}+�S�	����<���ny�Ok ���o��o����q������B*�S�ah�VS�γ�L��H�df4&`M����:���\aЙ��9T����h���li'��u��v��P���	��u3Tx^YT�9$�g&�C����2?�/�$��_�>q䍕����+��oxp:�H�4"�E�������%���>z���n�>�)p�8�\�{v�|2M�{YV*|j
H5඀�6������F��P� �T�Y�(�~��|>�2�/?i^�Ab��B�q����$dC���������:`�C(GC(�Ld�:�5K�w҇�R��DPdp	���C�,=��g��C��y�kO�������ف��v��6"a|t׮\��	�_
.GFF��g061���Id�%�.A�v©_��*<M�
L��QL��`TK�lq&��ߏlՏ�l9P��Ŏ� �ʡ ���	�-���^�&")6���{:J��Y�?"�L�
�G�3�H
�,�I�ͽM�a�ns��!�J��]����א���`����C����1���5��-�\w����2̸A;�x��.Z�ւkM��D��Mgʦ �#J�bx=(��Z5{3iM���&�V����Z5		��E�Cڑ? bİF!W���ńsZ���G��� ��f��6 b�Gw��(����� ������E��2�C��ي���vg��)�\�u?��4�f]}��J�>{i�J�nu8�����d��!P(�_&KT�s�UHsx�����-W<�)�Pq&���4��r�o߉?���bŲ��<qo>�}dO�B ��M��e#Ơ��&��!��â���2sr��
��:C�M��:h8iW1V�`��Fؒ��1���9��7Q��t+~X�-af�����~����*��U�������c����Hv�6�����u�2$)$����(�P@l�I�$�A��x�SS���8��a�:��ᛞDTs`�Q��h]��?�,ڥh06�+�����8��g�x?�Rv9�hk3��u���q��)Q����هD�<h��\�~�%��d�ġ�z&&�ǂA�=~/?����aۆ�ؼqF{��s�0��]�Q-��#ҽ�v���G�_�Q�X(0}� .��KDFG�D{�D���p��*r����b���Dc���K�{6[��jBEGQ'J����@@
���)8�#�������-$�a�;RX|�=�����h������>4�����HO"pf��(�>%���0�A4���P�dr5��6*%%�� _��Q�3[�+BQ�!�d�aq+lބ��=�Ěmb�)�������ǻ�A� Ba �+�;��ƪ�k�'�F��ç����98U�]��7�:���ϣjk�G2�btQ�M`b��L?V-��=�va��;e��5�^?ԇQ�-�N��\M]���MPh�/�@3����#d��|�q��ސ���4��/	(��֑ Ӌ�q-Pk~ԃa�ON���ã��&����_���zCi�y*�[WC)����@\�y}��GmЕ��a�MRA��q���X/9���*�f�U��#æ�l��D<���V�"4�H� ��fE�F�5����-��S�e���F[C۷�Ǿ}wa�������ƕ��J�P��GI��&�����_�D���kn��{��M����{��g���������_�y槿71�m"u���I���7M�\,�`w}y�~���a�m*�+KM��0 h��z�\��x�+bE#�[	��&�f�,t6��&����#h��#���K�ސ�Z?E��wW�����,��س������T͇�:p1�A�g��5Q�1�*&�i6�Vv*�1��[@��tʠ �
�&8"�T����&ej$z�6��m>V�߀�׊kL[{3����^���jU18<���>��+�Ǎ�!(��Q���3&"�W�pQ�D�(Q���oՒ��ͲU(��P(FsY���d�b(o�P8*�Jlꙝ�\��=tGP{���#V��4��	�7	�{��(g���RNrm���t�41�����@���8�� ^�D�%��G޽�qOL�@�9��}�����$干�j1��8��`�gE�
�~��P�I?��j�L�����ߧ�21���p9bE��ȃH4���r�\�� ��s�A0@�.�Q�|A9��5Ѓu�U�(�bW�P�x�3(�teR�Y8e��w��� �_���Qe}+H��Bz��jA�y|L�~��7�ȑ�于��OQ }�	�L~�y��{�E�V���>.7rJ@��C����	��i�����^�/��?c٢Ř8}�?�,�F�\�Sȡ�) ��Q��q$*��1�+,�e(��>�\Ck�@W2��paz�Ӣ�� ��0V�Q`蟏&y�4?:�q�����d3Bk7"��g�շ�w�óx��o��7^�?�C ���{��s_@d�b���{���w`�Bش��C���N��E�������N    IDAT�8��#J;=�J6*�S<}'_~��$��l���͛����Țm���j�@��j=�!N?�z���X?�I+w�ĭ�������&�{�*,[��tZn�<���%��m�ɟ��Zs�s��_��H,���7�1�kxo>�-\|��4�z�,�s'�>�E��v �W�;z'�{���Yٍ��e�>3��_~���-w���c�R�h��=s�s���Q�"��&.��r⨫ί�$d�F����a��{蹌�Lz�F����ރ�� �v`�A��)|��OP��E,X{�r�A4�B�L��D���Uc-� 7@ȿ}�n�0=��U���X��"�`��X>��v��mA:��aņ�ظk77�����	���x�[���?s�x�����5K�ۏ|A�����E[��0Հ@z������p��c8{�l��&�^����Jq���a�=wb�={��a�s�?�f�W���-���W4��u��ِ���+ƀ�݄`�NoS(zו���&[�'�٪Ք���<"��-�[
�T'�nh����šCq��a�������]���n@�sɖ��r.X�U2�j���r� ~��8 S�$���"���tS�+���~<T����u��ǒn�s��5q*Д��`d2�"v�H
]��o��oŶm��m�Rɲ�Y��K4�&��l�Y�e[���|�^����DS��p��?`�������+���W�[_���]G"ՈD��`H�ATAe�&I����R�����I��E�-7 -���
��7-���E����/���, 5���W*��0�*b��D��@Nr(���)R�4�?Ō�minD*�n�P3B�k�w��ʘ�d�^���E�[�(*��n�и<gޔt 2�j(�S�V\U����s�i��$h*��6��3���ǆ�[�a˭h�߉��8�����_��6��Ó�qcP���i�����:r�:��
U�c2aڧ�*u����'�Q�!H7���SG�lK1���k���?L#+j$C,�D8�ѱ'��8�4��s�������&\��-�Ä��jY�>�-W)͢;p�v�Պ��ԥ�V�B��ff��K�+�["9���>�H\����� Zeo�ZU�MD�4h��:��YRv�UP�W�Tx�1()$��D3P��B�%e``sb;R*��Y~>Q&G����*��|�Y�]1b�ȑŭ��С�"�3�0��[�jEE��0U
_Z���:Jl�9�
��&�N�^�ȗ�e0u�Z�姲\������3jJ~��ץ;�)�9嬡t��O��й��ǌ	<m�GD�Z����膒BKM	E�V��ʥ,j��m�oş��_a��e(�?��?}��Q������"n�1�LH�W�
�f�.a���q����:�:�h�D74i�2 5��Ր�V`��������9��[%ր��hx�s����x����~�>�zϧ�X�����F�r�������w155���hN7"H�J&8�u�~n����O?r���=6�c3ED�8�b7�ǁ�~ �_G�6;`�c�f���?Fr�vTBl\��4���p�:����8���c��,R�Il�wv~��@�
�^�"6��TM�Ͳ��X�>�M�\2�I�+� ���i����&t��B�����}����/"M>3�*[�����c'jN�B����sOA��5�V�\҅s�cx��P��q���c��=h]�j$� �U%|��`]�`+��b�+�M���Z�|�Z���|�\��Ӱϟ�R�	�ƶ6�������t����џ� _1��ݝ�64�Z1����s��8(�,ѤI�HŖ 0:̔
���Kx�_K�i�FU�����)pno�ҥ]X�m+�ߌl����i>tO=�c�>}R(0�iɄ�u�W��,��\���>659FXj�X�2a[�%��T���N"#J��=u"��4&FzP-�ᖕ�q������`Dc�̔P�|��U��҂)cxQ�9�U*��`��+}��ޗF_�=o�H�P ���\q���Tz5xͿ nn��2�� � ,��4Oܸ�� ��)����Q���q%�G���������=�3��~$��LuWTn�
8�P��y�APZ,���0uBb8*����s��r<*7���I���A�~�t7�loAkKZ�M�3mn�ݡ@Q�\*��-繦(3Z9��MG������&�?�����ǚ�����#�PD05�J7˖@7�)��wӈ���A�M@�9Ju�+
��:WBEN�r�1��7L��I�;�x��9�1�M�-��L���@/t�.	D^�l�M|6���#�գ�#�H�}~��|�����0Q�c�X�(o�X�H�#��Q+'"@1g�*GZ�����C��"#ވ��g�R�>�:�ķ����mǶ����{!�������P�p9��g022�bfZ�f�{����y���Qd-�D�uab�\srt"��$M�R�C.6�@-�ԠG¨tL���I�Z{2{��V�T�hD�E�K�~I��29gK�!�ʭ�����
�������%0u��� �j��u�hED�Y�=a�4�Po���k,u)
eY�
BW���k�ϢO�S4(����v@,e�`7wB�O�e���{Mg�:8h�`��`@C�f
$
��PWTˆ\��:�X�i��*z���Q5H۞ �ޖ����� H��O'"E$�i�:l�,Ϳp���(�=	rR�y�i�W� �ZↃXM���@��c�f�"y��Z=�*+�'Wt���|v}��|�/��^��~����̱<��+B��騕��228�b˶�����%V�^���8��������L�P�RIj5
��x8���{}���D��l�m�t"Q
A]�\f�p(�ؘ���f�"�:t��P@'�B(�ʵhz�����Dy`���	���GaZD�Xw������N;�`[�փk}���ފt2�u���)sc@Q�r;�]����bd2�x(�HYǥÇ��o~��~$�"j��W�?�*n�v$%�W�:��2�ũ�~��O=���#�ڀ�����G~���NLbh`H��T�A2J�r�"@�z&�
��j>��A�9zɦDbi�+u	W�Pp��#U� 5��5b�={��K_��UB�XGO��O��{�V-��ގ�x��1ئ��݇[���X��Z�2u7�VbH��*��Tɻ�+Ap(X���Oq���r�$�ŢHǢ��кc'�yQ�=Q�̑����7�J��j�`�B�L�	T\=�n�\��hUjx����&G�028$A��f�Y�� tj+`�T�#`�	h��x��,[�b�g������~x�RE��5�W-�Cߏ%K�!Mî�Rˣ�Qy65=(�Wz��������ܦ85��	L���V���5���Cw㮇�G(ـ\�B�@kU�G�!�n�\�y(���Jg$�A�n?�X��
�Qf�|Qi�z�a��Yi�u��ё��$?kok����&�X7�rO�R��2���Z�:�ս�4�4W5W7 wnN��+shP��v�le��>B�!�$�K���Zh�.��QlIϣ�L�Y^��8��YnT�}�Y�:K׫�:/����y��M���:�1H�%SC�f�����H�oۓ���K���^��	}�?�#�x��������7x���-�"�L�O4(Q0:�T��(���K�u-�bw��sv�&U_�(ʍ�b��7������Kl}J8T�f�7iP���k�b��I$�D�#1�1"�M{3��0I����D�Yh�Y*=�g������B	���,E>����@���JQ��5&/W��W��C��
�xڻ�R��l���g����8Elܴ�vlǂ�EG��yd��112 4�r����Je&F06t�W.ʦ��u��(���l�YH1a�m�6�ѝɆnWE�g*q_!�?h��0��z�0��D��t
�HX>?Ʒ������ɡ�kA����J��S��u�q���{h��"*׏;lz�	W���S�Z��V��F1Z\r����>'��U���T�P��V���)N��\<���(n<�I���72�ۈDR�����,U��B�� �禆h6����j(�p����J��P��8�����e���` W�B0��ل� ���������S�� �P�Ѐ�~�Y=���<��tm�)$�)�-�S9�f
�u����RQt#�<���⊡eo�#z�P�����k=ΰ�'��J�+"c�%���z����B����7�?����5+Wú|	�y7���ݡ����MA �CI
�)��L���*0Z�#W�෪h�i�����Дu�dk~�flLP�s[�1��=A#��M9#�j�r�}��_�I�kp�^|���?#dIǱr�>��GcA7��f191��'���9�y��I��b�%i���a�����Ѐߌ"[�!��(g�|�}����@S�
G�"�x!��_�e�ݨ��P�(`��/�쏟ǁ=�Kg!��a��;p��>��m��\�����Ұ4��"�L� '�<��TP�˂���z��!7��|�p��P>ۇҍ����o�ܛ/!Z)H�s������P���@���i�z��(\<��y��&�nY8{mՐ�5;o��]��Φ��C�H[g��p�6���4�k"<U�#
�������8��(�?�5�0�0��f,س[y���0.�} �}�t`ç� ˗����B�X�y�KAh�I�3�����(Z���|�'&E�� �x<*�����e�ĩ��}�74 �щ:��\�.^�����fFG�P)g��{!n�c���"Nr?,�%��*�YGcB��=}x�7p��B���7R�$fs��M�W���5�Ч�Þ�G���������R(�&�_��.J�m
�1"`�h�n�l�o ���%8@eIx�]ց*���3����\j������ҍ<;q
���km(���R�Kw��79+�aGX�n#��'���4j^�>wJË� ��M\m���[�
o�!�	V%=��v��P�f@��Je��*�E�,`�M��y�7�u2"���`�n�]�wSP1#ѿ'[�!��P�Щ�
����7���c߿p�w��7F�	A��&#�\�&���8��R���/7���ˉ����C�Gn27	QQC(>�e���L�f�+���?���3�0r䁠�@TS��73'�H�� ���F I�C��pJ`f�5�j@�Ot�0��G�B7�L86�-q� �I�(�PruA�ep8�6�V�Go(���(or�#l��a���b��X�i:�C��Tr�O��aL�@�g�ed2d��0����%�]@�f�gFP��=� %>��1@��p A?7(5�D����z*R@*3���UR
�ކ�H&M%�"�����?���s�ru��+�����Ҝ킇�x��f�6���n���!�Z�5�"hv=�:F4��9�D��ғ���@��_�����sSC��u��V%�����1�B�w�֒a9����~Pq�«�I3�5(��G!?�\����iI�mnI"l���+���JMqx�z����fIy�x�*��$A�_Ю��~D#qi�+�,�����&'�1:��U4�b�p������0��.������'q�
�����5��U���AQ~Ԡ� ��	�~<��R������%@����͡��W�~Z+ZE8yw(�Yزe��,Y��s���鳧��N)�P��t 茇� �B�[PZ+L�l��K�g?2�Gd(�r��Pૣ ]���B��4--f��(�Ő�Cȵ/@�ßGb������y�M|�k���q���^���?Ep��.D�"��q|p��qt/Z,�é설�2-ٲ�(�����ϰdשrAԈ#T�pn�;2�'�#(�\+����C_�+̿�>���M�ǆ�/���7p��p���aƂX��V�,�y'`�p��W4Vm�H6�P�,A.�-��,����qd�锜lp'�'��L"h&eS�����O~��{a+'=��k������}�yP1�A��i��ٳ���F�)��d3��+�Ƞ�%7`�]�ES@��ZUGE(o���K8Z��/�������Y᧞'�Ǚ�_Ʃg��u���BH$�,\�e�m�]@(	��ű_����+���߾���$;P�����l���Y�ՙ@����~I~��ގd<��LF�eHK�hm�m����~^�� �;Bǥ��r������_�˚Aw�|lݺ]K���c�U��b�S���X�P�.���^|���UIwO�E3��]�O��A���-+[��g�=��4±-�T�<�x_+!1k�j�Ք���`�.,o���������@m<��r�S^�({ k��P �^�kP�S;z�gA�3���x�F�Ź���Hx[J��\# sS���.�>����y�P~�2SQ����}.k�#��9}���*Y�ב'�M�>(#�SD��\O^-&m��ڪ�V'��u��ѵж�j���M|�J(������̿ג~�)�6뿪�������=��;{��R���G�""��F��%�(�\4����c
)R�����z��$g�޾:������bL��tCL�#wZq���:j�kz�RQ���,1$��	Zp��u"���4i��6�h���%�Kt �ѐĵ�A�k�0�Z �hy��au
*Ŋ��8w(`���f��x�g2��E#o4�W���+��:��|�SX�jVn؀��f�!MB�(4��LKSN+96��Z�I�����E\�~e�@]#_v�?K�T���W��CQ�B�"����c�Rd���2��e�sP���Cb�� ��n2�E�<��b�~�^q����&gtn�(�}W��]3s�~�ܢ�ӝ�c���y�
��C��~:�*P/B#�#C8��*5C��p-��WEI�����7ޡ�I� e������`�F�Ð{D�е���)���r(��/`��qe�F�pJ��O����'O�{�Blܴ--1�괫+�T������j�`�D
�=�x����
֭Y�;vn�ڵ�� eBr�����f2sM��ƅ����5d��v��D�Ahu:,�n�a�=[��-�Lu�X/~�����)��J��G�0����#�m�����j�Ǉ�����s��N	u�T>l��TK9Ac�mۆ��ɟc��E<yo��	X���2�9�Р�
"\���2�U˒hLM�iCǢX\�C��ʝȣ�|]��`,�CD�Kh6L�H�A�"	dAL�u"~�в�v��?5��C�����\��������U���
��Z*�^��g�0�=1�����0`�L�sY	a�#�N#K �	8�d�᪎��g��u�cא�
�}h-����_Ų=��h�S�(F����������
=�aَ�������;���uhxH��.q���;�KYJ8�������ԀX�I�~y��x�4�@�|�g��������G��ҰZ����=���?��m`���r�}���=s��q�[QL�p��0�9,^�[�ڍ+V�-�_�Y���r.qu�3�ז <gX̉�R�EO�2
�8���qᅟ@�ч���UE�w-����s��zp��_��;�b��Nl��{]��d'��84�	��9�=��� �(�#����+�p�C4�chmi�,�Y��/F*���>��ꀉ�y]0#I9WFG�148�|vSSC��{^(D˗wc��X�l������I!0��Й���KW��O��_��?�c� ]����*�qT�q��j��ý���%�<3�Ֆ��4�!Wh��k�eE-�)ne��6W�s�ļ���u���\p�21]��л��.���K����v��}B��	̳�ρ�K��Y$�͢GT�����m���2ޙ5��y�VA�.�R���g�l�ݤc�d4�#5`��%t,%b��o��Lѕ���~�{��#e    IDAT�����W�4*�Y��@�9[Q��C��Fv=�)�����'C�����9O}����������/-�����2�T��ؓ�A/vI��5!i�$��>�msib'O��OtT����;�{��Cn���sJ��E�����/`z��!D�E����79����!D11-��2!E��'��]e�Q�
Ѩ#��0�q,X���܂�����l��ڸ0>���v��؅��K�=�]�3
H
��)`�7i�9'x��oF~yN��dL\"�o���C*�U����uL��"�lB(�D�@��C);&���?�bU���P}'K&=�ə��̚>�>G4��UA1_�Ͳذ��'2�!O�Q6����J8PT-�n�$�"+џ+�EZ>�9=�Bu?���gϦ�W�����"𠢦C����J��>{:RsEMԱ����&{QW���jL"�r�Q�yE|����S�
��h8������85�j��"��mX�~�<v��CN��Bb7ZQ	�eZ����i;rǏ�M�f�r$�|��/��!�xс2�2���P��7�G��Ǎ8}�$�	�u=��ޅ��c.���I�)����ЖN 4�/�sm�=�.���a���C>�.sP*b՚$��6,^4���8p�":��L���`��\�FB�V{梨��ǋx���v�<���
�
vy�������L\<\�RR
9عT�Y��oߎ��ɟaقE8q�>�=87zd(�U�S�#�:b�ЇH'$�l��*C5ӹ<�
���J$��ɦ��H��Y��b�*�PP�ФX�J�-�F���ڽ�>��-ۀD��Q��O�ҿ=���u��(n��C��O��𲵢E�5~����`fJ9��#��7�Rb0��allLh�D����hlFc���|�2��/?�-8tB0j����K�5�>��S����3��Sx�߾��^|������p�oݷ킑nD�X��� �V�޽d1/�B0F�\ƉS'e0 ́�J��S��;�%?��)����8��(^�	��T`�M,�s�|��\����؈��q�٧@Sk��.�:�pa`��Hu�b�-�x�ri~MA��K�h�x��9��-	��M ��I�����`O�q��)\}��OE���҆�߂y����hL��ԏS����．����[w#�no���3�j`H���r����Q\�,Z�X$������q�b]�^܅֖&��7*�c�@@�������Ӣ���� J�r�qܸ~Y+��q�-X�r��$$�狈U���5�L̍���<��'��\��V,_-�� 
es(�F�՞������?�@$�|�� �b�x���>��g
���~E{�j��,��e�T&���zCpA�����U����,��n��:��,RͿ7��2v��`s�늂����z�9V`e�"�GYm$<��5����Ny�.p5w(�eS��	�ot��r�p�L�C� ��	�t~��#��;E��~��A@9�l]��Z��1�M� R�I[U�D�3�p�d�P�/��ѯ}2��4�ʧ���������׫�{1m���#����[D���=K�p-��trϭEB��{\�@ՠ���^&�����Ή���XSl���U��IA2�T��İ�"÷�H��C��B^�p|<�i𠫹�z	����n 0�N"0%(SOD���m���{q��7�s���N����� f*U��Ѓ^�%KD<�}A%�f��
�PHaT�of�����`�G,ê�+���-X�������\�P�$�iD��@��� �{�s��+jZ%�/\QZL<+Ij�j~�U$�:��?�2��%_��)�ae�z�zyn
(p�����L&�?�R�pz(��퐬,焷x����f1TU�$�p3��f��~n8��T��"����p�o7�L����D�ߵwV�Z��5Tb?5��py�s�ps��D�uDc�T}8z�~��QͨX{_�KSx�3��be7��q�o�\I�]Kd,��U��ת�l
F��11:�y��1C�ɠR�BS����֣��I��S��p��9ȭe�^�'ځ��8��޻�c��-0�N������cl:#��Em�m�
t������:���Fϵ)�K��,Q�o�UmcS ��tc�m�%c��wo�}��_q�cӶ�i"D�80�ل�eo(P��䈻+w�i����M�7hz�0Q�<���t�����L�*̈߼r�K,_ԅ����'�s���)��c�����И:��>���K4l�94�����To
���b0Uvd(��X��+�9E4i:���'E�T�&ݲ�O?�\+���W��w���/�_f�Tk�{~���Z��-.=ʮ�01AZȔXRK��܈P0"[H6���e������	��[�lnC�De<�����ǿg��ʌН�����/!<�5w3#���#'���>�7_~Z�C�l���o��6	5�[��������}�ҥ���)V�v��7n�Jo��y�1��tɆFh~*ơ���8�ӧ`��G�)	-o
6��~;����G�{5P�YL8�S?}����/_&D��3�22'�C�5���*�Pr7h_\PK�j)��_tS�qht5SBe:��'�a��E$&F���a~Đ0H�kV~�n�H��re���E��ҳ蘗�އέ��V��n�Gn
kn��T�ଡ�A�oxx-MX�n"�(���k�"���`ldX�\��i��$��h�X�H�Ù��ׯ�PP.�DK09v��(-��U�Va������h
l'(�/C�h�-M���5<��sx������+b
3.*yTKS�N��)����Ɲ>�p��uSĝ�e
=H���!�v�b}̡K�N��V�%!� �Mq�/�;��fc�&�*��|z�Ho��ߕ-�!x�ܬ�J�%y9���m�)���'�A��W𨮲�/7a7k�<��y���ͦw�x��&��b�t����JE�T��CY��S��\�*Am��Ɵ%�_b��aDQb�3�@��=��P�*cɅ�{%G�Hi����r(��H��?��*;�_�Ϫ����_���Ǿ~����VE����q��q�&7��*$>��M�]�+X��K�-ڔ��P��{�CU�1�H�����c�iF�"@&�H��z`V�_�
��4���d�(LMH��۝�ѦF��hf8.(f"�@#��"�llC��02�2�lX������cp��	A�g���܋��c�,V0�ω5oқ�g��7(���K"�Z�Ԋ6�!R e��P�.4ш���`˶�X�f�lL�rg'�s�,FGF$8��m�Pi�1p��._Eߵ��k��l
Ul�����N��h�44~ĵ:�VIhX�LS��N=���C�f˟G��RS�L
g����{�ө
���5���Q�F�v���-�m�[��1y�yC�J?VE^Yt���
���*� 0@a[�*!�`�j�n[���v��5���w��y��㷟�&t]��^�p�
�@t��Q���1	!"��Hhظi!�k海��3���QL(}#�h�:ʥ� j�B�i��hAg���F�:�x܏M��q���n�ab"�W^=�C�A0�ÞM9S��(֭^�ݷo��ŋa����!=~�3E��R�۽۶,C�)��\�?g���Eü��MG����g�bqw;J�:�=to�uV��n�Lԙ�k�PUF��C�t��+�D�b�F����@�7�p8)�8�L��>+*�L��\mL=OJ݌�l���+���W
}�g��|��$D�s���0dS@KR
lI��j�)���M��D�!E�P�Mnղ60��1Y�P@��M���*D��i�BQ�w���瀅݀ƍӧ��������l!��a�}�p��1ҫoA�!�![:mB�1ĮP���U���Fr��
%���Y��d��q�I����x��P�A�g!��Ԉ��2���)hM�F%>���U��;.��w�xN6�6n��=��{�CIg"vHH��Q�DP������|��0dirz
� �!3b���=i����U5\?y�>���O�-Č�<Ɲ2�o����g�\�	Г��$��{'�Ch[؎��w��X����
��5h!�I��T�A�\D���ZR��t�����X3[�R���d��qS3�_)b�^G�Z�����vlx�з��������^Ǐ���ճx��}�u�N�[Z12���T��%�t���(Md䌚��"[�ªXH6$�a�lܶI���^LMM���K4A#�C�r��,]C4�Ƣ�Ќ�"���q��%�l�Y���E.7���nټ�W�F4ڈ���\��(§�H *C�����O���WߐMA��er�Ѷ�CZŚFf�-)w�މ;�m�cf&��Egn�C���5�\��4�Ԗ�6W�N,V���
�F�#�r�ϋtc�7�T�:�}�
bs�u��K6�B�ɝ���z�(nP��\ 2`2h�����D�ԣ�o�Q�
�y�+�A9��G"��	+ښ��=15�5 �!�K���;�E���yS;Q�:�~���,��Z�rقR����_��l�a��>'��U.~����*U,Zz3���r,��`��>
~͍�����''�>x�����/]��Q�H��͕f$��'$���#��������ٝ�§qe��hxQ�ړ�SoS��~6ۀ�*�.�	6����P��@ov���.��)�Dc��S(MLˊU3t�\�wߍ�+W���H�~��H���16��T!�HC-�)�:vG����Ĥ4�}�Ӹ>��`.���r�g��3Ƭ-��8�C�
pҕ���#�����e��y�,Y��	��A��� �:3Y$�i����o&�+�1=zC�Wp������PP�`Qx)z�7��3QT��7q���-#�22�&�s�T�(j~���l�����3����$bq�q�a��t���|o�&n�;��-�s�`��xȰ�E`1�s9��w5$�< D��U�P�9u��`k�va��%)��!���o�������q �JR��2,KJ�̉���5\�CO߸P����4�{�ٌm[��������G02�CЌ"M�8��$`��@�}H�"��1��-�g�ύ�s^j֮�S+���kx��3�py��f�X�i�W�^�Ʈ��c���hJ�0>��Ϟ�Ώ S��g�Ocߝ�x��5��-������K3�$Raty5{۶.��6�b_��z�(�|x5�ap�$;�}�������d�k����&SK�ϩ�k&f7J^0ޜ�;�>��:�vXȢ��to��5�����X�|�����qԆ�P����<�\�AZME�P@e��)��"��o�>bIJM� �y̐>�s0A�%��}~,J$�B_qM�P��]�� �F5�g����:>|�5��,�����^����E�k�U���K|�uN�0A��XŜj�j@�\�&��I�œȄm:���)��x��2Ѓ��Ї�[�c�~�[���N��s���p��x�GO�Иۥ�[�c�ß���{Q�M梁�(�_X[� ����L��4�K%�I� 1e8i&���ۏ}�g��#̺b���}���_A����� �/�|����2c��t"��
��.L���Q�+�m�� ��`�]E�R�U`�EF��9�q��&´Y(RK1<���ʓY4�u�X�s`L�"[ʠ�ڀ�����44�W�}���_C�4����й�z����B�r��l6��%�n��ٌ��hnmB��nt,�/���Ȱ<wn[ZZ0==����T�hlL�}^7���
���tW�^����`zj�qH�`�kQn��v�^��X����)g+�C|�j>S��/��(�������K���#D�Y�����{�u�g��	7��h��s$� ��,��ɖ�Y�xg��fwkkw�5;[�מ�m��Ȓ5�H1�E�A  "��F��7�|���;�Ѥ��jm�����>�;��>���j���iX�q-���W�5��jC�{����=��w��_"a�K��j�I� �	U�Z^d���L�����u�(��!n6�}Cu�٘a3N��8@S=|>�^Y��]F�_ҪS�-��S�"]izб���U[��w�c�:,�Q�$� Z1]�ؖ�vD�c�@.?_K��؀�_��pW���y�Ϣ��y֥S4�Pד;�i��t5�&(3	U��r�Ԧ%�E��&�g#�!��y<�hI�/��,]�������T]�������?]@MQGq�6db��C�}�j������i5I_�4���d�a�Ca�mZ3/����G}p��H6�.�Ϝ`	�bK�ʩ. ��]*�w��M�5��9B�b�Z�$�,&H`R!;	-Z��7.�"��4D�Vjo��3կQ�K��*��H�2����uB/�1r���1�iI�7_*b�u���@v�
��Ą�"[*!���m4ѨU�ΑN���ʦ�k~��x��?Ǖ�`�I�>�4\4-��B]����˛����ȫ�䄉�	�.�&�J�����"S�=���'���+��T*�M[�å3��l4��ك�s�*��U���c�?�N���s
|R�<S:�t��������4���|�\�w��j���rc-G ��J�(ML�=9
�����.q$
'�=9��u�'�)�x:@]�ؑ�\��:~�ʁ�"�6WO�تNs��F֨�&�Ļ�0\t���ё��L��ü���%SM�+M��3ƞ��$YJ�7��p�I%�@O�d�P �ð�d�Ll�q%/����
^~�-|��&j43�d*�t��^��D��*�i���[��5�E�z��܉�����c׻��ח0Z��գF���U��Ž��έX�h:\��'����Soax�|�N ZWp��K���"Ho��?��K����-��e��{��a����w�]�ch�Mg�0�3�ź�@�������U�\9͚Z8L�j����dQ��?����y�
�>A�*|�;��k�ax�><����w�,��+Ш�iZ�M��9��:@�1A)Aá�K���[)���>�IA�s隀��z ����z
�1�,��¸�ˡ��|���¥tP�бcx���/����::�p�M���������z^1s`(�$v3%)i��Fr?�����_,K�ny��~3Yspb�;����<�6�P0k�F����Bj�u@����"�¡G���O?�'�
}h��uB���FX�ƪ�X��C*�'�r�l����X��N�(J"�v��h&���?�����
z���[HL����c�7h���
|�o��Fj�<�]��;`,\���E٦˛�Ww][����wR�|�݂���sŖ2���T020��pa���t�rt5˰Ν������Xy����s@�lxe/>�8��_¯"�7�M���}��� i�I�p�ʇ{�/@EOqj�B��r`���'d�@]�mmEi�5�2�$�-���k6a���<FG�8t�^z�y�=sa�D�(�Y�w�uV�ـ\�C�C!�
h*&t$��c�N��Ǟ�/+�iG��&��}�fޞ@{�J�ퟻ�.VY��k�zǽ��
��(k$�� ��Т��ue�&��I�~Mm�����`�g�O�d���2�W���ȡ�K�Ƒ���ߟ�L��\Y?q�f$�VT$S�h�m��j��3rK�I���(+c~�a�tqꬊ���Oi�ƯW�C����n�t�Ur5��{�8z�i�4ZM	���k~��d��d�lCl�#a1�v2�P���j��-�2�6��K��?���
B*�ԯ�Y�(E��������s���˿+}��ǋ[�O��2�o,�I�Q��>��h8��/��f�f��n]��9a�-�l馡뎡�\�����h�Sad��<ara��M���"�A�� �:��4��Y-�@���c�#���R��5�@�0�۱].7=�O�<{a:���    IDAT�֜]���~�N �����0$ze��m5�ԫh�k(��P��r^���Ч햋z�� -��8���$ёi���(c�2��xr�2��FgO@��
�)O1����f�20*5�/\@��@6�O&Q�lǌE�1�J��'�;�D���L��B�� ʵ&��.�Θ�9}��YLc��'����
�?�H�M*��	��H���.è�"KP��Ʉ�7�-|�ɏ�Ɖ�n'��W7Z���Q:��X�|�,[��N$4��\<}RF���.¼ūP������1��;�3�N������<W�RQ'>�+P`�(�)t�:ڴ E�B�v$��ɚc���e@�� C@��.�#Ʃ��P(#P@%�Dl���L�d���D�c�]��ZD�-���1�M5�V��hK�sFő�]����
<:��2)`��3ˮF���#���w�㉆:Qv��r:�6�F&P�1�##���4�;=��n؀k7/E&����?�k������#�Pg���b�Su�g��b�'ֱ��t3ð�t�æ�Kp��7#��q��a�~�0��qsR<��Ф3U�M7�ŭ�mAww����w�b�ۇ�%F�!�<r.�ٹ�^�M�����+�1:"��& ŵ���	L���{�bي��(���s�����5��!!�M���
e��W� �5�Ia2�#���+ #��:����D��~`[pkh�>�֮���w�n�:�:���C��1�r�E�`v1���NI��tJr
.T'Dh�d�ʤ�/_�\k6�ƾ&�`�q�v�:AA�����t��P��W�嫁T�O㭟�>�,�v�R�\=����L
�DV��Z�����*�H)� ��
���Hb���,������ZN��o��'�/��k2Di�"��{����E8�)K�X���}�1|��S�pTt'�В����ʤ`�b#�HRE��Hl�%�g������2�3�.܏O<��Oazʀ��зe3�}�@�,�K����/��Q,�v-�ݱ��h&���B{R�s�!���5M�߅�N �)o�Ь�Qo5�L��)�u.�a
3�I,Ԁ��T���z>��w���/~]�슃]/��'~�=�.���#k�Q�▚�L~&!:7���4N����*A%*�,�I۱��a�Ґ/f��ӆ�K`���d�tR	ǰo�<��/q��)o�&��lڼ�?pV�Y�t�]��8)g��%�)�(x��'��+� �Lbɒ%�'�e��"��By��\�6l޶y��CM�����ɡ�V�{�2x��_��1�Ln��,����Q���65{��?-�x����	��H�y�8.�<��7�R\?��3U�&뒎|b��&����:B�n&��U�����g�Ώ�)�@�G,��^�ٌR�P��baʹg��l������x��5 �)��be6�iMx��nk"�I!���=�l�hZ�X��k$��X�'N{�z'��
ʋ�!�w�p���_�:���b�8������u�NZʄ^��ZA��[]���Z�u#��zB��]
%JP=��PȾ��Vd>�Q�6$hS�[m����x����巒�m��9}����慺懒�#I&��R�YTs��=y�0C���,�i8�i)��h��jZh�>�s��j�/����>[�)ZJ3���i�ȅ��	��o@Dw���u���{Y]72���'� 4:L-�ka��>�a�W���:�%Z�;|��p|��_��"l�ph��;*]�\�@�m�H�b���{ς�E�Ӭ����jbtx�._ĕ�A��#8��ֲI�m4��hò��T���#7&��a���tr4R�JH1=9���k-�=�KמI��pQ�]�l�j���<B�	ز:r����)4��h�Ʈ����qj�����7w�o��6��5|?��?������Pm�I���Լl��MC�U�Ӑ�)"�C�Wp\0KW@�HW<H)�rX���I:hw�4rYh:�TF�Q,����v�6z�A�6�F�$��'���㣧peԖΑ�,�����h�t(Һ��f���h]}%�F*$m�ia�v0�c����(��.9�\St�:DW�ߗ|~�G��Ym
 (�5��oK����9�ft��ʵ�9�SfꟹaO1(P�*8G=�L���i�l�`�ҹ�u���fM�]��]	���̧-u��3*|'z^6*n>-@9Sx�����Tk-�q"�j�l�~�u�����@��;~�`���!G���_�����p�%�14)P	�1�� f�,a��p��u�)}�����e�H���VEB�Q(���~�2見����>���e�z� u�&�YӇ[oX��f����Ư�\@��@�,���uF��4�ys�^�3gM�ɓ����p�R�4�rx2�H���I��a)���iɱ��8k�\I��4�6���l��n�tv#5�q�VK���`p�@P��?��n�
�}�1�x�g8����b�!���LK ��Yt墦��e���1b1���!�3�c^�$�C9N�菣k��`�qP�(��t��1=���^=���r5���5`�z �G��E���O��C?�^)#�^Ģ[n��/�9��`^D��BIڂ���L%D�����`��6AA�0��|b�i���t����������ϣ+�!0].����ж�&)fX(��05�]��'��{O>�����'173�oFCOb��"5��>�ވAA��MN
��޿�|�D.N�Ź�{TO}�k
I�n{�7n����&�is 7%��ޡ���#��9���6��޻�%+�f:$������nqla�3;�,�x\Gg�����,XV-����c�!OC6�Eg�֫�OG��^�^¨�b��c�7���&l��x�G��'!T%&�%��1��,�h�у@�ɨ}�w�s"E��g����X����%�ܨcZ:��c��9X�i+V\�.�Ccu<p���!�����2ۤT0�y�Z���X�f-R�ǼW�˟Ji;=���?>�'}o���P���݇l�3�W^�|㘓�P,�X�������xZN`��6���S ^	bi���d6��i�{�%�C�G�������x�� p�0��ji��2�LgR�T#"�ןd6)΍���d�LN��:>֖E�&v�5j����ׯ�1}z�;���+�mL�w��E����V<}�t̥�Ȧ�x�:�)�>��Q��d,�A�ʬc�sP�iPᄖ�#��E?G������dX�|)��f���Sr�lOC��s;����}�IEd�,g��&22��t?W(}?�1�O�����a�������
�n�ֲ�<�5����i)֯>�4�
0�H�O?U���?M�DN�b��W(o��1IE���D����&1^_��}��?$P >	%d�冮�<|8��^�<�,�	�E�|�S���"��w�����]AC@O%Ӳgpj��T�\Qa?1�N<c�CW..W%�1ɓ���0�X��/@�M�mGQzȵ%�T�?���ԟ)�!�Z���o�
m]�Ξn)�&���&��YM�̩��|�d���c|��&��+`�v|q���/ ���e$Q@$Z 7�&�R>��q��A ��'Z����Vm^�6�G�qQ� �-i��ZHwuc<�1�l������|�}U�A�h�	�[�~�A|�K�!����3��Z�uԝʾ�1�h�Z�#s�0������z�(	����{�TP� l��(����a����i�c��Q�lN�9szq��b�ͷ��=�� 쉳�?s���C'pe�%Bc����7a�H&��P�Bd\G�[ѱ��:�F����a��%�mH&!�a(��\uj
h%���%k,��j�^qמݛ8Mr����i4�Z��Kf?�
�BKF�S�F��+A�g&�Ȧ�n�X���l8BA����+q�]���-+>�����R�פ#��CiTB\_"����@}����z2�K����=G1Q��@���q�]�
�LcОr�a�.�*��o���X��w�ٍ��&&j0��v�̆��yX�n�c�O����{��;tN���i0)
��!���3��}n��O���(~�� �|� l;]�H'�P�q��-�v�bt�3��O~�4��^_��g`��nsfgp��d��%���(�~�}��9H�0EX�Cj�?G{���Nrzxx�9NEAqq9�}(��[�<�T
m|��r���j���Q������5����m�&x���G���]�a���b�\S�
}������b�"�@%bI:�X�t�%)�ϯ48A�P����oh�+�Л�& �&�K���_6l�Y8�C�������~0����oƍ_�&2}�$���17�S(SKJ#%���^Q)x����^�:�^h(`#�d� 'w��W~�#4/�F�a��]�/Z����o0m���SEXQg�!n��x�%���C��лB"(���/b�歨�D��"�a�(=9i�U�%��q�Ϭ\\Ths�)�QH����}�q��Q=yX��FJ��Oc��p�~F�5�>�p����ﱇ�8u��߂ҽ� K�#LP���k�G�]<ݢ���(�4���ׄM^�|���B��rW�Q?��{��r�&��n���%dW��6��~����q��a�4�yh˴!�ts_G��BC��Q/Gg8��6�y6��`u@HM@Ҭ5��s�V$v�	tNoG{ofϿ+6nA�ҍ@������ǣ=���/Ӭ�Knܴ
�}��Z�F2�&EqP��r"+��c���=�7^yI�Ĝ�s�+�#�.ș�Ӱ���f���d�ô�%i�K��}��ܗ��,E��z#��l.�\.��.�9ً̘�s�%j��e���TdN��@��STB���@JC!Js�VSf��؇��i�*�X���^�<��n���G�XL�R�y>�3*�̫FW��D�҅�JE
hI�&-�^�$dJnN������t���2��( �Z�"Pg��ZP���	���V�[, ]���<��А���7�Ѱb�R,Z�K�/��U���=�{�p�ӼO���#W�8-n2\R�CA�P�A�s�+
#�lP����ލ��ط�]Ǚ�8v�g�f4��o�h|��F��.Q\����Q��?���}濫�
��1���#�:Ģ�-
�c"���V�N�wK[f"S� >+�������8�3/x%�W#�t�c.	�
��zR	�D�K��x�H���WȗT�'X.���B噘��}�YW�?a ��H*��>	<\%�W�əlZh�A�sfΚ�ޙ3���&�n2��ֳ`5�쿌�gN����ѡQ�DZ-M�C�b�J�I"G�E`��%�B����t��$�c�)H
0u	��@A"���4��իՀ�1,%���4`�
��p>���O.]ƅ
--9�Z��F��ғ%�Y�w=p�'��<��a߫��9V�$P�!���.#��1؉�7Q6�R�K����q�"%���*B��J�cp���F�J����%�tvR�]	�f��;((͘�fc��#�t�>�w�������3BJ'$�KKP��|�l�Vy���A�'=�Fb�1仸�(#@%�$���+����vtt��
W��MI��<�:q�@\�ɽ�{-r(��N��g��fx�X�Ǜ��/��ædS8!��+��I2A����`����k��0<�+�s�؎4⌡�� ^���+�.�9\�b��W?���/�- �l��v��;�bŒ9�������LެP���l��D�/_���*UG
v
"�!p&t ��p��u�a��A||�4^z�W8w�;цL�#pZȘ֮��;�	m]y?q/���ￌl�[��锏�K�q���b��98��O��+#.�y��k ���֭�q�mk�3���&�~k?~��i4Z�)^{Lq��8\*Nu���bfD
�N��5����|�:f��vdmM�<�H���|�bPP%(���k�����]�~��FG�G�s��+�	hO���Y��$3����ؒ�r�&�!�Qu�GG"�I�(�	
�!FiI�Y6�]@���4i������W�ظ����q����w�#�򈀂y۷�/}����r2�lҙ�H��PF巐�/֚��a!(�}�x-x�KҞC�Bg�߃������m����=w�η���`g�����@��/Wq�W��/������mވm�?�E7�@:�3���k�-�B''z�#��y��]��M-��̱V+7�>��Ob��~�i�8���	���� �IA�Z>p�0�?��Nƪm�Q��.`�r��6XZR�^����! (E9$�EI����d�Ϧ��#��Hr�'���a�?������{o�92���Ò�w��� Z�O��g��#?�>*CP,$�����#��5\u�j��y�s?I�S�I%�Ե�g��Ѩ5P���hQy��@ǌvt��ĜE��b�\�l�L	N+���~{�nД0��,֯[�{�k֯C&_R���aJ�HQu�͹N~rO>�(^}�y�p,Z��lz��D"��޶�$��U	񼾤���Cq.k��\�<�	�;R��idx��-��f0{�LlX�K����z�2f�J�"��b���.�0���/��1�1<|E�>o\��a��P� W�E�4�9*���x��W<F�U����#A4��t����\Չ���De��RK���ߣ�ac�Bi����PFA���J����,L���~&��`��f&�%5c@}����6#����������U,�5֐N(0OP Ծ��h�/8=G��0W,�0�1�/
��lPP���61�g���fa�c���3}���ݳH�ȟbRȧ����u�x(G9��O��*�+�~.l�">s,$�ԑ3.jbP ]�(hC�NU��&�<��ț�&gZv6]!W��(x��,e�%�}�{������1b����
a��a*E�S�a��)���g[~�Z���
� ��>-5'&022���1�i��.��w"�+���mc�j�eqCNs��&]�b{'�Ϝ���Q,���c��nm��q�_¥��08pCCC��z��2[��Y�%S2Ί_��C8<�2�7/7r~�t�8���=W��R*���`F>��@?�E�VC�i
��|�\wn��NL_�g���G�p��RHVo�b��a�ҵX�~�ݼkV.�������
g>����p�?��&��k�L��B�	r���+N�9*�x��Ql�Lz�	���+W	U|��ʔS��/^�;�µ7�@��>�^�����8��>t#��,�5��kH������y[�|6�F�n o5P`
*׳�DK�1��}���� �z\�at��eZ����88*��Nʤ +�X�;$��_@���+�fE?"�Ix6\8~,)�t��B��\B	���!�)IeG�ݵ&��"�e_�ҽX0w:���*$MS�ȩ亊�W��NB�Z5��ǻ1��$ƛ&^z�=�;=:�d3!V���?w#f�hCyx���8�&�7�&��`�$0���Y86�*=���!lڴ۶�Ʋ%`5���Gx��#i"����a�3l���p�u�p���#�Mb��O��S���2��n��v�%pÍ˰}��S8}�"~��(�<�0,�гrm|w�D>�[�],6�G���˯���uq��!.�U2 �W#g5�N�)��
 �h^t���=�_�.��j�D�@M����89m���'ЪW�>V�߀�~�7�u�zX/�_�>�(�����3��7�af6���vd���418�oV0l5����=AMA	3ry�X���4&`��r
*��t���%LOf���0h��C���̖�@�����ί��?�?���bg�ܾ۾�h3��$h����oI#`JRQ�HŠ��&�<�O�"�܃��Ц%pz�<��a����Jz$�B������=,�� �|;(khv�ҍ.��6�x����+e0w�&l����q���#SSB�B^&������I������K����i���<�9�Of    IDATx ���%����F�a�Xt����w� i��_�\�w��=�K4�Ŋ���y��З����C�l�	��fҮ��q}�tn!e��1�4<!�Z��.S�\��q��ڲ���1�����u4�/Ø^D����lFN�㹇��?�1���yga��uX�j+,N�*�24��W;=��B�Q���e+w�j����19W��'����t�H�݃��gb��5�[��|W����_>��N�!v���k�.�}��#� ���
x���T��95H���x��'���ɺ[�t��$��f!�Rf��E�L{$W@i�h��{?��+sf��`jORbe�v��h^���%l�zn�~3����6��x�ҍ-ޗY�p��ݻo��:>��n؍���:�S��W�;Y�c|�������ZZQ!�B�1N�U%q�ς;���1�MJN?Ȥ�#�ɤ�d��s�������֘��i9L�e+���@j7������E��D�5	�P٤�F6��zԡ>3�~�g2oA~�7�z�\S2�I��̅�8���Z��d���~1(�
�2P�a�>v��Ǉ�7�i���cw�E'CpbΗroQ�#�1���@��eCql��/]�Ȼ��T��Pě��~�)H�F~��bu>%�.�O�F&�z��ԍ�1�p�ȥ�@�Dw�`��z�����VQ�3e�w��������h�xVJ<�hAr�_o�T�vYe�jI��M��y��&]�ic@���Ș$$�f��q��EtvvK7��Uk4D�?Q�Q���.��8�ݤ{�4��
��SI/����8��qe��%�`�Jf҇<�lt�P�W� ��<r���h����e����t:%7_�Ѣ�)Ҧ������fvu`��E��Vĥc�pz�>�[-5ivDi��ك���5̸�z��]8yo�څ#�����sN�mڈ�W�o�l�#u�*���+�~�E\9~ZӅ���d�Ф8��d�Ӌ%�,#�!�'��p�Ǣꤊ�P8���(]�X�ۚ7�tD�$i�P�>�x�b�z�Nܰcf̞ǩ�|��݇���ޏ���y����E������#E.�m#iא!��YG��C"��H]�@`�s1긨2�X^KB��%�y$�ܜHHZ2����0W���\�T��3�0Q��r8�.?J�~6~���LG�b>�m�v4�&\�n-	,����ۯG.#}T�,x}�a��7*jB��}Q�����y�D�l"�����,궏��
&�m�������v��m;W#[0q��y<��8y��L�K��I�K&LXy�i����b�z����X�Z��lܺs#֭_�L.���x���p�����BHnn
���#�na��v�s����-�?s^c�U<vue�b�\�x�z�X�W��������������T0�'�/�̞�%_��w����Q�2����L�fN��M� �F�Z�wER����ȡ�S�Eb���e��PS4�0�t�FP��U�z�������WX�`>N�ڍ������9�B���LK%qMRGo:��LQy�'"q-�u6khq���h34}�"ڣ��F"�Q����q��A�0;S�5�"
�<�d�]��szw� ������w���cg�"�ގ��߂���M$�-�&DZOK������H��h_x`��ᑤ��q���qS�k�Bc�n�쁽x�o���aN�6�:�Rۿ������bK*=?@α1��.���`�3�K Zϲ����_ǲ�7��iE�ɴLI��'<3���֤n�<h�_��E���x�I������wc^�G·�d�Y�;���#?o`�͙���A|���p��c����}�=0,��(�H�`Rt�d���	���EW�ٲ�(��'5��a
�<�1�>̦\����K/���������K�Ga��@�����!�y�	�6n]�����܆���^7�>۰�4�_���K�4"��s�/bt�,T��tS�hř�g�I��T�Qo��/$�;�ݳf`֢%H���$�F&p��a&�i�2lk����K��m�$]��y@���U&JPF�Sg����ǫ��*��K�ʄ8�L��$�2s��5�����2 1U>�*�5����PK�:�|WZ�2��!�q�f�b���X�	Y�C$i!g��%����=�\��믽��{GPv	�b�0%g(�b��`��hZ�j��$׵�$�_&u\��!?�_��g��r�M���Ч�.���g�xS�C�Zvtt �L��j*�����+tU:I����B^dj���L �U���Qm����hg�_F���P��@e�������Q���"�% �U�\��������o`���e"$�fڔ3�M� W��҄��j�K|M�y=��?�w���B���7)Álm���ry��=���h.�DZWR�!*u�T�=$r����n�:I��f4f�L4e�����Оz(���A2��NY?}ě�R���Q'U<-P]�X�.4+��Z�B#�"R� S'��G�Q-*��ԂIx�|m��]�V�.��d��,Gbb��EC���M�F��3[@��I7P����Z��2ʕ�|�"�b./	��LAYb%L�;#��q�`Rf�9�%�+��Wn�f�#g2����!I�$(�2<�+ã/WP.Wа#M�x�+T�L��(�x����Z�=��u]�Eqޤ��!CP�@.�Do{�-�������S�|�82���"�"!0�)v�{�Æ�v"�|�l�'����#�q��i)�ް�W-ޕ�����n����9
w�	�Q�nR� �CCC��l!�d6��CLR�8������5Gڐۘr��t:vj�)V:ނ�Y>I���db�)ݹs'�m��g΄Ӛ@u�N~| G>ڇ><��:�>���`hH�5�%=2�a�L���݄٪!I�b�o�@3���b� ��YpXhkG�X� U^��PߩŽ�Gt��苋��ލ���Ǡ�"jn�����i�`�6l�"A>ӦѲ�2u����:�&���'J�4�W�\�֨� 7��@7��|��U6fz�i��Y�^���f�jM`��x��]���T�)mL�%�`�G��pS'��SM�A��xQn�m,��z������cl�͒<B�C2���'����k���!�2q��E���>�������{��~�R\�i-�͖��;�~�]������d;a�L�۔%��5+g��nCWg	.��'_ÉS#��H&K2��
zc �����\S�SA��3���������	��^V�j�w�ڰ���c�^x�e���44�馆B"�NC��tt���%�/0P'@*Ш]K�J���	і �r%�Je�c��b½`�s1�pŪa���(�L�-an�C8�$����݅�֭@��#�8��3��_�߰�FQ���ꝷ�o~���	$�$�����"�b����T�,ir�FQ/��"&���Q�3K����>�?����t����u�c�}�b���w:ň|y�F���x��?�[�?�B)����p˗���۶á+��� �$-�I�$B%Q��J0O7$�Vh��0��Id����I\>u���G8��Xb�hOkh�@i�R����E+����8�{�b�3�#��cٍ[����/\�ψ��׋����Id�"_�4�\F	�E��.I���мz������i!9:��={����?Nk�x?zn�`t`��y<�����?G&�aۭ��������hEMI*���
��\ĥ��8�S���IS�4�z�,ŴY�rY4�L��s ��J�f�x��&�b�r?.]<��D?j�AI6�9kV�Z�� ��P��4Ġ'b2#�
i��8s��}�Y���;R�/X�@�?���y��iRӋ}).��j�:��!�n�w(x�R��&�Ӫbt��aK��{֮���^	%��K
R9��>�9\�x/��:��y�;*
��I�l��.�G'�Z�$M���'���=_%��m7���N�����I��8Q�Nm�!�)���uk��V��<����R��z]��6��9���$���T��)�Ԝ�y��r�������31R����'q��q\�<(�7��F�h$���G*rgc�ɬk�c�捸��;�x��H��)����$mJNEI�R-[|#�e����'�l�ŵ��󷎏��c�V��oȂj�Z��Hk^x9T��k�@����@6=�P�����c���?IK�rzą�g/�ވ�f�dR "�pFa��7��)[<�d�w#'����O2�&"]��P�o_��������%���Ϥ-�~�7d&��dAZ\�����g�u��X�{���r"!��zu��j�jl�W��5���1��I��E��B$�e3�55�
()P��ӃL�ŹC'uvUH�i
5���A��xU@5-˃���l%2f����Ms�!AL�t��S�"n,��
��bXזP6�D��z>��m%��
�F�`�-�]YW�b>�kC߲UX�y�߀�+�A/�141���aq�Y��ci�=��v���~�&�N��a��Q9����Ph6blx��/]s1N��#�p
����DKm�-+�w)�7�6U�^"��@u+V��w�)�`Z�ح1L\������㣽GPih����t��-��YvT\F���݀�j@W�F)�[�����
erCI���J�vq��
�;��#��Ԃm�@�OW��H1G }�}�Y^ѧ'S�=���4E&n,>D�%�d�2�\�@gg
mmI���bUIK=qJ�e}���ν(%��ޘ�)��I�P�����Rɜ�7�#8��y�?zA� ��*ft�[=w�yzz��|eo�j/~��*mm3T�KW�H�KΰP�H1�4d̴l�Ǻn�m��㖍螖���+���C�/�w�`���B8�	`a_�ڹ}s;�XU|t� �;��:��{��ׇukWc��Yé��p��	|r�M[�+�&E|��Y�h3q��[p���l�����c�al�:ٙ0:G)װ���� D͜�ȏ���T��,'m	���ς�S?bm�|M&��T�Я�@�:*����G��¼�����sx�?�fT�X�ϡ�y�$u,���1ak:a�a��1��q�F�QE��L阝-`z�:&��P�u��j�[�ji!�M70'߆�"4OG3�E~�Z�=x�j���؉��������!a9(v�c����o~f�<���qM���K�\���x~(��a�L�uv�5b���8��C��Fg?�o��'9v=�aC����߆m_�Js���9�#�A��G'���^~�ad�	�Z�;��%,�n�|7\�ژ�b��뜶��æZd�*�윞2&[0�����n��l�h^�K?�!>�$�6��	Դ ���q���kt/_�)�c�?��gC޽�%�֡�����%��:6�)���j�!�S�1#���Q]e�(�.�(�$�ǰK�ى
*{�b�ŗ0t��i���G�M�r31v|�>�4����U\{�:|�ۿ�k6�95�M|���*ch��p��Ia����>M�Vgh�����t
텂$eW+�UǤ�0RR�$�E�K�nx��� ��K<�o`ƌ�X��.A��-�]��BX�������܅x��g��o�=�z�z�wIG�k�A����LX]�����Eܓy�MR��%9t�#p0�ܩ�<x�;�EK���7cݚ�
h�IG4�?�C�K_}:y�������w�S�a<�ء/�ڑN��HhR����%�� �P��L!)t���ߓ� ��:'��hw���U�Ť�2kN	WPSf	u-'�BI��Ο/r��h�m{GIB��f*:[0�51H�A#S�0Ӱ� �.
El`pX��_�I�ǆ;�̼f\3��q�4o��Ϟ=[�l�u�C��hY�h��ꩠ@���� �+�M�k��	�+�K�������?X�^�w���I���A�1-F�v�텛���x��!@=�ы59����[;�DB?��x���ߧ~]Pb��*�Y�����<�y���4�镣Ix�J�@�)��K���(�#�����&���*�L��iD
� ���t�q!,dL_�5�#ɜS��(�x�~�����H3��� D��p�m{����O5M30C0�ϼ¦�=���ĤkA�q�|��2|��l]]�r9��"�.D��#�h�<:����qe�څ��W���JڐZ�|�u�5Da��6��k�ը��QѼ"ʈNT�����,���4�L#N%��$�b�F��DH
����Xg`fK�_3sV���[�cٖ�0�9�t_J������Ñ��*�=X@zJ��'�sR¡�XOo/OP�R��Қ2�=M~&'�QyPO����4:�/+
z�W����%�>v�R)S��;����oD���h��0|�Ν8���c���Qc�X�#���y� tp+P`	(��&`����$��	5X��]��>Z!`˒�5#�4�l���%7���}���n#5i��R����$������Y�	Q�6�RĪ�.�q�����{n��z�
�3E`J�Ӳ��١g�L�3+�9���f?�"�"��ZN#�=���ًG���-,����;���-+ADz��1���>��0��(Q���c�"<����#e��2�޳Qțx�s�`��H$\<|O=�[��)�G>Z��:���aۖո��uH$l�NU��Jņ�Σk�L��%�*cߞ8r�$�䗦�Sp(��走n�b<x����j�D��7�؅W^���G2�)b5]����}�d"p��:�i.<Ԕ�$*�#0�?�]����>�4�h[��q+��Ѥ��w�|�����o�f�{�5<����a,�d��C_Q�h<��Qv���{��F���Mq(s،Bt�L��ГL���{��|� �Dȟ�c�gh�����b;z9�N�f:�;�#����E@���k�#|��s��2���qn��o"5,#���C��.ܨ��N�F]B����m��<N�=E	�MRK�U���^��a��>�������}6��d�Y�Ұ�m�v�����O~�_=�(R��o݌���E,�r�b�DQ�,%��S��rJ�~�f�L-X(E����N,���_I/�k?�;�}�t��(%54�m�
����A/]~�����>�<�ڬa,ں���+��	Sh0�C&(!<�z�*�XR�_~H�	_/�5����_5�t�nc��D�a�6r����g�G���p�}���>t��
�9��W��SO�'?�z�޶_����M�faP�'�	����)�2Ư�ܙ��Up�-� S�c�Z���8.\��f�!Tٞ�v��lV�4�f�"gN���L�Їu��
j�2*�10p����^�u�7a��e�<k�����D	��$����O��_a���[�9�N{����h[MyO���\N�2�;'
R�r�@�QUf���ΐ@��I��a���m�mX�b2�.����+O3�#�M�¼�����C����\)��Sٛ�ud���gjH&����'����.J�vd3y�yH��D�M"�gq�F�:�tZjaR�˝�B�cyBO���6nP�{�̍3�x�
�h����ݚ�y�3��);U�ߏ��R�ӌ�agRKŨ^�Р�nJ3��h\W"���I�)q|M�6�<	�FU�=���}R5!YmĠ@�O��':��0�\��������_lI:00�Zó� �x��0�����zAW�{m����RfhI?�!e�����5�+f�x�i@U�$�J���ATby#/P�&��Ò?0�P�e��%�_z2h�tC�	a�l{�H
�6�;��bV09A�2n#|�nh���ԬC~���O�S����lT��W�i�.�)��R��m_�$�I��=N�8g�@F��-C׭�!�� �A�g� LZ"d����\?p}/��.u������>)Ja��v���l��m���x�V�~�e�6%4=��`v]��Ʌ�Q���G9�-ctl\&�*�զ���k�x�S��I���({v�Au}n ;��<�
���x�s�.�ՊX�ykč    IDAT�M%�;c�mK@��4�1��	}M:�<�3�z�d�:l��v,\�Ll�t����	�~|���~����?\�i����!,�I:)C���s@t� �(-P�%#��dJ����UFt�����f��Bs�5j����T�V��i�W�P�u��6Vs#����'����#8p��-a��&�����)��	
�5��[B1P���@�e1T<����=G�t�b�f�@mIrR��_
b�!y�#�xAG|�O�{4�����3v��B��X�$��'[=W�Z�[oތk�]�ZyH2X8��eRX�8�4ET�cl�)JnB72�k�܍���7����
�.A�6,½wm��s0<<��_|{>8�j0���}q��.Fw 3@̿���u��I��j"aj�V��x7���D�6���Wv�a �D��m�w-�����7\��+�"�jBEgl�1�d8R
͆���A�?}	N�Zi���Lf�q��S��l\�7o�"!�C�ؿ��ͤei����Q˵�l�Nf9�W�ڮjdR��2
�QA������
W'F�)�5`q6'�x_:6�zM
'O�r�Z|���6�^���w�?��.\��DB
���M&hВ׶1j50Ns߁M�j�#Э���\3sy���@=�Q%(����	��>:a`N��3��RMf0�����>`�b ݅��ǅ����#�4�l�wތ{緑_�n2�����~(|x���Mg�W�x#���+�@�c�-G������ǿ�]�ڳ���t.^"nG}7�7�7Q�����8ξ��}�1�՛HdM�]�;��y,ڶzG�d?=��Fo�L�侌�Q{U�9�S��1h�L�ّp��������r�a�M�f �7�ǎ��C��_=U���~�~�!�F�r�&�,Z)4��B�y<�/\�(^3�SC%@6�}7�I�u�̜G�?������h;p���ŧ����}�sV�{:��
0c1p��]/���}�?�ֺ�ͷ�����0�&�)6h�е�H���Ȑ8�_Dӱq�m�Jn
��y�^8{�j�L��m��V�t��mՑ�e$�g+!�h6\4+��\��	jC�;��7l����#P@(��2fN�ˤ��e�k���g�{'O�ļ�����D)�2����*,,�	�YRD���2?acOip��Ơ�JC�x����-��[wތ5�� [�dx�����ӱ)-�m׮w�>,�!�j=r�s� &�R	e�ş�A�R)���N̚� �|Q��K[G�BF��dB�X����443��k?C1[x�)�!7-ݩ�Q�!��E@�P���C�["�
6�x]RY�0��sR{:Y'�AC����9�d���8�G�.Q"2br���	�[3���J/AM/��z,�Q�D>�;cG�x��-:��4~6W�n�c���/�WD-"sdd$���d�Lh�i]�?L����i��z�Ȫ�9/L�=M���fQ�$e0R�oP�9��<�e��t_�<u����`���{����O6ͫi��'a��=�WO#GTsA���w]��2�65�2l�pLÎ�T*RKXW�|� �����$���Dz^�l���A:�SZÌ�����д���&0A�
++��B��~/��Фm�w2?W�xvggD���9���j�xe�Ҷ�Ǐ�{�s�Jg���8p2�����Ar���S���uWuu7��}�E�A��M�&%J�Hzl�w|����:��u�a{�㝍���X_cˇ,[E��xS�-�$ �q�h�Y�uWV����evaͯ�-M;A��]W~�}��>}r�����@�-�F��͈],a�6�%C#�F!�jXdqAsB�U�wwS�&�x"��L�Ie���!}(7ЗL"ύ��-Y�4%���!�	���,���,ݰ��S
����$6*�B?z���(�qd�~ۻc��`��8Z���8��5�|-��q���N�0R	�Ve�B��w%[;%NUKG
ܠ)�@�@,�8��X�7X	n�k���'ܲyx�ع�6�/���2uf�)8x���蜦��73�cK3Ŷ�ۘ[D��X�J�4�)h�G��.��2]ĵ#*�-79A
z(6�(��@�}��ŧ6������g9��������E�07L��ǔϔ�@��+:�F��I��曗����ՋQ��':��g���Rhї<4�� p���j���:H-roϓzs�:i
q��6v߾w�\'�+���7���: �:��P@�D�<FNj��"3"�kK
���m]�tJ�M��;~Q��'C�����M�z�2��Pb�F˪(Ѣ�����&<�f����6�i��;C1��5Qp�Â�:�թy�/�0З��n�Yo�T��Xn#B�T-��e\[]���Z�q%Q���#���1t���)�g9G��h�R8�ύh�c�D�F��p6n���o�܂�;���?�S��*�{�x,�H<+���>�n��j���������➏|��i���f���ѱ��l$h
:L]���k�%{�v}�iv�D�H�M7�8�|����/��o<�QG�Ա��=��/��6n�Gz �
��"�8��s儗7O���<����|1@��P��m6m�1��]|�+�3~��kQ,�i���B��]hEL�fV�sǃ3>�C�|�^x׏��0�u=�|�3X{����B3�V��
+f�N۶�
YPz5R��'�J�����ۙdi#��1�}�i�|�U$��H�5h�=X�{'��W��؂a���w?�޿�*��+�rǭ���#���h���F�wVǕ����Z{��(�n��e�����<�#� �b����#C.9=�}�k�<��)k�=�>� �{�-���._?�[�߄����c����ZVL*�J�"�Sb�=9~�F1���=��W	~bb�N����@��>�8�+�LO>�� ��O�㙰��Ѕ+�i�f.a���.����⦵H�z��!��	8�����t�����Cx�ŗ��o�9M�֍H��#ic�P��s��[<�B)�
p"�t�r��hQSHh��2?�<�Vc������¶�w W���_&�
��������_y
ǎ�D�R6uc.'�O��6bQ�u��˗b�=�c��0������d��)���O����iZ��9���\!E�^q(����Q���L2�~>pY��FBX9 ���,R��lBB�	o��쬼"�D�I�k�����2Ǝ*
2�{��Uu��Bmw�wC��+��W��5*��8�
m?���R���Dc7��|1�bS��?�����8���7}�k_���+��������a����V�x�z>9�
����"��� �H,6�FD�_����(��D�^U�;M��eق""����Q���lgR	�X�ߏ|��Ջ�p��Y���ҿ/�}��	l�c��Y%�w���p��wQ�>�L�C˗J*f���+�=y�܇מ����*akm-
W��2F� 	�z>3��MP�ٽ�DK��ڢ
�`���|K�!��8,9
M��#\zVʓ8�4�)���) R�n�暂S����Aj
(4��\F�y����
p3:6L:sx��-	P��~���+A]�=�5!ɦs����$8_��>�.t8Y
7ǰ���Ǎ,�w����(�����e�G��Q���m���������,�
d2&�VS����I3Jq!�* �H��d�i�JH�5L� η� ��Z0Ry	@K��\9��4�UL��05�B�Nc�t^�!�M]�׆�fZ�I����ˤ�Xq3�L��L�Ƥ��(WZ0�iq�؎9V[4&����;"�W�x�M��W/�թ��N*��QHC��@Y�W^��%�A~	bB>�Oj�j^��л��G�v�	JQ���z�����������:��E�8��j@3�^A����b=�C��رq�C�p��_����b1dAm��f�Aٵ0�jK���HC`\[z��s��x��Y�*�أ����`:�и��a�����|M����ܴ6�6�|��u���W������,"���م��ʯ`h� AG3�7�k!dw6B��Ae��ȩM�@w�`A�����:h�O�ҁp��0��1Ԯ_BV7#�-Y��?���s�x
$�#�0��q���Sx��1u�8bI���b����{�@��a� F2���U6����G�������t�!8�� ��>�П�_��~�Zc��q-$3bC����=���?���44���O?��l��>�� �>��_N������rQ�/�+ʁ�hThY��J�������>��������=/9����ދ���[�z{/��O�����V����-�oC�����q\�<��W�p��5�\'�-��oh �>� ��n�{�P�)����^���}���$Ӕ�'`Yu�rC#bIE
������1q�2�e�
�P�Nc��ܲi3VߴN܇H�=���Z��IL�SX�_�|M�*�=s^�WH��?e��#�M��.N�?L&���)�1ec�l�
-3|/�r�-8�4k�^��]�܁͛v"�;,{�e3d���F�Ajcb�ͧ����Z(A�;m8v���&�z�N�a�Л�m;oǓ?�\׏�ٶ��L_���U(�(��,B{��	2D��}jn�����ex�1	4�b��e�����$v܁�NHA"O@�UF8A�N��@k;���MP�Oe�s�*nZW�i6�O5xR���PU�A��;o��G�����l�R������Ƕ|��yaG�{a�?���������Tԋ��Ր"�Bf:��ȔEQ2����'.6NtYa��|�p�
�ʹiI>�o
���f��,�j���	L���n6���3	��;�ތ�B�O�����֪B#�蛓��{n����t�J��Ӹz�8���6�N�Bk���T�B�oی�{nG���@2����_��_��2i��#֜��Xh�/N,A���?�oMAj���,�N��J�US�F@lЂ,��㤾�v�
r8@Φ��lTM��044�]F�����<xD��r�GGO#������z�j�����t��y�Fu�f4��	��	6�He�F�HA��#9��G��n8�{5�sR01	UX]a0]���˲TP)NB���!�^�4I�*�6�j�J+;��hpܖ�3������l_��I1@1'��s~�!'^	��2<J�g��MэT�ed3	��8U��4��I �����)ѕf� ��8�Q��MY ]
���eC�b����M���i���6�xJ���bt/!��N#��\���Q@�7N�����e��*�w���F�"���y�A�aȺbȵj��r}���G6(��n1�	�)�^BRJ瑄�� �7��kL�x�ǃ�M[6:�b�m��e��_��ں8{W�}����(�lZ3��ma�U�T�.Z���A�C�u��hu۲��}��XTȣ/�����"q=��6ƭ2�^[ЋA?�E�<F�����[�}�}ږm��Eu����U<���V�-�a�����_�E�2��Mmr�d9��S��4&�
2�z7%�Q�!����\<q��՗�ދ�c@א�v`F\�Z���p��Ob�C�@�ЏY�+x1�������_���CH�X������p��@6'�[����x햸�q_ac �j���
5 -���8^y�%<�ԷQ�>�l"-������� �������_�d�u��c�w���p�ƛ��{�ظA�nU8
��@x" �t�qK�lO�i�n��$�����"��o1�ȩ����;{q�{��z��)`�}wb��'�������������W��b�͋QX8��N��`zz�rV��>>_�-!4�|�n^���
BNTNR�c&�Ɍ��j�Yg&�u�d�A��W܄x��cb����G�De�*,�,��7�]�;�܍��l���!��W'r��D,L*�s���*�����SB7s%�1p���q]�45��λ�c��h���+h4Z���K���.�D��7*p�����wݎu7oC2[�!#�?1���H��p>參��ܳ��رӨ2Q[h:�&R�µ��e�^�ic��ex�����'~
�G��\oZ�{I�a^w��WJaS��ܩ³�{����V��9��p�0U�qp�� ǨT?��P�/u����Ĺ�C��0Gռ*�~E6�P,�Txgx�*}��-���s���;�B�iT#��'A=�����H���Le~?�3�{�\��ߪ>o4����R?~��O������?�Η�|�"�`�,iÄ�h�j��5t$rY�im�L�8r�8�S��f]�I16\����"F-Z%�a`#�c�2c��VA�^�}6iS�MKc(�G��8�;�V���ǈb�έ����$������c�Q;��,
�ËA'd8R@��5ذ�v�Gp��	��ƻ8w�
�M31�$���~�����9�0-�Y�.&�����S�j�bO��A�զY4�Z��@6�����D�%�.H�=�݇m;w`�%��p��!�]8)M��c�0Y��A
8��OqH�)9)DdZUhs ����E����u��.)�1�q�K�)(� �J��`rCA�k��G��5ܴB�-�qý1!7D�N�LL�D��@)�!R�#ְ
��;�lҾX��$�`I��B*�F�=�*�5�f!�x��@$>���h�llXvK��<�]ɑ`��%��/:&��}���-ЄBl�"��,
QAx(P�W۲�B�mwT�ɟ�2}��P��J�%�?�Mbv�(ᄜ��c#/�fYޫ�'$m�0)V�b>l�T����)�4D�x�(���Ix��A��l:�`�t"6�E$-����Z���]���ћp���w��<"B�g�8�K�v��YE�n`݆�����7�c�V��L~�{�~�mqM�Zh�DZ(�MT(��<�Y��&��4}z]C!a kr��2I�4���r(�-D�j&F���,@�H��%�Z�C��̙\k㝿����~��D2����x��'���;`�r��\[�+����>l){�hZ���]�=�SHes�tl���;��^<�����#��>��'�18������>�i	Tk��%��'��Ѷq����������}=X�c�>pVl���~v��-��X,�Dܬ��I��g#rc���W2����Sx����bE�|h�k3����\��#���{���O"�`^˅��`�<������ￎх޾I2�ق�&���i�Z+�'��G$'�!Sap��k�͢a���f^��t,%�v<��f�h�]ǥ}�<w��$��(V�w��g��!2���7��w���ԑ�̂��� 7���9��1An:�M��`�`�S�T.+�����Zzv}Vrdt�L!5�P�bh�nڸ	+7o���U�p�������֛�bv�:X+g3��M���ǟ��[� ��G��D��rF�7�6�����L$�G�a�r����Bu�0=M��~��д-��h���p��9Y�K�,>?�2��4�Uxn��f�k��ظ�Vdz�e����� ]�"�0���><}/��N���ZSޞג�?��@��]�s�6m���}~ⓟA�cbb��R�!�C�j���C=��7A��sq�Tׄ���N$6�h7���ϲY�޿ԙ����G��E�Lirz��9wΠq��6��!�%�9�VF5���_�:���
�#
Z���l�`a1�����h��) **�e�K�������)�g���������ۿ�g?x��G��v"��K3 y����x��7�v���w��|
�,7NV���)�@hr:(~lx��PS8]W��O�,��Hgk�Ѩ��X-$�r�zi=���5[D���@��`b�1"�/Ω�Y8�(���W������R��f����W.�����tW'��<Ŷ�I
�H��=Ĩ��G�U��h&IkR����@E�RЪ*XY���u�Z�H$9'�*9[%�!��"4��n�}<�;o���(�V	�����u=S    IDAT�� }�����)�D���A�-�'9�ؑ�\Ku�d9��hhu �m#���j
���F~0�baS��7�y83��I�/�nl
~��qG ����my���&����ꊪ	S�AB���"��rr1��3�����a�g	
�!����|-��p��xUu8v�J,,HӲ�e8I����SCU��|&�v}
�U��"���P�F�������7�L���8���/H}�i�g��U��'����Q�"�	"(<�I�c�K8yQ���`Ǡq��+��K"{P���� S�3��P��f��!���!d����&-�����~V]����o0Z���&&v��S�hG�?��	k֮.]�ī����}�Zu���Z��L�뼟��8��>Qw}$}�z����X)N��>ⴂ�ˊ�܇���95̸-�\6�hD�4�E=`I8�����지��%$�n1�~���z
�FE�BC���vap�
)y���e4jexß<�$����~X	�9���C��,"	f�k6yeWN����hLO�ɐ��ψ �d��ރ��n���s�(�-ɨ1��ً�q���p���q��^,�p3��,��ʢVkHN�֠]��2C�V�|nf�p�P�c;���|�PE:t�4託�(OL�2=���F����G0�n�7�G,�Fĉ ���&����Cb=�Bbx�4�CN�B�\��3�CO�w�>��$����+W�b9�h[R�Q�I�����t>/�4�T��铰���5'�ױp�F�nF�L�t�2�{�%���S�M]�n��G<��h�=�T<%�RV��ٙ*�*Ē���q.C�lG�6$�^�J����h_oC#�^��۶c��w�H��U�p��<��x��WP������a�J<��Oa������ͧ��qy���S*�8N0��^9��� <�d0�P~��PN6~:�Ç����\PG�6�h'Œt���6lڴ=��#�7|A��`n�� X�ƱO�W�Ĺ��G��rh�@�QA�MI�8Mh�:z�֯]��o�=��H3�j�(�PR:5��E�K�^P�W5lR����
��*����NE�X~���}�A�á`�ϳ��Ϲ��N�؂�a.7Km�y����E��$���5�����&�U�89�xV�ӏd��x������Ǡ4�ѽ�$��o��~�����V��$�(��Tr�B�!}�t���=��0	���1��R\q���"ŕ���M�Rh�B�,����2��_��Y���B�0�4c�3N�饎��-��6nr����@a�_���Rq�G���l
b�yLMfc@Ո�nh(zIu�	��<� &�f��Ou`�ٱg��,oN���υ�t�t��~���&|�rSIԜ�p�v�
�p� �b'�l۱>�	l۾C�h�f0s�.�>&H��g0U��j,&R�Z��&B�|H��!�nJSu�����ii+A�00C��eJTI
���V�v>�/l��Ʀ�w7B�M5������Dq��.K��1�qRL�h��I���Z �Ҳ8�nKz��1�<�*��`OQ�� d�"ŋM�;�u�ȞytǢ{'�t"��$M��Z���U�S� �C��"�G�� ���%��d󎅸�IzT�����g��� e&�}Q�B�/3;(�c� ׭�2I����biò+H%c�100$��1�8�S�qCa�|�Q��yJ�"z�@���s�BCțHLw6}r.4�pJ<��4�t�ᣇ�/��s�K[�[��պ��i5��ΠQ�A2a��O~O|��X�h1p�.��}�N�73�ri���P��lԃ�J�#pڝ���i:FS9�q�8dB�X�F`�DL�m���*�P�C��E�0�X�7(�3	�GG�����v�ťxiSW���6��v�,D5Z+�R"��k�!�ļ%���<��kv���N�����I5���m�b�u̌��:[�!��B��>����	��Zf��*X��%8�����tON,>-�C�C��ZB�L�b�A�@��R{�4�~�\�x�BA
t"_�z��
�j�l��)d�si��4l�6gḾW)�Ӯ¥��D�M������$�S��Q��7�	x���c2sF�U`���
����JXezn�M��N��~�{����;���_^~Ɉ�d��3���oB�zJ�vZ���+�)�E�Ȥ��2`ju\����;[�C2W(��#Y8�E���n�,ߺ��xv=�o|�i����ЬM+w�y�J<�ēر�d
��6-�Ӆ�/�V�p�&MQ��\$�̙k
橭��*~C�*�#�#QqPb^����o��&eS��ğT���)X��w�s;�lٍ����8<Y��t���~|���x��w$Č��^�j�U*��[MD\F���+V�b�֭x��DDϣ�p�p��@�Q5
߳	�'(��@OQ���\��Dt�ί�aV׹(L��VҮ��J�{�>v��{A,��RE�ь�~���92��%���+��_lc��_a*HN�"$)�����CL4�D�d*��d����>����d��/?��_}��w��)f�X&�E"�`�i��1�)t�N9,��DJM�y���"S7�*|Y`�N�)��) Ն�ӎ���h�P+�ѬU�	$ah�X�De�րS��o�HF�$74�w		Ac�cj���m9�����L:+nb���X��)�p�O��d�0�F!�.��9I&��b:��	%��jI�	�R�8�VZUqB�Im 0
��m�h�.�M7&r���ijرcz�غc����E�N�¹�Gp|���4--t61�unl
"L2���Lk�ѱ=��jЇ��i�M3����|_�lr=yi
�=l���P��n�a�nX�a�u(�����pS����ki
�/r�;�w*W">�d���"H|T9���t�[���c3��E�ijZd]˵c�0��-��I�
����Z���9	l5�&���%��g����nwP)7qmlB�jS�N~s�EO:��KF������$N�:/E���%���q��3�t�8��G��QwOd���j�%l��R�M��<؛X�|�.]�ёEb���b�|y����xQ�q�w
[��.�+TP��,X�кQ��9�W����ݜC�¦/��a�'�A���S����h@�%�IuO�U�<_v�9T�����n#R+�Z�D*�O~�s�̓Ob�Ћ�ɓ8����Ջ�&��R)���t0�QMI_?�E!�@���@"��ߤ�p�bé��H^�t���fC�˚y�8��bH�PHea�I败]��]wB�};0�DT�>�sY@dG~yL��`�k�Ḗ�?R�tr�9S��ƥg���C�`z��]0�/��5kցVhY ������;#T�P�R��I�)v��NJ+��13 K��DO��b���,�PUf4:��"����GZ��ϒ���;�t��Lm�k�6l:���>a/�5�9@�R�k߃'=Z��XLx��c�ي
���m2��CAD�'^������ k��E���_�g�����ó��8�֫�D�;R��~�Dѕ�s]<�Nz��n�Ǖ)dO�aQ��l�\��T���Ԍ�������h?��122 M���wR�qt=r
O��ׅ>�X�1�L�֯�g[o݉L��6�
��8?,6yQzLP�q�Y�v���}Z�q��9�:ga͜6�f�N�'#��LG���P��ϝŒ�����=زur�	�fO�&��*��c'N�� M�4l:�,4�z���	3�B!�X:�-[�IS����.������$œ�(xn�
�m2 	S�װp'�Aro��p`��	�Yr �5v�apn�9��|����� W#@��:A�>��������p�Ns��9��bR��ɡ\���e_�DE�����jn2��b27�qS�#���O���������/��� Փ'4�x"�L&Ğ{�̍s��O���V�0(��]aD��UY\���+��
��oL�gDHɹk��$���8c{h�jJ`��A�}�cj	˲X2�	�My&�&5�"���!��i��70�l�]�>��x
M���
�_�� b��&�?7Y�d��!|{*�P��σ�7j�)���X�^s�0��D� a�����m�n�>��۶JxY�9���9���0��� ��PSКK4&��$�l��oN��<�bNAnˁow��
�m�Qx�7�t�B�\|�_"���yI4�g�p�}�)�d�B�&�˃^
�.�񍈁�
��n�5,<e�T����ɩ\�����s��"����Ą�*XTh"�ǚJ&&em�Pt��X>�o%ò��Էq��|;-C�-Z<��|�>�R�X�m��pa'��eM��=��mWb���p�b���~|���!a�b�:,^���p��p�_&�Ͽ�N��]W"�T��Q��]���X�|��{'F�̙8{�����G����8y�
N�>�Dڔ	��*�"W��N޿�H�g�)0$c!Bw11�v�9����=�8��*�ix��:��9������\G�cwS0����L���c��W+h��ͤ�ēO�ǟD_:�����g����5A��-"G*F�j��v騆f#��|���]r�UnK���V[�۴U(P�(��Do2-I�z�Hj��QDn��;�nZ�D�,RYp6�G��]
i��pA��$ѓ-�ᐃF�:�wY�2������
�7�0��S{>��1U�K�k:m��&�ZCm�$�������OT\ݤ�!����>����zM��K}	�l4Us���ا�'icL�(��{L�h�9"ڒ ���E,�I!�a�B	I�T�Tۨf�D}�+��:��7m`#C�c�ό�'�Y���@�A���Ɗ���^G�m�E&�Wt.~�����8� ��|����gq��ah�'������$�������P��z��&M��%�EB�q1],���Z�E},�cxd K��b���y�n	�l7|���y�[x����)�u�͓>���ܓظe+R�>4�6��U"��L��R��`bݽo�X�
 ���s�T�5��D�(m�)�&u���{��]��;�g���]��m�hy��vl�t��B{�r�kg1/&MÃ�����^���gQ��a���
�we��k݀�0������ؾ�V<�ɟD,^@���^��	��*�*p�
��
U��t8�S�7֪τB^�36�9�T³�sP>{ʵ�w��Bܑ ^E���n�`~(��8�s���HA �s�ý]=G��㐇?'�U+�JB�v���=���!+�G��:��?Hd��c>�W^�?��c��p��~�����f�׾��w����=�"�'_PV��P�vs�YE��J�V�4���&�a�v8��{!AA��H�l�.TJEt��L�L�x.4ڝ�<����s�b�ЀEe~$�CmMm��z�@��c0��܊���<L:&m3�����8��z�y�(H��f�(*rD�L�9Yd
�O�Z�Q��7��H:sn̤;JO�M�BS�界G�u�V<���e���,�mU�)�p���;���tC��t3/Z"��9cS�����:4�.!mtHa�q�) <ӄ�L`��B�����*!V.����ɛb=�߰Ã�{�.���B�Am������Gy8�T�{z#�ΰUN#s(U0y��L�p<^�6�tDD�&V&>򼁳��c]�vZ�i>FFz�j�B�\�9������8|�,���>����Œ��8q��\�D2��K�xat���'�e�r�Z�ã#8r���̋�t��"��cb�
��,n�m�� N�:���;=���ŵP��K�`*H�5|��{�6t���;{S�0tSܼ�N�E����*�@�>�D^9~PHO�VW�e޽�x�4_�O�1Q����`�	�'��S�#:�-�J��� (� �{�ux�J@_'_�O��Z�K3h�Π���sO<�Ǟ�)���8��x�����0�t&yRkBG�G�e@Yو&��@<�|�@B�xl�}��8�(Z�J�
�uq?��z���D��u$��o2$�^3~
�L���mڊ��[��ʴ�Y��{��l��\�2T1
=^5��w,K
��9�qS�R�v6St�����7SI� ��1`��;r�;vEr=x&'&0{}R����V#���-�kרg��9�,�^}���/Sƶ#9�=Nf(�J��F�,�{r�c�pZ�2գg��N�T~Nʘ�)D���,�"��l6'~�n[�6�N��h�*�e�e�z:/�V�+ "D�y����3�4OZIs�c��'�٩7s:�#��]"%�!o��-�cm6��So�P.N�����UL^:�ZD<�@��06��7�B����I���(7P.�0v�ff�pe|3�r�0���<slx$��3)�C�X�b1�nق՛oE���jEp�����ؿo/*�1I�/���f�*|�ǰ��������J@�w�4��6��v�J�������(�e6A��F�M���<[��KW��/b@]A2�R�;-�k%4�M�;wa��[��Y -;YAi�I�2f�u|���A|�ￅ����li���r�S�E��׆F��V�`�m��Ǟ��\��C6�[1xl�I?��BݐG�� U�0+!rH]ì���M�c�A	�D8�k9O�������P�T�c�FC�8�^�Fj�ن�x��
��
�P�L�"�tn�h��#MA�ܕ�j8�t9��YLԣ��A��pS�����������1~������O�w�]�ݓ��
}R��J؎��Lٔ\P��B��Rl��8��sA��|\�w�'�|������6���.��Ч/9�>>Ŝ��=�v�J��A"�բ�2_�����Hy����7�c��Hj
�Ly>��mL�@S���S��Du�]uz������O�&���7�_n�?L�%QD�ʹh�)P��*Օ�nT�F&G�_	3"M���ߋM۶bxxN�.M��s����޾C��#�]��!](1�L�i1)�L�.�D�6�vK�/D�XXT��t��&']MA6��� ����eb�c�}��i�<D�=y�+\�B2t|��w�a�N�����M�cn�s�DWXZ���QAQ��>$i b�����cb'*7]U+�iZ��s�q[H$"H%��)�[�B�4^yu/��?!����k׭����q���c7�H�y$=RL�1�3�ذ�&�4����0ꖋ�_x����Q�m�Q�N`��EX�a5ff�8t�4<;%CTI�֘�����f��+cǶ-8���� �I��TR1ˡ����D(�iR��nA9ƨ�@��7)���A��Xh���񀕆7�	"L����>i��6'ğנ�!�<�6��5&�.
�5N����$Z�����Ѓ���,]���x���?B���R j���u������Ƥ�47KҦ���B���j�F�c��n`�j�as������X�z�II8��s
L-�����z��苖C���Hh�K��v^��TTCڈ#�%�:i��0�qY/v�!�*��B��w�"�+�;,��/A[FR��LCI�q�Y���G���~ij��q�TiQ�VJ��5q[�n�X��:�p��6�aR�	d�4�,Z�T*���,D�l
8��04ih|�{SId
y��gk��)�b��F�saq$�&�f�Ae�C ���ԭiЌ2y'�����(�O©��וMv�D�'=�+��)3.M�]��U*¯���a3�I!���5���6S�33+z1#H�.���Iz����U�-�133���W�l�%�q>����1�q>�s���;bix��$�Ƈ4D�/�>�C��ȱ��4��ē��Q��&�ԓ���G��x"��y�.[�E7�G2� �$P���̉�8q�Ʈ��l�2���}�]�y�d�HSRB_�&z��#Ё��*�Q�о��uPA�.S�@p��>    IDAT�J��*�H�z��vp��%<��8��i�s9ѥ��n�Q�B�6���n߽�l�)Mߤ���@4Cq���<�/������o�^QM�$�=���`�w)�$�X�|;w܊O=�9�	6��p�#�.�������,������*U(ۜk���T��y���D�����!�N�Y� y����8����RM��G\��P�M�����e.�!l
$?A�O@_
�A� ��h<�9+�3�4r�ZE5^:���Df�k
~��������w�}arl�vK�j#G�<m7����-�'"�dW8�C:\r���s'��Y|�M�<�������2\��5v�VS�CI'
C�3�+mW�MK�1P�+�c��Md|�@���a$n`PcH��V4�	������`��Z�@�aUf >@��툎��J��i�WW����tf*J �Ѯ2����N9�1�Z�s�~n��e�o쑊�}�fA
6m݆�Q8v��3�v�,�?��{��dM&G�I���ж���+��M�
��Kۄ�=��I�1A�D�"�F2������$2�h�����s�$q~C����+762��j
���°�i)A��ZЕ l &�+ XR3!AJ&�b�isMx�̞������U
z}z��O�صk��|�Wq��)q��Z�q�Vl�q���WQ,��{б�{�F� ����ߏ#��BT�qӚ5�5�|������i���Fi�ap$���>�9}�Ύ�jP�iµ[H�Z2Aaq��8nݹM��o���W�Ȥ�D�� ����,kJd�#� 
�,�׉lN�����������٫�UX؋�58��p�)@�/�R �
'g�kj��H8bJǦ�����IiR���.vܶ��뿉u�����w���󇨞8��A�k\=ɬ���tI�	��=��X%���vE��J��h�/�|Ӊ Ӊ`��`8_@6�iy��^A���^�L���Df�:�FF�2�9}�����a��%X6��X\�_D4�`"6�*3eX�L@�,�Xf&#�T{��E�XDifJ��j��Dmχa��j�p��q\?w�l�#CH�SB�#2�;Ћ�k� �U�����2]��esH�q!�`:�'�4�`c�y.�#�@��A,*� ��
��2�i9jDS�۬�0bq��M�&�u��a.JF��SzL5,L;>Jק�Vj�3�/a���C�f`�0�)�I�J3�g�iX�Xlfs�SI�	C��U'�ј��{&h��s�dR��R���tQ^��'��U��q�2�p#-4�������_�_1��Aɤ��2*�E	I������������U��ƍ)⴫n�Ȧ3X�hX�*��/K#B:c:�C�¥�Т�wP��������b��~K�/7nނ��oVMӪ#��)�ЈB.P'(Y}&���_	Rܷ� ��3Q�;��X4����
4�x�^x�%�8qRrn�H��X���٘��p��6lG.�/6��%�u�"z\D���~�kx�ͷP*��0��i�������?Ҁ���tq?�mچGeS0�r�C��4{�5����z��x���Q�ǅ�Ua/�1��`5�q@�R�f�����
"�Q���YA�BWP3��
v�
}L(@a�O�HLZd���Se����N`�!͝�q���&�NR��L��g�b�Z�=B"�A5�t&�����o^��Qy�?ǁ�C�����}�w���>N
M#%�I����Y�Q����$!pb!1;�B��XB1h&>����A^����D��Z������B��gH��ˌV��y%��i8b�{*%Sv��e�W��'����0%m6�01�vp�e��`2[Q18�7f�-B:���w�s=K��"T"=�y�0�LF���gN -��
:b�&��T&�T2� {�.�15qU��U�V��{�Ýw܃%�W��,�8uW/�áCG���{qu�,���
�L� )]}��-�8�c�Uۅ&�(Q��q�&�1`��<��PH+�
�}�
B�"U!���	��D���ps���M6������/D����?\?!_R/R��\��
�Rl/��I��i���4䱳� ��dSy
�y����D2����V��[o��S'ϢQo��w w�u6n܈W^y)��k�����ӧ1553����C���������=��S�x�z�xAD�C���Q��⥳�W�6"~R�(��P�xߴ�:��<{�3�p~��D��F��d�!�o��g��2GWMJ��PA3�&]a�ϩb8�g��{lwM����N&.����uha�\'!D.�D�K:�K(�G���jKQXN.y����k��Q��D�ncӖ������ؼ�V�?����?���E/�5����@&A!���dYN)N�q���O���w0ќ�dce���O��lyD�Ւ�i&��4���4���`$Ҙ��p�TAux��vc`�N��I��Ο;�O��MKcA�Oh/4wW��c:���6�Z.LZ
R�cFd&�C�9�8f�gK!9��!�(4II��8S���I�]����A�,D:�WR,�x��~Nћ�:��̈�|��D��|)�)�W>����"Ǥ��lDL��Q� Rq��v���I>5e�84�r�Ke�+W����-j��LZ�*W�����v�Vl3�M���s:d�畅߆o��qy߰v���X�FĞ����ք[oI�#�'K]&Mq��&<��2����S'��W���g�"��=����mچ���a�Q�O�nZ�O�����M������w���O?��%��]S�bb�jp��-Y"t�Kϣ83.�D�sC��/+�V���lq��Pf�]�A>��ڛ�b嚵H��`{Qx~\�5_��K��<v�)J�+�!�>�b@f��7�,W�u"��?1����x�������N�Q��!�ժcf�����p��X�q��ӒJ�Ld��&��XL|x�4������o����c�ǉF)�������N
^��,��غi>�����\��Zu��G��j@D�tp�<A*}��/�˨�+�'��*j�*Ε��3�{P�x�2��/<�d&���^����&��R�>6�
iW�'	��aPg�V�j�8o�@�Gh����KcNND���w�Fч��	���~2���L>��2����V�����Ǹ���|i������>�ݿ�6��մ$��ˣ������EN�%��Kl�C�;�,���\�N�p��
��
ꥒl�Qۆ�(w!3$<�*�~�<��G8�찅[���Vi ��/MA��bP��Ԣp��m�m�}T�t�qXt�ހ�2ue���+�k���p٥0�D6IqTjI�
�É��X�"w����-ƒ��1�:�����K�v�<�V�
ر�Vlټ��Q�Q�:��W������{q}�.ׅM7SM�~]��i#&�A�u�S$ڲD���F=����3�h�"(�ۨ�n0���P�e����C6�WB�@`:_����ڍ�;,�C'&Y3�D���9��:Q���9D�B�7D�4��S ��
�?|�a�r���|n����
�q�Í�{u��m6Q�{�.�Y�����i5m-<��n��<�M\�x^�۷o��U��������d��X�
'��ɓ?xϞ�x1<���(�r����� �-[�\6�����?�˗��'?���!�&�NC\�.\� ���GC�b�ݽ09U�z%B6��Q�+�
"���� �r��JP�ol�x��;D��ܔ?v��٠I�:�ær���!-�E!Ǘ�ݕ�<V ����l�m��"곓��ml޼���6���7��q���� �J��Lb(f�W7ЗN���~DQ�Ǣ�t�VS��3Z���b��=h0A��A��!�82S��~Z��G����x�*�zX��#X�'�e���K�9��S�$)��Ԫ��I�5Qt���@^
�*H8n�0a��ER�ӿ��)�w6MԐp\��~:-��)�M :�
�UL6W
6�����ϗ���-KL�U�&�0�t�J�,�J���b�͟eEJ��?��U�MG��g"�$�*�>&�zE~&��2
UNF�,U�/�|�jȤ�!���?A��
�/����Wh�JB�_"1N._�S_�}���4��d�����l���5���ӯc�=��~���<$k��P�-���x����l���#b��eB/��ĵ��~<00����۸z�*�)qB�L��H����D�r$������z�]G_�6n��5�O���r���Eh��\���
�$�ӓLM���'��(E��$Sُ���XB:� p���4/����NI�)�8���ʳD=g�h8�=w���r���� Q�?��ǏKS��׿�����f&�l�U#ER~'� nTћ��dQF���>��0�Qk��f�b�����g^�ȣ��"�d=��|�G �B��U��|~Ox���9��8��Y
�@C�S!� T����9y=���(}�� �뤚6����M�זBg9�����U�j���}H'h�.x2��ߤz{~+�^0�qS��Ya�w�X���������WΝ:w��LI�^ܻÀ����\��nX��E\X�	L-BC�۰�R(�"�kY(�Q��EF�ɉ5���D ��9�[SPf�-�]hLb/"�C�P���t�h���'eG�妅�mŨ��n��P#À�Ѧ �ⵘ�(7a�=[�Ӹ)rr������4��Cݰ����.��Vb�ƍX�d)FGG1�;$v�R���'-` Ӫ��j�Z�r���(M���g$�������TCn�x*'B;�@$̸4>iC��(s �)h��V���䕲���hh�k
�$�v��4���Hg�������^-oQvO���Ы>��s�	���',�i$�MAxu7����7Q~���;!��^ټ����c���4Fc��D&Ş=�JS��/��G$�{p`w�u7֯ۈ�|�+���q��W�X��~�Ӹz�2Ν� �7�?��_A_7������������l8�Ɍt��&�d� �-_*N��΋Ȧ�l�r���f"o�$C�rI�k-\��^{��&�񈠙rP�Մ�<C�Hw"�m�s'K��p	C͔M ��j����Ѐ��xP�׌�&̵�C����U�5f���{߸��I!{��Y�JN���شi~���7oƕ��ܗ��#OQ�/�G�ibTO`A<�B*��խB��t|\)Ma�Y���䈃z�.�r6'SX�Ρ'Q@�7`v4q<� ��M���q�M������_��|�`�Z�'�xq/�NN��������LlE�B!
kU��3��	�������J�N��擏�i.�pN^�l����Y�����::�iI=�X5���`Tp�^�o��l^�xB��j�q	
��� �J-��h�k#dǗ*��r�	��)=�)'��@�cRqz�-)��(��4>)�>��ʆ�A�d�h(D�%�jk"WNB�k��p��$��\��F� #�#w�M��?��>�]��F<���(yzV��������w�+���1�����ilV��?x��.]���kVa�ͫ1�xm�Å�Q�40:2��˖ː���K(�L��ڢ��A�LKz�ǂ��1==�KgO�ʅ3�ݦ��۶l����O��r�p;q�o���p����kq==��Do�)��:p�>~Ќ	%����g���j�8�"^z�nA�Nee�ҙ�8s��4��{6mفt��׹�����3Љ��\ǎ~����)��7Q�%Y�����)�J����ia��(V._ B�Gy1}+*��Z�Ja.��y�_�}v��",���5?�C�us]���2I{�y��s_��
)W�!�\��5��/A
$�R����nN������nh�X�7ԹP����@�26�k
�`ӑN徚�+�f2�7�qS��a!������><���^������s���)x��E,.7T8���Yx��OgUq&NDb]��N������§�z��f���D���jTt����FaD4	���>�DW@(M�h�
0�H�P��f�q�ܮy'(;1�5\m9(���$ꈠm�`pEx+���t����`l�)�U��BW���d���LH�z�q�z�߸�g�|r@R/_>���W���l�J,_���Z����������cxg�L���0�Y���q&�W6	�5��vm���o��n6�#�A9/���b˒���OqC�#����E���;HI; ����_�0mn}��Em] �'l
�	q����x���
���h�Y�T�w,:��,�L0��?�F�@
�`:�ܕx��BԀ��a�>v�ކM����W_���Ga�=����{�,[�O=�.]�$Z��+��_��'q��5��R���0SG6qM�x*���m�9s׮ψ5$�s;~=�86mڈ�|��?E��!���F׌Z��������ا�ɓ'��{�0[����H%��#J<z��Bw����~�f��㪼���v�Q�H��s�i��uQd��M�`}���w��u.�UwWuW�0�DN�9�	��$R�DJ^˖�g��Y�g��ږ�zm�)شlRzE�"%�"�� &��A�`r��]]�]{��������s�|8���ĤU�w���ܵ!~�
���<4^`8��@W��x�3a�:�rnZ����\��>�{���0q�^|�!�����Йɠ=�|3�6#���Lxɓ�u%�o���h.�\�"�>s�\�����#�!�'��Nfq*��ȻU̖�898��\	�ypݗ��>���.D=�dᙱQ��Y)a�5l�O�JsA�/C���VS�T��F��Z r�@�R(ʯ� RC��rf	0Ӆ�q�)�8��1�L��V�ȗ������jL��ЖN��Y"����'`!H��EK紈ve����8UKD�~+� ��Xv2E�sK�i�h�Q%��i�z�G�ҥ����M8U�#8�0�b F[PR��+msAc{���*��7w������[��$E)��N�)΁�z�*
�J���*3�`"�E�l��K7!m�g��w~�ן~��2^�G2K/�=_��\y���%�E����Gyt�<�8�#� ���V,�ʵ�K�p~x��Y���
�б�8?pc#C��0�a�_��A�ᓮ&�<�1���h
��2X�v5V�Z�h�U�C�zH�=7��4�j�6�r�ꐗ�#�bb����C�=�����.p���u�.9*Ǐ�³�܅��a1O`0#D;f&Q�łyI�x�5ذi�||DXh�J���+��n����x�'O��=�a27.�Ld4�����Յ�5`��ѰxQ�
��$BF'r��i9.(����'��K�g�,�<���\cOB:�nxB`/{I�m<=��\u���ݜHQ��I�
/�B�:�C,��$�����k8�_8?ZЌ4�s��lV��O���{.y-MK3�=�lHJB��O>�lk��h���C�o���-�Yç��{��7�u�̙��Oabt�j� ����m�4͎#�0=���5�@BfsY�N��W�%ԛ
��*���"P�=�R����#Q��z����p�b�M�:�~}]�mD���L�Y����c��P��)-+b���Qс\��<a~n��q�갫ʟY������-���⻫��w:�F��ꦁ��.�+��/^��TJ%�L���lz|D���/�ebYIJ���q�<v����}�P,��&�L�LY U� �a�j/�����Ϫj>�}�� P��sC�Hl�&�"+"/���n������5�>_�$c���aR��������s��b�����a� 8�-����S�����)Q��>'Ȓ��k^9�L�)±Ѝ:�mۀ-[.��O���;(�15�]�˗/��^�;�ޖ�ݸ�2�ر�����/wallB������X�h���F��{��_�#    IDAT�P��P#J�O�7�z�*l�p9���GQ*�{���<w�.֍<?�0��ĝH�bxu��y�!l$Kd�!��U	�4��p��W�W*�Vr���l��w̿=A�7������.�7�������c�ф|m����_���5�r�t�&�#���o�A�kV���Så6��.�mي���������0��}�4:Ba�e�������wf�&+%���bK�F1����@J�5j�5�#*��&��h���q���J��iL2g�X��n�_�2�߾X�v�����8��+�''��rH:5�5�D��J����I��'�ؒ"�����ê��3����^RV ��fK%L
(T���Ԉ�{R%1���k���둜� ���/<����AX�chK����.��b&�HDta �u����	��!hD#ؤ��q����`��&�uZSb�:���t���r�jMPX:$�;:����q�-� ��-"~'�����������3'9��i5L��S�Alj%)�.�2�f�y�&u��)R)�R!��~EC�*&FP�Ai?]�X�S�Ҏ-w܅[?|7ZZ�!{b �}�G8��K�YhZ	U;��VG��W~�\y�"z&M��op��s�870�#�ajb�ƪ�kpъe���A��e���� ����V
���yԪ%D	t�.� �G��:���LM����Ԅ�Vw���n�,[�f,���h#��les<7x��a��9x��rB�2���%L�n?�˨b���l�;�ݻ_��d�dZ�R����Hv��7�x6\~b���\:�fa����AgϜ�KϾ�������(�nZ��Ԇp0p�ۈ�eD#��$%��#�4��^��u��^�v�s���k�3��-R��FZ��@ů_�RR���C7�RA��6Jj��W���3Gm�p2 ��|!��?WI�e��a�Au
���>.�a�O�����Ш��K]�*���L5��5�{g�n��i��P��D
Kwv|�4[�>
~���C�߻��o~���k�9��!ڱq(A7b�"
�7���$S��!��m9�G�ƙ�U*��mȤxs�mS͑��^�}IIHYH6|Ǳ�\	8�N��X z�CB9�P� ����#芆�>��:�l���X��CG=��l���m[5��6Su���������%aki��ׁͦ@�!�KKk���`���h�b��SR�Y�	�NO�u肅+0��"ģ�-*�p��8x�?�CP'1J�BI�k�M K) vU�R�
����Uz�h
.&�D�dDQ\n"O!)�;1y�t�����/����� �5H�E��Ĥ���<`4�״����_w��9W��&ߧ
�(��)Z?^%�#D��c	u+���hO��#�uk�a�ʕ�?q��ƹlI�`[�l^��ӧ1BX�vR�h�zs/,�A,��5
K�-7�"~�O��i���t/����bѐ�('�q�:9�=o�]O��&�F7�)@�YÚ5��n�J�wvaz*�r���,����(��bbb
��}�@^s\T�*��؃���L��<4j��� ǆ�����o
��������.�?J��L;򯭹Ô�h.d>o�� �Y���e����}�]v)f�����.Fv=�n������Ӓn.�!R;��B(6/1Z�c�V�P)�f(�.3���)�>f6��ټkz%����F�3�V�(�,��*F[����"��������`�������0rYt4t�AtG"`�0��M��!#�l�+Ȃ�A@6�l�ؕѺ3"�Y�w��D��YMN`�PD��-Z��L[6������q���"9o��#xg�.<��F ;�D�E�.Q�ȗ+����q�#A�`M4X_¢��jT��B�i�!Rg^�j8*D+� ��4J����I����d��"m�u���ю�w݁����^������{�G��>rI��LL�#�i��9��f��X�*^+��+��7��2�Lrj����3�.IBw��{>�[?�)#i��6��οa��a��%�Be��"hzZj m� �1zTY��5+rB��K��M^��w�͓��v���UV͑Z�F`;Ԭ��9��0�z�c���P�"��8{{�~<�K�T+y,�׎����k��ŗm���H��D�ͦG���+�;�������ADt�^,$/�h��<���0�hт����CD�������`N�"-��c��'��/%C��-�DhL�C�Fz�ZHP�¡�F144�=Ͽ��G�b:?ǭ���B`3Xѡ�z�=0��46l؄�>q�)8�0$N�Ct���sY��U��!��9��ފ���P��tr� 
�
u ��#K�i �̹:�����kc���
80��L
Z�
�K�	.���y�&į����@�B���9��6�	�/B$~���C�'���2��o�-������g������_�ޱcG�;vD�W�Qk�����rЌ����t��&">E0�#n8,�~�Cn(:&gV��7h�� �\M�0",��)A����f° ���U��:�Ԁ���(��#��b �a���h`6A.���j���7���C(��;ܲVD��^R��j�؆eC��$gyޞ#���y�`�8&S|8�ʆ7����%�T".�G��G!7�r� ���.���%H$�Q��ϟE��C8z����V�2D�}c�wh�j~Xƹ�&��Z;�F�צ0�.ϗHA���Zm�>�ƇCӬ�ɤxv�9;5��m��B�m"��ȇ���.���T0��)�����_�~�����Z����E��B�s�Bٖ�X��{M�l�E���Zs�����V����A8��e���ۆ������l����-���&'��p�b�cf�B�ϝ���r�������\*��$,�CČa������%�@�� �$�;v����p8#�m��H��]o0�"t#f*��u�c4��$�2��\�ajz��S��.4���!t�]{�����?4��P�/i����bn𾡀�A3}�G
�7�O{�#�9����q􋦈��-�+B=T��
��,
�)9<7n܈~��t�*�yc~�������Й�#7���z�ͪ�
�"J��:��5r�Yo�H�:�'�M�ѦG��OG"^tF	(:����Ws��a�u䨏��"q���\s��Ȭ�X�恷������=r�b	���E���PP�K���t�ۡ���mhh��G\`�!.��hF��7�D� �X!���\�Bݙ(WQ���m��B�O���������9�)�$��׊�HR��t
��J���Ԅ�8|�I`������F3��梢k��(�4������1d���K\�0���b�����>}�rq��X��|^��0{�ZD.��xo0����ˋ_ke���զ��e��Z�~��*���%�O�i�Ԥ]�k��6��a�5��Ϟœ��]�&�#� �5nU,��,�zL�8��s��k�\.���.�wkY"�M�P�\F�0Q�Ϩ�`)����0::3�����/��`�ZE^r��I������o�Z.JC�N �^�w�u;�mߎh��Cz\P4��"�j( ��PH
7���$��r�ח�U�n�͆g!7�f1�FM�� ��y�8���q��w�����#�r1'ԡZizӸ���2��u����r�SV��,��p����^űc'�c�s�%�)!]Mco`�D	�D�vc���B�ւ��B��E#���쥰�6Q/���?����\.Q ��� zJ]i�j��tg�agB�b�R[z��HD5,���a��#KiղT�! -N������(�C�i2�)5e���o	K(���4OG��^�I-��PCiJ~���X<�X����ෲ��?�^���O���w�yg�r9q`F�Ќ$4N�M�����f��O+P��E%T_a���:�M�q�� ���X2n(��4���9�`&K�v����pa��$o1L�������s�BdV-�eF1�����C���Ѿ3���&��$��Z�p��m97	D	�� ���D$E��B��̀"r���C���3�E#A y��bV6b�T+�^qV����|
f�p��1�<u��d( É4Sb���CA��>R:�h.���jNt��_�Bd&���kbIZd���2�H8�x<)<]a3��G��Tj�����_V���=�}^��\���7o�ߏ�ą&�/����P0���D���B����uy���ϙE\>:T��tg�L�pUI����n`b|�,���L砎�69Ԧfg096�t�.�&��_���G,N{@G��gf�*4��&C�jWj��������(W�­a:G�������Fz���`0+b��*�9v<\��BLu���/��k�%��s*�����U:6����e@������ ����`��6t��M��j3绕���/*�O�=�|5�J���N�������Vc����o���F� ��-Gk*.\`n�k.��LT-LW*ȑW^��{�W'F�0�@O8����T�T<P�z� �L�*�d�"6�jsJ5��^�7�~�\�YD���~|����G��E�#��T)- ��L��s�a j@���V
eEɺ���I!��3��j	3���B��Y��1��
��l��1\w���r�J W¹���_����5���nH�oG8��$z	6��qv�����(�j����A�*US�]a�����/�qzte:�q�0[)��`�m���O}�%��f�� v~�_p���Q�Ag&"H�ZY��e�������C�=���/�D $�3Ѯh��0��F�
�cM�bh�h���gp�M����O>�'���0�Y
�p.ʲ(��5+BI���@r���2����d�+e�1CG�q0:9� ��� �ujAhg���mk���wc��UX�z⭽�:v�$�)�޽�� ��bb������qŕېl�ݠ�M��PK<4�oIu%���T��(�@�Ń��2G�M9�8XQ_�M5��R�BŪ���)�93�CG��\��p�dҭB�cFB�ay�I��i�u'q��-�l��hi떡�\�%?����@���8?8�7_�#�-��Ӓ'A�j9�ϲFjKhIk(Iz�Mw܍���d�RU^W"�~v
�#z��I�Ŀ�;|�f~����2��H�C͊B^DWZ��bT!e���<���,DT��V�zK���/�V�Qm����Ѐ\�a����Óؙ64؞��ù,���R�L|�tQUGmf�сғ��0�~��#�e"�L>�d>
~���oݏs]7���]۾�o?�����~��с��B@OHZc�Gss�{��͜����{B�5Z
V�o�<7�bu���I%R�@��}\d���I�
-��`�$iYj�%LB�4�J<N�qģę�ٚAz�t�[��[7�	�qj`��|8��!^(�p$�\������5��c9�*���o~a`�#n��a�t�FV`�**S��+���Z5���i�dZq��+�x�:D��U�/���S8}j���é���P�)�恩Ɂ��Ft��?[��.NCc�Yi�R�FӁ�!)�i�ʹ4?s+�!j
�X\�b�<�f׃��Ù6�����/��]���!��\�77d��kR��Pi���4�: �&Ľ�?��a��� ���_�����#I��v���%�S�!�fa;e�-	F�&Q��Ҁ3US5�eO��@�Z�N�9�m�j7܆ ��)�To�]:�u��)W���m��ӹ�H��!�P�h@�-�a�^���6��wRҤ�@�m#l��2Ř�C���T��H����Y܆��Nޗ��1i�|���ѐ�z�M��5����H��Q��>��\C�͒���6���%Q�&?���&�\�A�8+h"-I��֭Y��7�ĳ�������4d���Z"�j���JY(sDʞ���,���LPG�A;Su��Aqa@�j@C��b�r�-Y�:5�5Uf�4lTl�by����pӽ�C��W�v�~���������)�j�G�h�EБH"����=�B0G(�{�.�2���8[5H��b���c�Z���$r�J�"����&j��SGϦ-�큯�o��(�?y?����3'����U�E[8�y�$���G⊺D��D0�Md@5�E)���J�rXG�%#�k�Fϩ��Z�"UCjf1����Ǝ/> �C�f ����@��1��e$ctS�3	݌��\q�cފ
�"}òl��>r�k�Goy�K���M�M6���.#ب4a����,��܋��8`x���x�;߆56��iCV�@E��@8�B�����ֳ�e�,j�B>�C��D>�����aF�-Qb>��@4�C7]	1������B��M'y'1tnT��]�v�T)�yؒ�`åk�;o��͛���M�S�3��*[H�l;�*��YLM�թ����Aݍ�_Aw� Fd�R��N���B� ��!_,cbb#�c�t��*��F(������М�o��+����i�B�����+�AH������	����8x���E���N	��$*���LA�~d2A�Qn�~5v|�@��ٲз,ҳ*5i���xf�`��l�}�ۄ$�l��>�Ia�6_U1�:R#�y[@r���5�� ��^Y�*ʒ�����%i�M���U�J�y��O��,�Xo}�E�O��4L���;J�#C�|b���W��
��DD �L�L���43����9�u-����]׍����w����'�r�������v��w�v�FCXr^Rls��SK�/����^B�M�|vxTr�y��r�����
�*֚u	����!BZK0IH�R���*�x�Ḭ��wa^O.\���nt͟������ �&f�������W_���þ�0�-�B�=�-/3��.�"�?rͅi)�3¬"�d��+^&��P� �v
�Z;�����~nfv\t�}��ٵ z$%aTӧ0:<���Q�:=���#�
R`y<@��t��(�E"R	��j��EW��Ԗ��[h�
u��������C�D�W�^?�A/��4��o�(I���~X��\�%��M�ב�L�͢�y�x�}h.�����6�~�.�}ŝ�8����ƛ��0"���e�+5fST��0�(�IE�"=|�%[^
�E`'�\��)�2;��F�S�8}�iyˀ*^ct��Eh�*�L$C>��#�d*�.
���D�`��%şi��Jn�kFmI�*.!J��-&_�|����$����a�Տ9�!���ʵ邐n�@�P>�ﱼ����忏�����Z�k���ά.���
�i�J�G̡`��Uȿ��~�{��E�SC*n�Lą��o40Y�`�ja��SH)��@:D�B�F��f�qX1��LL3`�R�d���e�����:����YR�!7���w����v �p)
c�x�ɟ�͟<���0�\�@oOZ�[�I$�M�.S�P���HkFRv�ڰ!��6��Y��4��7���agz�Y:ZM!3аJ�-�1����p�}_@ۢ���ƣ�M��n9'֗u3
-Aʌ������ ������\�"�F��E~<)M��"�� 04:���ݏ��A�*Q
�-��b��p�g?�����	����ob��>h�i��3�B0ދF(*��	#b����)���ii�O ��eYA�o `�Á�)��,ڔ��8b\H5�(U-�l��\}Ͻ@$��o��O���!{�(�@	�#��E�f��F�h&j� l��2̰�rqP��$e��u"�,dPPKj��J�3Z�Q�L�=-�V`�Z����L�N'���'�ƫ���r� �і�!C���[�nE����P �~�c(D]8򎃑�?z�C�;��c��������� �ҷ�\6���@�v�F6_�I}݇��f})��N��[/`��\w�U�t�f�3���l����5H��}C�    IDAT�Bp:���w���C�-�̾FV%�j� ���
�Zmm,�{�}��h�/l�
� N�Y!A�dEbQ��||r$���JO����N9$@0"t91�,�L�K-O��b`���$�w���B!�婖c��^��<L�V�DO���q���U�IW�᢮���1��uI���{�?�Ȫ�p(�V���^�kp����*2?�TK��f�{��������|������������?��()$��T���<�q�.(ߋ^.v�r�����OO�?�fB&׊gG��p�9U����P}��V�U�*��@9��P3R����l%r:[��1D�),�h�nڌU+�c��%@4X%�a�P�ũ�!?s
��@>WƉ�8�#�Y�p���ך�˪V��dB���9����w��C?�Ln3�6���)��]�Xz�
,���X� ��*fg 8@ǿFaՊ0cQ$�t�I�\.br�4FΟ���n݀+�)�oSŇ�B�n@+���e�Bv��,�������NC���CPh��p'*Y��q�Pa3D����M�T�EP��s��_P�FsN��� ��ѹ��1i��rx?G���f� �>�ѷ�P5ըۂ��VUm2���V�%n~4�̸�7�C*EÂS����`*^�|δ���H��	�2�J"��X,:�:F3A� F�b1Z����1��y��baI�f�(���.h�44Q3#�!W�����e;IZ���������[Y6u
�v��i��{�Lx�Ԃ��+��MCA��s�!��M��>�[yj(��k*�?��G/�x�נ�<k�ɰ�:�]�P���˦�7���?���a8�7�oH�9�ǒ�4�1mۘ��2TF�a�-s�έ��È���f��x@����¦����`���
e�EB�
 �,�.= �C�B�w>n��˘��Z ����x��~��laX�l1�^{%�[�x�E��+*J�B`��R[x/����!k��
���7�Z����,j�2�c8v'�{F����eW�p����e��np�1~����?��[{P�M�g�",ߺ=+V#O#�����$�B�ܕ�����Y�Iu���'�1M���p!?6�w_ۃ�����@?2��}�m̻|n���ѷq+0����W8��+h&��X|�zl��^8єܷa���
5u[�"��q��V6z��X���(Z�-R��%���2J��Ǜ/<���Ym��و��æO|��}I��;���/���#H�D%��Vu�u�T���8��tk�R�7\� E�i�s�� @�RY�Dx�8䆃`�����$z�u����׬C�E�Mv��5p�X?~���x��P�
��3�;���V�w�PK��P���زKi	gT��J����x?�g8r���[H��݊�EM_g~��ѩ�[YX�]�ր�C*�"T�r�])bb���.��M7_�K/��S�I]opaC$��\6��?~���i|� ��&e�-92���с����D�B@:��fp�-7�3-�#<�Ԗ���L�:�aĒ*C�jâP�÷8\i�=��bf34(gF0��YZ|G!�>���{���%�B�z�ͿBD�ʬ��y����,�Rs��(9��j�s�i`2����ZD�j�Ĳ�L���*Bo�~/�B��=�W�I\��[FӴ$���'S���鮳�iZ�_����?|��W���?��Ɛ7U<�P�!B��|��	��|��SC涄^
�l�I=���%���iX\4
�ج���ڈr([64�&�l���B"~�����1o�rt��Ò�+�r�J9�R�	��'N���p��(���������l(Ju��2�rEd�U�*5� bѨpmJ�r
|��V�����1ano�q���w�"�0�o	֬�K�D:�D�E��cz�*���!�uӂ���F04pCC#8wn\a%��ݐX\r�A�D�5i�꺈��v1�X�U�ISJ���� �a"@�У��L&�h<.n���o���Yh�������M�P
�<n��}���J�zJs��Un��-����yA+�����D�����c������`����P�x�451���F
��2�tt�t��--��i0I���cffF�˪ �����==]�y�����3C��*�m�P�����
����Y��������5�BM�����K�xI����8x�8&�rҰS��y�F,Z���0�����x��#(+����l�%��C���b&��,^��9sV(|�Z��������^�:��gΡ.z��a"����M|�{֔���2��xCAs���n�}�Z#��u��!u=\HP���U�Ĉ�C��(������jەW��|����#G���"|�zv
���R���"7���6G��$�?��m��W�+�!ڎZ�Y�$�W�b� �X��VG|�b���o �e;�c�� ^��`��O �91������3w#�q-��KȓX�1Q�&5��"��PUȡ��8�s=A0��Z�<7$�$P*`��{xi�#>�R�b�cǗ��e����00�Ww>���1J�ϊvf�ƍ���a��-��,�.��f�wT�Vk #�V�Uˤ��c�/������<Ə��?݉c�<���P��x����/�-��"_~�J[����78��3p�HuF��q���:�RB'V���y@�$�ݠ�=B%�[,lU#E��f�����>�<�sȱ0{�~���� ��Y�y��m�������~�T'F���-��{1�*)����oO�[n���-��]'����H��NN�����9�c'��̙S�`��E%�岁�;��D&.Yn])t��a����[#���ã����[x�՗Q�O#��������æ�[I�Q���8|�,D$0�4�p�|���i<��#��?�D\9�� �f�h\�~�����Jw�ZD�$i4lni�M76j�����C�Ò&�.3�h�rX����p5.ټ�L��!YyuH� j��bO{��	�|�Q�{{/Fg&$�G%��t�C4č���Hk$
�\>=�����@&�P�n-�t�}}}��/g;�|��p�R�9"� �`���A9�9�seTЧ��5�^��Zy�EGӂ�_~�U詧)�h=b(�b�y����]�Lx��@C�̜�����x��R�&�+�F�\Hq��H#͔�~)�IP��<V.�$!�!UL�h4�T*���H���C���K����#/������O}�K���t��F"���P��lE=^���i�=���Uk�����!.6v9+
/`���!���z@��>	�j�:�R�JQ���>D�q�������k<�K�_�k��[�D[�������P���#Gql����R��C�V���XK,#�i���j%B��/U����$��˄2��Y0d���͈��xY�W{�!H}�4�1��-ƺ��b�5hIg��U�3��a�f�`Z����f'��̩~�>5(�7t��tS�)_(:
Е�m�&.*z�����*BU��˂%��2P����
��)���%2p{����+g����~��_�΃����GE=R(Q���;|BA��Z�߅B�чxX�ϒMᅔe����b�B٤�ZE*�Rҕ���zs�cf:+N=}=غu3�/����bGk�T�)���O"�l�%-@����:2�<xo��ż�PД&�C����Kc_����s�axp�5f8��[����]�F#��t:����ݯ"�bժ��tD{Z&w�������������0��y�D�
���FΏ���_���Goo7��<�{��l��� �9��9w
:^����똼�ﹰ��&�Rn��i^�����j���q�����N�l:)�c/W��2��)dg� ����߀�>�%�_�N�Iܹڑ��4�t�`���,
������"����0��&y�D*=d�U�n��[�򘨖1ͼ �inQ]�`a#����0�����.2�ob-��ǻ;��3��l"7�$.��j���O#�v�&]�g�^6R�nO��n�""�Eߒ)a(��W\Θ�	�\@��P>}/>����/�t�t�QO'qǗ��ŷ�$�P�?�'��8��N��Y44+�lƇ��{HS�k��fBܤ�.F	]U�r �	j�`"�FA")����K5�;��v>�7��!ZCu�:�gY��~����f �fKx���ƞ�Enrf&�M�݆����hd:�:G�`sc�4�[����p)�_C.
eKhB�D�vT�����OP>���gZ2�K>�w|�~P�3���qx�shXS�u�n�҃0{���/|�o�0�u�`o$�z.���az�<��38~�8���ܟ�tFj�El��擏���d+dZ�ȴ�!Ӿ �pN# ���g�����ό#p1\��c���MbI��2��]�U��8��wq��:�ԓOb�Ν�V@KKL����	1�P.D@��U���t��D3	��*��!��H�$BU��03�Zy��r�\�iZ�{�vš����LT���FǏ�����y�e�N�pV�K�4#�H�G4A9��;L��Z31$�:qQS���*��������:�k>V�t���IID�.*VY���AXr���'MsΊ�ۼK�D�j�.����O�����C,�mj�BB'�qB�Bj������� 򰍐�Ck`�Ho5��MᢑHMH2ol'�R�A�l�i{�F�9?��sI�4��I(�������|"��Y2��Pp����?E���=�o|�K۟||�Ν����މX4��ɢ@�>�ƜH�L�4��k�|��F�|��b�ᡉk,$'frsyc���\��ڈFtD#!���s]Dm��͊�A�V7�p�Hr;4P��t�u�����g�F�<��(�̠��70x���?���'012"N$%6e�B�8���Iǳ�hj��/���(�8>��N^�ρE����A���1�:B4�����n�%X�b-:�[aFB(���{Re,$��s��38�'��b�칹���PD
���e�1�8\5D�6j- ױ� ���.�eZ�K�� M��D�Lzn(��֯�w.�Z�u����`^3�zx��+���N�o"��׌B���柯Bt.l�����|^�*�%�lذ
���������^u�t���Ch>QE��,Ė�����~$R��bExۥB�V^���oE6;-f�2^}�ը��y�-��0�/�t�\u�X���c#xy�+83�ºUkq�UW���8xh����b�z���gv���3��[*��s�"4��݅n����$m����]�Q6�/��J�*�-[&)��������S��K�HD1��G^������GNJ0�K��5Tz�V&�4�u���)Ϳ�����rc�7�{�_lzo7	��������+���!�b�(�i����
i�m��E��ތ�� K,F�� ���� f�P�P�W0S.��b�С��h���'�F�9C�8��̡���0S���7�Zȳ6���0��a�J$ DC�)h�j�Vl��^d6oR���Ob��;���߃=�E<����^�[��;���%Z�6h	B��!l�DOЪtas�n�<b�V�sh	Q��I4��^*!�X(�>����_��珣3�"5`%b��ӟ��[�:�68�~�(^��h�Ƒ/e���+������v-\R&�w�ҡPS���C��w��b:/��߈G%UYl]e��a�dO��F�Ň���`-f 3�*�����}	˶� �I ga����x��'N����[p����;����m�6��W�]܌z�n��!BY.x-�
�9Q�`1BH�<���obr�ۈ2��']�Ě�n��_�2�yK��<���������3����u�tuc�������i���0`q`Ԅ��ū�_�+��F*�����]�\��ёqDL�F:���Q(� ��YC�e�fZ�}���E��M�#;=�Bn#���Śu#�l���x_�Jd.P������O`jj
7nBww�4�PC:i��l��pi��^�	�M��i���q��G�pE�h�=3�r~]ml��r�߸��n��O�0�a���Ϟ�c?�1�{�YO�++�5��0�4A(��LCG8B��:�F@��(5��
"&�Ie�0�b�9
���_�CiK��\ߺN��2\W�r�5R O�&foA�����wd2
i�'��r�I$��9_��{��2��&��e�CVt�#����"-�1��&�صr]�:�3�&�;;��ډ��y�B1�k����z���m��̔�g�->�&�P����H���C���O���7����z������[�<5d2�H%�Tj'c�9��϶�"���S����\p��=��
�,�`��*Ka��l�(��(��*b��)�7�֕:��
�i�VQ"�� �,^����X��5Wl���$Vnތp:��u��>��Ǐ���엤���,GƐhm�Ϡ@����̃.��X��S�=k*ҝi�
(tz]8��qɛ���GP$R`b"��W�d֮]+�[{{��b~
ÃgQ�'�F��p�(��10�/T�S\-�0e3���W^�
�͡ ذ`�e
�r�|Qq�!T4ٚ����(1�����R0�>�������>+/�z��l(�6Fd�����+����M�m���������*�LdRs4#��Ko�V�\��>�)���^~�%)���6��]��[��������"Ӗ���Wclr/<�FHQ(h�#:�.�t)V,[�_<�$���Cd�ڋ�f�%8?8�����a2�ظuҭQ��为ط�]�9u�hn���y������V�Z��}��B����nT-�)�7��H��x�hǎEOWz{`��G�����p��u�rP��{��I"h��m۶J������G�1� :�)i��V0��Ӽ�榽9���9���oք�Uſn��=$�5Hs�1����r�Y4�<��	�!7�v���e(��a���ۅ��!��"jpP�������t�zAg$.�ANm@B���u\��,�󤧾�%��No|Zҥ�RADRa-�p��4<H����Ѳ�J�}�/����⡿�o�u��Q���Z���_Dr�*Xf��_���,[o��x=�u��H��ɗgSL�7��*r�3]�SG��?�	�5�@]�C[w|��y/��W�:���g�����(�"��`�+pǗ����W�	F8�P ~(���@ݢ���/�3A�:$4�	@d=�E�I� �vQ<u/>�0^����ʈj5 żmW�{�G�%[�@�Vp��g���}gO@�+��o�n��"��+�t�d�D��3TC&ɲ
���K�&�b0�Dq �.����Ŀ��_�|��Z	���R0(C�G�w_��.���O��G~�����E�YA%@t�b���ľ4�t� �5i5��Y������x�]8s
��r36n�X��SS3��?r\(k֬A{G�N�lv�j�F��ᰢ�r[(P)E(�����9�H��j(`cXGX�/����.jQ����?~O=��[�l�0�ȼ�d8�ZϜ�����9��a�dJ���RIҡ) ���u)7���8ʹq,��"����]&�y�@��C
(��(7b�>�䣏ᙧ���s�ٌsx�KQn�Ct
��\����C�h*�'"�j.>x���A�����:��G�tU&�5�m{�4�����o"i����(2s~�3̣I"��k�l!���1ͨ�,�&bRz�������䓧��FÓ��Y:�UG^�٩5�-c�`ڔ�Y�b9���&,Y�R(�D��e\<�e�����j�P�#I�\�L�<�Ns(8��P�[���zO�����g�y��r�����4tv� ¦� ��:$�����)?�[�_R$<ڌM�\:,�7���䰣�\A�0#N,�P���i��/�0�C    IDAT�V*�.��q����n�q�:r�*��X�~zW�D���T:�j�6�V(`��0�'�p��)<t�6��NLchjR�H��-O��t�Q� <�XT���Y��|H��6JL�q�M�]�n�`XCK[
��.���˰x�B�f���������e&⭰� �'K��� lT12z##c<7"A9F$&���t9Ĩ�̐�gf�@��@�*�
�C�g�^�B�TF�T��$����Htn(0bQ�Zs<��o��]��UC��8�׈B� ���� �M���f�A�5MQ���s��^����m�����_5��.����y<��O��k�K�%�P�>|d�](�*��SO��l����N�W_�]�Ã)a<ܶ�����-0��?y�G8u��ń�o��Vz�w��R��իWb�ʅx��>D�V�Z�C����߻���+����Ȑ����u�s���zg^�L���-^�zE�ն_�E���߇��磯w�ߵc�3����;n��g�/_�P�.I"�5�^)���G��&D��� NY�uV��B�e���U�{j���恍�n�E�ᣌ~����\��x�<�n򉭺BQ/#����Mw܎�~�3X�r06�����'���!��j��mq�a�n���D�|���D�:H�����rE��f����Ӂ�F�p��Ъ6t�F+��S	t��}o-�#�J���кuн����ݻ���ob��Y٦_|�����=���5��a���#�4(�k˭<�Az�B��B\H�{�r��(t.�9�ݏ�?߉�/��ro��|�_��D��?���
kj�����W`�W���_�c�ŲS	���Ѡ����hI���'PN�HX�\�(a�&Ciw�����{����Ѧ���Hvu`�m�㊏}�ҵ@]��_݃G��8��-����z�m��_�HdPw�ؒ_-��TT
O�q���e*����(�!l�],NR.���H�|M�;t ��_�p� b�*L�+�c͝��H�<���wƁ矃5;�dZG��EVs�Y�w��%l��N؆	K#��!�!Ⱦ*����(��y#�C��;�v�jA������3B)J�X��"tu�ajz�R�|՚�x�KrK��úɥV!?�l�&�ACM�镫�!��@(L����QQ�,�(a�ϟ����s�|����t��dH��e�f��]�k��3�J\q�;'���_����5�ה)��rr��#:��Y�FQ-Lc��>ܱ�N�[1jn 5'���PtD��5ڟ�bfr?�I���q������C#ֆ QhRfy+M�R�RATL6�I�%R��^X�9�x��a��1C�Ykp��*�8�z�Π�N2	(�W����׋�HA�>��Z)��`F�.A�C��%�B��"sFF'�z|d�&?��֧d�E�3SӨȁ�t�{D'�,M���$���z$R-��̆�ڮҶ�|}d_���RW�����'3�oD����^O�[���}��O�z�����kݼa�$ҩ6D)���_��0<Il��!��M�r_Q�;��ÀT£l!(��E:�l�j��8�5��(r�Ѧw;�
�
�bZ�J����x��C�����܊D ��Kqqw�m���FgWV�^�֎v�/�Ώ���·�NM����A�V,���������F�7)@���9���N���*�4;l):�'��7>��K�.�����7�a����g�00xc�#"R��i�lMx�B�S��D�RG� 9��:����H:4�N:P�$3��E�|c�,[�J��l��8TC@��'l@R4!�'R���ǣ��t�_�G�����o�������
�Y���9G�R|���=���G|��y�>��y ��\[ނ[�hk;��+�����O��^xM�����2��O}��4�����rX�n�i�?7��VGH3pnp
��&��~�6lظ{�y{��&����W��m�1=1��^zY�k��g����������W\�}��b߾}X�nn�Їq��9���"���ق���FF���{03��!b7��ޝ�����a㽃Gq��	�_��m��̋(�+"p���M7\/�^xS33�K;��]�Y��������c�=���D�/7�>��kX�xx������ޛ�Ur��*H�c7�*\�W����R��39�t(0��V�
j4p�ͷ��~�׭E��i��أ8��sB���L��jh��W4�n3��|��`3�UD���*F�YL��D�C�p�E�<j��)�u=�ڣI�#�ŤB.�@�꫑�� �%h^��!��������e.+V_�;��Etn������E���/]K��]<��uլ�p"f|�Yi+ӓ�8~{~�L<�4����6}�l��}��,�N��:��c�����_|�����_F�W)��ƚ�Ϯ�J��:!s�G��JJ^��O�`�K$e��	<����w�#�0t�^��L��;��ރ��5�q�6��y���?���7��J��[o�G��O�t@���C��5n]��8 �5��%�u̥*��� �bL-*a��{�e�u^	�{_��*
�PD΁ H0�$�b�$Q�%K��=�5�ӳ��'٭e�mwKv۲�l%�b)f1 $Ad9�B�W�r���;��sO�#Eό��,���� T�z�s��};��|�0���?E��)�U�*"�mX��Ǳ�ޏ�����[����|���!���PF���ļy��o�.�z���ج�IMᄺAJX��Gx��>���O����;oÊU+e�����S8s�Z[RX�z9�aC�W��X�T�AD��H��>3>6*�6���|�hH�G�׮C��u� ����&����>::�'�x�>���d/]�h<�@8)�/ϰ߇X��\�$�f�=����]tN?�F&���t�E�!I�5�Uê�+p���΀�ԭ�:��q��$�5xM�8�o?�y�:tH�3�1��Z�*Ż�R4T�u��F+x.�Z2�#����"	�� n �tP�����*<m�̵J\C=y�mg$�[��ϳ@�gI�V��q��h�@@C@]�6P������$P�U��i�	� �{u��t�0E�`�@7v�u>���<�	��v���l�)��O.�k*���*���av��hk�+�_���5�/�>��]������\��F&Ep���{�~:�(P�b@��\ц���N &(��NA9�,b�����p��*J�� )W�d*�"
�II0ć#j��^�S,��栗��A4` �7�ұ(:�5�T�ŏG����Ձ��Vc�5�1cVZ�f ֖F�R���G��t��q�8y�.��h6� ��¨RH�+y��T�#mHٕ`��yW���P�'&� �>u2P���9s�p�\tu&�7j�,d&�q��i��c@MG ����
E���S���O[B�As$�9�^pA��<F\�Z	n��F�.B�R���OM
��+�**7��i
���&�Dw�� u���G�y�*;������m.�A�� i���Pp��Ӊ�.�}MH^��[EEq����|O>��x�0j�!��R̠#���oļ��x�]8y�"Z�{M�	����6�����cW���1]ǡoڄX���K�P(��&�r�Z�=u���u��.\�/<�
._��%��|�b�����\�z=n���{�$�޳����z�q�����Sط�0&G��m�L`��Ÿ�-"8����RR���ۋ�~��y͊sz�-7���o�sC�c��X�n޲�\�@@�jun�ce�LQUꍺ\�"�f5�Dl>_zё�}H��\+�I�P}��%�ɽH_�S [6n���Uq��GarL|�n��F|�_�⥋q�Cx�;���[��Z��Y�7���/Ղ�h�tQ�3�ߏ�ߏ\���zElK��"�����0���u,\$��E����
��E�I���H$��:tm�t͕�k�ݣ���/8s� �aɶ-���E�ʕ(�|���
� �!E��,?I$����A[cꓔ�%�� %v���o�8:�s�ᝧ�@��yt:ʊ74�|�6l}�W�5 ���� ��'��gP�JX�y#���/a�u
kU�,E�`�+��2
*��s�u%��%7�i�pD�����9��{x�'1#�C�ZC�gb������� �:N��9<����� ��`������{@{\���R�V��n��a[���UB�$��EC���[�����2|�r�8���?�{�R����Do6��'����H��k{�ȟ�)���B�V��qL�U$���C_���z3�l�"��xA~�J��8����&���v�M�����,����ҹ�у�+��9x�������"�����v���pu�
J�I��Md��Ϗ���k�J�\��$3 �A�!�'ط<�M���!<���̓O�R*c���$RF2�bq0����Lv��Bcd�ݥV!��;�D���c���Zb����!�U�ca�X�
kׯC"����	����*m��;���]�6]�p������8��08R��^sL��)��x}�|���~��2Mgm~~)�eoU����������[�k`�a(�<��yNT�D�=��
�e9�=�&?��7������� 3zIy]�[�ߌ�o���_1@�^a�O�\�H��	?�TB7�^K�T�y�x:����_҇~����/<�����K/�n��H�L���㱤�+y#r!K�G�0�2w�\_r�]��y�m/LKYw�A��%���]�	�}�m�\a
��FOiz�Vn��RW4 � � B1�b�0&���1���-N+��G߼y�F�%N'��0Q����"�p	'O��g0:1)��p(&��BY э�]&�1K��qi�jL��������5��)�6�d�OԪY��c�p�aG���e�>*�/vs�I!��#dz���#�v�7�^D�P>�k�Yqm��5�Y�z��R�����|��6P+8�2CP�H�
(�$���μ��z4 E��6�Ct�/��,ν���;F~�Ӆf��4���y�9�f���5�Л��𰫈�*X0.>�+��Ov����F��iT�R�!�y�6����m���0�՚PW�q?�:���޻��9���<�����6oY�oބD2�L&#���h
�C��d&�`%�;s挤33c��,�9ugΜCgW/n�m�hE^x�\$5����Yx衏�������a�d�<������������+�Fb�v�Z�B<����N6�ްu+Zҭx����H��D�k�]�������>dQUJ�2��_�Dc^�r�2<�)�@.]�k� #x��N����D��	���蟩i���@?����$v����G�ZB��P��pӦM���|�W,��{����K���G+i�������V�wt����C:s�����ؖ�&1I���<�C@�y�qw��at��h�ő����EZ�W`$A�M�q0��qO����������&��߲�}�sh]�ZhV�f�*�ڭԕ�{��p����X��zmR�b�
c�8�o��Y8#Ch�,TkL�.6oƶO}m�,PP<y���?����BׯÎ�~�[� �)Q��0l�9$�j�������u5�%E��,68�-\��7w>���~��X F��l��ŷn�]_�2B��A��Y<�O��[�?��K��l�a�7��� m�Bq+W8u�SO}Y��j5U��Β�v�E�`��G���|0H���;��5\:|;���GG���>��5C@����i�|� ��g_C��it�9�,��Pp��q���F�r�ݒx=�ϡd���Dd�����pp�;�"�׭7]�56��_!_�ٳ19�C��>,�?[tãW��������D�lU-��C�z�6�e��6���Ė��c��u���P�3��{pA	�4�0�s�Jp�c�>���	��V�Z=
��tZV�(C�Vm����� �o?ݰj����h
����F}������>q9" �8��0r-y���������S�v�!z��z��*^�h�� �oґG��Z�D�PR׵�nsO͕��e0�4��ʄ�i��z�C�\����9���UZ�*�ٜ#@�,Z�J��r��K��S��|��ZQ�m��v�n�eCYf��Ţ�X�f5V�]��H�a�R-ss�Q at����3[�+i�� F���@,��T������B��e�/�	��~��_~����mD8�
G�oKH���}L�Yή����Ǜ�N8���$��?V�m���e�4D��͂��Y@�m	���ͿpR�n ��F�,Z�h[�W�L����>t͙��7o��5+�ӞDK:�P[Z��|o1�s8}�,�*Ϝŉ��p��i���(�F��jUK6Mv�`���+��p�'U�zm�}��*咠܋�::�3�K<�)�,�'�/d0x�"Μ?�����h0���4�H��+�? �j�dSK��M�3���DSч� P���ρI��*�:lZ�|���Q���t"|8
�;N� Q䩻��c�������� (�Ů�V��묋]46]6S���5���{�w9�*J�*�(⚅s�/�:�Y�z�ry
�C2�io㓟�_��믿��'� ��#��e^��ی�ہ#G�
(��m�=��ϑ8�c�e�$Y̗p�-�"3�A�@�L�=3���.��}���}�]��ɝ��D������G?v7��}o��&3e�\��W���d��܃�<����M[�I��o�.t"�	bf�Ll��F�8���.�
y��j%lظ6l�1�ǿ�$c�Ln�Q)�xM�6&�}�����697U{M1� (��k�iR�s���İ��a
t	��$���4֯_�/���b�58��p�s��E�tG�h�������鴢zB;�0����jå�JE�����K��P>lH�>tDbh�����۳�BN&��8�lل����j��@��Q<�w����Dq+�]������Z�V�b�!@�ȑ��Y�kK
����t��L���#�����Çp��W`��"VȣP��]��M[p�g����� ���a��O�G�ލZ���˖�O<��1^�0Q,¢�z!Op��q�Ԫ�� �I�,��}�D�w��@nh�v���}o�'�mWR��^�}��H��(�p�2��?gv�B�8.�`�-�����[p�Z���ȗ�
H���)Eƒ�@�<���&�-�%�5,�Z�&b1�'�9u'v���S'�d3�FjN�����(��.\=z���_�����5
U$RX>W�%�'iI��i�������(UPΗҬ�
ۭ� ����p\B�2�Yd�y1�`�Hé�V&�L���m3��޿U枔k8w�^y�E��l@�@[:�E�����o��M����ڠ2O��'����@��?���󉟈�bժ5b*��ذD�� �8�P���ٳ�b�Z,A,َH�T#j;\4��\�2��
G�*�����/�)��D]UM6e�K�J󠦔�Ԅ{&����ʁ����z�Q�f�j�k���X���&Z���	��8��sO���<,����!�r�|>^�,�yn9S�9�We5��;�&��MY>���rl��e��y<D�M-�`����p,���0( �c(�
�&�A���vu`��~��t��--��\�A���L�i	���t�n%���P~��M��c�'R--_�eN�/VO����o_�������K/�W��n�, 9�eG_4��<7#	ϖB��p��S�bv��tTb��G3o�q���N	s���Z��|�-���!
�89`Jl�B&��H�+UP+`WʲhE�P��!�.#��� �3����m����AG0v��!d'�A]�q|������p��c�ٓ'p���C#(�-���P���P�&�E
sڑ�͑�Th�7I�I��M�N���j4�t2���4Rɘ��Vjy)�����<��*    IDAT�
�2�ѻVt��U�$��&��X���p!�Ő&��cE�V(�K<v5�Y�
;���#g5�gQ"3Kz,ǑL�IA3(��Kxt!���`h�&�̒���bRK��c��)M�MV�� �F�z�c���T'Յ��hL`�@/��ﾄ'�܉7vP��=���q���B�ٽ{��yL	�0����u�ؼ�&<t�>�<J���բ$mҧ{ݚ��1K�EGG[[Ba�����y�q��%��g�t̶߱m�x�g�HA�Қ��ի�u�ux��W��A^w�fب�ȑ#8~�tV�e��|��9X�bV	?{�eT��,^�k7`xx��څj]�Rȼj�J�?yo��W&�2��(�J'��-R���$fD^8�H ��Cy�5��5���<�Ͻ���k��@��<�h�,��i*�(d�$ (&d��D�/�/_�ڵkp��^|����{�.sQ�J$��GK8�xDy�S )@ֿD�o�QǤU@��u�!M�h�[E�Z�a9��>����D��4�&r��D�f	~?��mh��V��p3г ��q�}�i���`��YXv����ݿ�it,Z��re�m���#B�M�+"0�Z�5P�3
c����ԺSgӂ��@irC'����wd��͡R)cЩa����ӟG߲5*,����/_û�_G6�A�>���6�\�E:���c "��C1��M}�x�pBMDWeQ�Z��+����S+���\8���A��Fg$�`K
�7a�'>����B�� ���so�	��A(���5����<��4r%�����h�)�S5T+%������PR�H�29?5	Ѣ�$�*cp�1�a��`�����]����U������
���>�B]�<3����?�ٷv��.#�*�I*HM��
b��Ty*?L�NG�B��N2��X
����%�p+k_��C�����g^�MK�T�3z$�l�ҕh���/F�N��sO?#����	��K�]�;�c��-�'Ӓ�K: �Y���+̐I/���~�����'e�uq4�=�R��mTP+��0sF'n�~+֬߄3�I�����{q��^��+#a���	QT����ҹ�Q8	S��L��pD�?$}���@}�Y�z��O74p��
2�f=3�,a���ii��\U�-o+z�8-���*@̕"��Qgũ��@�-�N����#�[J�
W�\�xo�}�Tuf.��Æ*}	���&��İV�-x�Yo��>s0�C��x��8&ѽ�L�M�A��q���E�[�/ZF#m����lI���L4�7_��b�؁���������Gė���Ĉ����-�(x��w��%�%(�఩C�x��Qĩ.@�?�>P�YU�r8n������p,��ga\,��͠V��"(�q��� Ocɦ���{�j�j�G/��71r��W�Q��׻c`f,_���}812��abdW/]���0FGƑ)A3����(
Rz�YI��M�O���]�k��I�>&bሤ�ƨ{�(�Qȉ;�-��:.T����1��Hׄ

�����'I}��/�Q�©� .l^ǃv��B�+8��X,�T2�X2�`,"�łP��>T�^}�ڊj@$�� SX�<n͛��(��RO4(�������BM�RβX�����_��]oa��#��(�
����zP(�q��a�={3f�����ÊLtvt`�(�-:tG��P�����$��D������s8���Y�+Xn���nܸ	+�-�{�����w��̛?�7m�"bp��ٳ��x�����!ڰq�-[�KW.���Z������q�
�Y4�ի�adt�8>&d#��N�>->��BS`xYGw��G1t5���N�8���IU�QA��K[^o�#�qs*fS��>��5HS�`ڙ�y�$�]�zL�Hw�Z���ȅ�W�ܰ�]-!79*��2�6l�����j�r�ڷ?��?Ga�n��\,h���Vt�y�k�]47@�i`�T�8�Ιg@1��^*�-85!�E�BkP��[��ιx�+�6'�GɶP��;���\��ta��9��������/��?l`�k���;��3Ws�u�imkA�AD,��B�4��R�h}�����Z�=�zQ������ǎb��Q�-�JI&�?��;�������@������K��{�?�%��8:/C�� �TZB��D$�6P�Ov4٭��
k	))�$U�\Sy3�*�to�dQb�ʅ��_<���M$}��gl�w��o�u� ��&��)������0���p���E��7��C�fT
I�'ZC�ʚǉ��Ӓ�g��
,�l4<�Z������D�.��A\9��Ǐ�R�@hF'6|�a\��O�w�|i���㯿�N���H�dQF���A2�6�	���k,��pn����%-�4&��(���$��������4-^��k6bƢ�̰$y�8^��s8z�]ɍ u�=,_�w�}6_w=-*�̡���3�,`�������+����O?�L�$�bs�gPY��z%���Ɗ��q��`��U0Ci1������.zE� �ɇr�[�RI��P��U�����Τ�@��x�
��P�PĒ�����bT%�{M���
͍'|�6m��Sӆ@pJg��M2!cr�؁M���}I��n^��*�T���{���I5F<C��Q?� �~�j�r�<l$	���?>C�?6I��9�S�L4�dګ܎H�1e{ΫL��M�����Vl>�x��d*��	
~�����G�lq�h~����ر���/��@�n�ɱc�|�t�
��٬i�Dc�����h����ڽ����3���L8�S"2�fBG�;�� �Xp��8u��Q��p�
f�������P^t�I߼���b��q�i*�d��I�9�:�1X�<r�#(f��wm�C*��#K�	�	�q�����O?���V�~~'�?�$r�N!U��Q���4�Ӎ�e�ѿa=ƃ�L�~�.ab4��d��"J��@���T�2#1'5)��B	A1��H�����E��x�%��ꁀ�P1ݐcJI &-��&�:e�*�|M�7�2�Q�b�@�ud�)�4Џ����V0�ت�e�P����>]-8���礠a��p�%�%��H�.KAq\"wYۭj���(��lDeq5=�����\(�M���w�zm�ɚ'DJzao~�4eH'�*g����y�f��ݏ��$��2��$I��F'Gp�軸|�
j�:�͛�ukנ�%,ɘ�bV����Gp��y
�֯_�E���<�3r��;�����s�OmJ��<r���3sg����D\���~��~�Z���-���$�=�+�/���k֮DGgZ��L��A��q���n��H��D�̐��'������32�O������ʵ�{V<�?����qR�&���Uo�8;Z����&��*�?�Q6�	N��]���Q�c��
h 0	����
�FM@�,�֬[�/���`ݪU�D��׿����ٶ�S혙H�5� :R�K>3��ydje�vٖ�4q���3ה�Y�@G0"�����I�ԅ~%̤s\�X(ϙ��O=�^D�1q�"�����w��@��`�D�'����!>{F�uTm��]���i����lg��̼�9�P�@sJ ��綡�q���ȟ>���5A?*�(�>� ��� ��^TF����O`��I��&v8��fg7��]Hv�I��M<֊�^��z�I��Gl|�C�������=���e��Ρͩ!$!��֬Ń���aƆ�@������:��܉�䐀:��~��@���pJ����Dg��D Ezg0L;M���9�:��W�2T-SSE�9��\�o�D��MgN�89�R؏�܇z�T?�����y�)��E$�
"&{-����H�b�����+c*7�b.�sl5>"Dѽ�����!N>6���*E���$sܢhik���+�p�Z��Y�E!W�����ӝ��ؑ#B�`/�=e`�ʥ������ƛ�("��i)J�$���s2A���X�r����d���Ƞ^͉�i[ԇ�߀���.�턑/5$��B
�I>?g$j U��:�ù?q��1#�{<�R���FM	�>@7��ԑtN��o�0Moᚠ�C���'�͠@O��i��4��E��jJ\���Iȝ� ��,�*��F����Aیj@��J�qZ�� B��SsO�E��b�	���������4�4h�A.f�Ps����h5�W�f�<Gԓ�Ϡ6l�� I!w(�x,��Q*��"��Z��!���5�����HȬT����U��ޕ�8��ڎ+_�,��uc�a�Ð�z�͑���y�r�������P��oF�l�����y�����} >N��t$}>�iU�4�&�����^��\�=Ӭ�F�4M�g�͆�q܀a5�o��=����L������͚�7M��q8���3�!�4�N��+�_J���뚎��Q����rhU�������K�;f��07��ZR(��a�?B2�F*���K�E"S�
G1���{�܄ʅ�t�)�і�-!7�He�..&74��&r�Uw��֤y�]
�S��3���Z�Q��012���|NɈq_PF�V �?��~�~X�,��ǅ�^C�TDw�r���Đ��=�����Dń`ǏÕs����T������E����EMUr#i��D�&W��0�=���h6��I���-���$^�tp�T�2z��]� �g'��`J���:�M�X�q����Ґ7X�(`�Ӯ�ը��G-�C�V�M����f
±���S�MJ	�UD�G
>H��szR�;���)'S����k*�����M<i�Q���͋'z�aʥ떑n	c���M������8�]��B%�l)?�%}L��aɢ�X�p�p�9ɴ�� )G����p��q��I�<qZ6���MW�PoT]�LI	°�J�&&��P4 t2&`��f
j��O���P1v�UWV��X���#ŵ���En�t�j��:�D�p�gv�xO�Z��Fj��C��h��UK����ˤ�)��.����nc@4w��x�}��������@6=�#( �o(�Uq����@17.9��Z����ob˖-ȟ9���M?����F[��C1����tlª�r>��bE��!����M�z]��� ��Q�4��Ii�<��Qi�y��������V�P��;�>��|��ˉ�y!�-@�o&����A����ʻ\6��21$����B!���Eξ4h���F.\����?s�� R����8v|�3Xr�@[r�.����N����$�=A=���J!>�m��h�lEό^�����x��z�	%y��.�2i\Е�S@ޗ|l������}������&M%�b�羀�w���
��ַ(��
�WG��b��`��U��d-�����lV� K��y��W�uk�U��Z��r���������$�"VϘ�>�?Ɔ`W�k���NM���>����{�~�Q$ʓ�;%NE�'&A��N"W�H��gҮ������/X.4-h	#��#y�����#t�*,�	 ΩMw��^��e+�=o),3�R��Ç�Ó�>���K��v�iR �ޏރ�o��X
�bu�'nL�WP,OP�&0>:���x�?�MG �Қ�ƇTKh���vˍ��{10	�5����9�(�d�0�W�&Y܌�o�PR��ܣj`H��T,4��h;��l�k@I�*���T���k\��Ue��PT���\�b���9&zŰ�~��S��Ԑ�4P��kP�V$���ԏ�.ٗYlMY�*s� U?��I����
Ш={:oax�9QL.���o (Ng������$V��G��ֽ}�bI����_k=�T�MY:�I�g��3����DG������?W{���
��.��:�Zi��0z��m�����v����a�8�U��������َx�ѩ�5�?*����I�D�0�n�pL�a�YS��ͨ5!q�a��wmɍ7z��>���ϕ�!%�,�*�B�xa��p�������t�����3\Fg�	�`%�B�!qx��5\����ϴm;P�[j�Y�[V�T�e�y9�k�6	��麮� ��»@L˪��* XTR������{n֢<E���?`�|B,�,�tITw`Z����/QsSK�ڐjia�,t� �IA�r�+'U���|^���&& �0�͊����(&��$��5e��'E�Fᗌ��B�d4f�
8�bN �~Ľ��F��|f��1�&�����F �����| w��t���o��ۯcF��~ˏ(ǵ������Bz�l��ǐiT�w�>���k>E<��%r���C��Z���t$�x��!JL���i��L�)z�yd�m(����)ѵ���ny��}SD(�#��KzQaj$�D�o덚�/G�s�L��0i���c{Guk(�j�(.J��ǽҘ O�%ނh".y�}��Qb�U��Z=Cg����'�'��4n���T��C�(��@�9�k��f��DO0��f�dr��c8��������m����LȄ���r�(^�t��6)]��R�H]B|X�ą�wR�K*����Lg(R��獲����
�C=N	�iO��A����fX��X֙&����8W?����� ��D�����Md�"��I�ұb!+�n��'���O�x���Ǟ�iAWn}]��,L^O� �yc�S���Ħ͓`�'���5(���Q�Z�_��oc��u�dG�ډ���̬�����{�T>�mc�R���h���JI����ꆅ��� 
�;G�R� "*UhB�0L��R�Z
#ۚF����e+�֋�DGw�ģ����D����(�}��Ē�[�7o!b�v^�b(f���/@h���A5$�5CZp��F@%;�ɋp��q��~���ł0�ݟ���� ���`grx�����?��d�P)L'ퟋ��^�-i�/���y��ퟃh�S����{����?��k�<&\?}-�T���4���=o��o�-F�����(��b�ǆ{�/�"�C�}�y��+p��f��8�����ߋ��Ũ�zv}Rl�uDu�R�{��ü�<2\���prJ��b�
�P�58����h+�neP�Z�ۈe��	�g>��������^<��0��
J��B,�����臅�Y��fV,A�T��dN��������,{%��y�����p�Ձy�o�l,Z��������W%x���^Ʊ#�
)h m)?֮[���s6n�$��DS7 �H��S�i\�.]ď��/��O-oժUhmoJ����(2���
ٸ�歸�{��7G��b��xCR���e[�(���H9Ɖ���6O��^#8�ѝ}�<N��yS���o�͏�.�-�.�ɘ���Wq�X��:6�Q�KG�k<�ƘZ�������^jN;h��u���
y��a����6�Y��)�Q�Z���8��N?�F��[�ʿts�ݢ�Q���Bݜ��V����)KY��4}ԋ�j�`�nPm!�S���U�Μ�o������X���4(�f/�݆s}�R~��h,uvڶ�(\����;N����}1��&�4\�y�����)�t/>��&�H��$B˥�T��HG��a�A+�<��"�{�.�i�q�-���d�8r��Uǘ��*�/� �!�:�Gŉ+N>N� �J���nb�d)dڬb��Ƭ�1�W.P��&��	:��x1� PT_���������(��×�AC�z����C�h�E"�FKk�Q�<$7;��(.fP-0��P�	5 �`2&-������(.]Bf"'h����E�fa�y��[�7ԝDv���JDA:A���&�k�Up�c`xW E��uw�-��3Z�ʓ?Ʃ�^�s��&+7 +�D ���.�t�}�^�V�x���+Pp�l����{���M!l��?P 7��u     IDATX�q!���]����͖��=Ȏ�X�i��m}��u�*�=����HKB��)`�+E�gՕ{��Is�Ȗ煓��Z�
�Z����j�E��@�qQ�k�/�S�D�h
H�Q��7l����O�K����:���T�a�����z8�4TyS&�~���������9�L�P^��P�x_�\4y;��qH��TP<��6�fIg�Ŗ��s!�d�	��<ę����rIG���N-�Y6�G����3i�� ��i�|d�h�	7v_��ή��i'NL7��dP�}0�$`��F��*�&p�6TA4�D��D@J~
9�u�z�^ �:?*7@5���=M�Ҡ@[�6�i��<�iZ��W���AM8s���٥��˪���k���_�MlX�(�1�ҋ8�ȣhϕ��"F��(
N�Œ�C�Y��-z�)�߰j�H�t�)PԡH��X�/)��H��m�)���h�O%���{��F`�\4*ο�"���?Am�
Ba?&PE�m�e�Bl��~l����Q�G��������r�P�}"Wm+�E��8m'
�j����~���>�d����
������၇�;N��ןz
�����`���A���KV 50H�0s� z�z�hkG8�	�|t�PU]O�r�r�y�f�ˮ�P��W�:������#F���\B��37l��k6B��<�/���\9�_G�MW+]�;���.E��JӉ��;ٿ%�E�)j��p3NX*��,̪��2S��E\y�m�A[��@����Fx�*���#@�B�\|�)|�)8��1k(Zy4�Q�����7�{�*X��o��2؀��q��e�;s
����s'0::,�l�l,y�_�A*G�=���Y�럃�+Wc��h>�*���n�z�\8w���H�ٞ��E���~#-�[Q�O5)��j�Z��W�����=��eZ_���n��:������\�i=������IA�Bǡ�(p\6 T�j��(�F�7k���).�ZQ��~Y۽�N�4�����n��#�g�[�iF���¨�%�2T&	S��Zg*�F�*����ż���=���a���Pi�Yɪ�3�uNV��z�=%��RT���}��ғR���ʎT��hꢛ6����d��z/��U�u��Y˨�b9�Hsem�x� �j�M�[����������O���e3���z��ڢF�
s�'1U�lxa,V���)��I�θ�-gς��4)>�����L}�^�����"I��u;�p�<jW\X5��@�T!3]̨Q���7wu��gT�[vDH� �K:�2��U1w�m����]qz�7�0	ҵ�v��]	��u��t���'r�O1����U" a�K�܎|^	���?C1(R3DCa���N���>C;7vq� (\M&�D���ޅ(;U��Stl4Ш�β���$2���*��;��Ό��aph�/bd���
�~�P�b�F�S�u����E⁂\~���ud�1L�'��e&�t�.´�ǣ(���݂�?��X�y-&O���{^���o�~�,�\	�`��@r�b��gR��Á���SOc��{01:&"b���	$A�~�p�p�c���KP�{v�t�<��HJ_����S�7�B$�n��9������k��э��7����s�)nnC�.w�#���2��[櫕�k�8�n3��o�Lo�J	9�EI&;�$��T����0���^0�BM߿�}��~n�_U�;=)h^`�0�4���鍀�х� /OЭ�0���i��>4�)�y�d��Ug�롌�a����e�����Rԛ�)�`�sJ�ؐ���N�%M��h,���S���p*[l�AO��c�씪%Y�y�E��7����e�+?Y�U�K��������0}u�T�>�*4D�ȱ ( �7��F�fA��b� �1��x�o�՛��z�Q�n@���s��9E�&���������y�cu�U�_�\�M_e��6��RКC��Ǝ������_��Z��Pܵ�z��R�Z?�D#�.�g�c�.jj��nz�U9���	�p��ӳ��AHm25�S��u�?I5w�#M%��k�7m�J4�ؾ=��?�L�9�){f��*�/��7�~'��8
<�\#d󦑀7m�Ē�*U�NxH��VHټq&v�"���o�G~�X�"��	�����q�ßA��@��^£�������D���h]0N<������Պp,�H��XR%KH�2TP���AIw��L��
��u{��dϞ����9�T@��˶ߎ�~������P��o����m�?vn�B=b"<k�߀[�~ 3,@@�3��x�Q�͂SANJ��ٜ������h��:�Ba�/�� �wb�,�4���Z����t}h���0�w��Q��2Jf�.�޸��^��ο˜P�K��Pl�āx����ۯ��u�nN)��\�Z�H��eb�F��ٍ�����%��ҥ+8t�=?r��Q6ט"� ���X�v����ۻ`!�s�� �4����z�'���O��f�|�r��I�8���5�q�m�3Q�R̩hh
�j����t������H�N��Pu\s�A�����Ԥ�����������A�{�����UY����=gS�������\x?�G��(�����4V����hj��BV?w�:��p��+�{��&�
�8jP �C�Tִ�]����7!���׆��R�#�<��6���*5Q����'��jH��P*��t;:{�=����b���oan���#}�^]Y)��sݪn��U���ڎK���U���>��қ���>��\M�~�S�<ׯ�/ʟߔx�*:;~��^̪hP C�<�<�M]4����u#��:2��9Zr	uF-a��T��Օ��~^'�"H�)�R�W��y�Y�S�-��e���K
�-�A����/F$�P��ՍD*-�7���j�����P��`)2����'���W��D|�	
��( ���F���� �����%�bG�� �ڙ	42y����a�|:��Q���y���O}
��N�5�������'_Bu<+I�3V�Ċ����;n��� �~����|��I����>���A�xѰtC��J�\Aį���[ѡ�7�}�K����"(���
D�<��B��a�|MY��5��,�r����\ �(�#!��<��@�����f0 �ȫ�"���|C�_D�1�����Ң(,��V~�(��g9��`*�YX��gP������"R��	��W�ì�SL/=��I���,\��Dc�/m�ř4ʄG�=Ny�H�G]�w���T�iX:���(
��g��jM��x�T ~�η���hI�Q.�x��E\�:���V�Z[�`� ���%8����>|X�Q~�x"���}�ݏ��6��9ѻ�=}��ZZZ�7��,�#�0�b���A?z�lEֈp������?k�;��'�vT��:������u� O;�ρ>��t1u��ހ�W �����k���&���u�������/}����/�)�R��X�!?1*֝�n؀/}��XF�Pa��_�՗^AhlQ���5j.�1��D�ހ��ɘ\�ގ-����ʄ�#Ew,����qrig�*�}P��}�eV����?�L:�؎ې�u;0g�����c��}C�K�Z����H�[��7݊ͷ܆x{܀�tUv��4-�o�9y� "�"�\�
��EL/�|?{��8�ҋ2)�F��f�f���ϡu�r*cqa�>���j�C6b�mH�[��y���@zf7��r�lG�a����d�-׀�O�>F;k%p��E�I��|���;wo?�#dO���� ��wމ��<b��P��|�v~�xw��p�u[㘽q���ڭ��m�|yv�ZI��scHm��-��f�3�2�Q3���� 3!ct���1�� ʇ�E��y�E;Z��nfܲw�r���d'�O"T� �`�]�����o��h�ه�B����&�L�\��=x�>�8N�;��Kaٲe��|��#0�c2�ݝi�gFE���J
�g̝���`dd��C�<��I�&@����/��W�F{gl�z>6�"R�	I���|�)<��162���v��Z��ʆ���n��-�z�&��N�ڻQ��������뻩�M���Ҙ �fjJ�?y�4�	Sk���+}�t�0�����\�+k�.�����d��Kor����oR����K6\��O5�Z�~��$���i*�گ��@Ӕ�g��O�ÛT)a��^V�j[��J��p@�9�L��H�Y$�0�t\.K�C������֌�W��eThWDC5��N�/6x�y�ed�������3�6S��}�׿

ȃ��3�W�Q��8&���o�&�Yor'��/�4���;����.`��;�S����Os�y�z�f}��c�#�����$�c!.<<9^h�y|%�/�c�)�������Y�8J�n�]"���}��Kowr��E�����cIР6^]�)kPZx)0�tNL5��E�@'0��\\"<�*R�oiA{g��m���DDjSq9�P��\�`Ej
J\��ȧ|���"��'q�� �3y��݅��5a�y�%ń�(}( (��<<�E�S�l	1&��0]!�i1f!�ځͷ܌��߂��$rW/��^���_�Y�P0t/^�e�o��K������]8�g/�3*j<h��:�#p��&ZZ�b+�	A i6*�M�����SU��C�F��r>$gț���v����V��2%E���40��X]V��/e��^G��2<�HY�u��c��n����:��HI:�i�9��`��	��"A�k ����[�'�����EZ� �	�HugC�kU����N�X
LXs�� ���<M���mިT �������\O/[�eX(��C �s' Ϊ"���;o@�����O���A������gb����`@���><<�H8�r��=]�}�6��Ǒ͍Jz'�}{�c�ރ�#X�t�/��d�i~�f8����xe�DJ:v�,Z(����#ϳn���ص�y�[�o��u�1���(������Þ�H�E*���oƜ�3��o�#�7�[e��=�z�ղ�y�@oN���SM��k��04��9�@�_8�M��� X6u���m�5�`�AF�2ݱ�m)71���`����/|+V�Ʈ��+/�t� ��<�be���j�z�J6�:��
�Uf�z���P� Z�A��È� g�/ō���'gŀEOyr�9) J`@#�) ��7m��w�X�R:�t����+\޿��a��$f�Eߒ��b�g�F�nu��sd�9Sb�����,���<n��G ��d�N�Df�
ʣ�8��m��{I�����>��Y��~��йb%�*�=s���`��	�\��4�3ѱpZ�gß�IN��y}�I�To�~��&E ��,��k��/C�������GN���c(���so�c|�ru��7݌�~�s�b�_uP?~�~�[ؿ�e�R}�Xq�Mwva��h���x6/B��Ȑ�y����1TK��q�4I��1�!�ڊ�t�h��¢=�p��Q�z#��(��Ճ�6���m�?�ґs8�G��h���T"6�31瞻�_���G��=O�z��K��L���c8������*�~�v,]�B�P�=�N?!���s0wN��GŁ�a�q=�9�b��	��9Ѿ|�<&3C����6ZےX�bV�]���^�l�5(�*��[�ɰ� &�'�ܳ;�ԣ�`ltT��X<�:�Ř]-"6���7ݼ�޵-m(��:E'�����c�BmU�7,Յ�g4�%�1S����9w@��Y�8|�z-���~.�����l�1��U٥I97��.'�V�b"�G��SC�ן�j��k]�8u�뉌�^�ez�@��Q�L�ޅ����OB���H�g,����(=��[�������r�+u�Er����UcQj����6�[u�/	�3f��V[o���b����u]_���H�R�Z�V�Ga�C��t�+��֨Ioz��AS��B��	rP�P�l����ԏo.�������8Eң$-x�E��Y6|e����)g�#�|���H����B�Po3��K����\,Mo�
)R���h�"L���Ք@��5�џK7j�R��57�!�vvD	����ґF2�D��x>�W�l�ݢ !`�c�eԴ�*5��P� �+a��(2Y��]���(�>q��Vr�o�b�܄,2j&1F�Y�ry�
��*8�+ ܡ3@�F�f�h ��tϚ�޾nt����F�(!N�o��<�q*'��3g064��ȨP��]a�Vb� �aR�,��ܰ��D�O�&eBhoJϡA���x�'<^'�cv�^C~�4x#W]�<�d�Ѱ���a�kxI�ZtL�J5)P�!��
�u��;+�,��o���s�$���Ȫ� ۨc���D�A�!M�P�IA[[�8��i����m���N�ԓ*]�4���WT����N����}��D?l�������pC��kC��s��׫����ү\��W.^B>WE8ځKW�p��i�o޴m-X�p���]o����=�P0)�zOW��yW��|�z�Ә5k�p�_ߵ�%�����%�|a��p���ǳϽ,�$��uut�����z	��{���ur�<��'P*���щ�_z�RF&kVm��?45/��*N�>���n��&tu�㝽���{a��"�k�&7��Q��]iP��;�0��@�{�5,���5Y荛!N�ܼ��G�T��w��T���?��u��a�l^�_��ob��]<��^x���H֪(NL �� ��P���){4�@��Ć���"���D$�@��JZ1�h{,E��!.F��)��M���1P��0��a-��q"����^���u\=p ��J>��$�� 1c&��v̾f!��Z)�Ci�[���R�[B8A<�4
XC|����݇KgO�,W`��>8�T���PUN��.ÖO�*fr���_����?�Ń��T+���w��s��LT��,L�gV7V�Z�X2.�GN��N˺�7��a�m����ĉ�"ᨸX�<r
��C}h���h����@.���$�`ֆ-��D�¹�^���{�(���L�[�r���@D&�@"2�b�dQ"m�+ɶ�YϬ=ci<���3�G3{f�Yi$K+Y)�Q$0  �� �3Ѝ��Օ�M�����]��<�9����!�]]��{��}���G�x����阷n-��m�=嚍�O�ʥK������0"��q�_+�_ЧꏖL2��K'�loEk<�6-��~{���Fn��v$�^�Y�lKY�� .����߼�T� ˚@5dюY�>}�J8�n����:@$��zԽ���c��7���w�=��<����D~��s������BiY���{�`lx��J���K�Q����I���@��y-�ǡ�Mtw�a��U�s�J���64�t�
����U�S ȕ��]���嗐��@������ ���'F��ժ�Qm�'�1�wS�w�;�vn��ڱ1PM�G�l���n ��F���������y��I���!�����ԀhP�C��$>^�p�m��ړ40�6M�*@Lٞ@��)0�k^��6H�Y�t�&�ݫ�Zѣ߫�9��d:��.�	�c4����F�TF�T@��5�(�5��JЎq�4�����)�f�Rf�futO�F���O�YM�4,���Bn������Z��q����8�-�+�쟚`���K������D��+�����z��	}���=����&��Їț`���Hq��DA�$zIx2�(�����|��@�zᰘu�(nk &#w2�]�^�p��DP�I\U�M"�-�<}5�P���f    IDAT��4��9Z�gu�%6��D�H�LR\R�$BQ��ҙ"V���!�Bn�bcN��T�RAn����1+r�Ș�T��XT{7,9��_d��t��Ę�<H���>��\A��,aB�����7,�?� ��,\�H��f1-��l��b׆�pi�#c��z#7n�W(��9��䳑�ˇD�;� F�*'�g�M� R��*0�`҂��*�z��$�G�1���2ire��5G���z��U��t��s��3y���o��Qh,{z?��H9)�1�!`��YX�r���{����k�n�l��Y&�
E�E��W�ѷ?"�N
X����zԑ��|�6���{�K%�Vg��(����E�=��0���f*�<�+Ȓ��������ɞ�j
4}�B�i�I�u��B�q�g����?������004�H�u;$�D�tӺR�׊�������[�QdK�Ɇ�G�:�t2��w���U�g�;��?!:���F�Z 7@ȿ��� ������lq�{�ct4�l#�/�HboKK����v�?}�ul޴Ct??��0QAkk�W�GO�)O�9�i�l�|7�ww���sx��i
x�	�\�����|�y�x�Lm�j�����믻�5�~�/�V���a(�Ks�a�����	��ι�ܡ.�&�Nsȍ dXشf~�����W�z�>x��p�]F��G�ni�	4��s��&�P�GN�"���_CW8��`->?B�B��$�L��81T�N��X��dt��6U��A�%��܅�>
_�rA��=�W��]�/�G57����xw"��Q��Q�7omŢ�K	P�1>>�j���&���������B=�K�S$��p���!d���F�0�b���⥟�����g�x���#�������G�E��I$g�Ez���8�{W{�"��k:�� �l
�(�����Cj�����Oj$�dRU���
��t2t�9������>4s�Fht��U��;�����B~��1��h[����e�q���y�-ܼ~�rNb�O1Ր��$,H!��N[�L{��z�,���k���ȝ<���
�g3H�]�����Y@�(N|�ۨ�;�6��W��ё����C�S��n�4'(�
���+g��x��]8z��_<�=��Ђ��_�r�he� {fa������8�UC�Z�d
t��ɤ�Xȣ�C�0��A��L��)!d�HF�/c!�r	DO�����1��{7�����0�����Ƈ�0�8���+�)�vNC�����u�b��(��m����j
\ݒK���~�|Ҽ���r7�v0��v��C8�(F�5��Q���{�n\E�T@ȯ�Ā���ME �6H"XL��k�u�i�{d��F�?��@�)Z-'l��s��� 5MS����:^���o6Ԗ�`��Ȏ��A��l����nkoG��.��)�[r�"
�P���"u�}߼.$PΥ�ӑ�t�Tk��e3��n
�?ZӖU�c�K�5F���Xf�2����t��;nh��#������h���S������qt!r�L��d�H~ˢ�'� �qZi�]/�$$�P�$��#u�{��{iB%����ϲLѢp{���E�I��0����@�!jk�F�"��hX��=��a�����(�$�A��t�Q��`V�2^���*!w\>�CgR�1�ǉ����z  jg�0�lP�����+`v����{� p��;�����4iS*�ø�ўL'�>D�]2(B������D^����A��&�Jİ6D���<�+bp4'i�z(�����ĵS�zq��h�:_�7�Qy=u����X�ju�j"&9�&�F]t!Q��(�S3�Fr�4�Z� �7�ê����֢�a�Y��
n��
B{��y�x�]_�,>ߦߏ��1�@�f�z�SW� ��j�0,��-���e�-ad���+��>2YT�AnJ���� P@-u= 'R����3�]6��˨э��w��V�h�5&�=��1{�L�[��pb�^]����8N�-���
2=��ae�jAKK�4\d��Z�P����g���k
��	�3���ro�I�1��idqr�?��=>hs��!��4A���k��'��[}�)�GմM��<��`��t����S�¹8q�4>-��襟<�2t��M��J8���}�����Ec�G�2��Ts������c����@A���]'�"�����v�zKU��ֻ"�fQ�M�M�eU�-����+�_x��%l����'��D�,�^l޴���q��Q���8f�l��{6`ά����A�:s�FQ{X�CL�T4ӏ"[JS�(A,m�K�&���@�F~;�Ǧ��f�Ƹia���N��u�5�5�,6em��s��M�}^(�!?6��i��5k��_�2V�^���+����Q:�!��!qL3H�;*�P�S	&�����&R��%�V�c����8�8��E[�<��L���X��v��^���3Q���[{���@�<!�{A��V\�Q��ed�Z��U
EiR��	���a��`� �*�҂��n)�����ѐL������Q��Ĭ9X�䧰���ԩ�������C��A���q�ħ���[�8y�.\�(�yL���K�h�M�g��m,�M/��(�y�4���jK#Kظ�Quˢ%x�7����)(�G�u\<�.4��`LG����2{�6�{�0^~�U����ќ�ԃy,�TA��b%��vYKHv,d�,_��v܇���Ѹ5�ڵk0����[�q�z,�� ��	��{��F�A֨��O���QI�1���q�=�N�A�B�C��YZ�o�;tｻ.~���a˃;��ىZݑt���a�izz�a��n��U(K��D���jddׯ_Gnt�ZY��ޫ��:�̞����a��B׭�,�H�Q�R�RK���������=�E��i���Z��|f��epϦu�����6���*���L
x�҅JD�����|O6J�˽��l�4������XL��MSboo��<�Գ��j:�Z�c�J�ֻ�������`�LsZR	i��� U��@�ǟŽe�o9�x����8�ݼ?��,�As�Κ*׌F����#�,!���6˵� Z"�B��M�����f��t4t2MD�AC�\;+׮��u+��=պ��D	��i9ew��)�ȽT3�9C��N$�[�%�g���;����)�8�-�*�F�����ˤO�k��й�t#�~)��h�Ƕ�@@o�l������Q�s�!ޛ\FfVeˊpzB��:�n���o����n�R�{ѧ�9b]�=����i����¶͠m9��ٍ`P7�d'�T~����s4�X��5|pJ�ϩ���`؁�_�Yv�����h�D`ٚf�^�wW��IB8�.��2B�Y������&�&#�g���M� ����l#����g��>�2����`�������͚fϷ�99b
�W�ɦ�a���F�V��	��Rc��&PȗP.VP.��ޒ?��P!O�OY<��ڋ7� j��udq`s%	��]$��cN���/z^�DΓ��8 i,L��]�A�T�73l��/��Dz�"�޹[فy��A����An�XV�����u�����|��u�&ju����R$�U�
-��e���T/R����Мd���`�n����Q9�(�"�|p��pV5\\�4�ì(�&ؚYF�V@�i������t'� ���N��>�W-F�^�{�v���98Ն$OW4`�g��xUR�BQ�g!��
&j��X1U��Ѿ�9�@����(��A�k��� ��a��������n�uk�Z`����ཹQ�i�����4M����<�éIH��S��񽳑bX^�T ������������%����Y����~ܳe-�Λ�˗�����ji�Q^8Bh"�9	"[�t9���O^xe����������D��ȱ��?��b-�vy�r��x$ Z�[6K~�s�='���6�sz'N~xB�����s�@ݳ�-��Ud3I�s�FL�n�����ԩ��E��..bj
li_j�B��Ϋ$�&���������ۧ2B/�l������,x�%`�����P>�zM�G��$AZ�A�l9�b!�R�����[��e�Y�
�[����gqu�^�弄_1���4�FM�;Y�i]�P�/��ҎQQZ6`�I��>�dR�(��*�/-X�������(s�����Df�=��-��.��9�7�,����XD�mkw'�X�<8t�>�tUq�C#6�3�����cѢE�L�ϝ�믿��'OI�&h�}��0��k�0����p s2)d`
8P�=�N���?���7��껁��M\9~�i#�� ;!B��Q(���ø�{M(�rM&]�BΞ=W^����^c,7*���9s1c�,	�����☕NF��,I%�͵�^�xi�93��ӟ�k7 -��[���qd�^����*��جi������`��x��0>6��χh��p!������Sn���q�~��J5�i`�]k���1��ɋ�'Тӑ��H&�%����?dg�>0�W��-��z!_��J��r@�ўA�⥘�x���)��M�#�a��\�x	�O�B�XĪ5�����Hd[��7��}0�Y���ڍR��Z��7o.f̝�tG'��p��1|�����c���\��,i>�l�r���Z ��s�Q�+'���}�W���/K�4k�,��~f('P)��R���y�v|�G��ՍB��JM�Q4��Ƚym��2YC\7E���DSu��< �{֬)�^ã�{����x����] Fݖ�|��q|����7D�$����ân��%��)��$��RR���Z/e��q=�Cj*��H3F`WQʹ�
%����ӐƯ�f�pJ!�m����Vtd����J��7e��nw��
-�V�H�D1�L��g��wJ��{+�k$�&1O�B��e�^!�6�n���-�?�n
n��"Ξ�/�>]��QvwZ0�p�my�{�ϽǱ �y0��_д��=H��7�.�I�*��}� �?��s�����m�/A��S:�&�k\}��s5Ƕ�D��Z�f���6V`��z��P}h�����Y��P`�޽��ӧ�+��nq!s��_8��ە\K!7�ztt������,����2&�6Q+��^���Z�TE�j�V�n�^�Lf�RS�4P&�Ub͕���h�F5P�\AΧD���8�������U̱Xi�hC~X�
�2�rZ��p�D�dwD�
�"q,رO~�sX��^8�A��9����p��%L���WӐ꘎�V`�ʻP1���W��.A���.Ҥâ��ځHX�X�~�ڎ��"�]w78�6lM����
�ɽ����QaO�����x�^`Gߒ;�~�^Ǥ�i�TQ���`��ڬ������3��:2-Q�[��6�E�^�;/��s��/�D^�� c���������) e!����M&$��)��(LJ�2�� nYj��M@g��Z\i�����xz#a��5 ���}_6�ۜi>J�S��)x�w��mb��&�NҘZ*��q_�O�`�R[AÈ�䩋8{������F��u�:̜Չ�W��䉳����RTo�P�!ۚ����3o!��}�.�@E� :fveq��̝�)�n__�x��^�Ol-}h�dD;��Fp��r��?�>�\������܂uע&6Ϝ0�E�p��e�����kVaѢ�8~�$�� �~x6�D�&Bv���$Πw�u�lN�)���<�xǻy;E���ی�M�k�y�-�R 0�~�~:�UJ�3dj"'��U�V�s_�"6߽��A���gq�W����A�t�e�**�A��0���j:ZlI6�\ҙ=��ᴂ!\%�](C��/-��r�IjD��P�zG��^,�c�^��wp��)�Q��ét̙�z0�s7�qmp�JU������{����ܑ@ C�x��Aix��X}>����Q�_��B����d�~tGtL�����%���d����Ǳn�6�
�����탿^�Y��hv2�D�ԣQ;sWo�b�\����5�/�֭�q�]k�H$p��%��k^}�U�3\��n|��'�'�o~�CH2��( i�qG,�i� b��ruHG�|�:ܻ�!�'ʸr�<>|�F�n���dU0�("4�k��9w⽣g���������n�ӭ�ܵ�EI2��#�՜�4E��9�|�^��o؂`�®���J	mQ�Uׁ���930s�pbY���q��i��E��*Ղh.z�&̸�N_�H�tV�����&�� �rD1;���:��/��Dm��bi�͜������t?�;;�p�ܹf%R�(���;���/I�1u�ݝظyV��w,Z$����؁Sǵ�\�ټ�z����<���Y4��X�Z�h�J�8�,aA�,���<��#�螆�N�4�S�I�i����prK(������߼x�fM������<Z�W��<���a:��\h0j��7��{�����6�����m�s�gH��d(��%OIM/����<����f�}JVӣ�7�F#�Z<MM�I7$ H`F�
�c3�5�{�A{Q׈Bi;���C�i�g�5�UK0���s�Y@GW�=��v�@&3���x�~Q]K:q���E�Re������N����G����D��Y����ppھ�v}��@�oWk��\�AU���$�V��(�a�����Ij�V`�@���,�t$P���\T�h�*4h�'�OI�S	���t���dS���7m*B[,"���b��P-!`�H�R��c��/}�#o��ŷ�`��%�%��t_5vW�oي;7���sg�֮=8~��n�������	����aA��:츮AD��0Ȃ'�	wl�9�!s�<���l
�Qx�<ҏ<]�0�JE2D��f�<N���/B@"J!lQ+��(�N�r�|l\�LZ����>��\y��Q�D�cb���T��6����񂠂��6�˗]�	����wOKB\�	��_�&�#*��z�"�,&&�n�Bk�PdO���b����v�It���m����'�fV����Kۖ�4~��O	�s��M��W`Q��x./ǝt�����\�������=�x���6Ӫ���X�J�2��՗�D���`Ȕ�#�ў�#2�8������w��r9iJx�uw��=��h����p��i�:�[�a�:���q��	�MY�v#��*�~{?.\��T"�lk+�/���������K�!b9�HiQ�6;1�r�M�W���� 9/����aS8�l�.�Ռ�5�^?�Q��W9o����D�"�=qT x}�Q��Q-��b�J|��_��w�:8�}�=����� aT	��!Ņ>�B��Gk4"������i��Ⱪ)����09��D�`�		��`S� Su���0�!Ca܄�zG��NLX&Ο:���Q$b!��P�tzK��\�B�� 3+¬X��������k�b��̟�#E$SmÑ6m݊�|�w����#�舆���V�A�H���G"��A���,^,��Ё�( $h!��T1\3��3��sp���"G�i�Bg�4<���x�OH��↟�.@D��_����|��%�����o�y���3����"��p���UE�=���Q���`��Й�Q����0Jcp�i��ԧѽp=�W_c�p���g�[g�t7�,d�w��	�+9��
j[�j���k��]?�1�������eqx�$30�8Yj�1_�����H���O�>Z҈��$�8�3��nT�s2G{Q6C�U�����Dc��$�`����3���]���5����lb��� c�y\�|]D�ɖ4f̘���g���S'�aGA��y/eZ?���^�^��#�e̛�@��QEqb��A�/���[�ؓ�@6��    IDAT[W�'p�@�*�zj�d��l
<��h�Ri�y��-[�J���C�e�s�e<�[{<��0x��M��5�{=Z�:����q�������k*d�s��|߲?٪�a�%Y3nC ���'!.OU�����n*GFESস��09  �0a����+�se�2uK��b�»��2�!�EK�*m��bEK��c(�H]E[G<�	=� Z��_��O#�{�,s2,nO�h6Ls����Z��t]����Ғ�M���W�E�y[����w�С/K�i"���=Q#-q�R>�U�yD��nvR�S�����U�@V�
%����E($}����?d�({���dSP�e_�2 
"�-�S+	2H$�V�n��t�� ��6���~<��O#�g��\۷����-5(Z�`���P$�9�b��c�Vž}�p����j�[���!"i|�N�AR�BDθQL'#jqh��Yq�e1���}�P�+��kQ3��y��|t\�\�|���lv|}�z�tG�;q��4dci�m©ذ+q�C>tw&1�5��aa��\�����,��q�A��ɖ؎.M�/�G�>�ꞆU��k
����&�D�Y4av��F�4�9��yE���Om*S�������"�^A�\�z�k�z�ա(G�+y�*P�q�J����?�(��}p��G� �'WVrRQ.�a����dSbKz��	$b��;j����x�l̚ݍ��!�����(W,��5�lDL�G0�aÆX�q#^��>8zL��IUۼqڲ�=u�/^���z�@K[۷oA(���?��\#�nن9��ctt��D:�����^�=������8��U������j��ʰ�u�$PЅ���W��+�~��6Q������[��&^��bN�NP�릘�^�L ǆ���
����j�������K,[���A|��+x�������\[��i�p�!HBh�F�� �e�Ѥ4�h49�u�����ֵ�<^O��>�~"�Ċ�p>�C�i`���8��\Ku��cO���7�(��f#gi�1<��a����;�O��3�w�}x�������a���x`�}X�p�P8yۻg�������O!l芆7j���
�%���pP�8��:Se�n��Z�(�_��Dm�z��ۃ/cp,����x1��˖��'?���$�}�]���C"Ǽ�=����!.h�������_��S���l�鈛̋%�҅��X5���4�E	FF !G]W�j#�q�Ӵ!���O=���%x�ݣx}�.��2��F[{�.C"����d�H(�-�V
�ǆ�^�E4��k�޽���>�
�C$`"hU�4*�[���i@L��Y�)��4����p@-�Lպ8@��!DaX���g�`�>T�v�Mh1���P%(QS�T4�ew.��Uwb����#�^�(�t,�LW��v��v"�lC@cƌ9h��@,�ds��U�4�4�p)w�
O����g�����!T^Z��c(�O��͊;gc���x��Ǒ�d�-�Pi|r�)�n.ʽ�vrV��xEu3��[��'�<0������p�T`�T6��^�6�R]�n�Ç�v�5J|n�6�Fp�@�r (���4�w8��y�����4Ge�d�=h4B��T��L�EK����JH�E�q.T�a`�Z-4[�U43q�����U��Fn|��,����x�эزm��3��l���Sk������|�l
�R-�璭��_�US����������w�����":X{B~��q�q|9i#�Y<J+�B���R�#Y���ͪz����ɻ���c=Rn8��-NV/��M7{I3��Հ"q��؆�D_̚�l�S%F�!8�l؈'�)���~��DK��i�IGC�ҥ)�"�h�޻	5]Õk�p�V?��*"!�ljf5&:�D�Ԙѣ�0�L�x�j�����t�x��r�Q�$ϕJ=�7?��I���C%V�e���kA�f�h�da�x�z��G���z��#�_�g#���M4A�mH~|Å�-� , �|�DR�1��p#e�@�DTeK�̚P��ݳW��SsR4��|t��PK�YԵD�2�����B�&��9.��K�#��+,��HB;�tAcf5�I�c>I!�'x��'0<6���C�d���q� m�9�S���w��=�[�n����׏ ���.��޻.�����180�D�����
�Yx�,T�9q�ڴi�lۊ��x����Mv͚5�;O���_��r�ͨ���H"��;�������w5��ٶmzzz���wp�̇BM�r�F�_0'O���W�0զE��}���$:��Q���=�"�B�k
<A�w�<q����ys]���`i��*�w�CuN��@�/�\���hܼ
L��I����¿�
��X���8N��&~����*�>�N�H���H��(�z	������09Jr���wN�l��������@JL]H(u�u-�u�ɿ	z���:Q��rC���߇�ߏh:)#�\��<uX�R3�#�h8�{K(}5��|>'�ύ�7�������+/cll�f���?�u��#�H�Ұp��i|�{��+g�"h֑�}H�uL��)��4��t0�Q`o(}��9=�L� ��0�ֹ�݃��/c(W����lT��فx���o�ؑ��7����1������'ф��v����	N�:�� ���&f��#N'?��J=���Hy���%�z3qY��(6j�Y�����h��W�>�]{vctd@4:˖-�g�7����QP�:�ZR�����^zW�����x,����޵�0z��_~��;YBV�C
��[�0�rvu��~��j�ŀ�y��1�	�xm4H�S�S�t6����V�>T(&����h��wc�=��7؇]��R����uz��AϼŘ3{Z[��`�b�Z�RL��m� s��MI����Sp��r�O~�S�>}�XR&��^ͣV*��=�{6�-t���6���L	h��-�����N&�7�<�w�d�>r)�|3������_���I����ɵ���K5\����1�0C��b��"��q3�䞖C����;M_X��)�i��r45�R`��#T�S��e�&�hښ 6N�8U�ӌ#���kV*5�'��ZF޻�^���B�ʩi����
��L੧�=�6��}6�v�l�� h�"�+ �LE����#ݒ�I:��5_8u�WM�/q��xk�ۯ=�{o�����9��{_$C�%+���,T�O/���:�9���LZpү�����k.������_6�	�]X)/��5ģQ$	�|�!5�TKrp�լ:B6qn�O��3t-^����E,Y<o��\xkp�&��L��#�[>��>����B�����XҾ�d4P,Մ;IK՚�C�^C��/c�?��Xc�>�z�ϫ)7���W�}*����(��,H�
	�QM�I�W�~VU���nl�{�\���>��&n�;��ذ8����z Q�I8����6⑱1ܚ�b��!`���mW}��q	B"BF[AIC��Bը�A4jQ��!ɗ�\PC�6J'��sQ/B�G��dR�k]��(P�5��6o�|;]�k
�E���R����,�y+/�j��X<�g>�	�?��a���"�H6{&�'C��6m��]mǱC�1�?�J��ys���O}z����{�!�c�/�[��h�}�,Ғ��\C��CK:�9�� �L��o�3���+p����C~`�>�yo��t����;�b��.|��C�N}OK�,ú�kG��ϣ\�=�]kV��ҕairX�3�f�-��<�G�60W?�hM�ɧ�G�������|�<�'�{�Z��\x�E�$���D�����4J�F��5ܳm+~�w�֬j�������s4�^E��@6D4�-�Cw<��`I���~��Q�2w�Vz�r����T� ]�Tf�N2Y�+���w��",�����[��Z~��U�A��!����Y�ZA���`�isQ�pcl:��2�R���ʚ��ez{��SR��C�i[�݆�f������8p� F���9�RGP)�;BgDG:B�v�t����B�c�3>2!��dʯ]�P9����h�� '.�@�HQ�u
�u?֯߀�?�$����/��?�ĉS���|�3�����EC����"�<�"�i7bF4���$�~�F�ZA�NařL��"1#Q�Mc�:�3f`�㟂o�+��b�[{02:���$�oߊ?��?G8��T�j�� �G��Iܺы�����{�@�0�d,��[6�5w���%x�5d��5���94�डAe�ԅ�0ꕆ�=�������ǌ���>�H��َ2ˠ��T|��|�AU��N-��G?
��q�}�p��^z�T�%j��O�5!�1��.¢%+��1]���	݄Fu���ab�-��^G�	Ho�CMG�i��ʷ���Ż�ǩ'��	E.�?	��̚с��aݺ5ҐP|� ��b���*�<��&��X��M���v��[�?
LC��y���5��^¥�x��OB72]:�A�L��E��γ1S{��&�b���1\�:*T�N��8������&��<'��7�}���$��L���>Y���	�{Q{dX����~|x�F�r(���|r�5j�ղPkx�/�Ъh��7��8�;��fa,W�m2S��f^P��'A׾^��uAk�TK��T��p�⯚�_D��K�����'�ٽ{ן��f���$[�mkG4�Pn��w��d�)QN���L�òX�������<�.eo�D��(��q�"Aw'P(NH��cH'��f2�0ȫV�])�N�M�
ݬ#�C���_�y��W��MO>���38���8�򑓈�8^�ᴤ�X��߁k�"����C(r
��\g��	0
˯+jS�$�,��K#bB5?s]��'�V�6�-��$�M�Z�]�-nj/�M�q�kr-ZYm�3�c�l�w3�#8��Oq��[���C�h�=�D&F�"�e*�c�:��y��a�b`��J��:
���������s��G��rB���I�z��xM��Ių\�H@ZB��'u�����sVhF��Qb��o�Xd:��a��͝ ��7��������϶�-����k(W�Du<��ǐ/p��Q��#J�r(��"	`Q�t�g��?�DX��W{q��M�F�X�x��z�^��B~LhR��#�y��(*��5k�⎞9PB�ӯ��?��Wn������ �Ν+l>��]�?���	|��������o��J�$Ǜ��˗.����w��̝�U��D:�E>o����΍���Sȍ]T�N�y���;7��~��.Y�
�~�'y������
 ���)�����q����&��>u��{�P����8����6�����l�jX�"N�������u�
Z�qqm�:�I$|~�Laދ\���J �% Pr��4H'a �VX9�)���]��XԨ�Lv�� �HDt:�F1E^w��躲=���a��!�>e=��r��l��|q�P@���Z����8��6�nl��tvt#� W���ٳx����LL "jՅ:��ݪ�pH����DW��-愋NqU�F~��%�
��f�m�B|x��o��j���M��ٳz�%����4�4��f�q�a�:0<�Ç� 2��!�Xh�k�D13�D�i�F�]$�aR,�q��?(�&)6% �Y���O�������}{162��]�x�я���U��cϞ7q��Ui�99[�q3�������~���a�~h�l^�
�O��o����_G��X4�kUC
���ác$�C�Ib,�����&Ǡn��sN,X��Qc�)��%����Ǉr�B�b����uk����10>�_y	u�z�o[��4�B�c�W"��P4�PT,���Bd���܇=�a"��i�I �r[h���&FGr�v��n�4hN�F<�ij[6��3��{Z���*�[��ȿ�H!�J�	n��u��'�?��^M���=���\�GM�&�k����~v;���̼�dm���Qo!&"�H]輮��$����{N��Ƶ�nf�[ޣk�-k#�,�?I�����׍ l��e�7�~�9�����s�H�3��3>�é����{�v��L%�R~�\+�"*�l��3:���ܹ��L��33J5�{,����%{"B2�y>�I~-n�������E����g���ҋ?<\X�")�H����DZ|n��X���(�\��������l�0���Bɛ�_DOx񑷨�\5B�����<J��
�(�iI�-�A�g�(��,��(a3�ì#d�jR@DD�GagZ��S��g��������pn�n�}�%
���N��v/�~�s��w?~}��8�|�[�Q��z��rH
eҀ�G�i�!�2�K���c����(4��)���4��r.R^ߊ��������#V��T��z$��t�ع�����	������`�D�QD!�P�G�^>'ԅ	��LyP��(Y�U-ԅ#˦ �ւtKq��u4lz�pꠒ*��� Ͻ!�'�<Ǟ����HB|(�X<"�d/�C�m��v3B��K1�r׽kf�Im�)Lex�ӣz��łu�O��OW?*�"�a=��	�s��5�+Ģi�x���1of�d���sI&�2ps�b	]�ǣ�|ԛ��E�O+eC1L��fRHĢ���
�*�?4(�l"�B2�Q<R��)-
�y� &��J�lD�H�026,�⊾�	5K�+��P1�Ҁ�I�V�#��pP�T�&�C�M��̲�Wc�)�|3e�yd/��m�������m(�f�jl\z���M5j��l$�u��a5�����R	f����W�+_�7X�f9J�	{�5����C��������0�Y3B�� �vǖ�iⲤ��-��-|�#~�
�"jوƀ��>A��;B=Ą�ù�!���d����@1&_���"ۉF4�+�9��.82.�w�<�4��_BQ�ù\Kc�7n�����c��(l������;D�RD��K&�Vljhm����t�i�6�V��Z�ӑ�=�o���>LT��u��iܱ`1�nىH�h���I��j��u��9�޽[ҿ9���UtŢ�D�A=�_CȮ#�K�<,�����L*y�ҍi�T���u�<<��gP���+����octl��u��'×���������[����nn޼��� �L���w�_B�^ƴ�6ܿm3�Z��Ƒ����S����I���c~>�����9:,�>}�����4\Г�!.U�A��l ����\;�Q�-Ӥ�m�X�Qo+I��Ew�����`~/��<*FN�BaML	��]���ː��@:�)����B#���qmB���eS .y��d�\���.�m�r�Պ��d\�o�������+!���P�9�̔�U�^6�nj�*>��	���[��oO4��6�?��5������\#<j���xk��|>��D齩����^E�v��.󁀉�`�隫���c�M��{*��[�x_p:A�5�r^�l �?�=�����tU��K�-�h�G�q��	>vׯ_u��K��H%*#�����#�Ұv�b�߸��9(��*�X&�.���m
4�����IA<�z>�m�j�W��_D���������h����;�{s`g�aE9!�2��C��P�i�sp�+7��M;-���>�&��Tܓ+���-��8H����W���G��l�
9�H2��H�c�m3x�R�S��,U�50&¼Ye4�}'�E�����Nlڸ�h?ξ�g_�����d��qף����(~���p���:����$t�UV�J��ZUY���)7V���t�4E �I���2dlj�"��V��H�f�s�`�CA�ES�jI��f@P�P��:��ލذ�F����OQ�riH�ja�#ID�-"+�|�T�a��ӹ<
u�t�:�p�F�����    IDAT�]e�#�M!�I�ț�Y��FNpe�ba��!C�|�"�+�B�!QBj1jF�=d��Ơ��^�5�$����@x�S3Z�ъh+S	!䇥��)�/�r�����NZ�Ѻ�%�B���j�+�(��,�"ؚ4dg�<f��Ȩ�|tZH�*ʐ��&K�'����utŐ�#4ٌ��c���㔊MV�7�J%��O[Q�L8�*��g�/a~,$��i׿���|L�o�n�^�ތ�yMAsb|3Z�|n?ZLM
��Sӄ)z�wΉr�ŎY���J�9/[����kW���*~�����/����8��#q�
jRC����)��g�榕R5�~d���k� �>���ir)N���1b8�3�L}�2.���F��ј$��Y�а�44h�B9����J͏�֨b��5��g���}B,qϜ9'��Cl��r���k7p��	��Т�:"��[�\��w���w���倆Z'�a�M ���^�Q��E����i�u��H��Ƒ��P��c���x�c�SO=�� 2@Ϳ��B�E�k�S`�c���׿�u�=s^����!Б��Н�#�%�̚*"a]�uҧ\w'ʤtR�U�Yh�?۟���~�ڛx��}B%��ف'�|���_��7��������~ܻe#������l����Ͽ�r)�����vbݝK%T����@��Q���FA��t4�L2��2P�Tߖ���'��t���8��C���i	���7�A�^�FʹQ�lTM���
��z ��,�������ʫ/�P/��7��ino�����Ĝ�K�)H�h
 ����:sYGR���OM�U�O��7=%�#���_쌕��bY��s��Jr\U��WPˋ��'�һ<z6*^s ;-��&��z���B�[/���r?6Y|{?��j��}V^�n���æ���:D&�nގ��qm�����.��Y�Pk�G��&ܫ��w��r�Ǜ)���ǂ1ɜ�~�����L��F����Ð�����-����6w��%��A�C	+���M���NCrrZ�:�.�ӧ/��Pg�K�j��ޟh
����'i��p�t�O"�֯��)��.����g�����돾����M_o�]�`X�1s6�� �#"�Ff,]\��p����gբ��=Z���N)�qZ)���<�%�N�T@���ݠ�A��	>_��Fõ�5S�HՔ�B��S��]2�<u
�8�.��;�݁��\���ӧ�\f�F�@b�B�X{n�L�w�,zFP1}h���W�*]6�<OH� B�T�༹)���ӽ)��N����6<V��O�Sڞy4�.��Q����&_�Vv\��B���>�0ۼ�����'?��ѣH�ua�"�4��8cD�;Q�$q��Y\<sA��>MC�'��� @����	�CAqZ�m6S"%ｒH���Q����u��ɐT
��PW��soD����'��Q���1��C��{�a�#Q�-I�lh���b�#���L�M<�Up|U)2�{*�A	���b5k�eBƑ6�M���6C�O$ђ���
��\��c���i���Y޲�$���M�o����m9����z$}�K�
u�z���1sS �K�R����c���z���:͓O��=���L�_O���\�!�X��)��+��]n`ɲe��?�?�f�*\<s?�������0߯aA4��SG:`!�D(J�Š���"_PL�(]��t5"�RTQH�l
x΄>$�>08������Q8�8zKU����UQ#*��f��e�X��"���i0)\�h��o�Z/a��җ���������Qs'o�ᑲIn���.\���B	��q��1�[0K�w�ډ��*585K>��-2��� �=˰k(�K(������w�L�(�\B�ހ�T�d�|����'׮�ĩ�g��3
ȅ��A�x+���!�=�X ����L3b1tƢhdJ@5�NIjw'��}K��x!���F��y����q��������r�Ok�⡇����Wq��Y���	��O�vn����Ic���<'����1ٍ̚O~�a��s)���:.=��?��1��0Iֶњ����i&��!�Si�.��k?��A��)^�<�9��RKI9�}M�H�Xu6�o�����Lj-�-Ų��Q�,�~c�0P��*��ɎV,Y�
��,�� �̊Ͱ���)���N�R�: �Z�k����za�j���8�^�,tYR�܄r�$c���3'�hĵ����d���c��M��^�5'�~t����������7��~.�w���P��j�|����}���ђ?�ƞ�M�������7q�6��4e��;�)�]pG�zqmd�]tRo�&eR
��ؤ���8CaD�1q{�G��q����o���8��59��V�Қn�ZҾF�n!��h�2tv܁jM�i��<*-�$���'lN9�G�MA2�}6�m���p��?Uw�ʒ�Q���<��o?��]��w�����j�d�H4)\E�:��M��\WI���r(4�@ <<�����>��M���q�A3-eo�P�^zGZT{2�4�l h�r�c#H�1*Kp;�"��(��zPCk*����`���c@�5� ٲ1�PϤ0bk�g �����0V(
����%'�^AQ�G�$�b2�D�R��XP3N	�.!���j�����z,���Ѩ���V�w����uq��3����a��e�;����G�|�}$HE"�M�K��T�/����`ڊ%x��7qp�>
E8~]���!W3�f��؊>Dg�lZ2Ml�M�BYoz������D'�U��ܣ��n�l�os���4��&Ҽ�7������x��T���5� i:�u9��_[�WD@*aT�/���}ss`��DWZڪb^}v!dZ�	�=Z�z��:������y������8WP`�N����x��rݭT�/�u�ZQ��G}wC�M�M�fA�Ɉ<��ܨt��k�b#�E\5~�3��D���;�?������sJ���K�7�>�Y�S���)Z�e��w�����wFΟ�O��o0�w���"��p@
��K# .C�d��Ne�$P!NB
����z'��!�$v��M-�Yѣq �Fo���n�1�%�ЂՒPH���2�0���n�'0V��l��il��e���?�G}��{q�z�X�R�OAn�4E��rg/^�~�F��7�h��0�5��(j��H�"ZDQ�t
�i�`�ڕM�!;,@�%�
���"�х�W�q�r?���j#��w���~��xࡏ��g�����Qr�g��Sq�J]]�sTh��PB䜓1p�x03c��9�sf�s�{���x�il��1��"!!$!���ZR�:��U{W�;����j�w8����ju���{�7<a��]�H����2Q�r���/�շ��ml߾AvC}.�S	tF���h����Eh
v1]�K4��B��T|�����p�-�G�x���������Z�p�Ɵ���������>v�ڎ�V�UW_����'��,~��G��#�#��Fwg3n��:�\�[6���ݻ�L�r�({k��ܨ��ASC#�� "F�LFx(c<'ǒe�D�m ��I�+_B�(�i�Z�y)�'l<�]�a����40�4-�Aے�(4�����RYF+#�6P�P�X��E+�ڱѪf�Up{�T�C*WrQ+�����wISN�y�;#'!�*)M.N�-�����+{��u�	,Q^^��ʛF�7����dv�m2�lQ0���tǝ���Ş�B�A܉�v!����X�L�6���Sg#���kEU ��1�	��3�����k"%�_�^B~5YU� Ef��t�b_ ���E�Ĳ�ʡn��pi���"R��c����*B����;�mo�%����1�w4K��O)S*eY&B�0��jdO����S@��Ehl��!�/%�f��I#�$*�2��u/���5TVV�Q�U~'�}�S�1��?��x�g"/=��U۷m�N"�ZƱ2�uF$��k�C���N��`���E� ����k'��.���l�dOM�1��ry��T�!��P����E��z�3�F�V�����iB�C�D�UB�ύ���\�k򇑰��7�8U.a�*#CI��z��R.7Ɖ�5��2-�J#<D�m�u&��I�o��[�; �m�S�<����s�U"��eU���^8�s�&���$��ErV/[�o����q����F���#�͡���ZL�<80>�Xk���f4,��+/��M�l�����"�h"�E�*+�,x�5U
�$$�f�$��붱᳝]5��92���:&�
�67�w
'�:�����0wR0�8�D�N*��Q�[y)(�I���r+���x���8J�*�arJU��a�[AZ�~0��&�2�Va�v���C�];���~��Z�P�&����3����xd�K]�h�_MhPtzr���h*&חP!�,�ѷ�֜ȽP���c���)��-%:3�s��܊9�:?��;���t��u�hP�]�s��\�|
x��q�3yM��o�F�af���W��μ�\`�v<�G�=�Z�y4���_*���t}jŌ*�əq&F�cN,��W8m�(�TA.�ǯ�E	�v�/��G���J�%�8<5����'䧺
�8��,���=��0�IL�Y$����Y�P�����g�II\��*IQ@}z��=��W���G�#+����}�r5����"�hy|�QY��C�P���MS�R�bq�@��Zs+��`��!��/�Ţ�|���ӷ܂|:+��)D摰&�Zjk�09:���b��$ɯ��p�Rh	h��x�օh_���WFQ��,]���$����L�
Y14��W,ƍw܉C#i���c�].�tw����<���o`�����_xw�V��E�x�u����R)?��_ᙧ�E.�Ƃ�v�xՕX�ކ�^؀S����B���HQ�}���Y��%/��!X���>B%3ܟ�R���D�*y�Yț��V�[8gacL�9�b�-�g��n/^Bm-���"XS-��L��\ȋ�f��iP�ֶ�T6�M��U��V��[H�c/}��t��mQ�<�]5� �[�
��b��xq˘"�G�����q7�r�9��,rK��vl�N�މMNq��m��������78����ZS��pH�>�<>��j�\�̠|�4,��?�y���l,/p��9�~�cS?c�9��L!���a��R3d�Q�FUU<�
�(��ݖ�[��]b���T/�D%:й��Ȣ��e�=Z	-�hj�_�	?G/�pQ��'0��	�����h�`���;�@����~2)������|s}�^�k����H$��fQ����W#F�+P�z')��h��%�H&?��HaK��#�Ci�f�I�I4N�`�S�@�eARRp!�Be41�(��*C���/J�#xn�h4�˨�{P��6L�<R%����qx�ׂ�cu0�~L,L���qу�2$Z��,
�Q�(��(�&i�$3,��	�BH���ѨL
T Q����`� �D�y=^'n����%����
}j
olB����(�P���w	&=.��@��g]|"�A��x���1r|Px
t_�j>L��)C����ހ���C1���ro$k���� ��M)�D�[A[>�������܄^6v��Ί�Q��Yf�;M����2��L}x���7,C9J�l�8���$�4�S%�hX0��d��=V�s}e�BXq�c�r�YR��vΝJ��eo�r����l���;�B4v}�~��i��������)*�����] !�R�hNA�"Z8<�)�{g��}�1�Q���{�����x�����kGX����r9�=5!:]8��ϔݒ���eB��oɴ�E����tg,[�o��ױz�*`j��7a�����`��U@�K�u�r>C,=!cټ��4N|ء�)�%'�h�7����)=����G9e�h����G���PE�e�:Rpabz
��i�,��#	z�삡�a��8>3�)�#�,]`��ӳ����`(}�1�&Zn�\���jD�UŻ;�����;���]e4uTЙ�E�zUj[Q[[���fN��M��K�,�,�niB��G'����x!�(���E
����x�'խ�U�X�������^ܰQ�E
j��]B�U�IAC4($ݬ߇yg����.�����ޖ��<?��BZ�-��_��OL��>�������҈[n��������6��g?��}�Q��O]������T?�ѯ�a������W`~c3�x�y�>��� �Y�����ˮEG�*6��k�>_"�I�ɸhʆp�E���2ņ��Y%����2�s]��\��<!��$�0�*B55!�҈@u�߳O�2�qw�
�Y��m�Qkg�QW^�f[�N�O����X(�k��,
��o�h�����^�r�Ԟ����X�H{*ߗI������Z�*���S&��̍�|���$�N�ߙ&;��ğ���w�6�f���	!P���q�@��
��������c����|)l�4'�:����eϔbG�Y|`��+F�S�OLL`zrT9���=U�hR��480�Ç��X� �3	x�%D��ǀ���U��4���t����u��(�����s�~��B�_C�2�@uL���O���>�X���/=��ҳ/��p�ѫs9�c��P����!�R��펰=�d7Su�q��ƕK
�@WX.�h�K���%!Ԧ�qdq�q�Y��� ��
9��7�$	�I���,�>B�h�ľ6qq4b1s�(5~*��C\�ۏ�r��FK.�� ��� �"�fA���ZX���=T��!\�]N
��SZ��Hڱ'&L�4�"�2�4��@Q�t��<�:	*H8�Er�cow7���P��[o�r&��z.� +.���FLX>���x婧���g0~l@���������RYo���u�WN�
F�:{4?�B��h�ן�U�IjS [��0�f7T ��0lN��	�N�xnA��d��q쇵��rȹ��Q8�{�U��"Y�O5�꜄�.�� ��¤\9w����*N����zI`�U��e���U�r�����B@�5�U/TQ��>v�eC��9����K��ɀ�T��#�s-��]�s���ΞjH����7�0��"�u�Q��4�O�9�!�u�w��kй����%eg�Gv8[�|H�ȹ���)IM���RJ�|:�%����oc�j3��M��?G��C�����y⮅hM�Q���L��yՄ��#�)��"!�6r11cAE�]0cW�7X��� ʑJ�Y���F`Q/��fLfsx땍8�s�x��^�����zX���đBY17KʺBе0�y���­"�|L��چz�^{�����-8�ׇ��%��]�}$������0�>KW�C8��m���sOB�e�ҍ���\zS�]]826�=�"�g��h4���Fո`���E�[��f��	�����D����]�+Q�w�>�9���ʜ}��8���D�<6�y�o~�B��[H)��\�+?�E��ţϾ���>)��kq���|��������<я�߃�k���[o���4��*�f!��y���5�`Ac^�Y��F����F�B&�+V�қ������m���0�u;\�Èq_JO��'a�?��(�޳�,�"_)�&�L5��s�D�rzH�*Ӓ؛�t��X��ŋ7x{�N�X�=�Dň�Hm��@[�<D�� \D�۞���h��JǗ�V��U�n&�YAH�P��PA���1��Jgv����������͇�gB��)��P�mα9�r���������97�w��sc�驣
]s���[� ӕ�|/5m��I*Grz
�y���
�����{&�"�}:PgS"J�4��;b)=?��lɾ����<��	c����� �R|�#w*9#���2�s����r����	� �����%) �i*���9E���6��^
��    IDAT���]����r9D�[vZ�{�C�<F>�~а����(�Xe���f������w�o���t��`�!��"�Q�3<���7rYD\��JgbKm:U)'��'�Fπi�	�@��3���%�����L	(h�)�(� �(�)]9���8 ���c�<��<�P����|A̔-�(�_0p�("���F�`"H��h{-�K��J��I�IH�)FjJ�����b��i�|ꑜBL�8"���Yu^�����y;s�1&|H�89���ڊ�~�����1��]LB��nhF�EaɅ�!����M���X�2�x�������wXt�M�ɀ�f	�\Ei��?AT�jP�BDc�ysE������G��`I�Si�OU>�4I��Jϙ�I�;��D�v���8I���:ψt��$6�������t�f0��$�\Pf>�9��3�8Nq�A���(�T����m��j=�ѕ؆ �5��#P�b5b�ê*
ʪPf�m�����
��I���n�m�ν�A.��ԝg��/�"������	|�TAc�	��y \�T/�M�~>�rDQD�͝ו	��z��lnaF"�s�i����X�j4;ᐧh��i:8�ϖi�Eʹfӈ'�E��w�����ƚ�ˁ�1^{��?��L���(���xu�hI�Ϣ�x�8E!G�Tr���ĉ���ǧ	dB�-�s��1L^�+NԦOGF �B�E�w�%@{+̩���lz�iD�@D�K����"-m(��86=�����4e-	
E��G$E.����s�anmkÅ]��z��_ދmo�	�i
d��*�)��%��ǭмh1ι�&4�Z]��ګx�G?��K���l�0a��#�Ս}ã�}�c����(��t�w��^��Bj �4���.���3��F�*��g�ʣ��F������ec=.���Xv�%�F��i�<�6>�#��F�b���ĕ�}���Ϭ����iJ�R���C�X,�f�H-ΌoE%��;�����x��W%a��ݎO]}5�����a��a��&��<��(M�_����%4��(�����0���8��O�%�BR��Oy\ņ��aJ|d��F�4���s��"��L�(G��RIMǢ��ług���0^ۼE���	�	#`"RÂ�˅SP]�(�7Z���eJ��x{
�Ĝ�?�N�>�l,[��L���| � PҼ��T)�aBdʒ�'y��&��;=)�}�i"H��S[����.
d�|���!���r6r��'����� r�����/��s�?:t
�ñ�}�G>�F�R��ݯ&�R���:��&�3>�PR�!�eՔ_y@j�k��*�v�YR�Ї�$u����`���}�p ������e��/�f�e�aPP¢�)���F���O6j��S�]e���(�������Tz��ю���"G��q��xn�������.y���SƇHE��U��
��������d��|��O<x�[��ltt�'�ɉl�ˣ���IҠ�����p0�s��T�`�i�CXT�QD��\6-\n��dF&MOrx(�V��8_���Tf{t��+2��@����\����2�Y���Z��%�8�j~I��n&�BY�ȿ�|)�	PUp�BL�\mVF����**�7%x9���"0�|r|H̢��J.�`0,�?��K5'Yf���!�k:��7_�&� ���#=9!EFmG+Z��@��	�IBG�^jn{�yxc�x�i�y{;�&&�`���)v)]ȱ�Bzj��Q�EH���X���O�Cifɹv�DV'x�8�:�9��C�U��V��.�=rv���be;����ILf�`rL���_+Ȉ����Q1Y� TQ�~�HͮM����,�-�'e*wz��}��	ܨ���:a� J��_�O����x=h2��?$��eF��xZ%��q#,�V�N�S���Q�@����'dbSR� ;q
�&Dk�[��逸h�Z�����D}��1��"
l�N������I�hsD��p?7;i~�M�y�����ܢ@6b[��Q!R�D*�� N�n�4e��d193�Fow��V�jjF���l���èʧ�2�a�b�N�6���RE�i��?t���PH��ȍ��Xើ���)����R0�\0�TM-j/�����:ad2پO��+T�]i>���'Q۵P���tOOvh�v�eWફ�G�2*ϊz�J�C��*b�0�C��?�6<��\�2j=@gE��7�	nz�:�n�����&wh����;���aԄ�(�K�4-D��!�=�OǎC������>�=i���B<���p%�[ƢE�X��L46������ٳ_����������Du�/���\�/�k�����lG_y���>߿n+%~3]g��o�[����>���c��5Tᬳ��-��,�Z�VHSC�����طo?~{��u�q��n�U�]�֪:l|r=&�E[TGНCي����kp���E��K ���;0���(�A})�@1�2J��SF�((�kÂ�7�c#��d�"Y��}V*d\�\�2�D��G��A��3�s�988p
[�݅�����E�_D�ҍ`m�{���s*���bJRV?���S�Ye4��ZHltHSA|(�`7iD�ّ�WM
����l&ij)�߬�Gl��z6�w���Q~]���+�H������t�9�#�ߢ���Jȁ��W�Z���9���`n���ym���/�_onz�=����O�(DC	��!&��Vu�����خ����f$�G�{�q�V*�`�E�UzT�Q;[� �k�=��ɦ�E��L�~4Q���,i���9�W��XU��&'r�vn_	�=�B��u��G�P�xL���V�s�sR���چ�U�^[�[W�����L�?����'�ٷk�Ϗ�^>80$#μ��S��&�Ȇ�Н�9U�CJ&F�ɀ��T�=
3O>uS�)�V̱4��I�g�=t�B� 4�lT]Z˓���H����p,e�YS���1�n�c��Ű��#�8�ʀ���BQ`�`b"��2ƣ�eB�d�ir"x>��3Id���ILsL�T7�4�Ru[ݢ8���uc��#D9��������L.G*��MDu+��"@Gk��K�׮AT��2s�5?�
��ɣ'��?Џ���X�^8�m^z�I�{g'3	d(q��b�P���9R&.:FM�
�Q�g�^݋T6-v�9	ȓtG32q$e�&� 0�s�Ď���Hh#<�jP$}�6	/�,dv'hq�����,���u0����-1� 4�r�l'���e���s&tGF���'w��2b��,\>:��	��H�C�;���X�1.��<m���
(�w�j�$&�+ҮJ���ؘ;�1&�9�ۦb�;Ux[-�<v����l��8�n�e�1"8�����|&�F)Iy��x�p�Z
�O�z<�<K2�Wv�h�#�iŒ`s��os��A)Bh�4�zd���y�s�@P��p̐���0=%q-�P�g1�Cbr^#���8���~b�	x�Q��"T��H^�.�ww�����ΒbT�T��d-K���@�2�1r)���P�0~9	bQ	!��"YS�����ҫ��E�쏿�����AD�������m��b891�#'���!�8�����Dum&'��1"M�Wq
*+Dq���}�z/��y���p�s�������&�֍L���Ug�[�@��s%>�ؾO���P��g�b�T�	/)�މm��ݾ=H���y�AQ]��n��%KŘ�� �G�G�W\Xc$[Í��Ƌ^��`"R*��h`~,����2��֝��o�,"�z`�0���X��_b��n23�&�s�%X|�Ex{��Q�K�2�GC}�测;e��J6u��8FF�pp�!�����.Z��Ͽ �[;���c��1����54�x&��Ž���_A�W�I���H��������.&�y��[LN9=~Yl).�R *Pn���⇱�%PRƽR	y��\H�|�X��{��� ��G��E���*C����Žh�?��F�j�=!��q��9w{qX�{*&n��@[��!���GtP9�*Ƞ�l ؓC��>w���?�!sd�E��VB�a��ߟ~���g��l�w�r�89s>�5켯K�F�����˔ϥa��^ܰ���!LMMK��,�y_^Z4�4C�
.%ې@UQ0+;-�W9C�*�=�q���BIS6DTJrxЀ%�磻�] H�b^ɞ3?�u�����h����X�q�ힱ4�I��jĹd���55���e��\:�O�4.��<d�W�=��������{8���'E��5M�h�kۦ��x{��N����DSIbmU"!��MZt��#Y*
Ll�sV��v@�n���*bn&+xU3��0�zYH�C	B&�C`a��e�&{v�E�*>[J@�-ŉ��]v!����G�@��;���8QHa0��xހ���q�����S�n?4&8z@aHK�H�Ң<�M�{,Y(�&	�$�����=pGq� ��%�lJ@���Ug@ʘ�EA�4$Q:�P%&�-u��+p�y�`��y�"A^,�j��(v�ݍ�7�����k�<\p�Y�%8�}�v`rhD&yj#���dDu�����D-
#)�1�&X��l>�K��=�R��pC�5������{>��N�s
.S���(ƨ�d���i)��O�9��e��I���l�z�[Y�k~�h%��jnJ�R�;����@*s�5�ϮI��:�Mmd`ld嵼������O!%�� PE�(�Q0s�ј[��)�c[(�K����|�@�l�(���4����e���,Qo��q�)�=N�t��*!�/�#�P�/Mn$	b�w�S�D&�Q��Y�)a4V%����i�F����G��x<F�jc�I�ǃe���E�f�25�WV����?�{$���
��LL#I�P� �$7=�ϓ:�Z (P^�r�L�K���C>E/y�pL���LOJ�=�c�������|��b�2Bn�3�2�^9��	���N�H�H<��"�L�޲�}"�ώ� �H&�L0�����ٵ���*���h\瞍�ˮ��k�͐:����3dN��22ȸ�<a�5��K8r�(F�&�%_(@��������\���:��?���I��,��3��Wr����lk�S�=�M�nB2�F��FGPGODGG�O �T.\���߆�gʤ u�6���H�<������F��(�U(B�}��ځ��$r٢`�/��R�r�-�ꚇ�����а"O��~㒵�PW/�I?��O��/�S0Р�h�����-���40jW��o���l�nTb�{���>���q4�/� U=�xc�A<��zL�$���
|G��$�_*AU��\!�x2��/(��㱰���}.�.�E���8�w/2#Èj\�4�8�z���߁���/o���(��L0���b��)�HK�E�/_T�l�@6o,�뙰R�:�((Is�ui/�����0����"o�ļ-����(X҃���5�#�SS�2ƴ���1����h�DP�%����S۳� ���CJA¾U�sq2���s_���o .�7��H�s��"��ɸ�4��kG���<9<-;r&�D��3�S�oV�B�d� g��w�x~��ܳ���Q{��|�}?�(
��L�ܰ���&&�N)���9�+<���
��pA��̙�u��u��`�����VUazjL��AMC0��@����Z�%�4�a]8=�ϘPq�^B��\*�T�S�pEm]݈U�"W(��҄�L�e�4�
���j"�=Ö^�i�@�[8��m���}��7>��moo����x���N� ����fa��v�K ��ba�\��;�\�l�:����e���)��`�J��%;��t����&�ȥ��C�ۋ �REB��ˢĨ �>�%O3Y񜉪�:,�]�y-���򸐝�cxz{N�c8��tƀ+D������4!A�}����2�(��O�!?���`���X8cQgZ"�������e��'&It�%�(�B�D�"��"�W	WP4γb����؈3���5+���na	�LĎ];��{�c&��eX�r9���ߋ�#�*��4�ˋ����tF�%=Lʽ~IJT'ڶ�g��r�J�WV������{��	�LO�1;ɢk7"�JI��>����ɧ�I���Z�&�"5!�y�4G����������f�Tw2��c`��*�[�í)�^�|<��Դ�BDj�T�Ķ��Z��<�,V�nQ�I�'����C�P��TT�&Z-������s��I!13)�3'.��C�`���mw�,�өt\�G���g>����YSS#p�5��b�+6�1�V׏�x0�ں:I�x�C.2��&'�039��l�n�(Q�.�R��|A��3��&�
B��@���֎p$"�/!�ˈOOc��	dR�Y����������E����{yC��098�:�(IQ��݉���9fAl�N$1<<��1%a�sglhllDcs����b� f}d�$�F������d����Â���u�f��d��m>:��"�����zXL��sf�P��EI�8���Dpz8�4�9�̤h�"��Cw��er�������j�) _�<d]C���8��ڵ��z�z��u:u���1q�}��3�s��=����=z�d���e���EsW+*b�S��|QxK�|�h���`��8�� �����9V��MX�\��t
Qw	y>ou��&DW�#6þ?������`�����t
��u�.lۻ��4+'�a,Y��]v��k���m8|�O�T�Wx�"�
�z�~�z����J���x����!j��I���^O�:��&�����/���ݘH�����t����_��w���'�c�Ԕp��>� 7�4r2r�<�����-�A������_ƒ�y���v�*�Gf���8u`?��<<��4-:�/�5��ZW] *2�=���܂��(b�����㵤i#�^�K����P�g��ϙE�l���d��L8 .����i���Dm�<�L����)1��rȸ)k[��ѽh�ڻQQ��ٹ���.
�-�l�EU�.�j.|�i�)���ݖu�2QCcrk��9�U2��CJ�ԁ��s��
^Ć����L�4��>"2@j�������n���d\&�l\JG\�W�d��[om�c�>��'O(Cr�d͉Ա�.(��os+\�AE8�o��~����)TT���˙��(PxKU��"����B1��;�TPOr0�����P�PЋH4"�����SyH�{���e���l[�<�wuAD�((QR����b�����U��jV�h������'�m���Xyp0�q��;�~뭿�&g☎g����W|�����LDdq�v٬t��j�!
f!��ū��$�Ј�zQ:�V�䟼��D^�W��v�!"�X$I���N6���}O ZM-֜��]t!����n:_&���a�sh?��ÉSC�,!|Me2�f�1�%����
�R��VAF��p�!#E16)��t��x]�<��$�R�`R�r	�ԲgbW!$b�N��»�R0V$�|�@Q�_�DT���X�h$"2�өGF%v666c���X�d�[�Ka��qh��pEqбh���b�4P�t)
�����8E�ϧ�I��@��u--�;ϑe�B&>��cG����2�ǋy=�PY]-j	S�"�������'b�����C]K+Z���F<�9�5M��ĉ�A$f��{�҅�mhDSG����*B(���� 51)*,�xJ6&����݉�����l�k&�S����>d�)h�p����/�P�Q/]�U<A��CȦ��(�(�ڤ#��!�1�R�L�ap�$R�8<�XT�6b���hhm����gQ�N&0tr �G�H~-zӚ&���EUu�(N�x��>����\�䣦��zzP[_��UP�%�N�о}(dr§!���̂ŋPS[?[�2���    IDAT��wwbjzB�
&�--M�]��M����r>��xg�[8���d�
л�,��E��3�(fdI9����A"���;�%˖�w�2�56�Ae1#;�߇c�`z|M� �A�q��,q3�9��,�y�4?�<.D�l&�lR��<|U�\Შ����a5�sH�\p)���r!l���0�x�+�}H$a�(N�����0^Q��mW^�В��|(����<�����0o�ZL=��׏C'�1:=%�(,\t_P��eM�a<�iQ	��A��bA`�5��E+Q6K���b�J�beK.��@��l�HF*�q�gP}�y
�̆�O`���b>�^x«��ȩIl��.6o{��߁����Q4ży�y��1LLLI|Ҽ�Y�P����?��\ F���7z]����%��$L�{���;� RĳHmۂ��6`l�0̠�ȼ.��{Q�5�w�౧^���1��b��mY�i��@w:�,
�e���&�r�W��g��4�"�:U��<���w�g��w�ɰ���p��}�r`&� O@����#RonAe|
�n>d��(/��9�`�[�lN�[���Y��i�Rб�D>�>���Q��"	���vu`������P ͏#���G���-B���R�����s-
JfGc>�8ۑ��S�i%��ԕ^����	X!�s�SM6?�ß\I}��.��5���
D��P���fs��N�6NR͢I}���]�Ņ���D9��p
��=���	jQ��F&m�} ���Ɩ77�Y��R�/�}n4"��sR>;�S��S:t�8�Τ�f�]��L�!:�>�+�}�ͩ\�|4����#��� D3�
�p`6^a����p0 �b�Ɂ������V�p�aOz��7��hOG��ڧ=�((���߆��3�	���K�?��4q�@���ի7~cdh;�ZF�-2�Lj�����J1E�;�����d���rJ�E�YѓG�oꄳS�u)��`�C��~�Z<,D�S@�2��ѸLAV�B�� ��e�Z�kVb��3��٢4ǳ	�3i�G�q�812��'O���(��ދ��q�O��;�<���*��a��Ӛ<��Jj\G��n��5�{\�ΔD�T��AqQ,Ȧ���'�D����+�˛�ٞ,�`���(9y.�A�$ǎ� �,ĺ���ʕ����I��Gv�����_یR&/�WB_L͋$��0NB��Ls��d��T�DcW7�\p.��]#�;��ˆ���8�nڄ=��C"�~��
7|�6�uv��u�y˘�;ol�;��$���g_r	λ�rx�������]�����ʫ8r舂��A�:�l�;�\Է6##�KI19t
�6���{)��tR[g.��,[�
z��.
,LO�cϻ[���cz|RB�8��Kq�yH,��RA̿�ۋ��_���)�Q	��q�E���V� 71���ދ�7o��Go�}XԻ�_r��.�WWD1r Xd���3���;ȧs
Z�Ἃ/qc[�t��}�8vn݊7^~�x\�	��,Y�\~���x
�ѐ�#���g�C����+����^� �\u�t�b���`p�^x�9طW&,
V�^�+���.���n��ǇF�³���g��|����V\y�X��LBQ�4��$x��w��S���#�\�0���kp��磾�Qދ�tN�كM/m�{[�F��G4��c���^Y���"��^D]@�\F�0���/�!5L��J��.%����r����0N=8e�
xኄd
c%s�.�h�B��P�@�Y���@+TQ����a*C��t��@�2��I�ټ���cX��нe�/[��]�qӅ�GO ad1�N!���1����鶐�g�0F*��~�]�����ڊ`X
��1X�it��X��=v�D�b����|j�>O���ȓO�o���6E�y�:4�}Ǔعk?������z�#�B(�$Q������W�?����1��̄�}�#�7��XIE��C��K|�,�F�W��e@E08������6 �BeOZ׭E��)-�]��kOf���a�N%���e�Y���8�l	i�B��؝Dϼ.\w�5X�b%4ӃG{?�vl�+�@�OigV^|	���+p�2�F��1���#'-p���pA��'?
d��9@�,!��`f
0�LD�R
7��r����(�<(W�hl@��42�"A�Ač,��"UQ,Z�=˗��s>"Ս(�tX%�<av���_1�Pf��l%u��	�ʌ�}� O`�����E������䜝(OA@���b�{!��Q�SE���&?�:؝�uW�i<��dl�(�ŋC4�-V��<'��EQN��B�ȡ����q�^�����Ě��91�RT��	#�Gj������\����(�S|�mu>Y��2�6	��A^����J�d���#u�4	�"���
�
��
<V'��E8
*)U�����х��6i̱���(�����z��%�k������D��B����(��f��q��e�[�>uŃ��?�����Fΐ�Z0mo��R�	U�+R�,��$�}8��	1�j�x�( t����gB��eaQ�h)n��c.��%Z�����0�A,<�"\w�����p���������؄�����9�<1��v�Ʀ_��prl3�(QY[=@�F����j1;*/��|�I�(;ck8\eTD���!.bN�3��&�)�
�ü�V%1�|A�Z�<_�AJ�������QhliDc{3�OliBǼtut�ˎe����0���?�C��I7-�ܺ�#F0 �����
$�n�y�~�}�e���_s��+N&~��N����O=���!��>��_���?��%K���0�<t�SCX��cxቧq��Q�2,\܋[o�7��yxB:Jn>O�LG�����l��
�)��:|��?�gn����[s�d�����)���{����`Hu����ğ�s��^=�k��1����7ྟ������sK�|�O���t�8��fVʣ�M�͛��+��/�a2��y'n�����$�Kφ|{�݆��������(��Z.��*�v��t�*�6��]�B&��q�{�	?!��y������b�ڵ2����Naۦ�q���}{�G�ȣs�B�|���[PYW'�G�\K�ƿ���x��SY�X�+��w�}ꛛ%1�qn],a��	�����@� ��o�w~��1o�
�VgA+Y"���[��~�s�s@�5�]r���=Xv�J!�"Dҿ��`��������x٢������]wᲫ��5f�0f@��Ȟ���#�����2"��-*Zh�Q��QG�)'nE!�k� � T��D�N�,2H�4 ՟��E�M'� ���ga�U@�2�bPCj&	c�B�׋yU��z$[��۾,,�w�<(x](�#H�T��8�R��Sã����x��?"bfD.�E��7݂ɢ��{��B"��\�h0*�]Yꑳ1"�,�Ljx�<��^��2JK&GG�t�\�S'`���T��	W{�n��֜�q09��O`�ۯ![�ł�.D��Wah*��{�E�8c$��u�[z��:li[ȄWug�|��9E۽���I��� ����ȡcr#����Cp{�(��B�e��{�@��@ߓ��䦗P�M�~y;�׭F���p-f�^܄��O�`�d��aJ�0y�EJ�!Q��T�)"Z�pczzT&�qj�'<��8��Vx��eo	K�=���A�^��Ͼ���7J11�@q^�*
(T��nl��_�cr�԰0��7e�(����Y���F�dɴ��୩�Q´�#H�[fsL%�}X�t>��Y�y�� VۈBIC�Hh��NT����Q�NOfݹm؎�D���� �Ii[�xtH�{N���MI��g�.����k#�GT����Nؑ��WR�Ywz�x(ؑ���I�Åز��f<g��Q���S���i��?&��yM>l��I��e�M����8�n��8��Y��AӔ� ����|M��#U>�	SQ}�R8��F�>Dl��.����6RL��%����������
fAVYY)ƨ�W�� J�Re� ���Ԏ��
�c��8��#lOM+WDc�C����(������l~���Ϭ�{���ڵ��^b�i�C�(;Xs͋�t'�8��3�s:��a���klI,v��i�b�C�<^���6rR��Z*��Ӽ��\�HHC"�B�ST"w��W�c�u��;�����ط�^�Ǐ��Q�^��ŽXt����߉�'��[oc��m852��D)�O-D��V$4�inR��PRg19ά$�\�@k�+I��T����UF����bQ�\��R�U6�dFi�t�q����.�K��B���iw/��e�0o�|t�t�x��N�2yI����艓��C���8�k��tF]Q�q!�2�T�!i���I��\U������d"/���o����жj��iuу���{�~�;�8��ǋ��E�����K&B^u�`NN`�K�ȿ=���~W�ծ� ��~���ԗ� �Wܾ\d�Y�8x ��~<���07PYS����M|�O�D��V��\�t[���~�K<���8>,��˯�_��oc>u��Bp��P.f�啗���~�v�IM����/��op�gnU&�U�܅<v��	?��?`�;�%	hhnğ��p��	o4,��+#��w��?�����3H��({u\�m��}�b���(���o���~����yŚ5�����֬���l�L6
�oތ�����d�PƒU�q������n�r*u��R���� ~���#��{��2ڛp�gn�׾����*Ҭ����O�C<�����g�[o�7��-4�.Vf�"��\���~�����#�q�7����:�.�"Cd6xQ2Y#�����+lx��z�X�?���q��WKB,�������c��?>����X@��	@�?��@�>b�����,�Ζ���(n�"�(�V�&9�����en�іO�-�{��Ҁl,���Gz&	+i�Y�3Z�Z�RD�@�I�3/ɗK�zٴ.i>��:f��Q���=�B��SCcx���MO<��R�8c%n��N��x��qh�0j��1o�B4�v
�d��Wl���k�����͞�K��䔜J"5�$��E����#�c;tr
�6�n��+�����O��H�����+P{ɕ���b߮#0���~h�0�:�Q��<���ԏ�΂�T���@&��I��xf
��1g&Q�׏�瞃~�_����V�]w|RT�)�Z�,6����	TίC��E���Ao�}3BUд��p���y�GR��7�(,
x���������5�:��䤐�����8�~�E�{��BT/"W�a�g᦯|�E�ABF��y�e�OCe!	�R�9�r�,@H��sǢ�({Qe2���>Mi*Q��͉������������(R>F�y�MMbzb�Bm�Z���u8�s��9��Q.k��!��I�X`�ࡤ2�!7ȯ&���|�"����L
ܪ�����iYc'��pQ�H��g�� ,�	#R�(�?�p�}eyC؎m�*﩮�R��M�`P��YuCqdW��c%v^N��]�o�I��N�C��̴���,r��uE~V�4幢���z9�P�{�q�σ�W<?�ʨ��;�/Ǖ�A#)�YZIqU!�"�4�˙x�)RМD�'�J�H<$��G�*�S�dM���ʉ�DQ����}qTQ�`]M���ؽ�ښp�����|����k&���q�����Gy諯���WFFF�H��\ �͏�|�!�'����U0�0dሺ���)�(�Ġ�EI���.Dc���4q�%���֔�$��ʛЕ�x�e��Jvg�� �G����3�����.:��0�x�Q�m\���0b%7|%��]҃�3��b��؅ёI��Z� g�ěA�QY[-�4L*����Rw�[���kB��l�J+��\'�Z������CWW�hi3���x�?9>��qLL�`|b��T�)�t��M��5
h�m�¶N\y��8��Q��$It�H�h�A�ޏ81��050����pS;�D�+��R>��Rd7W�J��pӋ�6lQyZ	&U2J$�2λ�����еv5��%����x������###���yx�gP��(�$%�d��ƾ�[��~�7_�,���k!��n\��;`�(OʐS@�Hc��!���Ɠ�<�L��Hm���=�ܝw���E��b!���g����'~G�H�v�nğ�[��d5����(�9�|�u����.�����ݍo���⪛n�^x�6�QN&�w�V��?�έ;DR���w|㛸�s�G��Q��>)�L�x'���{���'�1EY麛o�_��t��Z�8zc&���������)��v�,����ߣw�Z�����Ȝ��W���w�@:,\6_��_��/|&!�R��`��=q?�����3ω�f}g'ο�J���o���E�ms/5L�������zF�!��S��]wg,SE�� cf/?��L
����B8��K�{�Ʋի��O�Z�=r���ƛoo����.Ɲ�܍ˮ�
�h�*��jaz�~���Cx��?<P�L��.��"�� :5�.(|�+� ,�/VI�
��%n��@ɢ;9an�� l�	#5��w���Ԁ��Q��C�Jݦ�jw 5� *J.h,j��P��d�@������h%�n�	��� u]H�Oc�����C(����¢����;���&v��7@KW7Z::P]U��?,16mf%i�|������@�d���,
��LW��,�2Ә~w+��w×H�,�w�B��t�+�|c��`��g�;mI�/<�g]������26�O*���i�@�Hy^�0�y A�I��Q�2N	�Q�"�G�a?����0�q#"���S�7�c��>��5��L�6����1y� �m1T����Ս�e+D�����ٓWE|?ey���7z
�S4%��2]yNC:��e194����p�m��?��"0�ʧ�(���Dl���-����F���I�����T~�(P�ԅϗ\�(0)MJ����-Z��-q=�珅e$OC*���oj�t	8>>���!C<�A]��s/9�\u/_=R�7�b��O�ZQۢr��v���l�0�
�"|).N�	����ν��g�Lŕ0��N�S�����]ez%��97��IR)G� �"%I�&tӹ��0�=~=^���q���@�nR7!�����PΪ��J����{μ���
�ߚ�����k�ei�PU�p����v(%���VÎ�� B&E �GNX�
��:p�H��z?	|�R
;�f$��H/��>��F�T��*U�<�81�&A��W�
S3�w����E��bCp��5�"�
䕮����%0NQ��Sj:�*X�?[�u"hViUCH-T�+���w��4e��o��H-│�l�o�^(�F{T:��̌��k�+�'��b�k�2ϛ��P����j�`�oA��R����4Gw�]��[o>�����O�|v���*�2��ő� �EYq_B��� �!D�#�W�ތV�,��+�6����B�@:;D�ŵ��F��.}@wct}����;��H�t���a��u�r�{d�M�SG�ࣗ�ħP��h�|�2v�cD�.MݝȲC�#V0�R��؋�߇ 9�E�w�U��zofu��BDn-ozv<���zL�<�fLP��J2�d��[2�oi��6�=���щ��.��،�4�2I�k:�5��7��*n�5�a��d�ᇛ�w�6\=ɖV��I������c����	ݲ��79
Ji��͕�ၯ�b�ŀT�����c���_�"f.^��D]�r������/���8,��Sn�����a�iB=�95
Y�����w��+����Ef1|�x<���З��QN��<�y�    IDATl3X)�;����=�wa0i�_V���zF
����G�~z���x���~#��;���X�t9���7Ea�����%P�$��G�������"�d��	X�䗰��'���e��b%��aצw��?� ��]���6}�Y�~���(����{���c�{�PQ]�yw/��'��)soU���:����c��E��{�(�o����0馛��Q�n��8l~���<Μ8.e�5O=���W!J �2��d'��/��}[�ȒT9�������?AyC���k��(��Ҍ�����&��"�^�h)��g1��[��X�������7������!q���`1�}�i�t�\�++���b�����������4��:<�8,^����j��O2�s�v�W_Ƒ�;PNJ�@�L����t�!ǞNF&�`h�H�����Ec�GMcX���< �\
��n/[��s~7��	�AJ+���%|�a�Afw�2�4j򕔮��LPu ��X����.[�����& ן���������lv!#N?�=�:s8s�F�Ĕ���,�nx�*;zt_"�t$r�RIYRKI^%=���TF����C��i���
��	xIX./|���j���̸J�g�^���
ܙA�n����"xӭ8?�S����Q__��Q�� �u�D��8	{��Fu�����Gʜt/�d\t�w�����ރ���p]���n!6�cW�E����� �Eώ�8��u�ZΣaX5�'��9����r��(`�G���(_ܣ�o�&�	�+PLN����I�X�>;���}��n��*�Ӓ�#��3p�cOc��� /�-{q��`4]@4;���c�@`)�[�3���Fg
\k��e�Ǜ�Y���T�A6���lЋ��z���&L�w��y|r�?���$���J���~��9X��a�:w�(�w\�=j%����0�]��tⱥs-�-RZ��f*�
d�\�[ܿ�E�hq4�Z_�o�8We�{����>�wՙ�"/�p����'�J񼈉%�Q�_��/��|�kJll]�J�j���(a�%KU�wfƨt��H����E��M��H�y���zqq/�%Q���}���<\�@��UM��Մ�4m���H(E�R8��ǏN
��2����D@��B�[ii��@R�����\yfi(ʳ�iY�du@��	�"?��W��
u��&U��
����?��s�ʊ-|��͝��A��*����%�%L�muQJG���%�^JG�A)y�� yӖ%�.䴠T� �/�N����'6���R�*��j���&�Φp��A�]��Xql���|�X��UGpd�vlz���w�t`�L74=������1�0�6q��$��H8^�e�,	C>?a�t�%����I��9ձH3������3N
1��1e�t�9e�b�:�+�}]��z-����իh�܊��6ƒ�[,H&p�q�T��7��7��B@.�d"��'O���mnF�r+bmm�u� ����Յ��-@�E�3�U�77�>Y q:��1E�Pi���/��w-�_~S�YL�- �4�x������HgP�0|���?�K��:.�v���mز�-|���7_E<�CըqX��'q�S�#X-
ELX�8�c���+8r�S$36�eո����藞E��񷇝p2�܌�^|	�?܊���.�.Z��O~���w4��l�W���G�����l������a,֬{��[��au�`¥`�a��w����^i�f�P^_������{ц��m��M|�c+�x�G�t�N����+0o�2�~�1L��E�ᢞ�`�j6��e|���tt�Ħz�|��� Sn�Mt��L���.ԫ��ހ�g�`(���	����'�p�}(6Bu�8.N%p��^����ā�B���a������|�����f���Y���G�?@2����ҥ+���g0{�<��[>��gNcë�	,�.� y��yx䙧0��;����(�U�Rx������_ęM�>L�q֬[�9w܁��Zqq�{58��vnǮ����!p�hP����`A����Y,F\�mhe�n3T`�$�����4j-�J §-XB��w�D�Q��ϛ��ؒ�ʏ�E�G,=�j��!N�T�:Dc���v���Z��e��Q7 Y-����ؽ�4*ƌƜ�Kw���׏�7LPP^SS��T��C7��,�4��W8MÃ"E��{��L-��y��!��a.]�7��Ŕ�I�Q�Ѓ0��22{��?� tAS���s�}.��9�8݌��$Bajj+����DU� �������W�v��Ȁ N2r�<|�����=0:���kz�p�U�s?PVR���^���3��"8��l�
k����P�p�I#(˱��{�2���X��"�Mh^Ѭ<>%��p��q�������*�G�(X��Y�L���=�����(��0.��
�N"�B��BZ�n�Q�U#�g���(�f�bc����U��h:c"ͯ�����d�>4̘��aܜ[q��
��p+=�B,3ԅ���ڼ�7����`�E0*��L�SD��T���LM���l��% w=݇�w���T�r
$��L��H�XPK�XqBTח"B*����Oe�#hg=�r�$Ē�%	�/����	�.C,�K.Ґ���C&�ɹ��W�(�_Nո6���L&J���kɭ�d^3*��������z�#5���I�E텒G����ԧ�@�zޢ�R�K�+@���5�&��*�Se�Ksfn�EU�~2WEhE���!#�x`u��E�S�]^��Y�|mǉ����/+�P�"���
��o�S|�|s��o��OW���|�UD�*���c��%��Nq�
���s����MTa��R�N#r���w��P�	\�j�x\��俑�g�r�.6� &����'�I�ql�t�?���}�����葇q�c�0~�v�bϛo��a���<a�o{`�aVT�3}B�G�tWv;�D.���l/L��@��� �� Ln��}��x�IX?�[�I����ō2�O�M�G#7a"f�t��i��N/y���J�c]mh�܌�/���s���?� [���&�n�ڕ�`��I�o�E �VE>GoOC	�;{q��)�;r}�W�i����.��58PQ|D�FF �aO�PTCz�s��[�硗U`���X��:L�?W� ae�Y��>��_~��m� �
�0�L��g~�0f�x�^�v����܄�_}�6����%r>q*��[��\_EA�.'���V���>Z�gO������X�U�>���z��.����.�8��_�%|�W&.o�/��y3o�F�+�C+���u�F���u���Gm�$���X��~T�E����2�C���F���+�l�7�e5ո��/`������p���ط�l|�g8w�H14�yK�b��k0m��b�E?=8���M��Wo����"�%(h?	��k�z�m��	��j@ǅ�ص�=ݻ��/����&M�]����+QY7L�UR�r�!;���.�8�D2�H�0�q�r�y�	���
��G+C�ęcG��������(ڍ�w/�}���I�X?�ʣ��)���غi�$E�A̹s�<�8&N�&<Z��?�uw`�Ʒ�qÛhj�7���[nª��Y7J�'����_��ݻp��B��l<)V����:0!��H��(�b�|��I�N�}10�t�b)�p2�d���t3KŁhH�b>AɁ���D�RW���Y�)�u��J�\w�������n�+���"�/[�@��F��C��_�%W.���J4Κ	o�p����E/�e�Dx�����<Z0��&K���8Q+A"�O9_q�N��큫�*|W�Q�~�L)��&���G�O�0���c8��D��
����h.*�\�֜����;8$^��h�(�e
(I�Q�zJ�v�X��̑�� �I��J�eM�:.��=�;�����\m��v�L��+�Ep�
������p_��OG}�C.z���zy�u���W��K�)��P���('�.�]잚�H�cѓ���[ ����kB��v��<	���Ae>S4�'c�#�c�\��p�����'�"��!��C����EZ�Ʉ�!�Nb	4�B�W�R�$kBGN3�rq���P{�dL�?#gވ�Z�8s�E�b~��xt���M��ew��E��	��d�,Hy��],8QL\�E�)�������b��������� �*�K�����S�{H�)��_�m��G�X�Ky"�%�^Q��{���
 �&��x��
-�����o��8DX�%HInW�.�Y�v���$��C����Ԩ�g*Qa�J��8Ld/�s�k��Ńv͵�����B11�zG('�6p}�Y-�1it��&Gi]�l]�%������'.Bu,�ڊ)��)��s�5�8����p�Ҵ��oA�oRE���^���|��w�.�2yu�E+�P����E>�R�{� \�W���b�6�.:O�@��;�`���		��E����2�N%��%��_����^8�Ǩ��1��
v,���Ǒno��>�t?c���E��I�s�#XA>�ߏ����e�6�����NƁ'Ҁڙ7a��w�ۀ��v��O��rkb��h���0���EYyn�!�5.02"dpE�"$��S9Q(`�P��E}m�L��7���	QSS#��ҥ���&=�2S��Fk�e�<y�:�s�DpL�h<�Ђ��ڰ�UaT}5ƌ�1cG�nD#���W���Ɋ��̩Ӹz��OA��($���BQ.�K

��>����%�i�lɜ�����u�r�\̻o&�z3
�W�L�G����_űC��ӛ��c�ͷⱯ�fς��f�it�?�ͯ��C;wc�{=�i��q#��Y�;V.�/��哈u\��=�HA~��ɬ�P�p,]��\�H]�=�f��Ɩw7���H )Â�˱辵3u8Onq!C��sضi#��!1r���4+׮��%��(�F&1-����6I���)�ъ�z����{�]��*׌B��~��1vl~]-MJ,��pۂ��w?z�d�|r���Dө����&�5_@Gw�1Sg`���1n�l�<v����+�N`��p��1��c(ibʌ�s�*�2B��~�g��Ʊ�{ĭ�ʅH���6`ѽ�1�
D���Z�LX�8��/ӊK��"K�p�p���X��>4N�$���K���{���!�&��Q?.�A�7^
HnXv6���Kؾ�m�߻=C)��~�0{�ݿV,W	��B�d��pg�C��S�c�X&2�1)��&0\���s#J�ZN�����!���±����3)Yvɔ֩T\��C&�FM�
�3�T�̡�r��,,F(�Aj�t�r�9���+� x�����~�~���'�����Q?u**'L��`�Z� ���!I�堀�|�c�ʚ��p�d�C�1�e�ڦ}h��>ۯ"�t	�T
��;i"^הi���^ę�~�+��Y��������Լ��ލ�d
�a���H�)�	̎(�R�h"���U�=��jL~']�:P��LI�Ќs���,�Ap�4�]��uPV$�@[���:���H�cG�5D�ׅ|0�@U����$�3��x��!�X�`�ii��4�O���3E�y
F���K�0�t��,b�8�&L�]�~�n_
�[�kF����;y�� B�<3#��ƒ��.2���o"�R8��~hg��$GC��a�.$]@�dCn��P6n4j'NB�P�{O�*���
y+������)̚=�.Dݰ1��RYN��r]�`^:��';����f�^�N�¬J?#5"��bg��:E�_׋�K��n;�t\�u�$���d�\u���w5ɓ�8CC�kςUq�K@�z�鸜ԋ{�^�6�t*��^�*@�=��E2���@�����2ڣ�l1���D�E�Qi�b[�J��<wQ�@���b1@�Ա���I�U�a'�D�ⴰt�D|��.�T�q-��*�)�,ײ�UQH.ǣX�)�bq����������h݁���B�����S|�ѕ�e��[o` [�)�bٹcǊc��W�3��}�3X�2�)����1�����K1E��xn�OF�*܄�v�Oj��Q�pds�LD� ���k��&ڏǑ�
->_>?MN����:��E��V2���"pľ�8�y3Z�생�i��i�V"�f%P��������q��q�	
r��ȧ-�����-]0j#�}{�@�Q��%����k*2������#Gb֬Y7i"F��
v�8��2�( ?5��Ֆ+8z�(��=�����b��d��e ��������m�%3~FM����ށ�# n�eaF-}}�>|[^'��L��N��M�SZ,�b���%J��D�sP�ޗ���o��ܽcg�DA���H�w����ع�=t��`0���W���'���)�ax�i��ZO���w���3g�V�Ϣf���rnZ�ވ_�p�x?����䡽8r`/�4R9��z,Z� n��N*����,-$�pf�>�<t�ͭ�Œ��{���q�Q=b$4��s��֋�q��~�:vT����G�ęX��>L�y���l.��`?2�8�s'�~vTB�8�%�g�Ca���!\U����qt_�����Ĺ��L�Z.?n��7�6O�߄���j+��߃S�@6G��0~�X��!Ԍ'���ѩ!\8q�vnG[s�P��θin��d�0�f�O���9��ϝE�P���Jܹ|%n�s*��p��i��^ƁO�����@*����W`��e���ɦ����	��{��J:��ƨ���h�=q��1� ��9l߼	m��Ț6,���3�b��3a��Щ�%�x�S\8|��+����J�
��ؐ��~�$��%�'��NA;�⊴!���b����v&?�H.
E�Y��|g@9����J�@Av2Y�R���	Ҫ��������`E���0l�}��ɀ�E��	?�o�3����gՈ�݁�7ފ�������@ye*���JW%}��
�%��V�
�%�t.-����%"�*x�ΞA��`�)=�	��	�n��Mmh����pFm#�e!勠u0��l����=fհ�)q��~"{@I����%ׂ2X*���D�00<R�F��gGqj�@[����30������r���'�#�ڇ��æ݀��E`�.(�}��fƋ#�>tiSF	�C�f�BR&��DA4K�I�"�֔���'���^�T��xfec�a��O`�ܥЃ� ��64�C4��W���&U��h,I�4ɰ�*�²`R�E�!f�X�Y����������)� 4l8,w�hʪ��Ay%���<��O��Q�p�w����ƎGB	
��pG(e� �(�y)8E��\�E���	��.[�k%�3^�ޯM����L$�8-��@
h�(q��tB��"��\uO�(i�nHRs��d�!B�#R��R��DM�<�ҹ�4f�e�ٔ��b-h�r��spm+=���Ic=�>�rѻ�Ef��w�8���I
����bV�LJD�@�(��P��(����l,�4C޳r�S�P)�JBk0'D_�@B�J^��E�Tj𲞓Ft�y���|0z5�Wt���oA��Ǌ���{r��g�}�lߺ�Ɂ���>�h%�**�c�s�"^��S�kc��u|=W�7��}��5�H����$��E��F�r*��Ȧ��dS������ -;�����K��ɏϘ@� �uX�r9֬���
>;��];Ѵg'r��7܀+V�l�bi|x`>;wLT�&;:~�,C::����xC@â�rԫ\ J7�8�6�nB�2LL;�gN��	c0r�(��B�r�����F^@65��`/����ĉS8��.5��ˍ��{��}&���t�H��9^CG.6�hD    IDATo�����LA����(�Ι�)7ϒn._�G/��v~�do�t��A�*���,���/��ƙ윣]�Y@�`��L�s��>�'�W0��܄��?���{����{�������B-�4f#��3S�x�S޶�L_6�X�Bݤi�i�L��&����"�����v���M�d�Dk0o�jL�3G@7�t_�:[����z�x�8�!�Y��n_O$�W��c���4�;���g�e��X:���������q�f������م��^q�a�����5�c�Y����Ѳ)4�=��{����p�X�����w���E��w����Kز�]�6��l�I��fb�cO!\3L�'��C��+8�w��/�bP�{g�r+�-^�q���]����c�����$��@��n��pU��{��L�v~���ڤ���Y�}���.̿k)BU����u9�j����l��C��T?�ogl�M��{V�~Dc��[����ID:��m�$<n򌙸1z�xY������m8�o7r=���SÐL)�P��BF<��$��ǌ]b�態��bd��(Rs�0׊aY�3G��E*�%��̯ +@Կ��tp2��l ����4	�s���ƤS�+E���:�"Q�g������5i�
 ��x���?܈�X?�L5`��/8��C*�E8R�h�^��FSv�,BB� �|��E"�H�%����B/�r�f B��A�����.8�|�a�C��=�v
Z������z� ��c�E��ˀ��d����@ͩi�;&M��j��Y������}���M���B�Ǐ
6�|�����	��Ah�T��o5p�B�>��W�p����v� B~f΂kƭH��(�4˔��<���R�~�N
��A2O��C�0��x#�@75�:p|�v4܉
#��
L�1b�L,Y�4*���~t��=;v �Ӆ�B�����(a*��LU�E)�r�N/9��9-�t
��ۇ�Ǐ��@B��r��!�3��7G����O��Q��gҳˋhYǎ����P[����QV^'kߣL��$�Ғ��d[Ph\���9#�y�E�!q	���s>�b[�:��|�F�)���s_*ԕQ�Kjb��l@���?]�P�	<C<���t7
L~甒�+����_���1�G�����|�x�tńb+��9�0d�r%�����-�y$�ޫ;�M�6��µ�V�m�ޱTN��`�<7���z*~O2褕7�)A�j�r�S�
���K� 9/%��cu�����4���ׄώ�(�j/�u�(X�s�e�_��^��}�_*/
��#���������';��Z�Ndu��C(\�p�\:쪑//I{�-�k�J.K�qM�_�C��\<XPpR��^�����h���/j�&w���L&-i'��R�䖃��
yx��<���2�r#��H���)�Q	�������Iυ���7��0Z�;���`��zBH�AĲ2�.�ۯ#�IK�9"�f��E
\|�VN���c6�q&L���G�q�H��{|~�������@o�z;%觩�2Ν����	��?t�#y>'���C��ÝK��7A�N�0�V�W��_yc�O���Q��П�g��Gϕ+��^/�R�D��z��Q"=�ZsQ%u��Aq�Fg�D��3�݉�s�@U�H39�#p��~'!4ݒR��f݄�<�`U%���1l�!ٽ>����,`썳q���3k��M}8�w7>��=$Cp����-���1̞7��(�f��N\9s����>	�J�r�"�}�ݘ�`)|ee��k����3ط�#���,�&���1So�ҕk$��� �2��q��>l��=���2���sp�"H&m����ִp���ܼ�C�k ������e���NP��N禋gO㵗_Dӹ���gmJ���[��+��U��>��<.�?��7���v-r-�S�-X�Uk���+�jÐIȁ=���_!��GA�yU���⁇qۢ������N���Yl|�Ut�\�[ӑ�$�{�]�q����8v�L��/�=��7��=۶��������>�(�h]	j����－�|f>-bP
y�P��c_��qeR@�y+���M�`�Ǜ��lEC�!=��+m"lZ��i@ЍaAB�&�NR�p��&:/RM���GR�.��C�u;�f^:�ir��'\g99O.�sb#�$^�Ld�!`8�Z�
*P��F?������#�L�#�!�t�W?��m� �}�1u�Y��οI�@"��P2%�%�>]L��Y�V�!^��%k�h�������g�D�L"��޽hڰZ_'\^Q�a��Ed�b�f�]�ys#���'�Ƥ��P��^pP��p�!y~WAQ=��N�G�8�����)��E+Ō��/��\8qg6��s�,�|�qc0v�*����@2���=h��m�[/ �`����mR����H�:��f���ҕ�6D����/=t3�D.&�����/�H��`9���Xk'voz'��w�����/��'�}�T
���ӟ��.D�{���^��
�^լ� ���cfe�ϋ��!��
�������z�ԁA+��BCvi7���P9z$*FL���7��~��KlTq+mi>��ͧ	�1|�p���t���H�����
'��_��Ȥ��xqR-}���̿P:��ћ�M@�lv	��DLM�TM�܃�����(z�&׋��_�z��gu�*�9]G
`M�4g '�@9唄�J�/�C��.=�NJ�}u2OȐ"����KR����7N�(�E�%�N�%�T�yf>�|a?H���2))�.�;)m�"$�@\�J4.U��!�����&��%f�lV(p.�rw�zc	���ѡL�5͕�P;|�'�u��$���(��a8�n�^�4��u]/����A����������" ���X���-�G���-���Ｘ��}�ブ�g�n)+S�성�����Q����q*.%���FFe%v/M��x�����&W�=��d�+�f�K 5z��]0���CIU(� ��8\�4B�a��t�8b���[���|tJ��֨�ˍ'�.3&��>:E*�r���IQ��I�M4�I	��\@$@�����!�C�b��\}Gn�t<���Z4����$� ZV!E��P��ƅ�B">���vt�wHo��n�N�f���3�?r�2-�e���q!���P��� �O؇pee�(����ml���P�����pұ��Wd<:;���L����*F�ł�������z�(ţN�q��Al~�e鎻h�)x0s�B<�ߕ��a.-�do� �mﾍ��^8�K��cf�������#T�����n�`6������������������W����� �� N܃7~��L K�Nw��Vދ���CèQr��fW��Gﾅ�[?R7���<�9w1�<��L�)֕k=����x�W����_^�'��5�_��pTMǬ<�ޅ���'>ݏP�ASyDk�c���j�CG+$9� ���#������G$�qb�,��;�?�_߁'T�P8 ��G�cx�ş`�';�bQ�?�����bͺ�1m�l�<�@w�y���>6��S�tQMK�7E�\��Z-�'�B&������s�gO���,)�|=�ƌ�ɉ����Ilx��蝍""�'L����l�Z<�ů�n�p)�n7�[�����?��h����`ᒻ��3_��	�$�@�t6�����7�@����A1@<O2��e�J�<��{�mh�ݶ�]��ס��	�upK�>n��n��Ĵ`p��צ8ld)�s��6�� h@m�p`�?Yb:T�t��/�4�艄08y��{.��~�6��\�t?��!��=��nXx
�0RZgڲ�Y��uY'����ӫ:���%�Hr\�*����"��D��Id��C�w���̚
�-���Yˀ�~d>�G>~N@��w*D}#L�% ��� wKB)�GI_�rkG�%�\E�R��Y��'Ӆ��'�ΞƩ_��©�p�)xƌ��+�_��Tql��T�h#��.��������s�*������;����3�.y�
�"L�ԥqR�KȤ���!Z�?A���ra�r>ٰG?�'օ�/�L[����"(p��˷нm��]�AO��kZ����GqR�%(�%73i<X.
.7rR���B]�A��pE���|�5��1��F�,ǇXl�=�H%z�� �P^OP�{�2�^D�(��q���-���s��`E��C���F�S*#.xg/N*yo	0(j�>�C�e��l��_��q��r~*O�j�yX�4-�J�����2��5/ �Xh�EPP�{R����}����A�8�I���?$���ё:�z�$�.M ش��MP�^���TZK��"m��9�9��(�����1�8���@Q���eV�;bj����-F�,
Z�z}C�7t���=�?�m��Y��
�ۓ�<�q�v!����0<���5�ɣ�et��`��.��v��a=t�|����������H������M�������۽gN2�����W)��HVu�ݼHri��K���ǋ�(���3HɒT�hE$]|ՅP��,�IJ�S��0�ؕ�C˦2,�D��n�b0���W%�#o"���[>�A]ЍJ��Z݅r���GG*�6�:�R>���������'�N9�\�,���̥e�T]��qQ�2Q�/��@ac:�{�h0��24�h@4D),b���1pa"��� ���%00�Do� RI+�|�� 
�yDuA+w&.�� ;@;�*���ӁFx����|3���[�a2|m<��HKV�M�[�V�U<՜����A�z#V<�߷FE�R9%q��a�������}��>�2&2.?f-\�����Z���*�|_�y����QH�����7��,��'��[/�+�������x��p��,�0�b9����˿���l�Т�O%�W�����O����e��,��G�g���������DK��ɣx�/�Ȏmr\(�K8n�Zt���1n��y�rj�vw`���H�LP��j``U�F��'�m�]pE��x2�8ux^{�|�*"AI�TT����},Xv/���n>��N���8qpj�+�%Fq������.B5�*0��A빓x�G����1lƴ��օ'��:���?�^b"?Ѕ�lī?�!:)��d�@�i�ҷ~Sf�
��g��.��?��_�ܱ#��Œ0!|��Ľ>�`m]QTd������cǇ��L��H��U��G��#_�&���D1���8<���s����E���NE����Jض��ױm����҄j�?-a0�� h��qu>j��8id�/ύS9ѹ�Z�BCإ�`�r�v �=�<�%�mɍ���x~�{G1��#�D�˚x�(Y���s��z��A�c.Fܻ=��!|��|��/�jo��꩓���0{�j�ꅂd8�0&L�dX�g�i"�1JD*4NB�0�䒠��`���O����л���3H��Q���v� Tt����}�d+R�&-Z�ʥ+�����l���,��E����Z,�XR.!IUU�@ph0Akj�a �<`���K8���pN�6�cW�Bp�#@�
�L�m�h���-��4���s���nÒ}���v�<OG
ѭ�N�v&��Ȱ�5���
00B^�|��ǰ�o����a��o��Aco��{��&�f��nd6mA�{��v�~Z!���$�&�@U^�B��H��ݪ��
B��ѕ��#À�à�C֭!PS�hCN���௨��*��J�$���.�����)>�Z,"k�+���ǟ!m���"�f3��>_P&�6�<n�@�2��#hJ#�މxG+��	�É2]����oQ�*B�|=Ӓ�a�Lf�E��:in�4'=��z���ĉ׮ڷ�6��%�S
j
4�pH������~���He��A���J���#�sӶ�K�P���e�G`������V�q��Q��m�tB�].M%�ۖ2�)�*�o^۲^�������VT^5��� XN[�dR&$�W�A�o�Zfs��#@�bk+|�}�e����M��w0�,s9ꆵ����a��T�txݾ�]��s�.l'�8 ��zZ7�+��u]��^��.<�ϗ7M�oVTte5�C����G����;NO�������������I�e��{B���yqN����ҖGR2�+���(�8
�hn�ZE���i�����,>K�!vԍ����a������i��D�ȣ�}";���,�ˑd�B��'D�.��� *8���_ބ��1��0��w�X'�Zi�'��F=�4c�n��AD�*�E�@�rI`T�Zp��'^⒤��J�TRx�\|�!ʢ!�E�}��,�Ҹ�qq`��"�� ��b(���@6ǖ��<Eq���V@��KJ'�����h���X�q#"�Tx��
O	ϔ��8.�Eh���P���5P�$B��é��7g.���q��p|L�5�g�9so>�Oػe+��}���z,}�!<���#\[x�JJ#�ہ�����*
�r%,L�e��iL�C�P�y�b��w���/�ܩcB�d�5_��?�͋��x8׀�K(��_�1zZ.K�'�
�#��g��;W�w$�Brit_8���_���?��}�p�~�<�0j���e)��\_7�o߂��,��L�D������`��%��h��������K��ԧQ� �!\]�g��q��{�}
�Y��������c���&giW�a��ux��/AF���S�+MX����s�&y�$9|���z�:ڢ��]��Þ�����<��+����T`ڜ;����@���DZ�F�3����sǎ"�M#���0z,����qۂ%�L�u����&l��O���L�u
V<��	d�`b��[�}����h�����Ǿ��"ıp`a��ͷ�k��7_D�[����=4#��?�E�WGc4�z�!��Z����	 E:-A/ן��CK0R�V�R�T��� .&Ӳ�Qr_��$�HB*VT#� }�BV뼧	�m��� |K��T�a��������ǯ���_�A������V����'Ҥ9����q�"�kbѶ�w(���N��Y��aM�!'j��p����Y���ӈʇEx�- ��/\B�����1h5~��?5w���
��d�/�Huee�6ɑVk7��,�dj���eH"�zH;�k0��|~�
��v";tNC9ƭ�Q���F�?���>@���u7#:�3\ܼNY,�A#! ��Y�u��i`1�I�l�p��x����娊jD��C�Kb��w�奟 �s>W��񦛰�����9� ˏ�;����{�4��ǩI�L���N��΋��t��nF�����GG�4��߃�l)CC�V�!?�ƍAø�VW��Dw�#�]#=�ם�*A��kJw��BW�$��@��K�z�U�|���ɮe�L�S�g|,8�6
l�t�#�z��+��i���}�o�.@@�m����w����R�s�@ "�\�x��[Q�&���<nRg����	t��\2Y������J�h�se�!I�4 �����G[h��E±�P;~<n��.ԍ��V�tj@�v&�B�TG�wH���#6�T)\� ���/4�\�SR)�xF�Zuu<\gsYIdv�:ܡ |��X��?ºZW�D��g���u�2]7a!NG����\Ü�>�L������~�54��-+�߂�����nW�-Ֆ)����|[��4M'|->8B⃌^~��r|h�%�,9z&kX^+h�3Ú[�V|����/��4,����B=��$�-��d:�P�C�H�)�	��x�ə    IDATY�7�R@���+a2�)��@x�D�T�+*��穱�J�c�or&�ٖ��u+���ꐛ\��	WƁ�` �� �.�#F!\[�p8����}ap�|��0L�ٚ�Ң2@S�U��p�[/����T(x��)�"�J7�ԁ�nf)��	��@\�f�T���2�P�A(��c	�DUZ�G�V���,���D<�B,�A��02]�S�D�����)��,bA��QrW�G����K���EJ�CqcUv�Ԋ�_�@A�77��O8�ŝl�������ٯᆅ�ħNF>��s'������Ʒa�~�3&j�OÓ��6�X	O4 (��࣍�ŗ?�7 �;�����U�`պ'P3vD$��O�������Wp��Iq���L�>_��a��7��O�Ddbh;���;��˗�V�}i���x�k������1���fly�W�R���;k��*n[z�Ѩ\�nÁ=ԇ�'���.�=�ryPC�ѧ��{�T� ^&В���O��W^��{�s������7�o~7-Y.�,��l�����m[�ya���s��U,�+��-�Ұs�w]�;����o�G��G�������w�`� �-�s�>��!���O��rI�(��j̻{z�K�W�!E@���Kg�� �B�ԥ�q3z��`���@�ǃ�]6❭��ʋ2=��I�5<�,��}/��
��E��n��M��s��+�87�U5X���X����܉��հ�qp������H6_D����A��z6O6�Z��1�eh�0eX��t!�9��� �ԡx�촫��uWB@e���GłOq�E0Z�,�t	>���29�a��\�[��[,r�^�EZv"��ԍ�K�������G�j8���<A&�^
;\����R��I�Up ��	�]r?Q��7��)~�G���^R�z��ݿ��� t��e�Q}�tT�}�)����±�8��s�t"2�
#��w����Q䙇�Ǩ�W�lFʳ]2lXr�"bV.�
W"z(^�P%���l1<���5�?ۍ�`���޳�+*F	(�x+.n�%:.�|rf�}�-ˁhl���@sr���l"�&@4p��ŷ�S�)K�o���+�����~���4n|[^�	�������M��~c�.� r���7߅��y4z��TQw��#�k�Uf�\�4јd��a��$=���sd�.$��K�;vFN�"i��J8�3��W���躅O��D�8�)��B8�I�Ҋ.��
��ҥhii�����Zx��h����	o0���Z�_�{�؎�KM�u���KMBB�0��L����	͇8��ee�%@�4"��JN1����_c^=������UX�^�ܴHIe��L͊����-�RR�g٢�ഐ�O�n��,V0qi�ݖ����2�֬��i���E�qf�,I��Ҳ���\
�\�S�ϣK��&����$�bc��O&k�d?�/ �����QW;o@jYs�	!��������/���oF׶������p{d&��It;Y�'��'�u�k���eͬU�J�_{��Ϡ�qĞ�tKL�zV]à�A9,Yd>��~��Q��_eՖ���d�I���u�A�tBx-W|?>�aE�wl��w�������e4]Ӳ�����d�a��9��MC3E��k�eh��2�b�4K��L+膦�.M�\��q�5��L��8���4C���[�5�mt�cܚ�pk�F&����^�-7i�9�F�u	ql��H�m�֝���B��X~��k��5��YféK��UW�/W�
9v�8&T<>�E�R��&q�����őN*�9�bJ]�j3Mdr��L��'�6}�v{	
�_
�����8�Ä�"(`q�����'�ʤ��-�X�(	��/�q�EK�0~<�/�.3�Tg�\����Bh�8q�����'�lŎOv�蹳H�M�6�����HD���\�P]E>���8���'soe�y��>{�3�S�\�<�!$�BBlI�eي�t'��޾�Wҹ�+��^Iܱ��Vd[��,����A�SAAQsթ3������ۧ �I���Wj�j:㷿�}��R	+�2f>J~���5�����,$�Y4Z�p�Ig�5'��e�qP�P������B�P�@��wq����I��r<N)CN\n�,��9�Ĉ۔�`�����p���/��g_��9s$|�ˎY=gN`�/~��7�.��/�����"NEL¥����=������hi��ES����	?��U��[��~��|�!�۲W.���/��1���x�G��1��M�Hm�Ҹq�~�W.bj��D���qS��~��wφ� �!��6|�}3>zgz�ۑ�u�0O��1�{e��`/����v���/0��)Z�H��.\�G^�!ѓ��7��Z�^�>�p���==}��{��w_��� �cb��e����8�g7J¡AP�ԋ?��K�q�+�2]����ob�淐���[�������쥫�P����ߋo�=�r-��%��|-x�Y�2�r,�;�X��?���8��Q�]�	S��cOc��K$���\Wvm~��مB*�D:�a�&��g_Ĥ�
�����!'�i;~��GX��A��}�i�]��z�~q spx�|�y��/aH؏-P�;$� `���cdY)�~D 脠�'�V��,F�;'	���Ċr}�@�@z��t����e���F�+α y�A�'�ۧ�P����@������E�QE�찉r��;����?E��Ey�o��U�{#�͇S^ǡ@��
�8��U��ƋB|�aF(ʈ���|z2�u]��F;��.���نh����'�b̓0&M,?��y���BK� �T���C��@}2ZXR�im)��x���S^/4IRo��63/�C�l_�Ye��`�?-�.��̆7a?�|����,X����^�$ld��w7���9T�k�Ұ�- JHҤ;�f׋$/����Ye+�L���cW	��4A�FiHƊ��;wa﫯 u��Fy���	����0r�R Q��1�y{��Ѥ[��̎��c�z�dR:�F��̭  0�Հ��FO>��T��R~�>If?TV�a�H3u�F��q�R�r�6����B�-jm�X��;

�4�R)fC�Y�J'q��5tv���GYE��b���D��0��C@�K��.t=�K�F��)ԅ��Ήd%�lS	w��a^_��Y�������;�)�ٜ��D;(�ݺ4���)��%/]~��(�1�?�,3ڋ)'+E[�E�,�>&"�0r��= @���h��Z�	\N�H��ӧ`�SOa�w�*Jc*�F2���h�������,!�0m�U��<^?)G��E>�lJ���Ajyj�����}:���Z
N?�a�B%�KdR^�!ҟ��]�qc����4�I�+�ǎlW�4b��bܢ�[��'巯��o���~��
\�$�m%�m��M��r�8V�c;��r���~���~���z�.�K2���tP?'Ms� �p� �:�R���SA�2螮k��K�-|�qEܴ5��X9��m�(h��k�fۖk���Fc讦��m�5��p+fM�|К�P��J�uXi����ʿ]�%�n<�>R�2醫���t�RSG�l�p��K�>��|���ۮM4"���uy��N����p\�Q�]ٶm�4F>����Bǔ1����v���k��i��RL1%���_� �D\����_b` �,-C92&�a�S���%8*�H!��"S0Qp�CLI�J�Q���DL����Fj��ǖ�+n"��*&[�&�Vz67���h�dk@�;G���7�y�w�IO�$�tH :r�U��*'*�������;۶��S��K�p0F�!C(4��V#vә�@ �bܧ@7i�3HWb�פ_w���f6+�6u�*7� ӞC*�=mG�MR��;������h�AM@���C�2%$Jз������X��)+2v�d��Ͻ0	[�y��b�^��(���'�:1c�j�z�E��{6��9�ӈ�?�w_�G�޲�dn0��IS���1�̾O9��O������G;�a���
t7_�O��G�����`���B�N�vm}�N#/�Df�Y����m.�Lq���~~�w�߸�L&'������og̀
�n�f������w���a��}�4jG�������M� �_Bˢ����3��O~�B"!$��aƜyx�{�b�z`�]���Ǳ��Wqh�$[���s�/���^�m��QB�r��]�I���?D	'XU��x��#�3:=�i)k��h������m�R�
�+����?����.5a^�<�D�|��6���T��?��K�`��O��@H�45+���x���ϝ�\�����8�=��O���Uu�S�����m8~�R	=u�Fcݓ��m���ŵd������������C�UVc���q�k�s�e�\	��Coo��o!�z�f��n�D4G@A3) � J��MP�N:����y-]Z��<����@���cJQ�H/�߳���%f*��[���;�˪@VbF;�����y�[�y����ɯ�?��H��+�F��1X��g1b�B�5����ͦ��w۲G{b������T�e�ϕi+ih<6D�E}A!C�zz�~yg6l��ފ��E`�04<��)wy�H]�韽�\w"͕��~��,**��QG^6�h�y�/��r:����"UEg�ĉ��a�+� ��W�qa�&X�|3���M��j�Z�C����I���6:[N�rt=n_��>(��d�� H�! ��
�K�Q
H_z���$�P!bl|�͎{x��ڟƑ�����_ �z�sf��a���0f�
��G��܆-�9�z3�2�nj���0A�,���bJ�Atd4�f��tf��60$|:2�bu�5y
�ƎEUm#B��:��2��s3Z�0��l�98�感S#����M�R򯽣--����)�I4V����T�ah��;�ƌ�lrU��>t}u�7m��O>BṡX '��!Ҙ�\νh0+@�{�=�ߧ�hRPs9�w�<b���T~l�0.�vˁ���y-ɨ�tb&E���#����YY}��h� �^~:0�f;�m�M%p�tܒ �-^�u�{�&O�W� sYun˴ ���ˉ��bvǦ&!�Q�<�-����%�s�P�����x��4���ĩ0��J�`�5�"2A���Q� �އk�Gׇ ��Gy��*5YiIv�EK <i&,Z����?,��������߼������>6�I�7��,�t�h�]9�v7��Z�U�����J[
kQ���������,ߗ�H�d����B�&U���&�x�-I���ɽ巊�/�L�7��ֿ)"�S��������I8�����K
wn�Z�ύ�PO�� ����*:;P��� ��y�`f'�υ*yE'q��w��j�戮�˗D�� tq#��<Y��v�:�Q�m���ߥ3 �d�X��I��t������xa��>	�s��]�=�ǓH���XP�û�8Y=�b�7y��4�իx}1�"����?k-[�A�őe�DQ?q"�?� �{��P��N�����D$5�P���fDk��PH������i��8{��h9-"v���h�i�B�c.sB���'`! ҡ�Jg&�Y4�ב�&�WD���{��+�:~��7���؂���h$���e~p��X0h�j u� ��ý #�����]��\��U�>��m��I��x��-�b���ȝ���5�5�ގ�k�a�s��лg�څ�vz-�헿��{�"�#4����x���c��e�.IF�l�tڱ�؎Dg���Be��Ø�r"5��9i&(�����ع�m�9y\�R&ka�̹x����ǡ@pb��[Id�Z��o~�\_���
B5MX�f�N�-P].X�{;q��8��~��:���r��������f��H|i��>.�Bn�!s"&�q�<����R1=�Z&.��
��݊������ĉ�s�=x�0���y�k׵�z�W����AE,�T�P���X&:�y�����q��x��ێ�hH�ǙKW�����B n:.����x=7�����@�,X��zZ�D��L��<�.������-ı���ͣ�ᱧ�ä;g �R�mN7�����p��	�P�(�����+cj��|m��g�f���@Y8,#��Z�z�1
�!��b�������oùq�~F6�Br@�Q�P�	��@�@�	�39B�7\)΋��Y��S�fe�n�**M�����,�{B�a�OY �6�{����(P�_��߇�X�s�H���r�%ϝ�O���D���3i7
K���,Y��t�x���A����F�Pޞ.�mL�[�)%׭׃��+E���ub ��8N��٫��G:�[��;�Lp�:���&���E�������@e%�r�ć�`����7�
:y��"�P�a&���Er�O��Xi)Jʆ ������i�����[_���� 6gP����s8��-t]>��э��b)���r�t�� �{�eR �>�7�Y��R�6�{>Tj#((ea-ǣ)lBsJd�������/P�lE	
�$P1z־��/Z-\����[��� *����ʔ�UD���s�%�̓f C�_�FW&�鄈��= G#��Ԣl�P��:�'MF��Z5�L&��5�-D�A��*���<�y��b�r^� ���Q��Db@��>t�
���$-�y�H45CmU-F���F"L{Z�K���"���5\ص��C���"86��K���� ۑ�!�wj
x=@U&���$�UK�4�����NA1�{���5�� �|M��!���s�Ԋ�/*^���`s@G�.J��@CR7p&����n��J0{�*<��(˴q�2�i��-2��D:
6�Y9N��,)��I��}R�
��H��I�6ܸֆx2���*DKJal\S4�[@(BY��F���x �{��4Guԇ�������7p��Gp��?l�sƋ�SW��w
��w�3ٗ���|3�k(d�JQ��̓���n&��);1�[���K+~���̑pqk�y1��f�s��@�X_)F���9&�
�bw��7E~x�s4$H��D�ܭ�^�Ű��A�[)�훡|��xm^^'_�u�{/~��`����&�*�"sdȅ�ߔA�g{㍰=[<��HwIa��ŵ�
O�*��nz����*�U�─���X��]�y�J���b=�M!K����Z���s�!JPp�Z�^����v�t�1�΋#�bxmIU��z���:�o��ȟ��,�Y��NA��Q���<4��e
Ш+0)����p�n�p4m�ᘒ�YF�Н���-�Ue6�ػf`��w�5-|��vl��6Zzz-���Hz�H��#I�u-�[_�d�(݃T`7j.n�ܬ�p!�%���� ˒b��!��kꨩ��0��:�GY6U�;h�V�Ơk�2�GE�?�M��<T��!��&ݙ���(Em�ű/^t�P���U$@�Y�v�`�5K�H+�ɮn�Z�˞yCg̀�fm��|~�2N�e%�HS�)�C�|�V���pԧh;�Dxz`ǻ��OP� ����UkQ?fu�2��ї{w���#�߇��
YK��M����G��q�#A9h�N��啿�90�P ��e PY�Y�b�ӄ�$|�D��:�ށc�If����UX��c�8�^���|��^���Slz�7p�򜥧��i������B�;�:y�;����c$�n@�l:r�X���b��Ep�"��EM��UUHґ��O|�EI�K˅��=��Z6��*�ƌ*�Ͼ�������Y����� �n���t�N3�����?�i����� ��Z������E��cxw�ho�, �'�B퐡x�[�a�]�d�"�Ѵ�s��?ڃ��@����d
�.[���!\V�x����������A,��    IDATx��员�����`�c��~��DHSS+�mcϫ�M���A5Ag:��?�h������4JЂ�ƫ�8���^,de���C^v^��rV��ε���<d�&���}���1v.)�.����D]W.L�Q���3Ö��>~��L��*^��?�����LCǍ��o=��kV�*/��|��aE+�ż0�5�u��k����	�b9�͇MV'ߜ¹m;`����'�k��u��ـ~���h?}�r?�Θ���@c��1 :)�F� � ����7ՐJ���c!~��W.���)v<��0z�ih!��m��@��y�V��j�X���Y�}(��:p���8w��8w60}=8���q���p�Y���(�?�EU�_M���]�:�ry�o�ub]0�������_��� *�7G���X���x%�%UB{�ڼ�����Z^��抖E�5�{��*�;�] �=�&��o��4ѭ%�Fa�;P;b�G�A���3���TǛMSN8H���WH�!Ґ����N0@� ?8�O��p��E�>s�/�GyU%�6�FMu=�˪EKPS_/@Z�J@��V|��_�Ԗ�.j#��M	����u��č	!��<Ƀ���. !@޿�)N��SlD�F�X�{׎h~��6�0��<� �t��(���3K��ʩ)e23!\$�ޔ�� .�38�Վ\I��=��_�>b�F�zJ�T±���AO�G޳
���t��	m˄�=�V�2q��N�7��p��%$hllDmm-2�,,��֢<��B$X�=�@{7Z��G���QQH	(��,��Dڴ�c�aԂE��L����IKO������&���e�5�&<0Y�J�]P��_��*r7��\t���J" 4�
�b��H(�`�*��_�)Soj%PaQ,>՞�]8��4�Tr�k�:Y@	Z����R�yϡء��V,�H�� I���?�a��@~�/�@($�w�fBڤ��HgK�@��GQ�,H[
A����;f��&C���"/A3���K&��f%]�z��B� "�����Vi{��N
r��Ò�]|N�T�Z�q�r+���@Wg⩌�̍`D@����
�{�	���]&�����M�C�B���r0��&��=ܓ�ʈ�n?�A�m���kK���H���Q����E�0s�b�3i|��lܴ���.���H��z�^#�
\3R/�a��A�ώ�a �!�0�oHA�d2�{/缚����� 3G`AK2:� T����;�g�@�]T+�:Ki��ާR7A�k��~5R�:��.�l��N�L٥�W�1�e���Z˺�������--���r"��K�c��'1t�=@�cW%�m;�6��e\<�F���x
	׏���._=,������&���2}��A"cc��u���!��s\�{�'�ûwbۆߢ��Ukn���ѷ�'�EØ	pä����i��9����/eRPQQ�@���!�s�L���n�����2>غ_���s��^ۀ?�;�܏ �eRYڒ��پ]���_�k.��c��w����!�G��b�G�W7��_��{�Gm��~�>}��
<���᮹�H�e�Eh��_��>��C� ���-�ʇ�c����Vt?�Dǥ���Wp���9}���7�n��g����O���Y(-���{;���w���W�������1�Ιx�?BYC���9��2�x�Kl{�7�j�&	�ɼ���z<��w0�޹И%�3��/����t��a����/�9KWa��G��V����y���.^���P�����FM
�[+�H|�\>�®��6mBd�5�g��6a�����\Z�
MG�d�aX��'�s.he��&�^�]&�d@�|��h�,1W���@�������ûm��Y��C�f �;&c����>[׹�kx��%Z|�|O7��+�d�#�{��@M���ȵ+BXR�D(a*�=����1CQ��+������5�Z<���sh��S�Ri��C��b�24�9Z�hi����/�Hu�~�(�͚����'�Os��$e?�3�V�ւ�^�Ԡw��L*�˗.��F�d��q���#F�y�8Ĵ B}i�?�)B�8b�QhMu~�<��S{T$�@_��ي�GJNB���y�ldK��("u%�-��$C E���"�����Vt*��Fo�\<sn:���R)����cזMh?}����p=�~�����,E��8��v	(�u�@�F
����D-�Nq�iæ
����l?�h���J&��` �����1t�m��e�GJ�j�B��$�ѱ���z��i�~�&-,BVaN8M�IKz?����	\�p_|ym7�zjJ˫PZR�Xi9J*��6���:_��v}�5���6Ƅ��������d�~�^�iR�p͒~�5LM��5�@R6�FC
�=�Z��T!ar���*Ndx�j������$_
 �J���|ٚlK�+��t$k)���P����H��0��UX��K(3Z�/�ݬ���bM�K|�Y_�(N�Ih�H�e��7C�Ϲ���ΝC<ǰa͢�`�M�M�W���	||�b(��P{���7��A��AIЅ�d�F���˙DǏ��EK�4�}����N����؜��q>�[B1%ŧ�Lz����g��7��d�-)RM���D8������9�x-z�h������,��a/*�9f���)���a(���$���Vi��!ca3ݼ�������J�S��E�;�`\�9N*�S�YRT�oiF�fB�*��G������N<<DI�Ύ"Hb��4EGl�8�c7� n8���UZNB�
��G�NK,_�1K����ĦL���ȅ.p�E�!�N"���1���P)��d
���
::zПȊ��"-)&]>�A�D�PFv�$y蟠�f41�P�G>'-�P�7-rjC*N���4���5���F�B��,*�(\�5W�7���#1e�|�M��tG'��ｻ篷!ZQ���t	0%��!,,ڹ��);�Uɏ�\�|(��W|fqz�'
���d7H'D�\�\z�V���ffcN�$	|"����Oa0�Ҡ��Y�z14�8�RWo�ϢF�+
��=.t��%�|e���ٖڄKJ����.L]��|Cf̄
B�(������[\=scGO@W�:���?�=K�)P w�"s�E܇>ز�m7t�g������g�G��H�f��+ٍOw���[7���I������y�$|���u�o�M-�Fk�8��:���@��ANڢ�h���/�]����xؠ��K����������D�a���a��u����s=x��2��*ߣ�x���s?�O�5Z�>S�>�:��o���kWQ_Q��^�]>�4�~X�Ǚ��\\;}����F���<a<�����] �������l��W��op����5}� ��7l�s��X��zTQc��1Ћ=������f6�hEz���<����0d�8����A�}8�lx�\:{R���ic�mS��� S�G&!�^�_u\��o����Aį� .~�y�x%5uphKH�u�U�ݶo��s4V�H���X��a<����#U��@N�6����;w�2�E%D�rYqq�s�Dh*+A��"l������N��K�t4=�?K���n�2:&ǖ�U:�B��f��!R�N3X��#����+`�;A���|%c�T ��;~���+��=(��`��1f��k�t,�(�8y	�Y�LW�>-�.@.�4�g�H$���x����8�u��}b苋S;�Vu-�=��	����Å�7���mH�u�_Ftx��V^C6�A.K_|#�l&/k����7����$6�ׇ��.�@	���3��A: �٭?�r:���y�\���J*�x���8��8�����t!���y�|^� 4�Z�����&܆1&�r-vu��������df��Uػ'�|!vѼvx^�{���َ@.���m�|M�'c�Oc⢥���1�߼���h�eeӂ�S(^�P�Ɠ��(hP�@�Й�)u����L��1u�R�\���&�1q@���>�J1��j��X��i�ɂ�� 'Y�BBu����"�I"�N���%?�%��]6l"�r�%��V�%R^�������ډ��}��~#|�Ku)P�H'w�)+u�G�L6��F0����:��bm7�q���"5M��xE{�F&E������A=#���P[�@DM�		h���u���X�s}�cF�I�Ŕp�5Lh0�����,Z��6��T���P<��u-A�
ҫO�>-9KcǍF]]���1G�<�����XxG��������w� �ij
��ߵК���d"�F`ⲕ_�{�wcw�8��䓓�����|vN>���B.+����bQ���E\�;�E���줫�u�Yp��T3�ų�táҝ��?i��+~���<��Myf�ID���>���l�xd7[!Wv�U����I2�w��E,�:��0��x�"�s�W^F��J@�����?-�+��x+��J����b�,�j�����(pS�e`�������P9`'<)�P��^���*PYU��2`�9�X�Ӟ����(�I%%�&(�ǫDG�tw��F[�_kG{{7�2Ș�v�H��IO�&S�
�I�$��~ٰ5+���QH�(da�
�Y|F�����ð|�2̞9}.����q����������0�6Ć��ox3P_����x�m݌s--��4"��2MYq!���]X����J�)���P6�^��#^�l0j����7�P�vqC!���E���#��I,09.ggW
(�&��X�ؕ)v��t5���W�*L>��]iQ�X�,�R$e�mv��pq ��ۧb��G0k�jh��RD��.t^:�Ϳ�9�7:��4�����+�5�ăO?-OfZ�&ۮ`߻���7�v�2t�/�Bʮ}�YL�w?�����L/>۽�6��Ζ�ʒ4g��i�|�q缅�ǤhB6����[?��Yp����K�(�M���W ZY)Ӷ\*����8���<x@:д���.V?���g�c��)t�����B{�9�L��R(�����~Sg�E��^6��@������V4�T#�ͣ+���U�=���aʒ�������_��W.c��)R^��A��Qx�?Dݰ������I��˟J��m�F#�>Ĳ���'���q��_}��xk�m߂��o�i/�Ri�7���ǌ����Rx���N��� ���Ο:.�%_u�Fᱧ��ܥ+�/)S�LV��߼Ǐ�Oܕz��¼�k���4f�ڟ��h� ��7��X�I:,���E�����2��ZV| �_�)��ٜ�sR�e3�B��(5D,6
<����������L��X%�z��_�n^d	P�)��gi`�-�X��@h{Bc��f��P";iF-[� �9�輁��3|�s�x��PU	�MȆ��ؖt}�?���2MI�K��(�8��'��aM��JKJ	D$�� �2qlT�:�:���M�`�w����+e�Dw�����֛Ht�I��HH��R�r�tK����V81�~"]R6�<[W:����H'�B=È%��>��r#�)�:��(?
���4&�vVQ�?�[������{�򉸜鼅g�ax�,�Ԅ�a�������Pz���6r<���	|�w��؉�˗��A
��O,u�(��r�q1v�����1j�y����B�����%4�����s�頷n$��`�*�;	 ݅$�4���J&�ǝ+V���Kk	�!�.��Eƴ���6�@��
Lz�׭/�I�ضc=":�ט�\:#�z�*������a��@��FJ�D����!���G�@���7l��-1:�`h��,dE3�u��Y�Vl�
M���(����D5�U����mP��/ԁj�W�g�娚m�����B9�:M�N4t�h
R>�2)|�ۉ��SV,ƌ�+Q:b8�p	4]�X_)�d�}B�{��[Ғ��a���=U�ɮ�ee��&�q�={V(WcƌBcc������@���B2� ���m=�8x�>A4ы��N��f��]�j�3c����i��S���������7�?<���?�l�;�7�0�����T������iE��ٛ���9U��JN�Q79餯0�ѳ�sLA�tù�:U'�B�°k/�\�!���������{���<yi��Iq�Q���`��'�/>FE႕�fG�Mf�Ȩ�WRp=�@ѻ^DS��Wba�O;�`0�H4z��_�ͪ�e�(�Y�����g8Jj@�ɘ���O�$�#�<���C(+�?~����[]W��!�������:=��c��i$�":����p35V��K_o�]}ho�BG{�P�K�R�DY�y���>�΄N5���!�a15��"��,��=�rⲡgM���C���%���sO��Ip��;_~>?��Q���W`��Y�M��t�)	�;с߾�w��-.�;�X$���a9��6$E�U;����s$�� �/��V�T�^芠l�/�)����Mm���'f��AP ʞUD���h ���*����2i�t5Y�P��\e.vz��򫆗LC��S��&Zݏ^ݏBeF�3�_���f�*7�!T�������
����=w̞���?�n$Ð�IΣ@������7���c��̱�f�x,zh�<�$��`f�0�N��7����O
p��s��b��I�^K^�n#���/>Ş7_E_�u��W�z��C��h�.[��Q�dZI:Mߍk8��a\��\��l�#�b���Bݩ�mDOW���������w��G(�Gb -�Ekפ��#$1���_|����F˙Ө*)�����~̘�H��F�����$��dvlx��øQ#��˫��K?��f"ZV.]�g�g�|yp?(�%���ի�5oV?�&M����*��w���ύ�ɮm�|�P@�wISf���5�a�P���H�u��{����x�\�����X�|5�Z��a���H�����Y��N|q��>yl�X	��;�<�ѷ�.�$3�F��+x�F'���yCkԩ�܃�>��1ca�C2+���77����0�zQϜ�|N˃�вLTE�h(���������+6rA%�%�L,E홇�y5x�bq�a3E�^�N>������J 6HbE�ܷ�	�4C5e|A7]�~~�	�1|��FM�IF��Ul��˸p�3O�����f��Б��$.�T	��6f�[?�l������<D��k�3ѹ1�V�9Bj��t1������C_oz]#��{���!��k`vv��_�
��R7����i��u�㸦�&6�����'f�+I��/�z�G~������ˎ66�GQ:�y帙EŸ�X��1�}�b�������8�������8�N� �	Ť5��l���]wLŤ�&Jӆ�z�-�ow��W���4ၜ����=yW/� kZ��α�4�|2�(�=lW��'͜�e�>�!ӧ�]{pm�.�ϜE��E��mTDƲ&�#g�l���<�H]��>j�|B:Z
Y�M��x S�/���Q��\e-˙`Z��R�����1m�u�4����h��H����xg�Ȧ�R\�ڊ��c��)V�l)�C1���D���t�:�l��8�e;.nٌ1>�1!���� �XS�f�Z�T(�x�����c�t+źH�.Z�:���
,22�)�%�z�d��	k,���j��}�o\�8�݆��!�`��P:|ɞ�Tt�kK6������|�o��|��`�y�u�ڗ4&~/M+ث����hnn�WM��cqH"3 >��\:r�%�օܱH���NT��=2$ź%މkZ��C)4>6dƌ�SV�{�����A��[��>�ͥd�r�L�L�ޒTW�nt��VYN%tN��&�B�V�RDqSvI�����TH�K��c� '.wtM<D�:w2�U ��_L���Q    IDAT`,�����_��
��̈́��˟�B-����E�l\��T�T!��/_�c�@�g��:���*���혎eY������0�)P���ܕk;���YvRn.�23ٔ�M��l���n6�I��-,��c�2�՜*0:$���(B�(�+�PY]���r���A*�
�ɋ�@Bl�
���T�Œs<�D_� z{���3��dZ�Z�2������l$� �!�I-��b�EF��#��Uԣ��H���W�t#P�!�����IE�a�K^�hC	Z�G�z7�^��a�c�㏡t�$��&S𕗢dD=�l��x����<~1���1)�~�@��	
�(�.(K;z���`A��}U�+ �V���a�e�Ѹ)�W���*�r�z��(�=ڳ	(���s���X�3\О�@n��G�]y�.���;���s�旲5�be���n�tܵr%&�{b�p�q�_��s?�����KW�b�\�c�L���>�1�����F(m��p�sl|���0�<�2�+�0{�r,}�;��� �kgO���W���[He�	̸�Y�B�Ɂ�3э���8�}}��tV&N������5�y�h	d��C��-������ųr=� �G����p�Ũ�m@6�B6ދ����h�V\o�(I�|���r��p����l�H,�x�5�;q?x�>�'t�k�ǽ��cɃ��n�ph��gp��Q|�m#�߲A #��HJ�G��.VQ��x?z;������w�;h�t^u�5s���{c'MEU]����lé#�a�;p��	9�Kk��<�v�5g�����J�M�Ǳk+�>$�h~T76c��:��4�>ݗD������G;w���p����t���h6R(��ۯ�(��?��;��+k�p��%��r%���2�}&o�����Ʒ�s�����2<�4���e"�P��"��I�v���u~8��[Hϸ��D�#�^9�H���$���*�Qu^H,��l��JS�e�m/u�dYă~�D����ƣy�"��Ɗ�Ȟ�G�������^9F��������4��p�����t�rࣣQ(��Ő7�a"#e��N�����	�N�C�4T	s�ӓ@t�P����p��y�fy ���?����p���QH��*F�=��A5R1TVT#���Z[���Ҳr��8�DKKĩ��*'�|nW�\�� �iᘸ�D�l8��o3qh��=�ƫ�{�����F��s�r
h�p��e�l�ca�F"(�Q�t{�@_G�����
&���hO� �~�4��k���ut�Ǒabm(���jIqEK�PX@��iw�h$��pi�&8ߜ@�S@�(�����[����S_)p��
�t�r�E|HD�8��od3�yp-�\���&؜�~�<�Leb�$ġ�է�u�믄�B1�y��|D�1��8ۥ��T��z_}��h^&L���Z	���i� P8�~������Ppa�F�@#K}��+^O�.zq"]<]������"O��<�=�~�+�ͳ�&mhlx���[b��A���T&o�!�d�h(��6`�\̦p��}� ��\�kV":�Yr`hgL�ED����N~��C�؂$s�"U���\��\�jz�.�{Y�v���\[[���:��e��a��*��A8ynOZ�uh�/"w���m�*!�CMI�$:p�M�7�	c->�0���Z{�w����򯪀�m㲅���Tba���m��q��U0��hT���R��ܠ����B�7��~W: L���I�Tɪ�#�6g(��}��.#Z]
t�Q�۱�5����z�P�j��뺖a��KN|�( ��dD,~�C����5[�=����������4�wK9�D9J^ �a2u�v\Q���_бG��{�u56���0�5E~��EvZs�y�a�/���a�����9�C�ڎ��m3c[�U�k���S�8�|��8i����u3C���Og�c���?M�rĊ����W���%�eӖKY�r�Ne�M��P���~q�A�O��Lо4-�3Y����y�KAD�*t�`��%~��D����1QP�D;�CG`䐡0�9�8w�V2��4��-E��IX��S��d.�f�z�o؎|o������F��38}���7aʢ���4�Ħ�	�:��ׇv��jc�ׁ�]jO�6��l��Ѣ{��٫<P���B���:�j��v5�T5�HR���{�#L�GJ�(\&�b����#	��M�[ֆƥ�E�Z
.yu_�NF4���E�O>�������`ܜ��xF�s��1y�kN
��v�*Ο:��a��X��#B��`�#03�8so��g8��G(�m���gއ�W��Ļ�AI]%�d�\���5����H���`�1n�L,X�n��>�**DSDَ��l�f��q#�{�ak!ԍ/�h3��GI}�t��L�O|���l�/���9	&͸C�M�?z��N��u;7��o��B2;��4��e=)��He%�_@.���W��mx���@�J�]s�ǒ���l�Ǵ�LG+���[�޼�DF(��ᣰ�ѧ0c�|D*�a0_�v�M(x��p��+jj���'���Q���[��tmNcϖ���'��1�q�p̚�sW�Ay]�7���|fw;vmy�?�}�=B1�2}�X�Q&�(-Ssy�6�~�!�q�v�*�+0d�h,_��ϺZ0���u����o��_�?�mMGM��~��X�B�˸���FA�_c�o~�+G>Gsi	J9ecB,��@�[(�Q�"b�%��F�}�`�W�5%#(W9",�>�و�I�IoqRP����gƤy�����&�:�sT	�w�AgLØ�ˀ!�d��{�Ǿ���.h�=�MMr3ح�ފ7�E����ۋ��.�|A���TU�#��"�]J�A"��"���<Z"�iv�������EcZ��ҊPUFΚ����ġ%D�g_z�]�@W;����O�P�	�\&��i�)k�Ҳ
�_i�.�r�9A�$���B��ј �!-�-r�9�\gbw8@C?|ѐ�	��B���ؑe�� � ��~h����|]]]�c0�"ѐ�N��'���4�.���H��/Q��ACY)��0�%���F�x��7�>D+���Ջ�1>�0*++ـ�<�kV�>�ѨPېL�>Ƶ�[��;�z�8�����Ҭ��s�)EQ��-����&��<��]�I��m�����̥���\�'.l�*��t����f�� f ��,L�XB5�rr�3��'�[��[�[�⫯��suʔ;PW�$��@ ����J�����"r�g����o��Jatd��)ᖷ�w�u�i� k�+d�]�VpPl�
+��N��.���<65���HB9n�O��E{)���`y�zPM4�����O!W]�ۗ/¤��`��BD�D	�z�O���DH��e:A*��RX�(�v�W�us�6Ud��r�POPYUG�v�me��l΀;e�@�ū0.^A���к��,�"֐3hMw�l���!9ቦ�w�Pu�C����p���59s��v�04of'X�5�2Cr�\���`����i��Cڵ��-�a�Ͳ���ڴ�%֕��:���MՉ��Y�����Y���L�>�#]׵5C35��k��w5�rm�pH�!����4*�r>�(���%���f�r���d}����Q�tW�&HYD��]��;K���w�s�1��ŸLIv��8�c�8�nS?˹.����<�����]�|v�P�-e��3|����{���Ŷm[�_�p#p|9���|X7{{}�ĉM/ج��jWO����g ��@HQ{�<:W�

Y$ҽ��2��K��|� ����E=detFNi��Dt)�.��
���Cg#eĭ�G����*�vȤFN�K$�䉷���$����/�s�4|�BY�G��*1n�X��oc�ih��5���Oqf�G�����/`��e@uG�'���ax3�>�J���~u[~�S9��וTT!��IC��\,�<��rIP�#r�2"�S�}/��$�0��sK"�`QN�+�Ϳ)�sq��<@�]���]���=gpM1�E%�,3���b��w�ʍ�YEP`"ak��uq�ڇq�c�1b�hU0uj9�~�|y�^}'�>) i������� �n��%�$d�9�/�Ư�w�p�.�$��c�cOで�A��-'XY��װ{��سm�=��}%�5���P3a���&�zn���;6l@W{'\=����Ī�Oc�]wA�rcv�C�a��r�+�y�|�񇈆#�ڌ��>�i�̓���Ca�fRp:���_�ȁ����%@3��ê��JʕϷ ���Á����-p�$�Y̸�~�z�qT�c�yȞ�]����?�����#��n���� ��0��<�_�2����Wp��Qqiڌg_�f�_
]��<G�|�W.��m���������	W�����sZ+�9��vnyG�G4#��/ŒU!�<L�����d��g��&��?�h4�q�o��G�@=�θ����H``�����?��$k#��PUS�������^8
h���}�-\��++���׍����9�����_>-���kyźF�~X��ޯ8�����k����Du�x��|��[/��hQ,d�錢��ػ=ս�0?/��.a"@�}�1m�C�>$]d��n�V
V.)nR����&����`!�l�7 	x�
�I���%���mJ��1?D��D�
7:3�P� 5��XD�s/@����*�L�[O8	�4�Ё(u���Ȃ�N+'N����aM~/�=�|N:�vN�0S��,����@��`�̳ڤ��o~�_<��}Y��J'1ޘ����`|<��ݏ�]�ڱ�[�UU �%��}"Jo�ژ�@�L����P-�r�!�+u<͘�� ������:wu��Ұ܂p�Y��R�V>H24�k.����^$�2�A��
f�^����P�H��#����E�?�#!4D�L�Ž��`8"t\��І��-ûH�9)��Z�U|���r6O�:��B��K�16a��!C��-����[o�2ه�%:�Z���N��]��(�}�9�בEc�bé �}���)��⟀Y���B5��Z<甭6uw�z��ZD��띅��*��l:=
H��h>��j8��A\6S���i�ҊT� ��hL��������i�FQU])��@�_ ��$:`�&����{���QW߄l�4t
���/'6D4g�<w��H~���-�����g�q.�m�����Ԑ;f~���G>���������x�.c���é����e�c��r�68c�޻�������q�	�b	��_�|6QoB�n��x�FL�C��b|Ua��M˲���:�����r9�G���Ly;����{}9�}�xw�ْ��/{�d�y�	>'�ss���� 2 &0�Y�DQ�
I{l�k�z�;[��vj������q�ǡdK�%&YI1�	�$"���7�s�=�ޭ���i�4�cUe�;U�*�7�{��{��}���9?;�'�n7)�7��F�}��xMԚ�+�C��S�	
�a]vݤ% ��I5y�L�o�]AG�J
��S8ԝ���݆��[1�޹7�	M��Co`�Ի����Fǆ��|���[���=�q������`��y�z|��/a���x5���Kx��X�q���"ٛ@��W���|�}z��x\�c��*Y%*��q���\ �m8��9� U�HF�h}<,:U��
(�|@�%pNQ�TԀ�,�{���Jԥx����R�R�~�b�&Ϡ��j��G`�$�KhK�*p]`��c�7q�'ƭ�|���A+�B���Z��E\z��������A����W�������с]d�E��i|���S���gP�+#��ǧ��u��ȗ1�i�r踀�r�4���w���?W�]w˝����2�B�Gr���Uh�=�^|�I�fct�ո�3�`̖)$�1��#�����p��W��d���Pp�����.�ۚ롵p	?������^�����ܲ��7�D:�z��;;��/=��_x�JU4<�o���� �v�9b
ozL\����&�z���T� ���Wpǃ�"o�0]�'�8�'��-�>�ڞ�l_����Î�!��'�d�8��<w�<�}=N���#�������;��l,~������E'@�}�ܴ���I�׮U�T.�#t4����[q��7P��qe���66qb����QG�V����O�.4	R�n��.�e�C�"�YQ�f�q��q���ΟG��#�~�Ow� ��к��	��ˌ�:Y�%%LDL ��(��J�U{͕n$;�a1-��Aʸ��X�����h@_�g�S�#ퟙyOc��e�疛���/ ǜټ�q�.��(��,"=j�b���&��U�s^w��߈�~���Pf��O�	V||q�3�v�h��bb�(�
��~������1��`���*� y�_�* �چ�v�[$�Fj,�ٽ'@PJm�V�)�>�R���C�.��H�6S̞�R��9P�{>�s���N�bY�P�����;qZ�]�?�Ժ��y�v�d�� ̊)�*�����0|K2"�g���m�T^~sO�޹�љ]�@��G-]6�Ϲྣ ۵t���N��c����E1�n��r ��7>�R����&��D$%N���1D�51q����d����H
1s8��ԇM7N���$���x��wE��}���P!%��N�⤊i�e���".��2N��Q$g���к\���Iܕ逪��v9p�u�s�&���x7��5ݒ����[���R}����\����5�!�!�����T���*�8v=x/v}�>���k���j�Ɔ�$N�xm�|�m�.�L������\F(֜̔�E�}�($(��� �~����ձd�@�m�WZ4,"zin�g/�x�m��+�HFۈFu�Z��.rR�f��urx��o��y��G]E�������+Н�I�������ȡ�ߨ�+1&�xN,����"�D����n��@� ��g�P�%��\1BU3�B�D����/% ��&ᤀN\����~-n��f���;�
&O�#��rZ�Z*��;yw��W�b�6\�xO��{h�]Ɩ�����0V����G���b��v�p������8�ԓ8�؏0~�q$]�  '��^��MHU�&%�3
�Y�� UEI���4dD�N�X '!���H<R�SWĖ.7�ժI�L±�Iz�V�FVɫԁ��S�YA���q����r@�\�±���@!��އ��G����шZ�$��k�����x�ﾃ����1�a�տ�C\}�m ?&|�N	��'��q���V[���G����؏��[�dTOM\~������'%�Fۮ���G�����笎EF���ܤ|�G^{���[��U[�i�7vD �S�ԫ8s� ^z�1��֛�����/��?���9h�K��������ơ�_@�0�D"���6㓏<�TO�̼M����8>|�(N}W�o�v����y��^�	u�8�� چC����sgD\X�;���������"�H�#C:��_{����a��)�n{]|�s����P�[�1U�f�ܣ���_{ED��d[��k7mG�P&xR{�\��g��h��x��V�bÖ�Z�
U�z�h�B���a��U�Ji����6c��m�(��7u\<}n� �jU��]��u����IӐ�&P����#����F��@�\��Ut���r��Q��d����F�U�-�����Ut<��s�N�v���IgO�̉��U;�\˒&�K.�1�b	,	
��,�д�hĄ�4��;��;��뙥��pz��o((8;@�
��ɠ�A��
4���4�=٠K�L�¢LLH�bԆݓ�X���:j�H��=#�    IDAT1��#�N,-��7���/
����x&�D��R��5�����h��H�t�0_��t2#z#��ua7�US�J�${]4n����TzԆ[��V�Ac~B��kX,FЩ=�^I�C�`�"��f��h2&`����C-_�|�w���Ь���/�5��D�����`7�6�COD�&-_�~>�24����ǔ�fcI�6*�~D²�aF'	�����f�z��Rz-����Bc��k�l�(6�!�����23�*�[�L
.up�zq�}�ᶇ?���(-�Q(���c1Q�$�,�;����SǏabrL>�\>�d:����Z���*��R'�T���Kx���e]lڸM�˨S�Y�/���
@�0�klӯ��3?z���JBc�3R_�3�l�-p������3��!e(��z�&���9T�P�3�`I�#ؐ�i��*�='���NX�/�u�+���P�F����q��w!�b���i���pH�v=ɧJe3H�S�GP�bJҕ��]����L
�T�ZY�H���y�����]�~� ��ρSK�A�z>:]3mdę��+
z�*2	 ���l,�Bs��a���γ#���vv��/�r��?�o
���G���ų����?����٧���� ;�[� %@ڿ�t�LmC�����#�k_�6s�����#_�i(���r%V�M8���1�zj����{ב��\������k&v�ތ]�� ����c�x�]��ؾ���ut���q�>��7�����Y���I$ҽ2¾|��:�.:v��ߏ�{��E���o�>���<Ⓔ�	ؑ�#-H�5b�1����p;�� �z[��$����
ܤ"t��"&��*yԴ(�_6EkJ�Ɵ���P�+t��͏%�ڔ�_�ЋLCr��$Y�~��E�3k�+�@u��ѡ&���z�f�������9�l�w��ob�7!�j^̂�q��rǟ�G��?|��w/50�~��;��M7�S��$���8��+x��'p��S��$���v���ې�| �^L�i`����~���Ʋ��;��o�>��L�u
�X,x�����O�0;�J�!���|���x���ct]+E�|����8w�X暹<n��A�5W�>�x�&&.H�ܹ���*�9�/\Ǝ���Ԡe�]��lfn�RE24芢����XR,�qajp�*���Q${m ���ƫ����8�V�<�u\|�y<�L��3�gb��.���}�Èo�F֮t@+�����|�Q���K�'��n�b���4jK7��Q�]9��
w�>�r�DHS�
��I�B��mx.��Tg�����C;&�|��j���1�X�u.�xrH碫x}fp�r��h����c2�<H��!y��M���,M�~~kS
Y���,��6����Î�+�B"�vI	1Ѝ&�@��Ж����R�Jw�fG�An�wh"��>����y�F���{Љ��e�X�rT��4R�m')��r�ZS(����5kW	�"b�&�q�01)��D�������^:syF8�����������z�j$�I,��T�*M�0�(��T&���j�W�U��ɉ�ü�:���}}�
� �B��H�F���^��6���{�P(�8�(��x�Q��7�|>��!�Xx�Z��#NLUϑF��r�.�� ��)�m��#��H2��RGka�5e�e'�c��2�q4�&��������@�ZY�x�k5$4`�w #�}��q�F��F�u�1�20	�%;�aT���E;ZMM�|����a�]Ǹ�A[���W�v�X,7[��؇�ҕN���qr|cc�:uH���8����$��`t�j�8(0ۂ M�-�2�&/���q*X�f2�^�VLD�r~�~�0PG��c���ԓ��2��r���}q�&����U�_1�P��˞*��6� �:��}��MjFd?�v"`H�Y`��� }��݁����c�9Pyh8U��W�t
���ݸ���d��A_�
Ĭ.OϠب ۛ����sܠ��d��[@�����s�u?;;-k�?_X\��hhh����|�.Q���Vq�`؛��Ff���W^C��!���Mј.�Y�ʳ���A[5�w�s�w�5��w�#?��ȏA�G�	�3<?'������/���JՍsAœ}Hd�R@�^��9��4�6Z�ȉ�*�t,�Y0�.�*K?r���$%dRR!(ࡼ���P
J����Xfw iDpU~k���X��Dq���2̖3�,�ݶ����w�p�u�;N�.�h�w>��J���cϝ��Cp/�����[���O�Lc��a��E5ӹ�C_�,�xn�W�<,��(��Դ�<H�i<N!�d���q�L���S�eA��t�YlrM�3^g��������l�R��:�^��Jp �]_�K�p�Ն*�yNvd��z�p����YX�]���_A�- ;�	��9�u��;�7�|
?{�	���;&��+����]l�����3vЙ:��^�������ʊO�q���q�]w�g�E�E��q��[x��Ob��9�L�/N?�������\���Ó��6�O�F�\�N�����q�> �B��PXı���S���ً��|;��7��C_�X��ZՅ����ԅ�(L\B�[��cG���~�t*
�ӂ�t�zGc)��l��"ҎR�h�h��˝�C��V�W��x�-_�a������?�h:��@��ӯ��W^A�� ��Ԫc�5���{>����%��׻U)`��8��8y�mI���&`3����?u��t�IIV ���L���K�QNg��]	k�tq�Q~�F�j��vD݋Rd�QrJ8��G�df����L�E���q��e&��$W�QM!U�!nwAN�����I���y��.:p�!5�t&k،(����7<�Ǫ�g�(��X�%���`�]î��i�=�N;� ��pm��Cn���nv�2 �/�tZ蓡3;�RxK��)q�2#��)ְb���� �����bvxy�(H��q�w�!��B��d�TJ K���uW	�ii�����Jk^��6������A�Y�G�[����sOgAd�;}64ē1�����L~�zS�&{�8V�`���p�Y��5� ����(���P)a|~3�"j�2:�u	��p���,z�(t�3�
���75<E�[^ߴ����.
z�=��MD�z,#=y���
�wꎋ��S��A6�$���VN���f7�N[\��6�>�:5�1fs�j��>l�q?"�>��R�?$� :51�S'Naav۶mU �`ș���FU(B���mܸ���h�S֘}���>�!�����d:ä�Ӱ$Z�~qhȸLxcO=���"�d#��Mix�+��+Q-AAh���{a�l�(�\�! �z����C�2�h�L=�ʢ���ދ�'t������c����Qy��	������"��-���=��K� >�?�J����/�����C:���c�J/�Kx������Ѿ<ߛAԎ�^W��bi�ss��BPPn)�3�<���h���ٮ��z��s�-D��w*BkGl�U�p�9m�k���ݶ��n���J�_�!?����o㗻g�ڿ����x��g�Xt2��f����B+zHWw�FīY�����E�!�8�� ���&�bW: �"((Q)�;���Gry�"�'��*Ш
(�J8]F<���jl��f\s�>��jL�~�N����0yi��c���q����}�-{�i���u%-6�n���A�?�7��ZJ	P~"IU�$2-�8��b�(�n�J_ �F�@ɡ��n�����A��8�H�%9�A�#�`
�N��b�' |�ٗ�<�y�qs�"�W*5[�w�3X�&]���v�oڏm�o�5�/nC�$`��_�b��I��G����j�'5 ��ͷ߅����PܶX����E���A���Q����=>n�y/��xV�_�����楳���ۇ03>&��}�t>��{�b���HPL(.*e�ON��Wߔi�Xڶ}I�ܱ�ZlڼM���8�vŗ�Ļ��o���"��x��^�[�@��b}}�sIt��v1v'�m������?�4&ZӹDH֑�؞�N��:�.��&�2y���DQN4�G��K���^o�G�@o?v�ދ|��mI���	g�;�K�.�1Ql%uvdx�7nƺ��ă���5P.�b~��.O�ZsE��Y���-����[�u:�X�'���c���}�7H$�@����B+���T�#�-y$��%r@�q��F���>� _�E�y�;b!i���4��B9x���u)�"7�ޠ��XXk��z��R��	�64��Y"�n�nWhS����J4�hۂ��ިק�Z��!����Ck�m�2Q�4B���}�����N�eʡ��_�$���RĶL�'�TSn�t�;� C
)�S]R���%�$ � O6$�$�}L�ϐ�5i��h�	EH4�3�xRD�3���A
T
�i�-Z��po0u�4�`!Y+�r��%�yt� �(�s�RN}�X4��Y�5E����qfv
s����T���)�Re�Ne�4m���V��E�k�A*O��r��
�����M�.���\��`2-����0�[g>�t���M/M�er���k-�"(Q�4����a��Ɯ�Ƹ_��V�U#���Oa���I&��1D�j1�Y��D���S����u�e�&$bI���W��	2��H ]k�ƫ`�1��M����<�{�]t�&֮]+���b�A��]�ڈ���z]̾~��)�J���Uɾ�޵�%��L�n*:Djn�P�_!���Q��A�W@����z�L%>Υ�f��T]L ��
�H��ߗ�R�Wl�9-�ML5���0������_E�-��zsUԚr�=�Ԍ�CӅA�5|,�?��*��X7���ό��:�91`�8�:�aFBW#�&(	�u�w�H��%�C�}�m؋���e؜�&kE�9s�����n��ݱ돇�}���cP��F��K��?��/����|��_\h���ydrQX�`��O�
+��whOƪ6�(j�1%<�lW�/�-TVh0):��(������Y@���Ho	��>�	�Y�5X�&��z-DPE����}56�܄l.���4�gΡ01�f���ebh�v�ذ��/��#Y�F�PE�fll֠En�h/�U+@#��+ʍj�X4�:Y�
���!�J��V�t�|tu�Y�p4R��^G�~옵�(چ��m=�LF�^�@����m�b,^c�Q��o˕��8k�]�!�I�K^s���e��4(�I윱k�l��
1bKX^2ߏ�ʕ��Mh�8������uL_Ǉ��z������"�͢`}}C��� 0�-g����&.c�R��
#5�a�
�e����F�t�bq�3��껤 rx����F�QԲ�M4�T�(�"��3�"���z�Y���"�+���/���l��@͈"7�Ck7b��X�i#�+'��t�]��]�����p���9��X�Ѳ���\�'��Q�AP�"�]gz��5�>�� A��*h��ˈWw��b\���)�fJ�p�]�-,�Ѩ�A�VB�mb�`)��H� L͒���g
oI͙�8&";�]�P�#�Ն8�Ph��K-���ur^�L��徼�j �� �0�*j�q^�ЗW:"�d����Q�g� F�<`ف�#w�s���E�i&��V	�O�� �^ڒ�5WzT�I8P �C��H��t"1�h���MG�l�u�142��h
Q�n$5LOO���s��t	���R:)F�VՇ���n��չk�x�^�ʻ�_�/���
F�E�5&M���=�I�N+�B�PXG�p�ʄ pK
�T��rb�U�E]�����T�ɢL2����Q�9��0I5* ~��B0�}�I���E��z�N��4�`�v�q]&���9�|���-����o 	z��ޙ���w[ܢ�>ĉ�eb�^���i\,Wю)�R~μ�Z�jq��nh;.tq��NH�x�Y�É����rQo6%y>�i���5��I����'S�Y̥��d�:��Y��BE�#"��4�ҁ�ns]��2.���Q���p�'��;��9Z(��,9:&.]ę3��,X5��dv	�� TUlL2���6���X�j���G�Fl ���L�	
H�>D3 ^�pR �w��������p�G?�=u�6sB��h��q=��<,�9)P��M?vC���:<�������<���b�>4��ʞ#�@�)��@{@��u�Ƌ20�&�?Ǉ�S8�.cx����_A~�p]��U8�_��W�U���˽!t�p�e�g�'T9RZ��F�.�N�VE�R�5H�5N)�jsr���m_��1�{�����{���s����y���F	c�"�C=Xy�3=ۮ���}_�ΒC�/]�����Ǡ���:���Q�����m?����l���ͥ*"�X��a$�Ym����P�2Qa=!��+�X!_���h�tV��!!A
�l<̵�$�0�uT�8�*����E��-�b&�,6�.��#�6:-K}�+���y�u\��$�+z0�v�T#}y$m�XM��\����)�<���d�U��@:���%�82���S�U�Q�}��",�$PHu'���f���6;^�t<�6����n ��X�fK�'��i����D��T�$r==��l���b|bL,��,�ɔ��cV����Sc�f�3tD4z���:qE�t�o��c�3��z���g)�B6b#a��lHaU3��������P+403W��B	N$�*_CO�C�J �-�]=���n����@�y^E#H�z���FOۗ���{���U���X(�A];u��L�Di/|�f���N�"�a�zզ�6ї�`EO�.�h7)7Qף��ep���F~��ȭY#��H��u����U����h]����?q
��y�y���(^��`�D�j:��J@�3,)�l:p�8�i�A�I�@���n�EJ�` ك�}+�E"p�1,�:"q�cq44Mh'F�V���~�� �H]�c;bʴ�:u�����.��p}WM�:�cRl�S��.2���;�a���7�ݎĤh�?�7P �xw+�N�[X��Ytr/�="�>��)~s,���W]��i`�"��A��;ɧ0.&�B6���,P�s�!�^�H�u�}Mz��^��;1�aRC��Ӫ;@+M�v�P*��1�}�T�\�Q�G�\���	kk&*a���r�#eȓb�k�Yr��>T^�+ֆ��	S�����Ua'�d�.JCF����][�B}?^g�HN�MU��V��0 �P�b�,T*K���̂�"1��fJ�
�2
��j��,x����pҪhsH7~eo/z�	���{mD:;��Ę�p��Q���q~vוIР��v����xҌ �[�J>��v�[�p] 'Ѽ�X�R�o�}n9��cq�3���]�Ф�ud
&z�@�kW&�
�0 E�$eM�T��K�ELp�n�~�3����0W���������f�Α#X�/`d�J�]/ֵ<{I��=�;4�pP��^��y�5;E�ʬ���,��&&/�����W�E*�#S��Iگ-׊V�ܣ�z醏���q���(����1�O)�%�Jn���]����>P���v�_�4W~?�Ίb���
B-_�S�ڑ�g=X��sX�wkNe��˖��l��-�۹�5[��_�X�=�"���(�Jd5���>H`�	��pіL+��͆��)�e�b���� sJ 5�te���k٠
AA����F�Y@2�C7�p�̸\t�CP0��q��4|�W��i�/��>ݵ�g}�_~�<�����O��7'?<���XX1�
�\�t( 'M-nآ�Wat��-��ǅA�'�lAGK��⯣��"�嘕߁[�©���<�-�Dۄ�Tk�`WDi� �Hz�    IDAT���R�B�c�7�t-h��mb"�lٹ	=Y�11�KA���E015�#��c(V�+����LC\4T*�R��|+a�;]��p���S���:0��Vb��B���ށ�p8vA�8t�chuT;&r�Vc���`Ǿ�%�'�a�*�E����c��9�ɤx�3��/WQ���S���so��X���Nq8;_J� �7�	vh�P��1����3y6Cƈ .E�+n%��L�5�%S5Z��!l�w;6޸��R��8�g�$�9��`��I��t-��f�����Η���XJ܂.;�4+��V��"�-��Q�d3@�!��L��;�,G"�Yp�Q��ǐ�M�EGP�☏&���ly�a�{�|V�$Zׇ�0���'�@W��	h�g�`Q=_B}�(�k��F��F7�Z�J�K��4�6E�L"5lF穮�L��LȢ:�Лm�&F��X׻z<�V�0�6�ܺ~o?J������ރ�8H����q��E�2O�z��C��@yAF���h;*E��t�-�J�z��&;�,�Y�v�e�^����"v�Y(��v��u���$9胰0����2���"���*��Q�F,ܤ,�09�<���kF��-U�
�Y�)M���M/�GХ:�\�B#�D���wb��k��e�IQ�W�`,��Q�c'��
X8q�� �g�*0�5q����>F7"N@���$вT1-�\ۗB����I�%�Gx�˄�B3bPa �\~=�G-d�RC� K�aA ZC{V-"IO �����tπ�B�T�*���:��b���r%:�uH�j��pG'8kB봔8�41�La8�C��i��_�s�d�\N�"������4�tce���4�|q�|E��0���Ѧ�$i�_Dk��ζD3�x�L�f�Tv�C�Al����-����
�,���%��@I&�ِr'!(P�0�:]����;&�"�[�����f����e���B�P���N�>�g�!���U� �������"jN�8��<�YNMO���j��0��8��LM�'�ņ�6	�=I}�� ���g�hYC�ZC��`��C�I�g�1%��Q���@��%m�^	
�u/k�`R����ax]x�`�&W2~,�(H���6,.���R
r�s��N��ۊ��ih�l���uQB�kѷ�:��lE2ӏ��)�/���=�%)��UJ�bm�T7ڜl�+�Ҡ��?���IЩ���D_h�l��qD�B`	���L�7����T搎w`F�
f�*�7f��c�m�-�n����߲�5�v�9D_������*�v�×��~�O=������c[㉬L
(�$�Nl���U�+�<X�a���t�X��ev0n���u�$W���E1AA���'Eĭ!�.R);��ցVYD�<Ҫ�TGC_"�xĔ�i�VG��H�h+�o�m����]k0��q���6_Ck�B������#oa�������'aIQ@�CM5�`DL�7;^�a�뉼O���#$y���6;�]�l	�Q�t�h���	2ِZ
4:*��ݷn�@��A'�ǖ}������n`U&a^���b�]Q����©��J�/����E�������/�TT�GC���[`�I@G�Ð�vG(Ci�Bo4��x)v��"����b��p��B�E�ic��F��#�j=��үa۽�=y��'࠭#7�z�JI
%�R@6���y\~�i,�| �3����e���|��.��p;l������Xۓ��XF�=ChE�X�����l���6iY
����moh��J�<z�ߎ�/|�e��G@ڜ���#G0��Q�OC�YBO��x��!���i��2��(N�D��{�T����GZ���:�D̴e�D�$������`ז�mZ`,Ά�~��z�ų0��Db�M�5; Z��g�<��N�D��H�$����������`-�(�ohp�)Ie�ǎ���e�<)F�Ge�Еy\����夏�x$�d[Nը��dؽ��?~���1X��O���Þ�e:&�91<��N!����%�f	P�L��f���C����)J����W#�m;��]��m`z
N� ���vqN�FɡQ�=�@�j ���9��ѷ`,N R,�/�2H�ND5M���|�aG��D�.�N/����+�GAW�P!h\h9���a�Or��nix]%/%�u�B�J�!�ʒ�X@#b�u ���2Q�v���C2ع�D`]r�5�;��G�{���q��)N|	C`��#�Huu�(bl��m�)eEв-�KXl6P�xz[��n�1/��-*@n(w�e�(�/����9Y0�mD���a&;]�m[ )�D���s�������e9���(���B�����^Ӻ���1ծc�����0�s��	��09����q�/. �Hb��-Y�Nҕ�>�� D��_�3ܦүt;�o���]�(�6CI��n��\��L��p҈�e�݈��eHPPib��70�ēHNO`E���
�J��!(X^�/Y����V���o��} ����͑��,KNz��&������Q�@�Zi>tf��j�ĸ�A�4�]���~�����"� D�����sU�z$Bt�]��6�[��\k�[!���K�'
�x�+�ƀe��u$tH�� >S�s������8ґ��teRp�>��H/��~�b~�������i��ԯ�J�/��cP��\�_ٳ�={������_|���
�����9���r ��iKB�
�),<�@�	9�A���s,��E
#υ�jJ��0|W���OO�E�VF��"Zo!cXHg�QmVQl����
7!�}�><��/ �fX�;��NM��t�cőR=�@?h�?���>���?��8E$�'*�9*̓X~r�����pk�r���"�+��d>���<蘱0=�^G��Y�	�-qv���q۰�(�G�v,�ڊ>�i��>ث�ѬϣR�G����&ڷi<MG�g�2���+�f��Z»O� /���Й��;�t���۔M���m�MI�@ڰ��ˤ�S�;9�n�qap�V�\��T+�B�Յ�������}�#�q3��Q��C�����EJ)���)%5���)��B���&�5�d���VS�&��l�G>�ae��(�ó%���M������Y����U��l4��\=ii�51��e�n�P�搽�d?� ���!85���������X|�,���q$Z-)`����Uo;��P��h��#4�Z-!�R�u��KD�K��fp���y�]�!>q[\U�:��yp}f�h��:���~`��@6+���K�^g�8<`҇���tY��kp���3�Ú��o�6E���({.����2DX<
M?(.ELiHG���^ ���?)hi0t��>SĈʡ��e�� 5���9QŝL ����fBt�K���P$+��@[v�Î-;�SG�]p��i�^���"v�M@$	��ξ�����D�����X�+���; ���71��K莟A��D��|
��h(�UW9�nl�+,����Y@0���2 ��fx$Aŏ�S�\P��$��@����gNŦ��nM}J������z�Z�dp�4�°vv�vH�!�)��L~�z1ҟ������l��)���<R"]��֢cW6Ŋt}v��6-�{��B0�{�`&G��b|a��R�EĪ��G� �t���d|�j�S�鈶��v���dtC��M�����$���4aV�p�0�Q�[ B��P�B�_(x}~���ً�&�Q`-|P(bڊ":�V~�6�<|qڲe�X���H�L˴�bW��T3�/�3�s��p�<��E���^5���~1Y���b���8���S56Cx�7�j����?zəqGڈ����� N
�� ��!��}6B�P��âf�^��`��p?�{^>1ǧe�!l��)�a�Z�x��W}ը��T�됽����Z�l~D2���āl�1cH�g�q��Ї��$��C#������r/�)V�6QTs��C�:����w�
�Uh���9���'1��hLP}�Qą�4�����������6lP�/��Ǡ�#��ʧ���?�ď��_|����b"��Í�9,Ak8"S�i�]:�!�8��F������:L:��oE0�h;t�u�F�>l��\O����z��gW�\�XQے��E���Z�H}�v�K���p�=ws�1{�$N��:f��D��!I";<��W�w�V��l�*��>����<���2"��)�v&�ueX���Ι �F]���Q[Fݮ��{�µ{����~���h�2AGD3��C&�"=K�ݙ���n����� �^t�`��1��Ә9q�B6S4#1̒��n#�e>��_úm��zǟ�1^�����t�&��a���AP������ۈvu�cq�G�e�!֬�nF:��S�|���F���:�N���xn���x,�MW�Ʀ]7��F�xX�id�D��f3'���n�o�(�#�J�}�-L=�4�W�Ft������c�S�L�����S�~
���Ek��bi��NUk�\��!���Y���cVE��Tǐ��k����6�AϮ��6mB'�A;���� �(P��u�2��̟>,.B[,�����7Ql�D\i7Qk{p)���rh�Ɠ�WY�
%��d
�xm����w4�#�6��H�
�����,4�y]w���(h6*0p�P�k��ꭈ���[���N��hbݖMX1��􎼅�㏢u��ꢲ�E
ŗ�+׏`AFۼ7X��� y��a�(!�K��]5-T�d�}eE�/�b��$H�^�i��6�%��Ba	iy2�W;_�ݖn�RWP	nâ5���Ŵ�����;{|и��Ln�v����z�7퓴���ǎ#�a7��:U��,tux�����b�-w*�ד'1��3(?��1mw�h&�ge >O��jD�����*��Jk��������)�T��➴�K���I(�T�	�o��Rӥ�Y6A�H
�	�M򝕸Y>j%�����Fν�oUH�|���ֆ.���R���6	��tq�i�M-X��\��bް�5#��R���R.22��-�fJE�֊px�6�n�E@v�	���~���z]D�l���ↆ�i"K#MG>��=Іrm��T�+//s^��hI���抝&��?邋����>�6�F�H�v^6�b"�wq�����K�w�k׭�0ӊ��I^s�����̃�G�'�f�&��&�%t�#�����}K�ނ�l��:iۈĢb^A�U���"��?x��I��.�Vm�.N��%7W�UG=�����^�)��r���ÂbzY�������q Vzy=4����]mSG�점�"���ؿ�֝@~�� �S�$� �ɫ��[�f���Pʴ��OR��������C���"fQ�'9�4}4N�d�gu6ə��O�~��sc��uIn�t���ק����P�מ��wh��֬	ƞ��*q���<�������n�<��3������С����Ih0�5H�%<lI�	�C�:N
��u��*���O�_a.�t���#��^g�+�S���`�EOWCưE���'�[⪱�y8_-c֊`��;��o�:��g���O<��7b����gP��pd}{wᆯ~�@��^z��8�؏�L�#� 7#��ݗ��������@�����4"��Z��\4t;o���X�}��9�'��m̜<���%��9��PFK�8�]sN���o~+�C�b�{�	������o��XE�N"v����e"�v5��'��n��<��?~o<�=�HPHJ1�Q��8=iR- �Ր7c�xN$%t�鞤�3E!m��c�^�\���WCM��t�a��
9�5����@��A� �r6�z;��a�(��O��{��\���O��[oR����cO���QD���D��cZob�k`��Qs*2y�����d
�&mmh�4
����"&�548��}��i�"I��1��tۮ���FM4�sh�{Y���W!�r�<�Fv�4�������(~�>���m��"&J�(�*���[�����u�!�49 |Ҋ���ӂ���ɨ]D[]�|����m���.�||Xj�B���f3�nz�|�׾��5�0q�4�������L���^��,��a��x��~�������=����-(A�PH��k��X�A��(<�Uh;�r ���_����C0���Oo�7��[�\����kY�Q��$T�  �ŵt��۽��_:�p2����D>�,՘�j.���o@�����<{�M�:����==���cpjeL4����pս�ƪ}��D�4��W^�ܻ��o�a�<��݈D��%����󣗊\@A
�ł���QJ�PP,������-Ƣ��kz��y������%Y¼�v�T� ��k^��V��4|�D X��Q���XB
RaC�#t�]'��	SX5�jM�	�9-��pG�;���ا�.z����G�HF�4J&9� �5�-�7J(�H��I'"�A��MޜLK���0�~l0q_c�{o�2��"�`"���xӱ���I��S[)����+l|rT�?�{3@��s��6%�N*�j*�Y��oFn�!�v�f�=�]}&�R)ؤZrH-M���!(�]����:kI�3��jj�m�B�����L
�yA�
�k!Vq0�ڛ8���P0�7a��}�B_S7o���D+Zb����`��`9�� E��5P�K��p2����j��KR��i�k&[�G�S1�n�+�ֶ]�䇡�I
��E�$E��']2y�d�%�] 
$(|փ�RZ���<�HDQ3��	�Ǆ��D�@j���0�ӟ����H8=����2��.C[9DPP�v���[���ֆw7~���/>�Ǔ�����
�{��ї^|����ߨ�j���wxj+�N��ȫ_��
7�л�^�R�s�҆ T �ő.��A�6��W*��U���XWC��E��G���FN�h"�x�!d�MPP�b,���}�sZ�o��2^{쇈��a#��9�D�̧3�n\����uo]8%����x�{�a��%ĵb����T�6Cc:�c'i������G� "�O�	=���_�<��ԃ0�2�?�:�����ؑc0��������M�!u-���̦m����>y?�t{�U<�W�w_8 ��D_,��a����8y����?��7�B��8��8��S�q��l�q�Jhfќ��i��i�ƒ�&�pd���A�t;��s�*�e4���\�@'��ۑ��Nۂg���H�Y��{��{f~���o�w��oPl���>��?� L�B���g^@��HV�½O��`Ns1Ѩ���Qo���<d"���c$��դ��	=�CA��ai��
�`��+����P���$zX7�""w#�:>�6N7�R j+F1�e6]���l@:��=��B��b8s�/���H��麘s+���Xpjhrm�y�tm)��f���aѪ���O��L<��m:hu5d����}Hk6��G�dZx�m�dÅ�D��M�z�^�޸�8��a�͟�%&&��/������{��3��GQx�q8g?�ta��B�\Xp�8����,EL*��5#0Q�e(��T�8���(3\����Bڔ�%��9,6@d�{P�"�r I=R��E��
�p��2�������3K�b�vCG3��]tP18-��ʛoA��;D0}~R���<ڧO��'����E�(r7⪻>�ܶk���={��ܱw�기��R��I�Dڕ�WN-]5M�3�"�^c�u�tOQkS(*�	������Vi��Q��8�,\Hyrdl�B$�>��(	C�h�:ݙh=I�%��	15�F�p��+H��N��O4*�$Nt���m�o�RoH6�b�&�4I��U�_7��nGtB
)�	$��.uR�(Z�Ņ��ql�8�c�s�Hm�
�%�	����R    IDAT|�|K\�4��MF"HP�F@������
"��=5@.��tIT�B�v-MĤ�WyEO���MPХ�m��fX��+�����0��N ًJ��f�� lIZ�mR	
�N��:�2(���t��{�����XĖ�J�eRХe�-�V�K�I�.C��w-�1��k(��
��]�"��p��;L-���Wr	�ςӡ%*O���Ꚑ>�!|��P���FM&���5�`�����^�&J�N�����{0z߽0�^�nn�Fg@��,�4?e.�^%��/���jR ��L�fi�ؤ5lӑ�C
B@�uI�HZ�`�[p_;��'&�#������x� ���5��^�u��Ϯ���Z��گ�4�/��cP�Q^�_�sW*S�g�{�s����w��d�Zaѣ�Jg�`�,��e�|��a'`�����e�Y<|�W1C�<t8n�=9 �z�jz�&��89�Аv	
��(�K�(1&��Q�[w\4zzp�g>��$z���ƁWpؒIc[4��#G�xv�M��~W���_�V^�hUp�	(�?u&��Y,q�[6���^+֭Ɔm[�693#�$��QEt$29X�$�d;����͛���~�5<�������C/אcg��*q������m�p7�f-����ĵ�y�$Q:}
 K@���~��8���.��p��������|�_~�[ס~�$������3����Ȉ�|j�r����-a�D�@�0Dg1�H!�4Y�T�b˄��ҙ+�L�k(��ч�	Ņ-�u�v$'�э$a�#�y+�w�D��m�ٲH�����W�7�X�V�G>�;�(p��ǰ��k�*��Mz�	#��<Z�j�Qj��|��]��^Mg`���bd2(�NW
�lTQoQ��M-����|� �>vɚ4���5L"��>�$b�f�p{��Ū���b�:	�A��n('��K�?�<f���@�KZXh50CދL�m)*[�M4E7@�$�Xj�({A�;�iN�6�]+s}��*s8�9%(8����?�����v�n�����n������]��_�W~���w��yt������;��)b��p��r�{̢Yh������%8לc��V�$�%vU�6�T���#K��t� U�XS��	���ky�|O��/�b���	˺�a!���a7���Ա���ׁ���;����1<
�����.�����q��a�ٶ��s��s/00,T1���8��3(�=�4��D�J�4v%QrUZd^�JCdY�/�9I����t
�Aإ_N���2�7���iS��!���1���Jʘ��+�V�Eî�L��%������\)�c���\�dR,.	&�;���F��0G�v�C��	8h@�T6���괐4u�c����C�]����P�1е�7Q��ޡ�Au�^<���R��І�tHW�J:�mh�ґ�)����V@��ꋟ�[��C������zS�l8�?>�������L�Ğ�=7v �I�ȑHC�p�j��F�V���O��?��.�wmo��U��J��,�Fi�r�ÜI�	& rnt�s�9��z�����Z�D�k�U] ��9�����>!��D��K�!��)��V���o?����J�b&�E0��2�'�Y�2��A����{��N�@6ٱVv��u�0�F�x�M@��9$�JnN��X���wp�'���)Y:-Mғ� ~�ۅ-E��L���m�T;�,4����^�E\��	
��&�3N:nk�$���i�ړT7_~vL�ה�c�ڀ�`!� �k�<� ��[�̼���1�/qP�6`��v���*���s���m1\�x�{#�0I�t�b�ֻ���SO��YO�T\u�,�b�9-��U���v��w���?����X~
�ʋ�U�v��/����^z��}�ƭ��\�jK6v��������^%�&���Xu�W:�\�ܘ(n��4�v"rm)@��Q���u�\P��e���IK���~�I8)�&�(yn��wta�ч��o��v��͋�1s�*Vv8�uL�O}��{3Uto���ۋ�G��Z�L�����'~�TnM#��f���XI�:��`�CG�}�44`�0;� ��-�R*r�.q��$�d�\�`�����_�?���Xe��p�fВ.G�&��B��J;{q���������y\��4�~�)������q)����l�Jlٻ��O���?|o<�S\��]�( ��L�	tl�G��4�����I	����9j���b��2fɗ�H͠ud �\ɐ��B-	��Ȭ^��;va��]H-�����oidz(_:��^|��:�:�-;�ӷp��?�ԛo���A��mc�0��0�*��|�A ��<,��B*��f�	��T�U-��h5)X֥ �}�W��љ�#
u�5}Ri��k1p`���>D)�9�3I AN�x��o������*j���*�B��G�FÌ��x�ʨTy��R&V����qU&��j�PJ��z+�� m$aEI$�%�ݽ�-�"�f��V|-�(ܼ��_y�/_��G��;�CӲy�g8���Q�p٤-t=N	(8���x �+O
����/���� �q�Ȣ7���U`]��[L`a*Q$ECQ�wR	�b;1)n��`���Iq�U�7���������W�r�aK�R8�+r�g:ڱ۞|+VZ�+�U��'��?�_p��q��>|�Ob`�nK��c8�_��/ ��AO����ɃW�T�	�m[V
�I�i�bׯŦI��o��)=�Eb����v�w�����oHm;d�w��E������"��,R�Ta͉@���I.��	
�6AY���u~ۀ���|��4,�J�(&�Q��F���f5�wq"A�©���[�CW~�L���2���=!��6���@�H��y�~�	K�m�E���)SL҇8�CȘ;!�8Q�b���$y&�p:(����� ڈx�F��q���P�r��2�<LNOI�3�x^����
�}�ŒԳ�����s@MԨ7�5㰹�y�H9��u��Uٕ�VM�~B�`�V�\?tD�BP��)v��'�uL�s7�4:�'�Րӹ�	x��	����w���I�mM�bة����;(>r�c�pg�s������I��Zw�-��Ro�Z� Z*�6P�90�oA��#�7��{4=D��P`��^�]l�z
%�?7)��Eh��V-SR��PъZUEl�W���%��L<�N|�[�<�]AW��T�E���4F�yC�Xq�Hc���>;|���u�)}���ד������Ug._��_{���~bl2956���2*�Rʳ���$�j����"ҿ�ĊDj��	�Ƈ� �\g�b�^�~$�6��N��d�2�ͤ�8t�	P��*�10������;x��HZ��
H�<�j���#����`)���Xz`?�G��n�xo��_��koI�9G�$�zhh��k��q�ǀu����"!�;©���'Z�џ_lj�0���x���7&O�G��'��H����$���1`�M#��l��_}�������ax��L̠4� v�ytt�[�'oc泏q��q���hMO��]��+�|��i9�1tt$ld4y�@@���8ID	G@�l��[�.�P' ���(&&C�2�4��nن�>��]���+�%)��f�sL�]Ԧ�Qv��y�h:1�+�{�M��-`0��af��n՛�jU��d#�ᘍl�#S�:S;�&�l
���+�Y�UPv}4�D�<�H��-����k �D����څ�}���^����Rn�$*��9tI
Q�y�˗0��;(���<=�#����(�����t� tZۇi��8���YŊ�E�p�]�;�<��DM���!�)hz
��5��������M�E�� ��m���r�
��@2��f��������#٪�#㠃��PK8	`KuW۠�k�kv�dJ��L|1������P��BO���<�S�I�jOM	X����;�'Q���^r�V�ZX��4 
j�]Ǔ�R�8�������/��VBC"	�ũ�7��жH��E������~���U�N#4-��_������7Gq��q���@�/�ѫ�q�q�Q>}K8������苎b��Gu4	�D�yS&1́B�ũJ���S�X����L����/�H`���B��LUT	��"mv��I��'��cw'�l��@�@nK�ZI#cq.S�f3�$�J�'�B_.�<)��w|V�$�EXh61[���pQ'�_h�������ˡGD��H���#�d����Ź�x-�Az�����-R�sBP��Q@ )r��V�M����d��&o�lF{�RT�Y��->�q^�\G^ӶfN@uhL���S�ȌPM蘤�f�0V?���� Hw�i�%A�������ꛮYb�s�v��G�| �Y,��Ѐl_4C��P��[�F8�Ѐ�T
�j�／�����Mt6�HFMe�{��!��,N���M#j��vR���_H,��L�X�A�b}���_�-�f�B�FB�^�N��#��w,��w���!X��3D�%�$;Hܶ�Hc�@�ۚ�b1������
(�'0�5J'O^ ���4���h}r
�/<�h�rfMX��na�2���9hK��)pw���܆]��ֱ��%��量_���_�Y_�������?>vsc#Ә�)b�Z�{��c�ve��(r�cwb�S��
=3ݖ�7��&�Ξ��A+�>ra�l�*�X:�Ug�>	(Xh��Vhb6��]��w���{6���i��t���w��/�������Hm��>���x���ŉ�~���/���L�`�A���!l?x[�솝ψ������z��l6/��e#0,q�p:;���W�ťw^�+�(]Agh��E��� �Гhvj��=�uT�����q���cӞ�p�{�tnQ�!-%r=�e�V�إ����Wq��I�'oA�z�2��"fӔ��N�B7�]82I�c���L���i40Y*���֗&�⧯��$E�G�l�fA�����*@�C�\Bev'>���u�.��V�K^]���f>z7��xg>��z}�;���`���d��"�h����F�F����L'����P��f�+�i�VPa�Bj.�֚���G�r��v"�ه��R�؉����g�X�?;�f�'M���d�V"��W/@�{~�}\}�E�M0�k��4�P�PԦ*��+�����6�7҅��Ip��",����m����@�Q��w�B���w��ӿ6���W0~�z�b��n`�2���M�Nc/a��i|���0��G�.r���B�ߙ�as��É�~�Ů�2��!N#�0��ň:�kՆ�
8H����&�)�Pt vY`����k2lKWl��H�y{�pۂS��+���G�>��ؙ��BZq�I	a�Mz�&���n��{���G���o�J�bP��^(��+ǀ��Mwm���a�~	���ￋ��*Y�
5EOL&�M�,X��c�d/^��P3�ۥM�͗ᔚ��+��	��e�$'�g&��N%��I�&v��QB��$�sL��i�E�_��DOr5I�Zt�!�-�v��ב>��7�G��$:;ЕN�&�{i�Ck����51W�c�V�{&Sch�J����	3�ޯ���݁��3� ��-�s$�-T�/�ѝ�aIl����ҨZC	&������-��}����f�_q�R�X�^TE�b����<K��^z���p5����`���k�`巿�̡�l/ZFR�.�E*�VQ��}S Dr;������"(hO�b͍�zy��� ^Óο����P�p��,�J3ǎ��S�Df|D@A�z'�Q�iC�E;'.q��L�b�P������;�U'���Hh���1]�N-ѝ?�Ϭ�z�'
*SEd�`�K	Ns�BVM
����.�s	[� M(�H�i�J�uz3ǓunŠ��ە�J�q�b���EiV��Me�!�
���n"�k��V�:���_Bx�RZ��&k2)�{1t�?�s��6n�����/�4�|���z�(�,x��.���?;vl���n�N	(��6�a9�)�l�1�@���� ��;:r���?9���.Q?K�@&���K�K��P��0�N�#���~.�B:�7���0]i`��PLw�o�6���'�n�N��z`��V�/c��%��.ܳk?�%��U�\����K��4�n��NAo��>��K�.�L�eː쇕v����X�R�G�k*�ޞA�RP6^m`�ݛ���$Hky�5����E06�Xp����3"�п<��\�j>'�r���La��wa���\=�ή)x�H�M��Z����Y�\���Qd�V�����nVQ0� ���Fg"!»�	��@h���uܪ1MQ���p�`�H�E%Gr99�V��A�]�h��(��p���F�p��{�z:���#ؽ:$3X(TP�����O�8��7�by���{��<&�n5���O�@��D��òll�#X[G͌p�4��jA�MC����3�Jj_zҁ�Տ�����V<H�I��>?�µ��L�ܪ��5tu��v�}�2�]@����N��/_@����R�a�H2����\���F	U�C�NQy���GЌ8�L�-���Q�lJz@G6/������=�����.\;wŏϠx�f����ʕ�~7�n���U@:�B����1s�>{�yx׮��Y��dl4`RG�[Vf�yK�Z��CU:�� .~T�H��%�aA�����
�],�cM�!aDj�%�kU��u��!IL�m��	����{I�A.�|��y�˖$���LH7Þ���dj)���ۇ-�|���kV�,U�h�M���K5�Kutv ���UԋS�97�� 3�ٳ�ѝ�ź�S+�����Ft���i �DT9���\I�d�FPC9�B�aSwE�R�(\�֛�17lK��tݑ"��~�+��f'\ٯ��阋�]|K��pYPѩG���eԨh���"늀D�̰�,�����u`yO�Lf���Ѣ��@9�0W�cv��j�U���*��� px-x_4O݉Nt�:��wH �4�\�O��"*�~�Y��=��!Á�Y��r�o[�~q��N�'�9⤀�@�<	��@<���b�@�NگM����>�Y
��V�������~�{�8��|/�ZB�T6�6��sUx r�����n�Q�i���1 UWM<(r�v���k��D~8sCC��L
�bSo��&�������6�,
�c���מ�87_��K��rbS��v��?񯡾���NE����<S �=yT߫�u����6x9��SA�b>���mX�Ѓ���~���vB���q���!1wg�oJs���!�K~ח��i)w�	I�tC
#4��!=S��
�����%�*26�1Q+�VPF0؃������av���AX;�UՊr�������+E3���>����}񹗆o\E��X��Ro	�=>U�N�M��.rq�;b�F�
VJ,rD[I���Y�W�|7�U�&���6ɤ��bN G��&2?]$����B��v�
���"t�uk���A�;x�6oB.߅ tahMg�ѬjH:�p2��uf ���k�c��G��=T.]�Sm�n��g`��ɸ�A��f:�ҡ1l�E���zY'#~��[�K��j�N��w����{���s�#9W�So��U�7��ۄ�0�h�$a2a�"�m�tN�����$���'���y��[X(W1]o
pa��+P�9�ɳ����l4��A�.>���)�{'�)$�y�IU�n�1V��t�,���T�kc��� �&f=�r���qYv&��K���Mc�U�ő�~�j��Бz��`�]�r�&�.����G���3�ΟB��M8�*|rnsݘl�V���h�Bt3?�	,K䰢�_@��.�c(�:?��򂄉QW�\����B�P��������#a�}�ֽr�    IDAT��k���Ƈ�C057�0k[g1�b%�����}{�+���)|����<}w�r��e�'�_'	G��U�TK(z54bљ:�I5��:���V�P�����W�2���<�l߇-��>0ԃ�g�`��a�MC+��zMD�H.[���бq���}�p���p��_B��K��g�2�$iCQ$���Λ:�Yh����uI���i���J #���%��qTN�II)W������*��,:��U(��Ch��&�-��CY_&+>�n�D��샸0X�hĢBᆋ�'���6�M'wH��Tuu]��ȯY��E���LF���p�E�-f���f�ߋvln��G���8������m��K'�������T�6טŹt�ؤږ8f$�h�ّO�np:�� ,�˅*�*�<6<���j��"���H�1$M:X[�h��N
�ZI�2��J)gA�>�,|[�,�R�J������6ɚA5�pˆ�J	Ջ6�< �����Y^�)k)�IUC��ɡa$�p#\�>���B�����Ʌr���wc`�Zt��!�ׇl2�\�?5���rA�zU�w�!|��1�^B(�b)�|���S۵I���"��Z��7�28�i%�d�F�πc%`E:��� m&��:��$h|a��8�s�G��\�4��}[�k��2����D�0)�r4w��{�	.<�q&P���~�۝u��e��<�5:��(K{	��3�h�ew� ]NCO:�t�������ϟ�5r+Ly�QS ��!gy�mi������ޠ��\S�d%�ŵ*���iB���`�z�	��f�h_b�]�����������ç��Q�4�r)d�n�҇֯��MϳQ��Q;E�O���d��I A�8Qzs���L(� �禈���A�1)x4�:�E�&��9���30�򫈮^F�+"i��R�d����`p ��Y������m��r*��U�_����^;������~�O��3O?�EP:t;	�}���=��d�O�$7�6���C���M�$"��#�
����>�:���X�qC�$ig�i��Z���#(H�j��&(H��8]d�Y)Z�����9����Ǒ_�U��ܮ,B��K[�ɡl�)���a���
�0
�^���_���HU[pZ�����>���0���Y�n]Cub�Fi?�᪔Qr嫉4j�K���l��Q8y͓'��s���/#�ұ��Yj�HG��`N�\��$�dV�k.{��¯g>�|�<��9�z�94?�7�;sr�f��+�4DP����t�����f���4�"2fA$�_�4 �R�5 s���:i���9v;��V7kL�K��/��F�9�)�ٝ�����{q�c�cՊU>xso����	�i�:���\dc���x�(�n�p�!�Xq�B]|��T
5#ĕ�	������H��@��-t�t�j�_���=���~I?0~�^|�;ǐ�5��:A��[����%,�����G�;߉�Sg��O�a�c���BqA�b�"hN:�����hi͐�Ҙ���&	��w��ȧ���V ݥKR˷��'�s��T@��g}�c���ШU1Y+��N!�z-69����E���2
/>�s����%<��|~�h�=R�y��b�ݦ��+�4����UlwFUwT�C�.��b_��P�􁶈<�-�T.���T�?�w�˟�U�֤(5CK���)1b
�tb�ˡ8���\s�^��2<�UU:�tY�,ќh�]�{r��
�+��p�c~�� �zavt�n��J��(~�1�>���8�ЅE�l���ZZ��@��$̑����rBj��@l����l���hR�՗C5�#�N����>��c*2��ӑ�0*��P
Ja����4<4�M���,M6�5eIOD����^�R�fG'a��%}��`���=Ol~H�Jd����-Y�t�R�]���X)��HY	8����[���q��2��b`�0��^d���)L�O���Oq��q�ZD�
aP�p�a�}G�e�}H�96pB`|�K������jV��>�e�6��H�SH�c��,�	g��owЕ+X{�%��Tu�E��fU]:��S�j��hRO!/�uLJW�N¢6�v�Z�@���p�C�Մ�ϻƽ�"-����!X�
+���B�ʢ%�����ZA�(�E�A`(�7�k��;����˴��/��5�fI�G�����1��D:����d���co��S?Et�V��i9��ښ���R�QE�����FdH���$�zT\�(�T<Ӊݍ$'��5ḩ�������tG_M��05N�h�a��!!� �g+z:*�,�u ��ǂ&�41�Ԥ�Te�=䋉� �2|qr�$Z
��0U��$C����<K��[�1�Dȗ���]���=�F	�d =b������%�X{����Iz͆��n���J��e�_���^;���W���O>����ǻ���Z-	�8���{Z�i+.��Xض�k�L
���ce���X����F�J�V]Ѵc#�H� �	C��=�k�n�%E�	�&��i�с�i�g�X�|����kq�{��u{��D��[H�2������g%��
�[ &�O>����P:w?BFSٖ��J-n�=t}9��-r�];��sg�]EstvM8e�"֮B׾�Xq`�������}|��C��D?S��HAα��I����=CW��[��I�y��7��]�0�-�4+�(���|%�<�0�v�R�y����7��]F�׀M�Ƿ�S�N�� ��0D�ka�Z<il޲��ѼX:��������	XV&����#�
���G����`�,�u�drJ��p������uX�]�h\|�i4><�dmFƂ�Ia��	k�UE�z"0&(跳��AL�NHAW'}hf��s2&f�)����*P4B���X�q|������.`vW�x��^Efd�QA�I-�L&��t'�y�1l~�~��œ����*�A�t$H�	�t�����t����B��I'��|	ϕ"��m���¢��u�C@��z��|��R�N���µ�~�2��L �b9��؁�۷K�Z�) ��L����Z��.6y|��e,��^r�r��N	�f<��P3^ט
 ��(B*���%b�/6�p�h�˧����>,�����-����G��Z��+�AM��,H#���vQ��H��T��%( �%5'�𷻑�3}A\�����^gU�ˡ�����Q��Ѣ2߅��6�o���Z�,�ʚ�\O\����s�^�.�`��v�-���ъFs�	��.�$Y�S���Ϯ�<&�s�V������Ffy�V	p��9���7p����)���6�²5C�w�(�6L\����~S�i�X��]�p����$*3����9�kV���R�So��'їa�����e��L^�f�ܷ�iz�I�۵}��)a��dYb� ^�3����5��*�o76��wݽ���r�׮�ԉ�q��O03r�j=CK0�7v<p?����F\�G@��g���1���p�^B�룗�/�l�3D �`r��)=*�A�-տ]�������@�A �لLI�}�*��(��n���$E�N;��s*���jl�3<��1�4mX���}Q�r(�6�&�(���f�߅�A,���a��E��2.��p�nm�׺��u���&�#�NW��FPRh/m�衫_���a�?Gt�<���F�z�.nO�˰Xs�X���W�M<dL�?Ca�-:d��wQ/�Fb{q��嶭(�d6�S��P ���︇�[Tuo�� n\�(4N�ܑ��wr֮F#�G�47����t-�\+�q��q�,N�X���P���DE�SI�!�@�}l��
�V�g@�d���D�.\���/���i�Et�t�ic�Y\i�!\ڇ��cp랿K���/��_Bi��}��A�Wy����nN�\���o���_|�>:q"[*֐��`'S0����wʅ�DD�R*Vѐ�{���e�Cl�Ð1��i�7Uu�X��0i[p,S�'����#�N�[�^�!�D[JCC_w'2I�r�`z���n�k�j؃(6826�=8�ek�`x��#ՕG"eB'������Q=s�sL�!�'�4S����\l�1"���{��퇁�� �LL`�����)�������A)&r�n��|@��̎�������+�F��Ǽ
2��Zt`
`�t���ʨ�tTBu'��Vg��UŶ2���J�#jFw��C�^���e@���O1�ʫ�._@�ׄ���CĴ4"��rq���b�E�V��}�D^��a��6�Y&�:�H��HjEd&��jN
5��\qi4}�vF�
��K@�Ы�����]�v���䧘|������0I�'0Ria���O�>ҁ�9�(d
�-D��҅�4V��S�k��"Jl&���l�Vܽ� Ç�@�;
���Q?y���jn&	s�Z�v@��m06P(b���x穟�z�z|ݶ�����89��`'��:��\�B��B�*����ć_{��O,"g�0��ʆ��{�`ɮ�X��n��\�ē��3Ә.��E��@�A4>��S���Dx���cHի��@��K���h]���]mx�����+$�U���t�Ä����f��ʙ�$֢͒%,�*�Hz����p�!|ZB1�SK��+d8�j�{�BC�f�<��mwH�������E���Y�	?�bA�^�K���@�.Y^��� �7���u�ٲΦa��<P*#E��5�n�&g�c���s�'��x������1��!܈)��(�yy�Q�mx˰d�6XkV =�'�8����C<s��[Ȥmt���P��4,Z]Y�B���b�V��M�H�3��y�>�\��]D~a�ƒݻ��o���~���/q�_bI��nU,U9��$�����L�Z���g�����"�FmUSQ�h�ؘ��^��_�I&p�׿��M�c�!�W�4�S���+?�=�����ķ�㑣�^�FM��VY,��������'?Aw��n���1( %ˤ>��3�,��E$V���ݡ�-� �,�z�* 	�jל�c�^�\�
_��pR�.̖'�`�#����]Q|-�
��4���	�U:��S��a,��#p���t��[�H�\������⤥쁥_�ר}ZY��gN:�Zl[Ka�����2� �I~wC+-
��]�S��u�#�?�����ߔ����ZM���v���%��/v�U�3��3S���-w���s'��^���/l�ڱI2�C�(^��p�,�����	�����Up�y4B���i�A��|jEt�MT�{�\T@�;�4Qx��%L\�Ȏ�'�>�@(ϟ��/��:���� U8{/�����H�+�:\J&���P��b��Q��������uo��%��_����"U�M-��o|�؟�ɟ�O���:��t:+��f8�����py*��Iq�rCi[�޹��I�������G
�H1��׽nK�hp�M�k�����Gב��ۨ!�nc�G1НG.�Q*�<WNr�7�05LT�]�}Z������]�1�j5t��
±˘;}�gN��P��ar����0-�"�� �5�w�:�o����	�Nc��UL^��K��o�RhC�@-D�hL� ���G��r�b	9�(�f�9y�Ldd����2)�]#����u��ag�d^\th��;��!��L
Q.��q����_{�����-���^ƜZ�D�:Z����B���T�$�lԍ�/<�C�g�@D�y�f�A�f#�7�hX6�V�T�T
ٵ�]���A�2�z<���D�QAm�j���{���y}�=̼�2O!�*��Q'Qŭj�0B�%xR-j5���X��F�L��_��$�n�I�K"�崠��NU�	�26��F)4�r�><���-k�	\���7^ǭ�OH��u+���!`�~��_F�������p���a,̠ˀ�=0W#of�-�!d��7� 6�Y-[8����*�5TZ4%�,��#u�>�(�|6t�N=}З�����q��ߨ,q�%�Hvz
�Na����IX�s�F���6u,�nӶ�c��_(n�:�o��.CqW� �5g"�f��Z�P�$"���N���E��3���í7P���-M[����B��Zv���Rn{��4�1%�-$l��Yt?��K���UT9r��ݎZ�m��G�.�T���ވ��&`p@%��jh���x�<���#Q*�7
�e�0�HM:9�,Ф����2դ�"�;t��]��J�oePNfнs2;v ����X��K���!��""��	u�6<xs�M��bk�MuO�"����\6 ;�o��O�4�{���M
����#���ǐ�_��O?���c��!t� ��&�đL���i��u~�!�ݽv��Μå�>��yX�~6��	t�a��e�����K�����g��9�]�..b�lƲe@g&N��Ͽ,��7�6z(���N�µ��kX�b%�+��t����_<�����VE���B�v��������I5ǿ��#�c�2V$���r�@�^�AA�H�j���JE7@G_zz�Q^�GirJ蔫�{�O��v�sO�]��!ň�&9䵤�RG��*,��C����N�B̸b�m��B���߇!����M{=*7(��S��dq���,Y;�J9��
9ܶt��'���.���q�>����Xu�0��40ر�	Eر=���8��cȳ�.���n�/�	Hy�+'2D�t�&�NP��+A���_'nO�.�h��q����B�Pwc9�w�۽)N��� Yڒ� 3����I��t�:,�WJ% �Iq�X +QqCȃFP@+Z�O�p��ӅD%ˮ)7�5M(րs�0��;h�ހ�6�4XI�^	Jc���9t��v=�X���_U��_����S;~����_��~���Լ��ՃL6�$��)G�(�!a���h昔B�5����ﺝ�H@�N%-�����w]�;Y��_�q �Z�D�2�t�"�BoT��<��SH'-��:�&P����G52P�m$��q׶�ؼg6�ۃ���҅g�1{�,�N�@��%��)��5ƥ(4
H_`GUu�(0�CG+�m�z�7mF��Up`d��5~�)Bi�aW\�&��]�����kb�j�V9ڳ����	B�l'Y��/y>�L�ݳ�� ��2]"�+�M�A�y��"��(B��\|�)>8��Fi����s����y�
��5�[-4
E�>��;��+�%5`iWy�KG&��[O�$��I�`�8W)�o�6���o�7�,@�¢�U)䋳�g�Y:Iw�.̢��	N����0���J
�|+DZ��	�4D@O*���.t%����	U*�F`��.&�E���t���?�m����-L���@t�7~�<�0�̄�I���38���b��e�V�dGi�F�ݜ���g�q��Wp��I8��\�`����A_�9�+z�GM9���}{���[�t��^�Zu�< ��]��q$�ޘ� ޛ�����L2��]�p�Ï����Dz`���B��4��>u�����''���ѣE��t����'+M
5 �&'\eS
\��
PPn>���]�� f��Cɡ�M%�d;2�ذ��eh�����4���	�J%4����(�:��o"��K�P�V���.�M�{��NLV��S�ӌE�r�f�.
d��#ը_gV;�����P��8����l%:�V�X������YT�fP��ꍫh޼���i c��)�6i��H����m���p]|�tI�|4�R"&��=�s�*��X�J�0ˣ#�q���V���K6o�1؍�p�}h�:�G�����0}�2�3������1�?�[��p�2�%��b��H;9��5<��?����X�i���5V�r%���/��9:�RQ����t5U2ɏ�s�p�A�������8�SW    IDAT2�W~�4���'H&�>x���7a�^���,�}�E,�ǶGH#���<>��j��:��]��Sz�Ƙ4�V�]�q�S�8��x�g���u�Q�9�0��rS�>���� [�G&"=R����)(�b@��D忔��<�wq�T"����ϚI�(�0R,a������(P��AV�1<Ї|2!�7�q�����1�q����)X��<
�wH�0�y�9����
��BN�I{��7�.���%\��*�X�ɉ콪���w��B�D}��V������Jo���W�@j���)	�OMZƺ�e��t,�?�ͅv�$C��5Sk�`��{B)��@�k���8�[Rq�D�:E�5%�Hi������@L���c���q��YRq�7o@�� �= �7�$����O�M��::��5]��P�M���U�yl����$�cM�`���ye�#\F�p{�gF ��Z�7:�����<"���t�Š�K�[�����пm�����?к��*�ӯ�C_���'|���e�SO���<��O���n�r��t �ɠ��[xu>��Ů��T���N��O܎[Wōr!�]L�?�(�£	]�����ܴ��*��:�`0����&�h�l�t��Jp4_8wi��>���b��rK��d`/Y�5[�b���aǽ���M/]�ĩ���CL�=	�QD�НN*{ 7@ȿ΀�^v_l)�)Tm�.Ne�q4�]�ذ���aٞ�X�i��,M�du��9��9��％��G49�^vB#M@AW&!f��^TH�""��"�@�;f"��woŪ}�X�J����!Caj�0eT�R��OT����j�oࣿ�1n��:z%d�� /\l�H�0$]��j�^��|�����_KkX� ��A�$Ô<iZpx�����i��8�����'��P�%]��{��!8�h�t�.��4��~�| m�2��,�k��8U��:�?�S]&)V��<���h��3�e�Mch�w��9����}9K(��+L�R29,��lz�(�׮��S}��3�s}x�*,Y��e�-�к4���(\����("˃o�8]	5��$:�4��$Z����ۺ�]}����f�2��E�Y����"&��)����&���٦�f߀tw�}�Q���8�.U4ȡNg���_D��g(}~���r����F� Z�C��O:֋	���c��%�FD���5"C������~��D�@��`/V޷�͠�nZ� .�0R<��@�&` Ƃ�� ����c��i$�s��6e�`�*�K�Ƭb�:p�Q�]�S�H!��S��ր�$<�׮Y6ꆎ�i��#�q:7lH�#w?�P��ǭ��$%4fFќ�B&��'ӿ0��ZEƶ%@D�|�hWIG ^�X�(bU����ɳ��t�~U�:�j�!�>�0�Π~�*N��n�8& m���c����U�'���bg�{���:n|�	&�� ��ax�*��6f�'P
�X�y���oc��ݘ�po>�
�}~��N<���.���-��'������O��K�C$ڂ��QSk��?t�s�A����F���|/���h^�'a`�Ç�����w�-k�a��2l߲f����>��ūHrE�w���A���x����]d���p��Wq�Oa��q��>�],��@�pu7_z	��AznJl3�v7:�3�Qh�|fĎT��i�E�PU�M~�w���ץ�#�>����-W0^�·5$��b�sL:�U==Ț,�I�����/�����׸����tw�w۽H�{o\��;MkbՁV�u�����HZn�p�	�c+ZqR��_��qBu��I+�-h�{��PDp�k���
f�]����6}��S0C��y�8I�3F�Ni,ؿh	�&��|�s�a[J.�Z#�f�h�D塴K8m����)]������}�Ѕ�.�q�Z�d�� n�Ѿ���:���n8K���u@���l�pu���t���f�G&�Fw:�OGB�J�4� 1�7�٬0�l��C\Ꞁ��5��$���l�
-�a6<NH]4�摈8|��f�Dѯ�FknO���Cߖm?7�m��k��?ai����A�?z�����'��������ꅱ-�K6B�\��]��h�.L�h�N�e���ы���`�D��e*@(������t.j]C�RA�\��l�Ţ1D,%�.�0��'�u��
Hh�&�DDQ'���+�����w=� �>p=kW�7R\�(0}��N����h�O �38*@��[)�+�e���¹'}�v�)LU4��$�n߂���݇��k�t�h����/�q��y�y�5�|�u��*H��J"���$��-iS)�i��t�#�f`��Df�FXݝ��E�R:Sd21��@�tQ����`�=waۮ�p���������|=:��%9I7h�H���$rz���'1'Hk�Z!r���\���t��'M86�):892A�.�0�j�ta��X���*ꭦX�z���*r���ѵd ����la��UX� �V�ﾇ���C��943(�3E���t�Rϑۺ1���BE!b�- �f"�KR�U�TP�%(�h�? >�ڴ���Y2)�ݳ�6�#�JY�X98(^�,�'
�X�~�3W�+U�4��UTP[B�B옷tX��#��t])K��O�D-G�Fd[�)����La^@L�Z ���_��4z����Ʋ{�����M��c��1B/�:�� ����Ξ���S�ܼ���(:l��d����p]
��	��aU@��;)0�)�6���f���!H���x��k��=���3ڳC��@����,`�`;YX�ل[)�V/I���w@���7�ŭ 1;%"�94(��$D¢��. Wu�\������Lq����'��O�F����>nن�Ga����"���ç���*���*s��`��<��!n�<��RE.�����A:�����J�뜮Th�,ReD�m=��`�c���CGeB��+�⭟��W.����o=����>4jZHe`���'1{�.� ��]���,
�3�U8)��D�Ka�c��#O���^̌L�⧧126�#�yC�	X��ګx�?�Gؕ"����	��Z���c�Q�����w�Į��}DsU���O�{	��4�I�:���!�u;`:x��g�>��W��t��)�Ng�M�;��#y�v��Oٔ�|L�;�g���7�}ù4���q���#��w�����IL��*j��@b|��Tq�)xIGU���@|H+Z�m` ��p
��k����%2�b���x�"tK{dSbyW7�R)�}3��Ɩ�L��5e�	�@Y�t��뇟Hç��$x_ق�N��F����;�b;��'����V��Lt�ͪ!@R���HB,%D�Фͮ8yp���paT��N8�r�K��F��1�:�X��e�&����{��o��q찓��|�Q`�p>�)N
,�J�SۢeEV�������a�m(��B�5��2뇔Nb/+	��P�<�h>�Up�4��6m���N.�.���0<W6�B�
��h�@����jNS��P�zZ������=X�,_�N=V�G>�D�)q;k.�%,�
���]9,ݽ=�n{�^���΍#_e��5(�*��?�k���������.������0f��ՋTGN6/��pZ �����R��aKv��@��^Q�ܦ������c�s�L�a�
E��j�Q�j&�N��H;�0d�i:}4�p����<T���ۂ��y۾�mh�L�%�0��d�TB���B	Z�G�'e#��x�<�<f.\EN����P`R`����맺ѹj��!�ފ��C��
�\��޾n���=s�����������,��������7�/mY6ܖ'�ȴ"�4��o���ՓG2\tt���f�jnMN�U�����p�����w�%�ϯ�������i(��< 8��A	���֎�_N�y6Z>�!ГL�7�C�v�VZB's:3�R	���Q�b�TE��q�\A�I�ѝE+��Q�i�U�"Q�ѓ�D���ͣ�4�g�X��.<�裲Q���.��J���-͊���q���"}��KF���{ti3
,�ua0Ӂ.;��B�&q�M���Pd�X����J�Z������y������-޵K@Jm����~TK�����;'��!Y��ު@�]L�fP]�upI;��4�-��%��!�^�G
��B���r�
!�����*�B�Qh��ݸ��$��z��5�_��3H���;_��:MO� �L�� 	0��(��V�%�6�[v����������Z�w(1'�E�� 9�����]�y�I���w׵[�-k�@�3=���s�
S�p�0vn����9on\u�͙-��`*�/^x׾��
�4��Y��ҕ��E�tr�ܗ�qW�]� ўO&�����ȘЗ�3����p-����]H�u �ޅ������֠w��\e|��S|�c;:������0c�|�w|���|	M0U-��4%v��l({@��F�4"yO�>�R_���6�q�ZU�\ܞ�H�T�c`�j,�x:W�:{�.�Y0�hE���|�R	�K��jȏ`ǋ���ǟ V� k�d�b�I�Ч��c�k�k<�$��gN�G�X��҅��6�����7 ?4�w��v��2�q��6n|�!���'`��_(
�\5����]�Е�(�
8w�8.>
�Z�D�:RӺ�����ᛏ�n��R��#�vf���
�~�}|�u�N�@+E�P�T�����rj�N�Ǌ;����G8�ë�v����<B���]k��o~��7!�t�����W`�]G�SÊ�f�li��0�0P]� 3zI6Y���~V������>��>��Dgw
K���|��Q~�=���GXW.!��rr�	�r�P�����'���+���e�q�@�!��x�ѩJ&�������Q@>$���꼖ړq ��I�����h�T��H�9���!��K:V�0�1L/bb<����A��XL��Ħ�N}�24�
*��I��6�6H5Ò�,C]�#�4q��^N�A�1�W0��C�aBKY�Q%�n�	�UG�6�f1��BW�!.��K�T5�:ߢ?K\�e��g*T���<���j��P���{R�}�/Q�qo��WE���!
��tob¹)�],�P�P,�5������
v\=���Y�?�ī5�}�c��.ǈ�L<����)���^��`S�|���MO SW�05P�� �ɥ����C����1�qٙ��ьޛnB�Mkߊ͘�ﵮ���K���S��)���{��3��⏟�������:\O�K#�ځtKV�#�m�<=:4��"$��Z��>=h����1���	Ac����eqj
�ܔ,�ՒS�JđN%Йɠ-�`���cHU�ٺ�=ǆs��{�`�ݸ��B�ƛ�TŰǯ�
���Y-:qA���+��ὗ^���;�D�#ޛ�4S,����Y7`�ʵ\��-�)���p���=y^�� f-\���A�*J�N���/p��Oqi�^$�e�h��f���>�bc!�`Tr8&�@��ѿpں���NgH�m#O����#����vwc��X�j9�����a볿�=5��]�%l�f(����(���$�,�t^hh�,�%RH��,>|�TFS5�1<�Gn������B�7�`���z?2^��HVČ���������s�x�r�(ϼ�6�m}�SG����OX�,�=S���*c�f���;��DF�������)T�V�ʑOT+(:�� �H�8�"�z�p�F���#Hvv�ϻ�>7�JEc$m����Ϣp�jgO����4߫!W.��
4���'B������n*�UY�d�����0�N�jM	�yCN��d�aƺ��������U�;}
g¹�q��~� �f��-��w߇�7o�՜J5�y����ү�BQ6�l"�C�X ��"^��)Д� �, �k����?c����	���P�Pdc����݉��-�Y��=�-,X�R&��{�ᥗ%��G��Xx�"��g/����@��\����˵�>l����ZQ'N$���A=`�`j2�wRH1�:k�ـ������c��dv:#�����8"���Z��d����o���ϑ�<�C_�j�Z�V`2����)�,�Be)�n�B�A�Ԇyw߃;R�K���������/ Y�a[�{�7p�w���7�t�
�2d1C�^X=,�v��3O���=�K�N���sh�ދu܋˖�f�1g �H�4�b	�kcس������ǯ#�Wj.<�Nc�3a�k�\���wa/\���<�=o����(<�Eۚ��'1�{P�����o��\��t�X�։�-��S�1��MH�X�8Mj�����]����µ��Ü�:���a5�y�������`+�;`]A2���C�,�$��k�WD�)T����9���K��g��E���f�K��k�ϒH*�_U'�$�{���3R3}R]�����꺝�vA8�B�W�sE��2'��˱�T!lRݒ�"�UH6x��u�~��G�_�$jR�ؓ�z�&@YK�8''��4�H��f+�,���P	��a����ї� _%��Pw-�^&2gKC���w����F��@c⚆�x!M�Ei��z}A4��$����5��/5u���Z�}��+�u�&be�>G��L�.0i��	��}�
��4,�y��~9x���
5�e�Ȓ�T.��1f�ɧ�Z�$�k��8�ʴ��%�a���V@��l��)�gA4�X�����t˸�L�ښA瀞пf�;�ٳ��ֹ�̟���sS�<��J��K?�y���?��<��x��M�����VhDt	2��<�/�;���0��"��M���k�Y�����*π�?��UW�b�E)��DЊ�)�&&��*O�H��-=�-h�����1���4���+���V�\w�?�0�ݱzG��X���N\��H�*:���z~�.���oqz��h'�.9,�T�+�Ʋ;�����.R� ����N���=8v� .�>-£��i��l߼o�)��\<��l��W_F���:�*޶E�A�c�,�&*^����e�\���cX��Tt�a^����@��\���RE^"�Xږ��2��[�+��Yt�*�>��RD��/n��:�i��Z22���h�b"�s��Si)��*8_�ĵ��LJf�Đ�Yh]�+�χ�+���^���k(���X����Aj�th=-0�)�3)hN��~��zSǏ��9���H��C�J�Z}�A
��4x��1�ēh���Iˊ���qyLY�{'+5L�J�84��fl؀��,[
�J>u
���a��LN�����o�3�.U�.,8.]����1���0�\F��dc+��9ד�4"g<�Y�D)y��d�4��.O����)�bd� NK5?B�承�b���Nl����}�*���x�4��?��T�S.�<��s�7�a��uX�q#���D�x�����/���!9���v��KN�I�q<W
n���Uʱe0]��
�BB��h-&���"sJ�F�N�鎁j��1����9s0g��Xt��蟿 ����K����~���,����?a���.��g/���܌�[C<��!A�Fj]��p���̑�׿�����#툅�|��X́�7n�7l��}�-�2�H&������RAܐ�H��|$k��#��T�_EW"�8�
؆F\5ib��ŵ�\c"�|/D̈�C˞8w�y'���_ݽ'�������3OC�=n�c�2l|�[��>t��DN�łE��J�AE�!�q���CC�6z�Y̜;�9��Ɔ��r��>��O����^x	�}��gs]��q�t�x��/q�����7��⳧_��/�����:��Ý?�>�޷	W�����������e�M�13ü�n45�P���W܀w�}�<��V�vV����    IDATe\���zG_~-~�2��zn�я`̞�ʮ}8���Ȝ9��r6Aȴ�%�D,h��Q�꽔eV0�<�_���k�\�ql�]��C�X���LX
�lM��hMJ��D܆FKVa������r�腚����7RT���h�LXg����U�'�B�kd(�;����11��4�6Ɠ�N�
���c�
�R�����A���߹G�y�I�F}
Q��UtbD�t�gR��� �Qr~������}3��y|��و�؈�`SMJ-��9	i���m�����4��Dŏ!�E��=��rJH��企� tN7�h�p�V���+�fj�5���i�_�c�nhk���^�PPsTS �X�gY'�|-�$�	�"oE��P��#D�ɨ ����elxNucn�����j
V�}?9c��i}KN�+������sS�O:L����]h~���������Ȳ�g�nnF���m�.Pn,.Jb����F.�x��2�b}l(M��*�v�cZ.@�Y��DLe4��u_e��Bc�#��ʂ
s�i�lDf��D)b[�v��k�MD��&���i�Ji
�������P��<񜶐�*`"?%��D<��&:�8��Sl}�Y������1#(�ʱ.�y�1�����q��	>| WϞ�ؕ��)��E�je�}㎻�Ě���p��ݯP�p�&�QIgP&����+�"i��s�=�9�yTP$Rb_�
jY6�?]m�&eȏ�pj
g�{���)�G����C\��D�������
i3��D�x\eZjZ:�!R-Y�&KU�p��a�Qb�� �J*��O|w���@OpmW��Y��s�t�8M��6����s�U�����8���8��f���H6s���hUDfⴤ��RhQ��i�:i63�$Z�i�c����p;..K��\�q�	���b�w�-?{B<�O�݅＃����4r�[A����~,Y�e7o�̅�(�@u�N���Ȝ9��J�(B9pqFHY�V�xӣh��h�'�FEj��RT�<�Z���j.'ӂr�C�R�넘�>a������5�W�����\B��$�''�+Vj1XM��t C��(��ͯa�?�'x�.�J�b#^�'��#.l�V"}"��]o �M�M�RJq棘V�euH�i��&J�m�q�������X��nd�"jk��J��Ma�{���W^C&����w�=:��Ν�ޗ�ǡ͛��I�Q$��a�)D�X�hdC-� ��/��R��I��@K��ZY�DGkU�f��o=�������R�YI�&��[�<W0�Nȅ?��3|���tp�v���0�`D�jd�4Og�D �(,�GQ�xD�9CG���x�/{�|\������o1|�8%e��­�z+Xl�;���}�ΞAWK===h��Ŭ���2o�]�@�E�c�0��:p'���6��޽hɦ0c�|�Y��i3qz�|�܋��b�ơ��~�	��"z�0R.����?�:��D1�ܺo��i�8���w�<�񝇱��{p��a|��ft%��;0����P�t����Gv���"�q#��G�P�7�����`����=�5�+b�_|_�Ҏ]8��-d.]D/�(��0͑��>)"u��np!�%Ȍ��*d���ܰn������Os�?ll%�B��U
� BH��Љ8�UNT
���	WZ�@h@RhK��}S�-b*d��*ѢA}�S�(��#\\N�|������L�\@�/����­IP�+��:jLe�\
d��ե� ���zː,>V��"�D �i�4$����rqۖ D�N��s2)(��VC��<�8�=���ص�L4��q���`РͽH&��h�Q?>|_�ӌ#pk_�<W�D�y�T?ȉ"�$�Yh��!,:���x;�K�k�*Ζ
�X�0�\��4���-�H3+'�d�!i���K�g|!)H��eZ(�,�����x�A�����Y��0�ti��Lx�F��L��U����w�aڪ��]q�����������*��-�ۨp�����S����p��y��z�Lg`�S�����E�)�u�t
��֘��A-Dr�ԋ8nܮ�F��$�u�t�$���� "�(Ӌ�>��c'l$���8!R5Y��N#D�J�|c����w`���ü��a�-��a�W�=;�rك�B8�B�B�����C���gq��בr�h�q<ǌ*^���y �?�8Z�.F17���!�5!ݒ�P>C�\B�TF��`��9��@5���-l�ݯP=w���$G�Gs��r</��?B� �ދ6܆���!�א����oպ�hjo��*.�>+������FU�8��G���g�<�V�0���g�����NR��,��)�����A����7a&,Ʊh��x�Ôb�(�n����4w.��7?����n��p��Q�B󊵘{�F`�<%2��c{V�P*���`�˿���b9�p��w5��u:e�!��r�	�D��z�NI,��l[
o�G�zL6e��E�����B��-ǲ�]�!ȍa�+/�����]R>�\ϫ���HC�V߿	�ل,C�N�ƹ?��`�.t�H2��1����J%
e%V�x0A�7݂�T21[l_�*��j$l���B���J�����&y�B��uX���^C{Z�5�RS��^�1��V�����.�q*|g��wq�W����r���@�M����"G�Kc��Z
����  ��t!�����,��B�����+��j�����:���N��g ��8h��0� ���g"��o>��i���ۏϞ{���Ę���h�c]/���bS"���^����֐�CX<�<D��+J;P�C�Ɯҳg㞟�s7=�)89A��$}�kU�ot#ARmԜ0��������/���cf&�DX�yn=d�5	7}���f��E�/�9��֩c���̍7b�wÌ�7�9��y �������+���;0w�q�<��.:�h2�(f_-��Ѻt)f-_%�8q�������G�������ۡ�.��c٦��j���.>z�e��{��5d�4A��Ս�:�'��9��˗a����w�L����pf��'�5�6݃ŷ߉������m�58��-E-��ȩ��r��RE����o����̙�8�2V,]���ND�8�sN�ډt,D��ظvop�0μ��c���e�I��p��5Anf�0u�������S��z��8j��x�~��"� "�U��NE5z�m+:e6�7-;!E��7�C������/6,�ia�}��#�_�o
�Y򆢊Q�'a���IIq�nLJ��Ur��'�=��)w	��8�j�������I�N��r�!�8�~��L�i��=>Iz���V����C��yF\��%�F��J�����O����4P{�{)T��c��%��<�f���!nR�!��&��)1�HR��� ��ԫ�?�7h���H�ьԱl�嘩�p��������H���Fd�0ah812�3��(�ю�b:��&-h��0k����"PjP��*�W���o ���[�7�L9qJ�͵�Ǜ�X���sw�T�������vL[�
��Vm��f��i���:�ϓ�?���Wzm6Ͽ��������C��$V�Ґ��4�F,N�����2�,������_ryqSD�Dȍ U��Bo�$h2MUQ䑯:m
�
ż��Œ�x*C&��t���rh<t�Z��2��&̹�a�����]�
��N�@�J��(�h�$�5����k@�:>�9|��F���%�C��F�7��mAo}�	L۰*��X�	��@����%`?aHc�1�U\�����������T��/~NN	�]!�`�8�Z�HJ���p�U�$��j������>�o��p�7}�1,��f)�.|�۞y���������N��B����k�dcI4��HYuے�jŔ��8S�GD�����*\{E$��"�.	��ηp�/� ����!z�=��	z:��w�=h[y�҂��.�������a�Bt�6�x�em�a�1��L��b��g\F�b�	7^�(��q�-m��8���}W{lH#�ᚏ����[n�����u��[��%Nl~��(�uSD���jTn�¢{���xm=��u�n������r)RG�Ř���U�+e�8)�+��X��c	�$�Ҽd�8����H[�Ŗ$0�� D{�J@_�Ky��!Z"�D �)�Q��\~(��i���Յr��P:|T��s\U�ԭ�6�I�uˤ0��V��\M�k��PX�ԑCR��0�8��h_��W�C���ΒIL�X@ك4�-�Yq�.�����b�{��ױ�P9~X�7�>d�j-2�zJ+K&�;!���3�����U�Z���n%��q����!O �:�x�q>�� �g���ѓ���э�+�`��;�Dv�,���.�v
��W�����G��
����"j#I_����%���f��FҐ�X�������Zs�7o��{D�E@����p��Q$2I�̞����`v�!�ʨ����G��r%N3$�>{6��E�a��������C8�.�8.���{��ʵ�aE>{�5l�)�k.�S,h55�a����&�"�܂���?�XK/rW�c��Y�\�"����nD�9��x�vmôӰ���Ե�ˣ<:&�'D��^	��_��7�ނS�N��o?�e�WCom�J�2��� E���n�:�ko��ʁ��6t��fת�k.4ڐq
��jZb6�XRB����rbq�_�/�n�������������9�!�Nw5VqB��oQ�b�:eZ���*�
�NH�#�����_�Y�54u�[��d1I!5_tU���m�m����^��z]����C��v��)Y*�Դ>�̂��!M�SY2V2���Qő����3Q�e��u�bn��
T�4���z���0����\SSE*X\��~О�ҤQ��ʘ�z�����=�Q��l�"��՟��L&ЗlF��D2�6��"�*��0��/�%�e�B�)���5��3
K�V���y�U�d~�NS�SbE�5��5�l�@K�F�n�U�(��j��V���&�1��+=l�8�_*����IzI�Y���4Yg�0��Hژ��*� �혾f5����ܞ5�ɦ�?7�J���?�6��z���w���w�l�gN�jK0Oqq;�����0��~ h�:ǆ
��Hn��p,�E�k�G���޼\T�
�QT�zl;|�Z%z�;\��0�̎�-n�3�A:2a�ʈs�<��l©b�P�XC�m������o�;v�G��v�<�N1.���tS���� �W� ����u|g3>{�)T.\D�e�=�,&*\;���n�Ɵ<��������_.�;	E�,�(Ȣط����!�����}������h��'G�����v�M�8n���o �9ˆ�ъ�s�􎍸�M�fR���f���_K��?�V?t7I�>��<�
� U� f�."�V�M��*b�̴��N#��D�ˆ-��K�UvI�)�ra
�~E�"g��Y=��;:�`a�)����/����
E��I���Ө<�e+Va�!���M����ž��3�n[�%��/vc�K���`t�ɍ��q.�D�	������Nл� ��iPl�cq�|d)$�xA�'7/�B!��DS:nو���;�����<���'O��4�1^���9����MX��=h�hCx�,.��܏?E_��DP���pb&�I�
�ӊ��=��}%�X3���O�Ţ3�&��B-3!v��J�H�3L�Z௺�������(��a��q�+ynU��`��Qa���Hϛt��;y��^@a�>�0�Mز����s�W�J��=Nȇ%m"��7\�G�mf�(����SdB�b���N̽�~$7���PBL]���GN"f$��7=3{��&LFe��)�(]����z
'�-�	t�-h�#�	�Sx]*�i4zyK�Z$H�WM��|%T��7釞�Ե�,b��ⶴc�#�A��#�԰�ݏp���`��(��xyA��(�Z�}���7�sh7�_ñ��`A��5����s[������<^�4�PӒ�aa1���$y�]����v�xǽ��A)��ղ�� EJ�9uJ��EJ�����[����$ �F��J	�SD���P��Y����g=�3����:�ٲ�?�ZB��3C8�l��ũ�����ǆ�C��K��vKy�*21� /Ǐ��7^G&���>�� N��(�(�� ��+���'���OP���[n����0�x�m�3���+.^!�މ�߆s�(�CZ���%�N����c�L�]6���n�L�M�`�b�k�dS�"V�"85Opq���J&'�רO���ujSg�Ӻ7�l��Fʖ����B�Tń���4��Y�� ��?��(,�E2��P�*���j
Ho���I���2^�,,Y_�g����_k
�l����`Ɗ�hZ�
��b,���$�]݇���O
�X⦚4�:���q<f�ƫ�
伨h@e�T���[�O��'"\>�E>/)z�xVq��������;��������H���,zZ����%�#B�z�/���i�+�����l�!d�����y��@̇8=��$�q5E�[(yU��@�ę��CA���PY���E�g:�*'2����I�%':��p6�O�P79��)z7�5,���*�T6�����ƜIx�)t.^��%�veg�~23c��?e���iR)�h�>&0f`�>��k��i�{��	J�~��_�̍��oi����i��<\��ז�\-����_:����!:�p����X��F�+&���i7Z����=t��Z���P����Za�J��Z��I\4I�)��P*�ິ�Rc/.��к�"�@Ž�v� ϧ�ȄI�H%�w,D�h�>Z��"�8�y�Z�uM��6��Rؕ�B�T@���X�TF����e�-����p�1r�8�my#{v�ej)�G�lB�ɰ���e˱�;��Y�;�Cￍ���g�!^#�f!��.V�X)���CX���a��%(�1z���9���ő/0�4�t�,��ftvC����ځw~�+\�|�bmt�Y����,�(F$J��&z��85�h�>�׬����q�ڛ��F^-c�˿�_~	����������ﾋ�����S��'�`�;���'�Bttɚ	��u!��ƎH�x�1xz���8�r�)Q�h��\hL6L>�+,���-l����_�L���#�ǧ~cd7�^����>s��}��=|�kVlX�M?zV6�k;?�����������F�0qCg�:�U����\�95 ���QiM4�%E�'%Zf�vBB��+W������� ;~������}�HA�H����A,�[���� �[?��_�}���U-�� ����1z��e���c�Z¤WEEcA M#� 	��F{<�&�ylB#��]�֘�e����Nt<�=��q�8^����߿�˟oG�2�����`R
T�[����b�=w�]�B��0�s;�.�ˏDxO�r6��h6�L�T%w�Z$BdZ��A-]C��qJ��%������O���ø�����~�ß�FO{�Pp>o���X[���\�N���ޝ�=�n� Ad�|g���j
tPBH�S�i!��5���j>>�<sr�G��/�D)���{7���vA����>�n݊�B��/�Űg4��hBǭ�`�?Q��Hg6��7$�H�e��z�k��x���lԔp� A�a��ȅ�0P�	Ⱥ�x�g���� �tt�J�0�j�ډ�P�Ditm���X����#���p���p��\��T&���3��;C�'���_je��5���>��D��$t�� ��	���y�P�mt/���a�����(��)F5��#G���{x�*V�\���-��"�ZQE��+ؾu+�ډ��N&!"    IDAT̍1a�S��d��z+:gNGS� ��ju/_�G��OP>v�TAh<i�s,�tE�C9G|�l$nX{�z��`�����ْ�������w�_U%|��p?5ޥ�W�EMe�
wt&���D�)��㈞S�����_���ݻqq�~�\�7
W���$��ymק ���A��V��$4�I�"����P-�B�MAr`�^�.6���S�B6�\�8N�K�4���;� ��8P��_+Q!׋�+���)�B�t�oV
��n9��5<��;N��]�2��8�jaA���d+��w���G�i!����s��B�v���W�&t̋����qi�C�I�$�놸�e-�>��p}��kE�WE�03�H����H��S��,��vD�I1CȈ!�H"�J��W���\N_�	�tk��0KR�hM�*-�)���+���I���}��X�����ݓl�}�u��#����_����� �.إR�	�܊ׯA�̦�wӚi�#�^��p�HM��u���0�
.�#]��0�0�6��'W{ �KD�q���o��4�X[I��^k�g��g�QzM�#4"	�V��sK�����~=&S�W��A�FQ��j����dGҍ�u���= ��wB#�Kc�n���t�0MI���oG�Z�"�s-#"<F����D<L�E~�g�C��9s�0�ǈ��f�i����]�n�B�ւ�����E�75C� 6@ɿP�5��L#��bq����R�DZ�|I�0�����x�
P�[+�Q*L�?wv���k8�����;��
ʅ�4S�
��H��LZ�Փm��>����8�,�T*���9�2q-1�=�FҲM/L�G�G��V�x��I=s�R<��c���ܧ[���~���Ø:h*{h��������f��w?��[� )S���&�@F��
F��E${��_�5V|��@SGwm�;�<�+�w V)��6JnN,?�Ń?�n~�4�f!��9�ܼv�C@����cd:G�2Z�AS_O����v�\�˖`ẵ�N�QO3	�\��O>��_���+��O~��wފ�<�^z����
"��bhV}�`��M���L:[�iz&�)���s�4:�1�����k8�rZ��:.�BL��� �C�7��'��vA�>|�-��\ǃ>���7
"um�x���W��M���= ;�c�˯���-p/\A��,�)Ds�b��(!������Z�����쁀y�2�|�K�v��j���6!~�:�|�a`F�x���N����ľ��bbh�}��~���_��;p�.���?���l�`�aZ�0}��{
ḙ'���?�1V.�TPe
.�q,�5I�B{�ӂZ`�B��^���4�����w߸h�៿�3���3�mE�X@�)��'{�D�9���S̸e#����Õ��<ӢK⫞�i��	��U�j����K�T�@	&�n�+���զ� "P.�3ET�+�G�������X��ۆ*E�e~�E�ӎ�\Y���Ƙ�np���qꝷ�^�cV*�����reV�+B�S�o
���H�z}Y��r�͋�=m9�Qe�D�fmKW���o =3�;|�'Nar�^`xfmRt>�X��l��~f��	�����o�z`f��X$s�S��2A^˞�mHL���LS�`E��J�Z	�}0�a���6��p�H'����L&�|�
L''�NJ�ׄ��Ξ:��g�IN�X�v=��Z�T�t�	\<��Q�^C��UT��C���.����b!�R/B�R�Ӵ���A��iX�t��F��FP���s��.��ٳB�ioi��,Z� M��$�R���M�̹�B٩!�`V|�y���>�e�Wa��	I���`|�KP�p�Xi� VV��_��(ǀ\&��M������B ��YiX��'*m]8g
,S�2��k���+t]��,���J�a��@��."Ulȓ	
�=�}�nŵ���$.p��V:�Ui��J(��;���F�ߘ&p����|C.A�a���u�	�s�1}�����y��f�o�4U���V� Q�*�)9���M�j��i���<ϕ�`"�7�lG���zN�*>F��Q-�Hd08�d����v5����{||���&��J��ɉ	4�I�ut	�U�US�j����fL�P���_�I�m[6-��LRYJSl��8Q�3���s�����J�8b60���ť}_H�ŐB�Ⱦ��RLFTiv�!58鹳�1���L�rR��p���c3E�7�^�ĳk�ks�%J���1'E >/B��ǥ�I6�G;�M��wƾ�:���t��MA>�����}7X�����o�D��t+K�u#��(;r�J؟��Q(l��Z��%��%��c��ۣ�I_ޙl���_!�HdlU�|	���i�mJ�#]�?!�u�(��f�S#G��F創0�^�����u�����Z���]g��'��.WT]�4��,k�e���h2�h&i�F).��(�!�NK@q�a{��*�{c8���| ����@l�CM��@aB��5&��a&�gM�M�0,���af\��8�V6�j\��&��HA.E��¯�Q.$u�M�Lh�'��x���Q)�0<<������ȣP��a�Ƿ&	gR#Ye�~Ǒ��J�$MAñ(e�&3Bk*��aC+�`���"�2�]R}��:��y��O���=��c��s����/�G,�[�rB�q��=����Y�k���x�U8g/!AT�� V��5=�W����x@n���>�;/=�k�v�*M�k�
��G���<��_�oߍtW8yX�4�~�x͇����곛&��:b�Q���
M��_�%w݃���G��S8����V]$l��i��<Μ:�r��%7.�O��l{�U�޲vq
�ܚ^��!�-Zm�Z��iےI�� ׎�������2�(U���(�*�v)ꣳ�f��E>0p��q��}O<	mZ�$_<n���7,��N>�w���^G�@7��o���p/��'�<�S�nF��l]��q<̚H�a+-���օt��Dc'�cj;�VB�:V=�f�D�n!E��0�&�c�E7���[�z�Z�������v��.&�'1w�r�}�tQ$�L`��a߽�wnC��Z1d+�u�:�ZL�a)F4MCE��bPC)�I�1Ӌ9���n�F�fcZ���	�.�w{,.�N�&J�m�V���M��X8�Q�xFv@02"NI��$"3@�� �oZ���Z��|�ܮ](m��!�R��0�H���1�leO+�=4)R"A�,��H"ľ�7��ӆ%|��cL��G߭w �z�ӯ
VZ&�U�r���U���q�\ݼW�m��O�r�b�"��.�O�|��"�-P1 �4*��Ā`��9��7:�q'~.�ǨGf�Rt��`�
� ��0FE��E��C�R���7�7���IYۿ׶l�w�f�!�C,G���3,)��=%�d㧇�2�	%�g�t_��S��O�m��օZ[;J���<���Ke��*�h?{�2��f,\��s�"��H��S( 76�k��bt�:�Ed[H���c� NG��7Nb˹�P���V�֪��Ír�1º��$<�L��<��l)15��h0���x^���"�7���4z{��-d��zF&'qmr9�LL�5L���*<3���iho�P�b�� q��\D�L���,6~�\�eK�TGoAϝ�]3 �Ѯ�RQM�XH�Oݮ��E��e��#ӃR	Q�"M��� �&��sm�5���V��t�	F�4*�r��
L;&��c#C�x������Ӓّ���M6L"�he�*�X(��8�ձȯ��6� �����)w���-�-��I���*5x��Z[��׍�����h�ߏ��X�[u�&�W6'��8�u�%�ٓ�qLNN"��#��*�,��'&r�=�B	-B_��X���-Br�L ��B�mPUӐJe���e	��CO��Hi���v��b�F�o�bYM��$�]}jCW��2D@�jl���B٣ӺY�����ɇp�^D�E��P�՚��@%�P���NCj�`�,���� �G.فDO)#N��&��p�Ww����ʈ���;�u�=q�R�V.���(���tt���{��]��*�_���Ŧ`j�ʜ �Y.����@�����tQ�s1���U����2,D��g\o
��:�Ʃ�f�/��R�7��d�o����c����H������R��j�16�n�x��T�uT�sq��#i1T��P&
MLԳ����6���]7���S
�R񤲧b�h�ܡ�Sh9�������WHn��3 �Yk�g�s�����}�4���@�w����ƀ'9�-�d�Z�Xl<��p
�P�Z�"R;$�X�P�T,�q��e\<����!_���m
��e�y��QV�T�zS�׏�bڒ6�[�7�⤈��"ź�k�E(��a�w���~�8�ql�G�v�0����"�J�Ȍ�e�L�,]�y�X�ɻ������q�[ω���^5�!iH������.V<��Յ���і?����1q�<2�'��'�5�b��������~�w`�/��S�H �������H��D��B9���q#����H�0H��]��3ǎ���Kho����`vu+4K`H��K{���{����#U�!ˆ�EtA���$Z�2�[F�&̌7n�d�*�1�ՠg3R܌�\�V(_����daX(�&�;��w?�y�I$�~��ѽé� 7�P����ع��<q�o��~���S{��[��5��C�\A����Z���(��,�ŉ�u�YgϪ���+�YĊ�L�D���f �Vm����a��RO�Y�}�@S����;ph�~��tΟ��6b`�b�+�>�'�}���h<t�w�/�ӈ�ٴ�d��X�Ң��]Ҡ}��A��;6�"@S�$Iv�ZD�A���N��k��b1�z�����m��
\�&
�
'�1t�23����SK0�SY�]���G!���VKr݉خ�D�<��M�N`A�F��<�d,�`��|h�#����\�,6���v�.\�삅��i@k�RN��!�S��K�;�:5�����o/�+�����ҁ��JS�r�L�m=�G8���ZA��"� ���u\����k[���u��c�)ރ��sۭ��~+@1k���>,ǖ�-���[;������Lm݊��mh�E�F�f��o���u�N�=,h����3jɦ��+��ˆ�N��L�>��b���(��9�)��*2��ؑ��N�$U�2ע0���Q�<"ېB�1mh�&�M��-�lҢ ��~Tk��[�d��DQ'��7�r���-�\jNE��h6yԲOk��R�ĝ���[9@_K��ײ	��5��sN�US�򚥅dͅ_v$Q�9�FoGbto����d�P�Y��^7HEQ}<CC��/���;�m)+��s(��kj
q�&��n��S��S�XP�b����j�"
�)ъd[�d$5�o_D�S�Ԫ"mnkG��Y���y��Ab8�*Lbjb��	��2�%&	,����F���&]@"��Q5�F�ҨC�n�����S�f��QÞ�n��E�u��ւ��4�bk�^)g=:��,ґ�[�K!R�Sy	B*m��ӂ�C�����8)Dh�Ǆ���ҁ��陆�9�5�u-uԞj��:��&�EB��:�w����ƁI���4D���1$����uJ(w��"�	����񏶢t�"R�3��-B,4DᤀYsж�&`�<55a#B��yu�<�e<����l���%4�z��iEc��`�s=��H=��:LK�r�s��w�^��_���g=��cS�;K��3?p�}&o��H�X%@]�lÝ���\������T�h�%Vr
P�.D�d�.�e3�d
������ҀE-/Nި�xVjoQz�k�XW���-������7�_
x��Y�ס���ho��8��,>����*R=��ɡJ7e�N���D���&$�\,����C������tE���7!)7\�H�!*�tR�rőCN�&.f".�D����R�c�7��Fkk�ZڑJ�d\��J����A�1(� ��듅r���/�ܹ�6���I�牢Q�E�:�"�:� A?�*�{]-�+	9���m�ഠ5a�1ċ$J9t���Ϟ�ᢇ\������/�5�]C��C�(k����=�d'��Fq��~|��K���6dj>Rud̉(BG5���嫱�އ1��v]�>�Gb��i�_����c���ϛ�u�܆��WPɋ��C8������{��%Xn(�d������H�]��C�����q�?��ߋ�'���8�{�4,6�u�]{�H�Jn�}��[��Ⱦ��X�D�92�g>U<�&�4�K&�X�2��c^�B�$�l����֌LN�q��q�޻WRPŊ�r)�8�2�1����/�M�?�kWC���'�(�������ɖ�����Ŝ��n�޷�`���z}D�|~b���o���u+U5��u�6Gn��;�6O�в8u�dE��(�@G�a�+G3��(�5�3)T�6b}݂8U''$��X���(�Htu���S�Jn��Q��"�Аp��2���%D��*�f�Y�0%E�b�r��4�U��#��Ys�%&)�PM�y����,�����on´�Hw�P�T�TK�[�I�cN��%�;���߀w�8Z#IrY��JҔDcO^K�gI��U�1i�&��Aj&�U���!D\ב�mx_���϶"lnF���Hgq�1(Tʘ��Į����'�Vʒ���'��"�H����e���H�� �nA��#H�ZC����TP�{�����h�I���sC]��u=b�V�3����2 �r�I%�eq~�*p�F>�XD�ݾ�N42��ŗh�2�`�G����fF�w��&���v����DÕ*.���{�RxH�'{oc�y��=g_�~o���;���$E�H��hK�$;v<��N$�I A�A~�_��3A~L��'��X�[^)�%q)����ޫ��k�u�s�~����m҆�8t �h���������y�%����\\kH�X�_���3�A������!�	`LM��%W�Jz�k�b� ��r"���Y��Q�C�s��	Rǒzk��*�i�D�S���l��
�˓fN#���6��+Y�m� q��+nP�a@�Mb�-��\�E��g�E�4`ӕ,�La�')ܖ�H���u�0��4����h����pw�Q�CT�YD�=����P�`�Wy�*�l! �I�g��X�+��$�5f(��6��ݯ"HRl�G؍R�cL�zt�r!�F��L�c�&��T�ͣ@��Q�� ���Hg�.�3b�[�>l
�H��r����LG4V:��$�ƍ�3G@���=����[\w%�E�x�ˠR�E��T}�Ʀ@�$�X�G�j>�:mt���$�0�	o�:�N�s�	�ǎ�8|Z���ZOT�ǁ��p���$I���3�PhD,�e�H����P&|�{�i֝M�(�UU`F��	�+`�)�ױ����=���HI� \ga�l�"���:��[xs���
�x*����?�)hGʆ��q\�!<���5B!���t�rC�i�8�"�NT����R�v��^����{��լ��cSO����H���4��{Na�R\��X��f�D�_Mf\O9<�$p.n>L�Y����z�0���=��M���7m"����G���F֐_e��y�K�+&�q!dLP���'�����ƍB6�,�����K�hJ� spqА��Iq�i i���'xvͼ��L'��H6x��ibL�
����:�ͥ�X��X�׫�{�L�i#	y 8h7ۘ�_A	Ր�]M$&���tT&>2!����[�FX__Ǖ�W�}c[�=q��Nt��+M����ў�L���?���/�v$�ѷl�l�\�Ǧ �a���vRXY�x�be�K!    IDATo���Up��3�ү�
=z�Bu���DjS!���rbZ�]�k�~���Y�]B��J��<D)��A�&��[N����?�n�[��na����1�FK��`�S���������?���z���i���	WN!�t6`8��X3��M�O݂�?�i4�[x������b��%z�J����8��i���ؾ�ݍu�}�9l��:�^_�`9H�7&7;���0uSP�I�5��ag���p{������è�Z�z��|�%9<D]� �}zj"+,D�����\]�-<������G�q�]\x�����R�~�O��t��~��-� q�W�:<��(�$>݊SN�h�>��U�0����O�K5���r�������`��11F��NZ�#((�}��܏#�H3���,ms�0`:*��6�p�F�R�TeN���T0^�ÉKlh���)��@��)����*��Vwr���'_���a?ΐ�[�����'?��-�.(�IF'��)�w�����������{�{�,��.\��Y�}�j��#��)���%�,Ie�{�uMq7!���mP�MB��P�,4\Ol`�Q��90��8*0"�#�aA`�{J�c2`:&l������%��!��C�yD�X\r�%?��˙��1E]t���_�U �40%�Zޜ�S�A��"`��y�R��O����L�:�zUR`ݷ߀�{��:�����X�P4Iĺ�Jp≮Ti
�
�ŉ�+�Y�c3�qbZB�����4��6#�0�����L���mcm���3�a0��ư�~>E���h��r�!��%���r���k-�b9�x���	G2�=��B�TPX&D�A��\,)��N��5=&3.tdA ;�%�j��Dӭ�Y����[v�1�{�mI�'#��Bmjh�*jvEhD�ͦ �شe�L��4��&VW�y�Kh���
}�q������_����v�Q�0����7�$��(��^R{���8q�A� ɖ��^	���r���`DW�.l�F�p�Aq�E�o�L)�j�)�R<��yg�i�B3�@���|���)NK>l
f���%cO�`%(+���ǜZ+���`��j 6�V$�ace�6�Q��g]�s�|Ptb>�a c�d��Z��v�-MA0.ЛD�Rk�i�Y[�Ih��[c�+�ؿ�� Y8D<���gMNz�*:�s0�)K�:�����q$:9�|܊�f���S�3V��� c6\L�����u����i%u	B���F}VB��-�:s���{M"
C,���SY@ڜ�� ��tpd]ƽ��(�A�<�Z��pE'=�'��4�#3�K�;�D�����_�}��������<)vK���Y��i0����4,Q�L���A��t����'*�e�J�D�y�H�)�d��e/�^�t�3��CVS����Co���(=��MF
�E�]N����̤����|֌̬��d���Bf��)�9eS7��Y �G�Q��C^ ����CD�&K��4`L�dSP�@G�@����J���c��J�JJE�6�M)�յВ-�F��f��h4Z�]��BIU����I[�3�)`2/�p:�B���5\�r��t�l�=i�dR`
�C8�<T� �I�`Г�r�𽻦��ic>��Nz��,y9��<ƴa<�1�<��k8��i���z�m���C{&��N��L�	�7/c��Y��U\�k<��&R#���h�Io�(��������Ν�	Wq�����(v�ˤ���y|��sx���ŵ7�@ޟ
�En?�'i�xW���~�ZaB3mL4S�FެI�k����7��� sLj]����Ã~���i�:y�\?y
?���5,��U�
!$?��ElEzK7���6v'���m��iI^?����S[��8iHY��2I�#Ls4:s�����l��S���F�!��L�P4^��h�`g��4�+4uO�$��(׳$'��@���Ȱ�<4%�Vի��
.��<�,I���u��³��	�i�� �tz`q�{۝Nq}4�n�a��i��@qk�U��IRB$��Ae?=�tр:j�]>�6rS��4���X,;���NPpS4��@#Q�(ޱc�?��㧰r�6����!r"�{[���b��l�;k�΢%�
Ł�pA1l�JO��JlG��f����Ha'��e�Q�,�l	�sư��gehX:�:Z~E,�đH�ey�#HsL��"ƀD)�5$���Ǥ/i�VabδpȯKZ��*6,�$ ��V"��;��Ԗܤ�p�tC�qE�Rn3��kx�5�����`v����M��}�HeB4ݺ&V�N:�E�i�$�8w��ې�6I'�U>�:'1j����5n�P�b��!A6Lla >�����=�Q��0��8��]��W��.E��8!n�zp�[aZ6)iMR+b��I��2��,K&6R�
%pv�~(��* �z^���12"��6�49+x��q
C�z�A
&4,�Z�86�iJ�f;��Ǣε���R��ڢG�?�Wt���|�M'>��B>��Nt�,�`i�/>��yX8�������Ɵ<�΍��1\F��H>l
h^!SZg�l�kj��;&Փ�'	s�(����i��BM��T\����F8HBhlh���	�!i���N�W�?g,������uLQ�#�<�vU�+�~���\a�ũk���~��C�tI�d���g���J[��@j����2���Y��I^���<�|��X�N���jh��B ;��?�T���!m�q��é����^���x�G�@��?��w��ɾ�Z�u�W���lȹ0��i�2D#>��L���VS[�8�P�99���Py��eJW6
�K��0���,���"��K�e��Ɯ���u[Q�C���5	MJ��.�����M��8�L/�]��r�!�$=請8��,�}�Y�����?��?��`�?���!�?Ӗp��N1e3@kJ�Q(F�;F�0+�y0I��^"�%��P�W�L�,�_3-�,���5����7;�R�0�;5ZS!3z�_i
J.�~�r�N^}?��4�~g�$nD*9)(8~��|3<��$9� �z����ѱ�z_꾩��"UI��wlfQ6N
�P��?jR�[c!XS�Z�� ��Z�Jw�{��k�G@!Q��B�3�Z��i.qRS�n0< 
�d��zsJ�Dbv�76�cc�����{0�A�GY�I�U�")>�j��M�'���s����<45s��C�����
p��� q�!LmL`#�V���q�}����C8Tk
��ï?�����b{s;ۛ�� �t"�
n����$���Ww�԰0�8��8��#��3X>z��X��)������ml^x�o���w�Ĵׇ_ �F^1w�L����Q��I7y�;�-�r�|�O_�SyPƵӉEl$M]6?�s�	���I�`0����l��oz�$��R�p+pjU	��#\?�Cw:�
��3Y,�#����<��N-9�|�F���"���_�r�ЬKj��&�V����'�?]j���8����%[��x�m(`����5
�B���zդ��)A���2�4.�(u*�ֆ�5R�,Sq<O���;��tj���[-�5_֞%X�q:�,��5-��BG۴Q�-��� MèH0�S��x*��PROU�*�~�%��*��ňiI�8�D
�¢PI�/G���^O�(;�`�	�&��\��D����j�3P�T���tM*�mr�)��@�<��ElA�aT����$�@��
u�@�t�d���'Ƽ�_�HO�ЋiH9��}Ḝ��MNu����JӃ��"�9�8�m(Eg"����I'�Y�?ģAQ���`��PDK�x"�y�	��qA����e!�t��.<)pbh)�	\��&y��H�T�HeB`Ccc@r�FZ%�8���+��<͢S@��&&2˒U"�ԝ��#	FbNHF$2�����h,�~vu���%o���$�B�RdD�x��B]>?�OWh�˹G�E�$Bͩ0HiI�9#)4����(�)`؝�&�⺤�Yg1�����!w�F�ZS�lvw�=Yo=���
����H�&��u�0@͆$�7]mZrG���,v�~#Gl8 ��n������W~�;	b��]\��?Ee}���2�hqrK9SqQ��Di�cT�xE������'E=�|���3!�L[&q���W]��HB�4�*]���ϴu�+P�����Rה.3�Ь���,�, �4-i<�g>+���,7d�1ϔB�����j9e�i�`(qI�.�p5�(�mҫ��\Z���y��H��e�üa�QG��F8�p��6bN�N3=kg��_���e��{�}��p���T���hm.���\[�q"(�Vǖ��Ϯ��%hQ�+�9��\�<�c	mT��g���v.!��2�q�`+`�+7d���~�Ty��C��Z���iK��Ċn�ƌ��qy���,g�d���_�vbH(*� %���aJ��{><@����sw��{��[Gϼ�oRPVػ�ȸ7�o&���Qu�"s��H�m����@`��g\8U��|&��ɗ+��
Wo_�vn������k�?�"��\%`+�]~�_{]銉���D�?�d��58~�����������'ګ
l��td6��]� teB�i�@,�gM�
S��(�ՆSiX\0�=Jd���B��؊��03�4�wM��LI)�Q�Ѽɱ��7�V~�*�e��Fqj(Q�LMB8V�b�И�;�1��}��_�@���no�^��ْ�@�]e"��%�'=0����,�"��b��t�{��%C��:>��1���8A�X`�CQW�FXY]�\���vz�,aDI��d���]���˅(q���xn��!�&b��rEG����a���Y;�����es�f�@��n�+��?�"����c#��pd����DH/dN^��ƙ�E$ѫXm~R&1,���<����/�����D]�,QW�#}�@�1Ed�͝v����5���FCl����1IBA�[�,��2h���(?o���\
w"Z��$Eǫ��P�I �J�����a6�#S� dSI��!�Ϟ �i��J=k�{�3���)��T��BK	��zT�$�~A�rA��ذ��!X+4T�M��=�F��	�V=t�)v�c�,{�Z��ج�����,�s�L�$��^i*E[U7dRP�ttLm:vH���	2t�p�(�q?a$�I���c�Rs�K�,�0[<���8�B�Ȧ�4<��S|OG��fM�V&����8���x$�L|�G�J,Y��N�\�Bg��Z�����1P�E��8L�������M����/T߇������Id�2�G���r���p��hU*�s��d|N؄����\��������C�7�~[3�B����f��i$M���`��T�i.*�-�(�&CRVs��Ӷ�)��bL�,:5����'Zt̖�D�S)�8���2�Q�禤XK�$ۖ�]w4���X�d���K!��"P Zu<�~-..ˤ@>��0�b��Eo:FFD���pY�$�yƍ�f��W�E�6lg�d�g>�W�>ߙ��|7��S�cQQ�g�`�����Δ{n�AW�������4m�~Y�c\��-��2�ӀI8�9�㔣��ԧj��y�A���@����(�|i8���n����>�_�G��=@/��!��ѷ����&�W������#)�q<�T�?�A"�_��KZ��Q��uM���1�_ˇ����uw<���>�̊�=i�i4 ���<SU�!_�nG���$l�Ԗ�����эfN}�>��2-(Mhڠ\���u��ĩ�*PW0dgIϊ���Nm��v��F��RK")�eme�j�<���ǲk�Dݖ�Dͮ�7����h�	��aj�Mp��G���::�'�o�)~��g�'0�>tѻ��f�EqgT{�LTU��sP��ʆM�h�=K���ؐJ��ӄ -X��34D��}��2���%����T� �5��*u	�$G��M�)�ۂ��g�8d���rZ@�6���m���(Brj�������,ƈZ8��ch�uϻ��S���@�������A��8�Ȋ|δ��i���i�O;R��N�М	��yd�H�� 5:B�jz-GyQ�*WG=�LM'N�в_�A%�\X��1E��q�e��ɴ4e��8�@��f��]�f��6Y	�n*��o���⫈ց;:���4�L�����E��n�|�r��4���|1�P�Ĩ+v�05M/iHE��^5��=l44]��3OԲu����L�D�����q�GQ�j&����TIVh�a��ۡe��ͦyN
hMMC'pso��w@��9�I(|�-T�uA��g�r��D��˔���s*��	��������ױ�����{C&}rB��;��&%��<8�����C�zp�A'v���;sԃ�1_�d�l�SDCTm_��QDMG�l�FǋZ�"�'&�+�<O��lb�P^��E�GiGh�NV*�@
�x2�3+�����T��,0��q��Nb�I".:u_%2�J��(�)*�nn��y��i$W��E
�8�BӲ�	ɲ\� %�s,�̑�Q$661�L2�Z���ma�Q�������Qi��X6v=\��Ew<�렆�O��bS�4:͐`H1!i�|���V��q)F� �m�B[��J���j��"Ė�b[���B��`��Pln :>s�H�$�=M6��D�'(�bR�ƄOե��l�I�erX�l� +1j2z�\~ݗdR��1Ź��}JG/�d�"h\9�%J!��A�T�\\>JO����j�̹>�\U-�Ţ�ڡ��A�C�eљ(M0�S�|�D�4T(����\¤�E�\ƴ�z���1F�/�;봠%��	����Ρ�qud&��d#&/����P��Ji�Ȧ�-�D�x��u�*lIs�Aɢ�3Lǒ���vU�'&j�� ��š�bc{�ť���������<'E�nOE�۰l,i�,_�.��3 ��=6B���+�jf��Dϐ:�d�%��ds�l��ft#�0q\�D�Ѥ��%�t�FB���\��e�AMG���ôU�s6l�z�m���)��%��A� A�6�`C���Y�ZA*N��8�$�h"N
�N+�ְ�vD�$mף�;�{��b}kS�!=K��*j���]�����7��ʵ8�ǔ"5`������<j�,("����n1�Q��	��lĉ���C������*VV	}��`��._�,y8�Vq�MBXZ����#9�IE�Z�S�,`���3��a���Ff�A:���p�l�~�Q��X����/�Ʒ���[o�*L�T�e�%(T�$���V���ץ㌙�F��3I��F�acӤ�S��T`ZL9)�8���SS�ͦ�	ȾO�UN�J�,��9W����&�%�uǌ5��:4���nR�G�T�j�b�c�k �RD��؄���<Z����F� ����ĕX$2@xHp�V�G�/h�l��1��/r���Юy��*.������ˋ��������㏝�g���Fk/��_�o��yE4����P˩�O������Ҁ\�Nαa�g�O Y~R��e:M���)ݾh�m�)Wle�0��s����)4�i�#�����VD1j��y�d�$1<� y�����GIX���m�0���TS~�Z&WHFh��?<�~�Cک`퓏�y������s��'^(��巿QS��+�����b�
�������%)�j3
x\Nˋ<a�ቡ�i�k��r�:ۅ�4�3v��/�6Y[���7�EL��l��Y�ORC�a�D�OCu��������jJ}ii�'��d�@�]}_i�#�����4�s3�9#+l�O��|G���p��z�PQ��������;NX���hZ��[r���TbhZ�OMװLM�����c9�3ޓ<
s��Y�e���Yjd=R="�v^n�e�<�̬Ra�kE�{E����$�#�eR���0�<<�SP-�_���]"������{    IDATG�Q�,V)��k�A������u���'��-E���Jg񘗃2-�`��7R�X\���JV��r<��0���������"CIX�k���Nc� �V�2,�ELt�q1��!|@m����;g��Pb�E�H}c0�Wn	lL�gG�40�Rq���Z"땋�iх@	Ʌ#�bVDz�j�4Ö����,�9��K�t� -����E���i�T��|�B�Y��T��|�>9-�3i��K6*5��*"M�~0�v� {����n�IJ"��]�MQU8I���I�z�T�5�ɔ�	"�E�ut���1��,��e!��	_��>U�3��#�ϒ��<4KK�
텟-�����'&ϕ��u_G("&&D����hps��眹��ؠ���YXi��+���c�E$�O7�M�L�e#���l�4Xl��\�S��6�L��ؘ/'A� (ڦ���Q6���a�a��u/r�5	�u�:�݊/i�D��p7��9pش��6�"�,*YN&K�TB���g�t%U�s��������,�j*h�C	��b3	�4jRXa�1��mC\���b�U�w>G���:��n���U����:L����GU�4K J� y�JsKQ۫�su?�$���������Y�M�/��&*k!�\Lh �����;m��
NmS��x'�� ��]L��`�T�~�l
]ՙ���PMa���H��ћ��T��l�N����4B�yI��>(�&��{J7�>w���� 9@ƿ2:K��:�[Z���a�;y虚=p��\۸*����&�Q_���_A7�;���\�!�rd�)m�gf ^���2�(by>�:�YfSF��آj6�q��HM=����S8|�=h/�J����jEMO��h��;v�u�
v֯b�ں�|�U�h��P�X�	2p��"Òfb�֔=Ӣ{��"(���j�Ï��_�e`�
��ы���?E���er�}ףΊ���,A�b�t��)b_�����O�ǳ��Dq6]�����t� ���"`�n��t��`,�M�t�$a���-�T$5���!�P9�FO�f
��/���D�G}��c�t3�9�?WX!���aY|����f��h)��0��NB��X����1ui셦%:$�{�:�rr���э-8�!:q�V�`>���&Xjב��m����҆��zL7M���~��G�]��o�%^��߇>�ˌ���y��@�/���3��@��x�Q��ͅ��)?�R�a���X�S<Ϻ������^(���Tv�t�w��|W9���S~Z�{�g3Z��X����U20�t̳=��#�l�ݒƝ{q��M��ɔO��Kt ܓS�#�ƕ��{E�������^4���u��'���t������D�oJ��ڜO?C���?�����E�_{�Ƿ���mL~5��uvע}`)���*�-h>�!:��ub:� �R�	�+3�<�x��`<��UP�&�,�Vu�b1��Z��x����&ů&�i�e9\
Q�5i�yWG�(�Gc�Q"\@L6m�rN���X&Z.st)B�v,G�m;c���Nɉ%/UBt�D�7v�#�mC�L�%��L�1�d��i���֒kQH�0w2Nd�&�Hڀ�c<!����D�&��P�N:H�*hb�(hk�)WB�,�*�F����Pm��Z��J]�;-���3'���1���u��8�0	7�t��9�A?u�O��S9=�AW7)h
��`:��B�r��lc���R����z3tǻ	�����M.��A��'�&�a��E]߿A��R�ʦU�R��{��R�s��5���� ����b�n�P	-��=_�ci����E�k!:��7ֱ?�#�ea�ME��9�Ut��ΐ��NUZc����	�9�~!��X5	���]k`k<�^� /�K3I�1��[��h/�b�=/���VS��Y��z{{b�p�t��MF2��Wđj΄�FQ6K���KaW��T�X�$��-y�������y�����;�h��3�3��c�p�К��4juE_��t	q�>��&iv�����C���T��I6B�І�<|�\�V�0L���ّ��)X�h)�t��H�K숡k�K��ԯ#l��/,��[������X�&r:���$T6�B�(�0��@�����pcO<��4[("Z,�{�c+R��0	/�E�j�(2.S2�����O�%���q�`�*~�<�i� ��<��������-w����Y\��H�x�q�qo�� ��v.���?����0�5CGU�<��:ZD�e�[rtIM��hE�#��J��,��^A���+Ԕ�%���׌�a��ܩ[q�����auVa�t���t��+E���?Dxp���Wp��ױ��;H�z��C,X:"�2U<����C�R�	��V9b��T7���0|w|��c��x�{x���!�q��!X�yT[(4�H�T�\���;�ܗ-�FH� 9��� [��mIpm\���U.�lY�^M��i��)f&8ع�qw_i0\�r$9���XES�lKD~Bl
D�&)M 8sJ|�}f� n��>�&Si
������h�/ð\��FA$k����Կ�la��a�ᷛ����X�0�~'����I�PH�o����~o���I�e�<M����������b�O��<��y,?�ǟ�
�z�F���x�_��X=���a8�s�u��ѐ�����9>&ÉP�igΦ�l�&,��� ��NN�T�#Y�b��p�� q0T�Ͱ8��OM�h6�|&��Z�M[���^�ayaA�	a@�L(��f�f�P�6��[[��5�:�琟O�#�f�p�k�R�P7�(z#���������)�;��~��?�~�;�~*���O�['���������7^Xy��W�ˍ��1�|�y�Z��Ƃ��3\g��q2��sL%�X����) /��Z�\�D@�]��%�P:��1�x�DFfI�E��?b8R�_��n�J�v��'BJ�v:�O�4Hӈ�90X(���؟k1���[X�VP�l85f���q0��ca�B�)�d�D2)0CMuT�����)޻�R6��R���g�1k
z3����_�|)�#h�>�O��d��rf�	�QCsa�WU�c %b5��Ý����H�,V��K��y�BUӄ�NdTo�Q�.&i��l�zġ4��� *�cW������:��2�����a��h�,��l�ʡ�CXl�����cw�:�d�A8�zo;��X�q?̠�!|@�xDGрx=t�`�!C�r�>�9�+"�%YP�q��p�E� Uä`�B7G?L�jM�	�:/c�z���C�`����u��}9,���e�PoÃL���M�h�͂��j�J�c�� ֢r��ؓm�j��x���|X&���a��f�g�،b�s�О���������X�!Nd�cl����ɥ!H� �~;�q�����!������.;�3��	��y3oy�px#�/�̈́��AG.>�����Y�POε�aH�u��>�z�TW����p]_�V���a~F򘈚��L��>.��6�;�������?a�o�q$��"��6�NE�v9-p�\(yb�H�`�%�,�ś��+�YB��q��a���1���[o��I�ܼ�Q�*en
Mƣ�8��~KK"d�1�
��/`��]���/�j�R�LtǕ���d���S�2��!���0�Ep�G�8�p��Q4���Q#r|x����C�ⶇ���@{A��'����_��5�lT�=ȇ%���F��9���s�v�=��Բu�aH=d���KG&lJ�ɦL~�\'�_�{�\�&��dZ�ncw0����9~V�?��Oc�λ���e��*l�(0e�f[R��F���:���{\��7�7�������PIb�,�R&�f��Tt]L���J��L5l�$N|�k��;�^���b������>� 0�
4��Ddn<DQʠ+�Q3�ٔi��x�O7���[o�څsТ	\�a���7���VV`�:��M�mIML@[�&���,6.|�,�����By]�H����̒��@�Q�02�Ѩ �]g���<��S	�X�/.��z/��̭��U2{"�������1GN��5��&L�� Z�+� �2�UD^i���c���0z�m�n�a!	ᇻг �V`/�q-�0h�P��.,�}N�� �k'o�0�������`�����a��i���a�w��&mH�6�iD���8�Flo����F�.vn�#��Q�T�F��KKj_΋$bt��I���-� a�ib S,�{-�Mߓ�)���"߅mU`[Uؚ.t�A}a�%,;���%�q����D�HSL�h�Ɯ/�n{x�[����������҃��̣������q֏?m
>λ���گ��;k_�׿�/^��+O�Ӏ�Dx�'<_ߧX�S�	_�7r!0{�46,t
��ZV	$���>�T|�r�׉�ѻڴA�·�r��@^_�ד�Rj�a���p������KcX׊ƨ$SI�4�H�^��7d��b�HFZvs�6=��@}e	f��@'�	�or���70>�"� ���x<����#�D2�K��~RZs�-T	��Y��E!��;��p�X6!��L���a�^z�%���"*m4��h���Hr�����i��Cw}�h�E�B-�`�(0���)��Ukb�����\��g�4U<����j9!Z�?�w#i��x��)�l�9_��܉�X��$���4e>�z��}���0ھ.�t�Ȑma��E�\��lwI�O�_�e�ŋjg�p,�`9���l�H��j
���ϟp�lA�����$:ߞǩ3O`��{p��;�e�(g%��\:	�[{$6���)�&8����g�{����Y7�aǱLld�6���w�s�z^FVx�%�AݲŪ�¢�v�00��0�=\Kb\e���
�y�	�x�!4�|WhW�I�鈉�4߼ͶX�y�#�_��w�ƥ�����h�h)R	}r�F���9�������uY�qĆ�"Wrˉl���#"ȵ&М���}��<�w�A^F��e/h�j±��?ˀE$��N^`���+o������o��l��4Dՠ�!t5��
]8�tu�U��;5#���=�3�g�:\��ش0jw�=
�����Ѽ�8�!&��00O0&"��^�Е�re~G�����$�@���������6��1�'����X܂t����1LG���6iK�)�i�o&*fC@�)r�Ǻ��Sw��/�"��9���c�F4dx&�A"��NE��h�`9,U#OF��a:���ɵ+8����՗ѻp~6�Bœb�t2Yo����k���t�Q�6H4M�|ez���L�3�݉O|��d�aaIh�CJ���:)� �^`�����R��*�4�����?���;��ʫ��2�ⶶ%A�ak��U���@��Mth�Z�`S�/����c�g�,� ���{����˸�����3@g��@j!!'T�k�����%Y
CLp�����c��y�Z�V��SAZ�'N�ȩ[Q]X��|��+���q�՗�֫/"�G�m�7a:�4<g���'�Bi1D�E�
j�c#)�J`;��*m��4ΚTLm��u:�Qm,��ӟ�m�?�S�"��S�B��#\�p	��}T5��1���~�u��)/C&W�~5�P���c�ҫ�}�y���Oz@�������0B���#c�3O¸��YTi���RdϿ���-������s���*��6�P%��*.�;N='#t��p��YܸzU&:�W/`w�*֎������5�,����p:<�����o��c�����S���eY���6�7��%��MF��#+k��W�-���c��u�z����Ṷ.��� Բ��-B$b~�f��R���?�K����|��Q��|��X=��{��o��������o��?m
��[�������9��������?x�}���UKD���w��P��=iJ���/�F�ze��X1T@�Xorq�'�`(}�-���E\�%ј1�S�3Ŏ�v�KڡX�#&�9���p�8!����)�Qn��@(t�Z8y�6���ðu���vZ��B$O�ny���w0����Ɔ$_�pq�- =);Q�q)c>���W�FA�K��l�J7�YH�D�vL�NT��`�T�0C�YX8y��&�������PF�1����>�`��֡�V��,���x������"��B3MP�2��(����vI/	C%6�J�(bL
#$(����W�ud:�QR��S�p�SO�O?oqQ��뛸tႌt���K���+x���i���'�ѻ����e���s��֛����~W�=��{�i1��h���HwQ�W�o3Q����*N�{)R8V����0
"�i�K�ø�O��_�e臏�h����⥳��<��4�{��X?���NW�'����Uq����[x�G/`��7�v���r�,6w�d���Dؠ=��\T��@���n��#Vo f2�[��na#��6Vz�;���#؍'b�����OBY���<6az��e�C|�������y�}�.��tЅ�fB1h��0E"\D��zR�<���9�k�x��<�����z�����G~���ԟB��O��lr~�.6j!�3;��D�i�����=�~pg_����<&�Q�T�p#�d�
�L���,j'>��'���~��T����S�"?u+��<�G��#�`���R��y"{�\s�˵�Fci
��E�Ӏ]#��W\��l��k�1z�e\��p��Xf�OZ	�٢���aK&����i����������r_ �2-����9��>�5����d��"�	�ݗ6��.f�ݺ����^�l��e!�|�=�]���?���ob޵�ɇ����Q�J�~�ڝ�X��_� ��Ie�'nA�K�c��3�N����#O�<p�|λ�PlP�T�2u�t.��� Z��t5UB�#(��ѻ|/�����_D���պ��� {���L�$�֨aY�$<��au��~͟}h�{}�����x��}�A4?�L
"���	��\���Hő�>�Q�=>Mtwn`{}]���g��xͪ��\�o�n�q���8r�]�v���h,�E�^�4�����|I4D��°i���D���t�	)5l"���'��r��2 ���CK�R\\:o	߈.N��SHb��������ȭ�"�+9q�*�'*��t���6�on
uةxbQΰ0Nx-<��g*�c��%�V��I��FϽ���}����H�����R��V���0��p�Zށ����� ~�<�����q��;����<u15x4��5`���s���N�f���+x��ױq�";;�n_G����>��|�i���pk"��c:�Ε�ؼ�>�lS�e��:�d�A�"��-��醸r:2�5�(L�x�8��~j�G �-S�	��ob��T*.�K��,.�#͌�ft��"k�B�Q/h� �{�(���\��Q�5�8s�:���N�WƉ����i����Ӧ����z�G?Z����_����ַ�� ����J��J�.���0r�3x�+�u�.YF�J;-Snb"�a��B����88�ݫA�>�o�*j](%2�u0�s��P$H�m0Fӯ`�Y��� �t(D&�=S
���jHӭJ�r�C��ة�a�U���k��L
�,�F]Bt�q��h;���{ﾅs?z^}[�'�R0�a����"M]D�2m�*q�V^�"�&Үƍ̮��eY>6�t����n�#_zw}�� 0�%f�'%���u\߼�
*�G��Шaues�*�/,I�i���1�p�� �;�1.=�=8�`��4���ŵdH1˂P���_\��t0���}+��;!��h`���p��Ob�{a�upasׯ���s��{��8s��W���y�����N�8�{�M��to^{g_|�kWmoÜNP���"�ҒV�n�Q!A��*�d�@�����-T��    IDAT�v�Ũ�����_���G��	��=Y���l��G��zd�V��b:����������s��&S� ��+�x�\� �d�ȨcUt�2DQ9��]U�x���P7,�Wr#��@G�I�#���t�v�9��1L�5�DS��pj�ZZ��U�Q��N�.��1���QLGB!k ���M�8�6�]T�q��%���HiML+^��Z�G���Ͽc�`&R��׎���Ƨ��"�5�3�b}kW��:��+��T�Ž� �(Dխ`qn�F&y�Y��� �h��=�]���^��H�f����Ɯa�e�" ���*V�@4�q��!�L����14>q�G� �܆q�c�`������$E�y�u*��}䕮�S66�	U��zJ�LQ�$ΟG����{�U��-4�>�u	����B��:_ �$�>�r#d` u�}�:z����Sx�羆;�����-���(��ڱ\	��t:;�=r=���8E���F!M÷L	�_ƅ翇����0�r�)�*�A��1�F���HEμr�����;�0�CN�:������/|ͣ�bG��L�d��X:|
,�B���#�;�$��4
l���<N�+2���ҋ�ѿ�Cl��'h�!�v3#N""e��!��Ja���5��%T~�kX��W o	�q��������v,<���#��UL��N�!�>³��Q�2�	�#lo�c����^��,��ݬ�Ѯ���h.���۰|�$,��S�m��p�I��x�G/��?�(�JS�38-��1�[�X�<���<�g+�Y����YR:T��˙-�HJB�#�E�������O�s�VD����
>MaD�h��5!5F2ũ7[��5i
���!�I��j�@�{š�)M���/b�;���X6s�.�}~R�m���?��/>�y;�Z1,T2Zw���?�������#����W���S���L�f�!ba����iL8v�����w���oc��U�]�;R��g��O}���Jt.�bEl�w^F<كVPt��Tވ�O���bf	eC�f�z�7XX:v
G�z ��adyqlcx��`w�7.�03TM�t�%0�6�dA�9�&�8G%�`C���{�}U7��`큇�������m������//�Ӧ���ϯ{������_~����׿�ߏ&��.��뭖�� �H�E�Kڏp�x�a@��.��,!eT��mf	�<PX�s���e9��]Pa>jlM�qLĦ|�(��x��X�ka�3QI����aZ�G"�MLi�h{�=��?�3x��O!5�x��EAǽV�����}O��Z1y���|�vvq�'��ҫ/��+/�K8�����[�� QXL*j)�A&��V���8��E�a@\�����/��ß��_�"n���*6v�1�3%O���q��{�X<��@*�f���k��X8�����.�o��o��\C�����D���~Lb���3�����I�5Q��p0b��ٵ�q�'�ࡧ���m���x�s7n�������C*C���s�4��F���Q;�`�9�����G`��^8�׾����&���,r����By(��P�dI�l�N�LR�	8�-���B,�����e���WQ,����>��*@��b�/4��$[&���s�a2�"i��h�lB����	�y������0�tN8A�2�Tx�|�p(��cF�>�A18ͱ�t]��*t�� w��/�>v��2�<ۆ���
H��/�.c~u�FC�-�?]��I��6�Q<���&ƽ}�MK�����g��o���4D�c�T��JX�e��ӕ_��Ҡ�>�Q�(��.��#X}���_Ƹ�������P�^��6�UO�C��!BK�8�G�-��HX߼�8cq��K.�����7q��]0���byK �-˖<tW��D=�.W, ��瘘9�ʃb�� �܅If�zw,E���fî�p|���!F,`�j긞	v�P%�2��V�
 �.��g���󨏺��J(���$4d�
��!�Z�q�^In��D �	wq���C?�s����5L�������lYD�j]K�J��C�*z��"=�A�1*z�J����g�����m,@G�D6�2�P�fv^�H ����?q^�X7г\��~��������8A/,Pk/��7�f���n(F�X1�S�D���و�!����'��U}xLw��x���w��D�.�����ɧK25��y]�2L���u��&�?�U�}�k@}'��{����z�	��'=��A;Y�xt8z�TϑjD)�!U#t77�y�*��]FgE�٪�֨��:X:r�n�K��
�1�N;u7�h&�4�{�����}�� ��Al	y`2�d���*�Ss�3��e&�|f�@��|J����<������1�zߣ�#��pmE�%jMw�8�hD�4�Q_��Z��AA�'{1A�}�f�+KRN��g8 ^{����%�v�	�x(�
=�l�?���O��@��ovX����~��B1��-�=�է����Łk�܀ZK�Y����CE�׮\��H�,S���� ���|��x�'Q[\EaՄ)�GҖw�ཷ_D��ҧ���	���lҦɠP*dŒ�D��"7}t�ڭ��j�`<��$6������&�h��\�HJh �-ەf�5)�Y�^ʍ }0�s�����x	N>��N?8t��p������x�~�|<����W�����W����?]Z���0-L�^�\�#V�DI(:6|�����^1r�i����ʩsn����$J��(�Ҥݝ���c,���}c��0`��6��^o���ɣ,��H3���(1��s���T��~UG{`_ɀU��n�������y�'�c��6Aچ��(�jvU�"R�6�Cʑ���oPS����l����/+N;$Im`W+�Z�$�+���S	$�"iCEf��(����r� |�Mwޅ����>�$z��K�e2�Η$$�@�ZE<�H�ʭT@3�n&>�!?9�ӯ�7NEm�:�b:�:��i��	/��4����:��J�t�(6�U��@â���#����1�s7�0Ŋ�Ԥp��x2�x"Fz���zMx��qCd"d�m�*�W�Aow/Pn�|����.�������P锡Q��BP
=�Fy��4l�ˬ#�@#7�I�8-�5e+�m~�x����Q(bn��ٕU�t��r�G_o7���+IFJK,��?�|�2ff��߃��F�K�n�ڑ#8���?rX^B{S�?�J�b ��,pR0�|�y�`�y@�i6f�-4�Y����b�݇��r�^,�5��S.ۍ,�F�GO��FMuK��T��"|G�xh�+�x�m���=�uyMD���S	��kE3a�L%+_�Z(��� �cm�0N����G���F�\.�I�V,ӅlOo;�)�t6#����*`��j�
��	 H��y6n c��9sW��G�PD�G�UQ�{��'(Դ��ߠ}��gQϮ,�P��Շ��q�Ͼ����Xt��b��3�$S��.�4s����$O�q���*��:f�q���a�� �^�gN����5�ϜD�0�t˅M�w��PHo�7A����-;N�y��(wu#طc~��@4�k�
-E��K8pÆxO�.�rT�Cʣx�iZ���I�_d���'`�m��懧�K]<�.z[u��*��T�Ùf�#�b�X��?�3���B�@�L�Cz�N����w߃�FS +�a�B���3i'�!Kx��I�K��)!b`��T,�32�g�����ϝG�RD���*�fM\�h+�B�]R���BcR'��= OW�t���:����
U����5��4ҙn�,�E3���j�V^�vQ�N���CQd
��ײ�F����_�'o����,C��(/� ]���L��8��"~���3����5\y�7���F�o���=�FPu�h�<��2�t
�m����^a��UW�������<ʅEx�z��0Z����$�o܎xn F$%E'�$qX"(`���k�����_D���t�dS�}e魲X�s]�{�B*�|��꿣��y�k& �R������B{%�l6�6b��=�ӽ0�YD�Y�ј�h	ڤ��P�RAr�x�	(H�a�Qqʑ�H	�d��)D<��NN�C��w1���p��:��i5�!�
[(9:�]qt�s'��{�N�b)ԛ��m�������~���|�At=����|�C�VB�!"���+X�[�����e��,�p��Ih���'ž��C�{ .4}�H��/\��3��-O#�h�%�	uL�Cv�h��RL�Hge�7��o���.��nT]��5	�)����bQ]]i	�c0,O/�k���&�ʺ�� ��ɥ*�<��y���;�bxߞ�9���[�]�Ӵ���_��/�QO��GYo���7~��O��̥k;�q	n�NLF��x�=;]�������X��r'����wz�K��."c�,Z�����xx����nv�$4���c���K�Zi��X��EAeU܇�zV�a#*����$��=�w�jGpuyV<���Qt����B�΁��S�f���&-*Dq��R~U
�l2���^� _�Û8��˸t�X�R!0�����<�u.d�}�P�����D+��
Mqj)�Br�f���m_{ �^��l
B4�#���Z�uv�(�a)�L[�Ubѩ��&>�	j5�����8���X9wZ�ֶ��ሚbB�ƫ\��YRh�v���=�
l��L�~{��"�㸒_���ҴZ�����(쨍X<"�d)N6ɣ�C��08n�r�jUy�1l_�Tč#���k��'o���WC�h�a���g��3VҴ�ђ�QF��>l'�{�4�=����؝��o}G���]G��@__���bP�]�ڇ��&~��n���(W�VX���VQ�~s���ￃ���fe�C�&�2�v�u��J�����P΅C�����{�w۝XI'qri3�"��G12<���n��t��vxQ�h��w^2i>��2��4�\\��(b��i|��_#r�:r��k��4^���Y�K /�CE��X��57M����<D�oo��=��K5_�{*KF��I� ~v�zQAfwXr<T��F����K�.�=3Н�`"�TƩ߽��/>��	��8L�B�FLw0� g۰�) -�{��1�&jF��2�?��w]�h�:�.��%D)�5��Ȧ�.6�eN���%P{D[s�b�ڨ�H�1�MɊ�ȕE4O��қ��Z���^F*n��(�"X�D]�o5T$W�斨��4�]}�������#���KK�8v,VY��5+7�v�UG{��k����B[9�T�5�I���Б-�q�՗q����r�Z��р��Ě���:�zf�Qg/�,���#�m`��ɿ��Ǿ���c�Ҁ�IS��h�Uה:2%�n�*5�� #S+��X�V�k�ڞ�Ek���G�Ɠ?�w�2ZC&H!�eM�x��E��8	�)D�=��o��Iqtapٕ�O�jc{w��?7C��,ܷ��	��̢�Z^Can�7PX��P����[@*i��'��cd�&7�F"7݉�5"D��Ħ�^�����k/�Z�C*�FZ&�~Y���De�t܈��;��3�!u�:��LT�n�{C��h
�	�N3�P@���Ll�'��N��%%��M8	ޔ3�E���J��z�MP@Ma2=�U�B�c�HӇ���q������[�H�H����5PH���{���~`�6�"t�� ��5L?�.��[dM��B���o݌e
"FL &�s��G�\Ei���J�K��U_�x���Ï<�]��B$݃��Zr^��i\:�>��k���a#���ם�*�l�(��챡i�пn����A��L&5s�>VE䗗�2���b��
�.9+�^Ğ"�?�,���S��̻�40y�6�۰F&�k���i�:U`|	��@��pѿȧ\:{6�w?���������4���Ww*#��,dl;"��C�/wRM�C���9�kw��|"�����1-�4S���3
ک�Bb����,~Y�V�U�X�ږt�wR+-���"�5�u4\R\,��{`d��@� ��$]��lD��4��USi�m[1��UV�r�`Ja�RE�Z�SO<�Va���N���ΝA��#Iy�B�j�-r!K!��E�3Z^ �"uՖ���n{�q8�f*�E߃��w3���]$#�B�m-;�"�c�.�e�t��Դ� �B�բ𮻝(���p�ŧp��WИ��" �bh' �0�(���M�>�cd�O�B�Ѐ���=��.��S���8�&'6b��8�j�C(Jf��6b�i�p��Ht{<�r����cuu�x;׍�\[��7��+����*�t����N������v�LYf�>��a)��#�78�[p��W~�=��o��hbhx@��;S����w�U��8�/��
'�%�ѣѭ@�����9|���P�x�jQ\�$y� W3����fa�I�/�n��UE�p���c��#��V�1\,��ulغ�=C�R�S��N���/RN$�c!ȥ��] ������U��Fr)�n\�+���?�H!/�7]	m}	���,x�I�f�Yp��5_�B���~����%��ߎ�3���b��uŁK	��`��	�t�� �����	y����%i6�"6z�q�f���ϟ��������HPCL\A���E��-D�G��6�O�cz��X/�m��{�Q�[7Ë%QgV�E���h�
�-8�'J�5R"X���p/���tw%0�^HZM�RD�J;��� ���a�B�co#�XA:&>��-�T[>VHY�i)��V*,�}�?t'��ɿAn���8��5w6ա��	9�\RIin�@n5�>'I��.�b�,�<�N��n2s�x���O�~��[CFRkh��H�"'3s[҈`�ꅨ&R�ڲw��_�o�n���hf��Is98��U;��f��5(oA��,3�!O�I�&�O�'�̈��������\�ë�ă�R�D}�8H�Lq����@;t �����y����x�Ct��bݾ�h�z�`fC��BѡUp�����e\�x�s���
q��d�36�	6�A4�XQɶ�xFIԺJ�6o��uy�(��@��d�],Iyl���L$��&�I�MG���~ ��N6� ��]��y������ظ� �D7|-
͎�2�I��ϗu˩E��P�0>����q�*U�!�F
B�;��n��;���s/����\�#���&�1��.��п�^`��@��I���1�����w� g41z�6dy֎�Xipa�Ҙ<c�m4����Mյ2*�JkT�y�,L�D�Ľ܍M��B������Y�	
�O��0Z5��Iゟ�t��A��2���v���п~4'�������|����9D}�9quW��}pS�_&[�TǱ�~�k��"�&��ه��<gt����Ѵ��Y'��\_��/����{��G�o����杷��_��j*u$�����n�v9!���ɩv�ړ�}{,̃���X���e���R�D�����6x<Иl̎2�Z��R�"!GV,�]؝+��Q����y�ܖ� ��ة6�U�#�Yl��6��؀��n	���*I��t�Xh1>�e�HS����H�@�T���<"z��D�+�p�������!�[��]�8�'(�N(9�S��3���o!;hx�3�h8	l<t�w�Z6���K��z�˸��BҨ��&�R(�B��	D�JdY1�K��y�B�"�p��ec쉲X2���;x��Ob��1ěu�ۼsR�D�-��6����j����ѧE�e�{�^������8�8-���}��;(��:����0��W�����{K�)�d!h�a[(U�������vL��`<���'�ڏ�ųg��V��<n�^)��S*�Χgz0�`c�oǑ���S���{d�\����"���N����u�i�!    IDAT3'4"Uv�-	(��ju�:Q/¡���4����p���,���BQ������
�� �H�q����q��=��#��N�ɥ�����cG�����.��vȅV��]���q(�ĀN"��Њ+���g0���h^��4m�@lYy��������Td�C]:ua�&�y �|��	\/����C
��������xo	G@�]��'7��C��1���O̅(1�V�`6��a��_��_���g`4�H��t	��Q�0�F(�Ť��1%0M��Lx�#H����B��_B�"�}0�(T����F.�c�!LH�Y���/j#��w��8(�JB1	]�z�!#
�*������/@����ӑim����&\����I�eG����������ķ�
�-��R�}�l:6��^NY���mzI'����r�*���D��̠�c?�1���2��Yt�.��Be=���T�q2G���Xj��1y�װ�Y �CX�z��Q��Lz�#��:H�c��^�
���z�~p�3��^E�RV���$Ҏ-�s���{8����ԑ\X�Pa�e�.�Dڌ I���B�w7&��/���*���Q|��Qd��0v�>��)4mGt�v�ʉ���4ȭ��˘��PS��2,�)�,���W%�v��fLl�%Ŷ��Y��P��;��X��Ƈo����u��О���LQ�Շgj�S��?+�n~����[�E��*P@�h1�ۼ����e�iE`<�9%aɁȄ�\,���-b}�r*#�6��)��8����IA R@�����w�/����a��@D�B3|���r�Bs4��Gn�Zߌ�p�gWg����8��/�*X�'��x�Ν�6��#y6�d��|��1���\@���XDiyQ@A1?��lw�{�9���
t3ӈ�w�(.]��s��z	�Q��7���ئαYұ����76��8��bp|�����E��ç�d(@�t�3Ӱ���Hf�d��ӢÕ�kf"9')6�8���p��_#s����=�?�G7�O��5������T_��/����{�������?_��>�7�JEI��/� �);�����E��K�0E�tq�5������wbv����Å-+�#ٮ�ј����*���7��tX����&E�c�@=0�9I����0�����-[p��ate���L�Y5B� _�cOFed�(Du��`���|?ߗC p���-#�ν�2�N��^��
(�f�<(��`QAF���i��Z��*�����Ǝ�E�v���ۡA�Si$�!h{M3�&Ǵt^���d�Ka�<\��HOJ�����R�K�� S=�f�����f��=�����"��No&mA:��&E ߇,��X�y�$��p�c�l݆K�5�V˘ؾ�B��n�R��$Nz���Ӑ�U�]n�<�حdq"Ţc�!�Ģ��K�g������s� �v�j	��B��p��λ)B�}V4T�����Ƈ���o�	ܾ!����Y���<�,�T��AL	�R��g[��(:��Ǵ���y��O�����s8��oP��p�m�C
��`������|��ioAtё)��ͻ��ڀ�ذp���n5��)� �dG���`��߻���ٽ��!8���b��� ��X=wǞ��>>�D��Oz���8�m�#�.9�P�)jvZ�v�Ǯǿ#b7���DDP.]���3�.�%Q��渁S*)�4�&]Q�dC{�"�*%��z�i�"QΟ�ٟ=����@kmZl`��8ud>I2��c��ҎU���F�t+�`d+��#{�X�E�9]=0�)���e�D�J�d�R�LR.�Ͳ�|I�o n+8cC���|1�|� �	�A��h:�����B��q��qeh��Y�(�jXgRq�&qk�6*��}�	L~ ���P�M�L�M�ҍ�>��ZY79���v����e�7��cjp�
�`.�k`�wp�7�@��)�X�6K�EMP���
�Erc�z�V�6c�c���{D-��JɅI�4�nC��#�MT���h1����*$ˣ������ �R��U����.$(Vj�����ß����<(��yh�}�,Y+��Xa����w��ە��ٓ�p�DrY��ٍj2+��]}60�8%E9&�'Nxn�
�X�0���2*�<�fE�C��PYg���۱a���t�i=��E,�9]"+���ñ߿&� ny���X��?���Yi��U�鏧+��~���5��bZ�.����j�6���-{�rRpC�õ���I����B�ה�\<���i8��D:$E�B֑�b�,��/���{��UGD���|˗��=����B��n`d������M ����|o?�=��5L܃����kj��!)��[�1�/QZZ�Tf���W�$ٻV^A<����b۲h2T�z.������+玠��	,�����Й��.C<�yU��#��!@3h��d04���w(X+y�4H�����������!E=[$�3��5��@�C�r>�+�x�i���~ ��������_5�����7��+P�e]�/�y���_<u���>�i{M��2��:���",ȸ�0}��z��m��\44�ewE��Mvi�����.��XT6�6EA��d<*�F��.y(I���X�(�I�.CE���Z�#p�0�G�۶a� ���݇]`jjJ����ݠ*>:˒��O`�!;�<���jY-�^XɣY������-,��{��O?��������rة����[]�x-e�@�H�{�N����:4�i�Nm@�+-^��y�x����L��.�m�MidiBs�S
�B���\S7Tӓ��b(��Y[�闟�ٗ�F��ǈT���O�"'�mqC�h�خ��1k���2��m��o�9��-��)�d��s/6o�* �E�� �X0	
�cM=�L4$?��I���,\	29�˹�)P�P�����?c��t���	�j*"���BVW�re3���B�����71x�0��8*0ЕFW6s�J�ɦڡ4
L)����10P�����b;_�	 7o��I��x�N>��}�b�RLf�N*Z�i�%k��7r��n*���N�z��&ħ6 76
Oh=w����
�N�'� q펝�PE�-���8��:zrI��&�4�?|�1���a�,#��U2�@M��R6"�k�@���t�Z�Xw�>�z�OaM�j��$R��k�
=t��S\q�?K^7C�:D;5�cN���
��%Tٌp=��1�I7˯��?��g�`�StG!ftq� /�0�!m�H�� �FЕ郵�vt�u/b�v`���0Lh�`;(WjH��E�H:�g���ivK�5B��A��*��4Wؙ�¾G�r�O ƴ�O?����
�#�"S/c0����(z��f�D_P=�]���}��/�
�B��Oŀa��8V��2	����d�fB;�s�Ƚ�����ZX�[�2��֍J�{����G���ȹu荢�7AW��EV���u���#H�؍]����U#�|�	��ݶ#NnN��JN�mk4nޟ?�8eM+��weu	n�E<�@wW���̛��;?�G�3���d�Z:�*uɬP�[=�=n����&������>�KǎBK%0�c��A��jq�(i���7�:<�&����G%�:�%�F+�E��S[wb��}�c]�(B�j���sm�0:������Q\���݄��>��MNT��D?)&��И�b����ѭ����Lto
�Gw�
F�v!��Z�x���ml�u�C������"�I!�`8GlB!�x��
DI:�f_y��bu8:]�\���5��j_
#? ������ ݚZ6?\�����x�?'��<c�v�͘L
he��N
�,�s�@y��F�"6��eT+�����u��n���4<=z��o N햯��O��8�H8���@9.*����\��d�V&0<���A�t�P��at
�6?{]lg���
�V�A^;ؐ̀���܏����ıg�R���a➽?t�����g6��Z.W��/�S}�+P������6oL\<���gΟ���f���－��DH��o��Cq|��0;��Y+|�"(�q&}� �"�k���ɩm��m�G�Q�C�¨�e���&|��2�p�(П�o][w�^�y�]�^oڈ�-��E`sdki�$"�Nw-�bJހ& �=g�9����V�(2ʹዥ&�iF���7C�������o���)X՚�����NX����z9�=9�C3��T�9�lۇ��}(3�`�$&wm��M�:��'��E	� ]&h!ɂ�C���(�~W:"n�C��#�n%��f����ǵwނ�VBJ�ON{��x����6�s�0lT�Ou�g��{�8�Z���Y���p���```@�Cv����x�r�Ș��k�9(��XY\�Hwo��\��:���|��ӈߘC���#v���KA 'V1��K�CQ�ѵy�݋��VcYx����r��MN6GᲩ��-�nP��_�v)t&o�颲X@�PF�^ �p4Dk�^x�E�K���Jg���Z�W���C�L��B`�P���u�g�~t�~�b��#�~Z6�@G�P�0��h{:��kF��ǐ7�F"ŵ\rC�i>���⢈K�FC�}��,�����s�}��/_Bҭ��h1�H�683���&FM�%(fz��1r��`���aFKe�.����L1�`��s�.�xl�h�ض揥۹�-v�<,��P��������|g~�K���@0s�q�;N��m��%�l�2Y�`�����w>���{Q�%0zh1�=�DhXh��b�K3��n�HG1�e��ET*�<ݤ�P�r��V���5n�X9Z������˿{�R��.�!���f����Az^��Z!�H���C�_bd�]p#94�H���#��)��F�I�A�2�	��t3���kֱ0=/�3��P?l=@8sG�#�{�y�X�",�&�E�YP�x	�	%��LT�Id�Ė�?��}w��G�/6���L���,[�$��Wg߿y��q�[t���B�R�����
��F�����Kￅw���.]�0��jY��֔$�~N
��{�0�?���Hç��;���I�z�1�{�I�5'�2Af·~+PP��RC�I��5	���ex�5�]��$b�ظm/�hN,I)�g3�ܝ�G@ْp0�c{�T�f(@]4FbP ^�
Ԥ@}杽���@�Z�

:���\f�ڔ���Ɲٰ�C��MQ�"�rw�h

ꍚ���I��-',�9g��18��=��W_G��DQ���2�]�C���y�~D�~��"��A`������w~�X�5�߷}�=}�6T����7(�\u�����2�媜���U��~	�����ƭ�d�XIiԑ������\�����[	
㤀{���&���M��^M��І�Нn��p��Q�M��C��BIJgH�+�P�s�Q2H������T`�^�p���1��3��
��#����ƿ�sC���[��Jȯ@��u����]�z����W�M[[B��������Z!}��6t=�cIO����,� ��KG�r)$G´"��F����UH-l�@&�ar�Q�������ђ�#2�f��R3Dd|c�B)ӅU3��۱q�nq��K��Y���%M��Kn��GΠ�)�����``my	�ss�j�%4[�Q��rn/���b���VV��%&����S�����<�Һ��?�̶}����Kch�6L�KP�۬ j�Ȧٹ��%��)�ءkW�j��N�T%��V��z����h�� |L��>~�'8��3�א����GƢ�URv?�)���0#(��T#��Az�a,;	T#�l�S�h���N&L)U��P-K	A��4ڬU%߂>�&V��8;'4 +� Ց�F��8��sx��?�y�*z�5Ф6�5��8��	�P��2X+����{߼��$��qD{�a>ҩ��&����MA�eZ�B�[���BĂ�ݙ]�^��y�@b��h�6},~�6N>�+X���_�w,]GI��&��
p�h��"�9���{����Շ��	d֏�]����$���r_ޜf���>� qn�`[�L6nܸ�����]�G"g"�0���x�N���k�2�hi3���R�C��5�C���Xw�Èm�c`�\�]}�uɟH�B�PRc~�\�mko�mR���Bhw�lGD��LV�V���P�]oW7Rn7�|�~���7�1��Ҕ����-G�H>r�����Ȉ۴ه�Ν�aٯ��bF"�Lo����U��#��e��S��*�2j6��,�kF&ͶP��1;��|���|4�.[C�Yŕ����G���A���k�XiԱ��Ī���&�Q��v=���߅X�8t=�Z݇i�+>.bO��	 P��V�X��sk��;Xp4,�-�T���S6�@o*,���_�'����e	���>�+;`�O.7�u8e��R%����Fz�AL��u����Z�"�����R0̮�&�,B�v3�3�=�s��@p��3�����E�2�bwL������?�=�gN`�nx��aӎ�L!���T7��d}C��6�3
���+��x]��0y`?��Xav� ����w9)���jZ[VQY]E�H��Uq�)�`[���`Flزw�'V4!{�kb�2 1����x�-�+sH9��U��"��VKiY�ͯm��=��ǭ�া����k��=��ɦP?Ó;��q��8b��Z8e@PP�n��0ڠ�E]��s�������XQD<���1���xTi
P��4DJ&P�M`������a�{�tM�@DK��GG��?���26܃�G��}+*:��Q����䒔tl�Cc��VE��B�
�\�� ��-;�bh���n��4͇��D��\�tk�gdR@P���9�% VBc�-��,w2���G�iL���P�(Z4�
uVˋ��3���$"�Ҟ��&)�lvq��Jx'-I�k>N��,f�{�Vº;va�pƦ�Q����H�.o>�W��˺�_���׮��8s�{˟���UZ��4����Q�<�D�).:��/��m��4DK(+\<���ϳ����BE��r�X���mM��dL�)2�z.��=�5Q�1p�6}�$ƾJZ��f���>\�?ۍ�;�i�6�qq�HY�$J�E�\�.�Mq����0�t���-Ȇx��%�\.פ;4��0� ~�"�O|��4�t�4�Ng��Ό`�QBvת\�#S��s;�����rش� r���ᵍ�4��i�)�L�)��m�P��[%+:'�k��_�ՙ�v�˄W��7ib4���ŇO��O���*���IkL؜�(�vR��PG�T��a��&v���"�nDBz�f���%��������ۮS���[�>d%�Z6UU�b(P~v��3(��p�:r�1L�eq��7��O�D��i�Z�Lޥ�� ��)�]�,���yıv� �̳q'���B�2SihZ],'%���4$�=���c+�?>��]�iX�����%����]w1V?z^|����E��0�\q��`/����&;��bj0�G1|�0���zF��܀�����@o�[8��������R ��'T�8�R[���<�\�&��#H�؈�%䏾�7��Q;s]����e�4S��@�T�0}��TcI4G1|����<�F�ɞA����IQx��L�e�Jf�@ho��擋�d�r�ތ����-�������bI��^����~�S���G���<�Ű�4���1�!bt�Xv,x�"��"y�n�x5\\Z��NH������E��cm��,� 
��D���"��Ŷg9�z�Z���dD�qD�1t;r��_|�/<���4�fsnha�^A�:WMM�ƕ��JԆ66��}��ݲ��)d2�[&3��h5�����n!��
��yϊ*����E��    IDATXx���XXXBh���F�
��Vq���̋�!���dX�c�cLk]�,_�R�&���24��5Al�m���70z�=�)5Q�q
kI��;�h��#?iv��=|�HV�,�eV!�!)΁f�*��Օ���v� 	q�7p�����S�\�j�S��u4t'�a�_��o>��� ���q���p��i�l�,��E)���z�dۤ��� f1��u����&>��	�kE���YP*�#��W�j|�fLm����X�Ugg���V��,k���z���;4kHGx�U���������j��3Ǧσ��`�L�Ln�+�:A���V�o�=��J
}H>#��R�5�覦 ��H�)���hCH��*��J��M�aU�9��W^Ax�cI��X���d�P�ۑ|���V���mY�[	��Ƒ����~���uL�߅�G�1�n*�J`B;Q�W*a�4��,�T�%���|N�����l߄э[�� ��p}�wf�za3WO������
=��u7݇�s��W�T�9�f ^f�S��G���F��	hQ�N�-��V�
���R��S0L��C������#M�Rp`}�{�9̾��g�}�Edݦ��]c�^K�|�%�W��˺�_�����͝=�O�>��]YA�pgΣ���RCy-�c�����\��j��ږj�92���@��H���tD��iyg��p'�	<b�D͈�5���נc���
�4��b��;q���#�رc��MD�i��4���mPp��ȼy��o(�6t�J�~�	���T(�V\E�b}�����1w�7�#�sM)P�i:)A(��LjV��V�vߎz�(*����E���A'���	�:�8VdA�����U"<��*��MP�@�j��Ρ����$vy�J��3�X�����ȟ:�X�G��՟mӎ�֡��u�#&��A׮�hnF%�C��	OLH�y�9tD"*Rp�!��&��dD$�9���8�������I�m�'�ݛ�a��Q���G����\$8�Y����΢���,2|��50���n�3���)�6N��(��9�|�.5�h�o߲�>
��
B�M�bffe���iyȢ�湓��ҳp�|��h���E�"��jI���PaN��:�ێ��8r6"5�׭�vL���=�s(Q�^���7���79i{��T+M����k(���@�ãx����� �MD$7��PD��w9Ʀ���z"sr�kr+�l?��cH$�r��q�3qq[	�oc��ތ�P�ZR�*P �cŢi(,�1���
Sj)�k�bM���8���P��r�'4�6�Z&za�ײՔ�xձ�NmE��� s�0�Uk��8����^D�1����#�Ts�j@��[�nu�S�$(���Τ�L�`�
�q�������o_�̳�(���$�m�X�ױ�7Qg~�I]��_s˃6:����C�����F�H�H���=�C�Wж�B��MO��w����m��Fw�ե<��V`�"���I±�_��_���<��y$��4(�&�B�,ſԑ��<� ��^d�ݎ]���w��B-D�Az'�$u�)ɆQ�6����4;0+�@%�yfJ���Dee�+E$��e�"̽��[8���w�4}N���7��,�^�D����|#?
dG�|W�}7Ο��֭X`� �5ރ����-]}�($�!���5\<s��U�z���q�򊸩Mlچ���!��P��:�m\���'5�����T��Hڞ��"�@7�t�Q��N����־|�s��[�EZ!����\u�+���}�ܾ_
c���=��o�pR�q
|�Tv$3����p�n�@�r�M�j�����+/���59�CФ������ޛDr�^�����ꞎH�V� '����~���em���c�ڼa�e_����f�x�F�l�X�[��$M��F��i��M[�02�	f*߈KN�_��L_:�f�"fC,I�.*&�˶k!WQ�lP�/s;�D�atj�L
4;�j��@5�hXB{�B~Y���N\ėΈJ���AA�e(8���~�9�Z	������}��7�P������U+~5)����������s������Gʫp�`��ԯ�H"$7{�^�C0��@�pc ��W\u���In	�Ph;rƴ����yܒ�p�;/�tR	�[�5���1A4�Q����s=Hmݍ��q�H��ئ���� j�&���l�Se�VPpˤ@�96(�.]�\\��)����/�Q\]D\k`�'�¥����fg%�(^gW��L2rf�,)Rd�8h�2�H�3}�ATr���Ә��6�{��qL��RbӪ��u帣�J������Xe�>�v�V�UĒi$�6r���'�����	��}���􁈼g&�:m�*�����������؋j��R]ܲ��ɡE��l2-��"t�v�%��̓7�C��Z�X-T�1���4�22صc
��G���	�Ǐ�;��c����!v��n�jYpƧлs/��-�o؆���r��WV�}�"/�|�Ʊ�?[nj�W�Ϯ��l/��13���:��:"N��[Bx�.�����=��G?D��5��bj�G���	�lG��Cp���Y����Huw�V+��Sw�|��{{(�̝��mm��J0���aq~׮���J}9��C,D���ÿ|uZ��*)X�웵d��"Y@�X GD6n�W}|̡u�]͊Ij'M(�6(�`1-<�v��߂�AՁ=L����mˋ+�[^�$?�C��B���T.C74�@�n�5}�3�D�b^?�Z̆;�	��Gם_��Z���&0�⿡�!�Ri���5䤡Cq!R�,�������$�}��X^Y���2�	G"�-� ��^���!�8�^��?{C@A>�0�Q��&\�C����][���C,;
��4��N'#}�m�,:�Ϲeu��[�+ۂq6:L�O�au�Ev
�])D[M�Wq�׿§o�suI�6�b�)�G��
�s"��B,�u!�g?�=�-��=�O�Z��ڈ4��Ƣ�e�)P��G�U�~fA$�� G�E]L�XE2�/Y514q��7�a�B�v�I^4]����i��n����3,p�gq���ٲ�oGk`��I��.��25_@'��뢼��O?����e!�
������¢LIڶ� ��~�����\���r
�{�YZ����Da�*bF�� (�&�U�5��\m{a��[@���1Pp�AL�9��k٘ڱ[�V���3�D�)�*�UxAA�R�	-A��ġG���hV��sR�Ĥ��u"H5]���x���Ob��V��u]�zu�@�/����H~ ��ۀd
���F�����q���OP��}��w�aķoE��E%��4*���t*7��=Y[\E}��j�i�U�YP�����
�>������>�QXč�'(Ы�4�c�D{���~���u׶�nO
B=.����]2�)KN"ʢ���ڊ ʾ�n�Y��	
hM�a�⾉H���}7~����;va��~Xc�@A��\"�|��@��u�����F�/|���g�VWМ��>F��"Z�z�&�AwCNh�Aa���%�/�1��|��r�<��h�a�H�6p<ۘ�`��Фդ��3���f%K�j�,S���F�����zw�kdٮ.�9�ϥD�&U�r�u�v5��˾E�Ǯ3EF�7�133�b����jML�FQ�|g_}��<�@@S��'(�HD%T�<��;���H�܇R�U���{В.w�ӝQ�Ba�SG��)OY���S�y
&GS�a�ve��*R��L�T�U�Q9����O���i8%NtH�x&���:��|r̈́O�Ez�mh�o@�I�{b}�������E2GXw�;�$�v�:B�v�u�c�p��'�P�b�^���ׯ���00���M�X>�.����Q9s
٦�8��-�[�g�-��K�A<���F$7�5���{�Y��_\vt��T�8d��@�v��@��������*nܘA�oYp�&2^�=)x��#�Bo�s0cZ�ĚL�$(P�
�j��#�� �]��'ѿq�}B�"��Nw��Ӯ67K�Y:�g3y/ӧ]X=�QWP*Ր�J`��t;!V�~����p?9�X�[�+��D�e+�16AD������ݎԎ���߄h�Zf�jS4��,�X\�5�I���p��ͮ���o��R����<WVE���T|�S}�=�~��(_:�n��9�v7���6��-�PG�I�Q���B���,���C4�D���lV
���~�39�L�ؑ�.�a5}����4I]wCe7�/t�\��*�L^�/�v���������_E*��t���t��Z�4;�и��_C�6ab�Hm݋��$����#pN	����������>�.����czzVܝ���Ұ�&
'��ܳOc��{����	Lg�M�c��i�+n\��Ն����-[����1v�^T"I,����t�B:�B"E�.+Jƭ��[:ܷ�<�".e�+�{̀�ɹ����$�Y���_���ڵKD �\�R��.��8b�8��4����o��U1��˸x�8z''���;��u>�S�,25m	(����5�h��X��C�PB�Z�����x�@��& ����̀�ڜ0x	��wgp��7P�O(ठ
BRPG��H�SW���t��[�筓���9e
[�v����M;�m�=HtI�1]�,+��Om�1A�C���,ˁ�0���!��}+(� c;Hс��9L���'�a@�a,�չPӁJ.l�@�����A�Erv�\�Z����|R4C['��� ����g{P7�p�t�ak�L
H*�X�Y@~qY�:]�8!Y�G�^���:i��a�6֌(���r�WO��r~cE@A"��e4��>$��L?;#��Ѧ�J�ol3�6��A�A�j*�a2���riM��{(�a�%�X�)�l�Y���g ^j��+/��[Oˤ@@�����}��ۯ@�\ �������s�M���߉V���]U��O��V�!(P���e"f�0�8i�b�͌��#I1��+�(������E�h#Avv�Y�.<
��n�z�����<�j�P"{h����;�������@�g }CC���!�K�v�!Shձ"m�����	�ZN��Ce("����9�"��n�
eR��xg_})	 ڀ��'�r��)�G�H<�FŊ"�}[v(h&3߶��~�%tww	8�W�Ӫ׫Jx������Z��� ��@��D&�Cw:�3(|�*>��ϐ?qN�E4�������#�䛞O
<|�E��!�{�p�/U�гON`�D
�T�|l5��N8�M0���0�֢��n��#
�+��>���9���2�19��c���o~���ӈ�*H�J���"Q�K�p��֙��߸	�m{�ߊ��V8RT���:����{�X���L�9�R{�}����&٤���,�Vl�Ǚ`�A~$H0�3�dd� � A��� �x��vd˒,�&i�ŝ�}���nխ����{�r(#���.Z$���~���{���&&$]w��sT�|�y��O}^t38��q]&�P�{������#�y���o�D-a`ٮv�{N�y��A*�b��`P��-Σ���P���:����C��[�F��4C�8�s�8���mn����$��s��X sm�D&�D
VWW��j�����������D���aS@���7K�Rh@�P�LM~�Ә>{��>g�a$�q�1�'��]/�P��G� �cM t6��B��먁���!����a��D�Sp4SZ��'��������s�2 1bS �uEC�
���]S�pv�3/`�{��A}��P�z�rU��Z��j�:�|*@A�hCax"(ѱ�,�F�k���6�;;�=l�~�j`&�~�m4���6��Y���h1:�TR �%���cj
�gϡz�YT��;{@�i��"�:�R��7#7��+4�����D����h4�����<_�B�x��x�7?G��E��̇83��{�S��h�T�0BX����O�Ǟo�mjM&�3\J���+Yb�+�%��Ɨ�h,�F�1"Ry�i��%��q
B�bΆ���՟�7���al�`�f��a(�uT�UJ%�NQ���ܳ8����4}��{�\���fq��o3�؎�	f��Dn&�)���tG��P�2߇�m����^g咉0�0���#l�3�Z�)H���L"�$�C�˷��6P��~�i�/?;�
�y���暡]��ݢ�����}���=��)�ty?6�p�8N>�m�')`�m�	xBJ&)/���O���J��|��[��-8��D7��2��k6�ٵ+X��;.}�z�6h�L������t���/�t���Iql��h������/�T�-{OF��g��{����.,�$T/�0��a�i��B?d����2�A
��;��6p��a?�$�s{�X(�f���jz��.��u��<64��hE,`V"���G�4]��S��/���s�k��C�TA������o�C��)pJE�犩�nS@j%
-�)(�S����c����BM��NKS��9�/1�����c��u��Yo}���K�c������5��?��ի�n"i�d���ō����-�vN
"�t��.��!�{xI�B�XNMR0,��(�'����xz���$zQ�������4f�z�^�.�=����3X8��;eV�v~�s�+0v��#�����k�8(�z}ܻ{�kh�w:�.984Y�ƥwp����o�Bߎ�{��?%N%�L�W2R<�8E���@��I�Ǧ#̡#�[��'۵06QϽ��DW�!�9/J�q�#/������q��
�8Eu�����*��Z���_�ҏ�ᵻp��L�mݔ"���$A��0�^6��0�䳘�5|�x���}p��1�U�P���\Ҝ��(F3A�	��KwY�Ɨ�Ut����%H����,���$N-�`�o�?�cķo�ʄ\���) ��B�5[l�a����s0��@:6��4	�\G��R���R���a��#E��A�u�E�,�4�b��r�[�*.jUz�F����?ǽ�ސ"��1�[E5�`�6~�L�es`���:��	�R�0���<jӳ�Mq�����F(i�3_ڧ���7��@�Bڧ����jH!�®^+`����U<~�g�ʀ��`CX��H���6��H��!R���45+� SO>cq	^�klF8]�����8a�=j�7�a�s�I��έZ�����f�nq�C�B����&V�S����W��_�@�����jSu��6�(d�[�v�,����Ȏ�Ɲ�@�^Ȇ�H����Rt�k�b	����Wcy !)C�`"�U�24�T�(D������:i�y����bϠ��G�B���p�-L�L�XE/L�F&9C���Pu:���V��`������Ax�)SP�D��Hp�ڐ�҉vCٵ#�^�+
�~-����4�u�.�P6�p���Ƈ�D����6�p a��%�j��!eC�5��|���ػc'���_E��h�:�Q>%%�IΤ�Y�U�{ٹ��� u7_҈��A�O�1��a[(	ܾ�+����	���B@x0�퐡\,��V�e��<����B?rV����>�g�xF��S���%���v��Y�H��`�#��a�'M�E����h�VP+[H
$X�s �����@����D�1fS��]e���ħｉ���j����,�G�!6{��pr��h0-æ_�Kޥ��&Y��|�1�&��sZ"=l
������� ��T�DB������9�z2���)�%h,��I��CZES$�f;$�g��/|��~��MT��B�Y�(u�T���0�x�{ I�"H��06���.����!�ܑ���|8r �N �h�^6�    IDAT(�� � �8���ow��n���D���vc+n��^�S���~��T65�Pպ�ܿ���{0I��Uئ.�\K��$�҇�p�G�vez	s��[����;�.fm}q���K�5�V���Q�M]��Bh~��'C��[o`�ݟ ���?{�u��6�J������]#��7�����ͯ�n?�m߾�_�ܽ�GD
v����&�VG�ֹo�0��D�T�#��p�� !���,�x���䠈W+�r�l
55qՐ�^�#��PK
BSE`����X��P�10L�U��:���|�����fqKRhO�.�0�� ����IS0*Xei���e���m���[c������q,U4�z�/�y�}h���1t��dr�0 &�D�tĉ�S@�Kp�
G�CݳA�*S���EY��Q���v�^�_�1I���_p}�`����Ȱ�j���&8��똬PTB�Wp��?�������^�Z��->U]>N�yȇb�F�	mi	�O=�3����-\]~�Bu�O=��)���Z�*�^�͋?]�Σ�^�9we��m�|��������&LX�á��?�K\��?���,�w6���!��-G
��6��7@[S�/,I>���0�Ze$���%�T��RW@acJq����W����s�b���N;[m):�j��7�?����X~�m�+׉�t핦@w]��P��K�SDע=�`�
��'���a ����8������8&��W��������n��(J./�?�����b���Vu1Q5Ѿ}	+o���w߁�X����HJ�>����!'�@)�P�Lϡt���0��W�@V��R�E  @߿��(hj�2\Z]2�dgd<*~6#�~�@2����?�����(A��1�Ѹ���#�}̰�-�UY��d��d()&M6}�5W<�{�tmD�`�w~�^�rB�a���2��@�Zm��f!���L���h�$��L�'��t����%^ �3������*:�~���u�>�:�4�+t�;Y���`������CD���g0v�9L=�<
���Smx� !�3�Ltl
�+���H�#-/ �DЦ�	�D]Xd��eS`ۆ$�o_���o����0�P���#MϚ�鈀وG����3�jj
��#b[|�W�3K�	��L@H���2a���1e��6���/��9�����(��
��&~�+��ś�_�1hB��N��a���Ӕ��Ϝ��?��a�z�?���}���"s]�e`v;I�����&�x��4
��7����h`smJ�32F�������0C������:�Rm�]�f�r�YaS����GX���:������3��8wi��QS �WB��n�'v����]��_�)��W��Ët�9|'�z	��E��еM�I�!fD_6��0��`���2R/�)0r�=����g6��*��&��{�O?Eecer�
��i@��س��y�\�x3�.�`m������J��(={�ϝ��� h���T~�Eld���r����}l�-M�����s�"�5�;w�~绘�w�₩8LN� Ýuܿ�9��2Jv���"�Vжe����
�w�vc�æ�H��}�Q��Ïh�HS�����vS 墉j���)H����Ψ)��H$M��(F
lO��;oa���0��̓G���S0��L��/�����\"~�r�4�����_��l�ۏ>����+���5�d�1W���h
��(0f^ y�#M�$/`WD!��<��*�k�F}Dqʊ
�n%q�S��:4EH��C�x����Kai:�����r��~�5�c3���D��X<pӋ�(T�(VKpY܎�NĪ���)� �X�����\_�q��3��V2��3�93��?���}�h�k0y(m��ZB�;��\��!�����uT��{��}��s���f06� �|VK��Dn��ܦ�P.�XX�%:���'�#%����l�Qc�c�^�`���
�h]�W������{0]���ڏ�M����80f�BA_ՠ�L�~�)<��>�|r��q���š��p4K,M��jlFE�d�609�i(k+����R��������ށ�e�p4Lfn��/��ޛ(56a�#X�/)~�Z5w�-7/tڑ�!Q0��. �݃��'P'�bf������#Z�;i�ϼЮ����.�a�1㯑���u�^���M�������~�?��?|�VS�N%�(C��P.J�U�����;Ȓ �U8��c��WP9r��Z�­V������!�M�@6�4Bd��[">|�x�3�i��#�|���8�,�5˟��_���/>���AIݵ!���-�}:T�U���`VH gv��^���v�±I�Tթ�0�l%��U+Ћ&26����-iw�8e� S���H!H_��L]L�����6/��CM7�0(MQD�B�a�.�<\��0�0�R4��~�����e�K"�M���G���[D�Z�3H!b^	=�wpV@LTg�N!�?��o�xC�a 3�Q!�eu���h~�1��e��D����RH���}��!b~��.<�fg�R���W1~�)�U�G�P*����I#b�#)Gg��#�$�{�<k�[����04��@��ۿx�{��2J�����cRo�%C������T@�%���b	���GO���7�L�c��2��V�sS	��"��/�6d|4ڻQ�b�Mr؉�RS�1x�@���x���ĕ7�+��
�n��w����%��ip��l�p��2��O��?�GP�|���u\~�H,G�{��CG(Q|�T��#�E�z�������:�=e���46�Z5%����9,<���,�B�� d�ύό�6��Go�����UT��D�rQ+	4�И�@��Ȭcw���H�����n�y�Ï��Gh�.}�A�X���A�:�"��KV� ��ʖ�M
��B9��G� ŲH#%��5 ���:�uM��L�?�͟���?�X{%������"�hs���w��[��|H��S۾���7~������i���>�S?x��� �A2Вy<y�%�*"�~ ��Gs{��6��M�>��ns��-�Й'P���]N[��!����&���ҙY�S��:��e��L��9
�1�� �x��4��=GQ�/ J���r7�r Z-�(�s�A[4�A�t!��w-IU?����BM��Ƈo na��Q�?}��C��=�����k.��>�\�mV.}����\���޶��=���K�>XE�
��v�f�� v�!��+�m81.��do@^eĨmL�O����my 	�QT�	�	ĬNm��]%C/
�S,�㠩������A��9\X����Gyr���������X%J���IrjN�%8�y@S`�X硿�`k{ۃ6f�<1;�l�.���лq��GԤw5'c��<�*�$�3���&&E��,��tbk�m2�U�ƪ(�]Tke8�|-rX��]R�s'!2Hs���>6��H�� ʎ��j���ʇ������뗐vzB�b�D>i�kb���>l��ݧE=�����?�pg��ǭ.�<�������̅��X��9uL�S��^�����~#�I9�i��Rzg���9v>���/@__Cax'��B]��)��|� B4ma?�}G�x�%�=�"2݁�ER�KQ���.H:�x�>4�2)6���)e�w��1�����43E�ğl�q��l.��{o��[oap�J}n����,S����I�t�Աv�޼��`����Ss(?�ï|��Ax��شpϘ�\��j1GԄ�4q�H:w�����I+�҈���1���l�����
���S	[˖@k�P��|B��zv[�\g�ɳ���%EX��p��<i.'�a�S�� �,?�kG;J������֒��<{	-�"�~�L�S�*�ĝ&L-��˸����^���2ҁ��f�NT8���f��)(���"R5��91z|��*�O���?�wП]��'2��PS.]̂H���`UK����)S�Ք�ky���~�g2$J���Ür��A���js��*���ݿ��CG����y��觉��A2�f(�L���B���M�+���＆P5�Z�Ba�\�i��t�~f����2��D
�0�Q4~~D�Z�-�Y�=�5�"ݼ�n��&vn\��m���3�/��s<2w���h&��(�G�75���ZF:7�c��� (ֱ���֖�.��0�`�:\Á�蒻!�i����.��E$��?�T�#Z~�k！�/>F�� F{����%��VP48v�ᢡhp�ā�����j�������{Hu��E����a$n4�Ŭ	&ʻ�즎DW+�M	�l7��}�?��~gccdJ�ؔ�Ʊ����9ǭ�%4���C�::f����E|�Ώ�m����Y�a�Sd��
�Dx'p���%<���&����݆AqD"�;^���<�}����,|�F?�� !Zy�V�`��a]e>��P�|�8�yԞ1s���a�
��lÛ7q����`��=�J$��}]�U'�q�w��W_�����&l6�����9~���(�M���O��o����g �
d�4�_�4���}I`&ʿ���^sJ0D�o��].�.��(�� �����{wnI�
�Vƫ1�6��;;0R:����>&�:ຒ�\�������{05��UBѸ#o4U�{�"J<?-�����%�*|�x?IH&i�^��jC�U�
n}��As�Nc��3��-��{�c�0����S�A
~S+�5�n�-;kW/�'��W��;h���2�.]F��c�;](P` --S%�z�l���8#�x��#�(&�M�-/6ƪUL�ב��t��������XR���@A�
=�]=��ǁL���i�hp�����g���/�ep����>�;�{�'�R,�*�����d$ʋ�D&�����r��	{��`��as{�A��p�`�y���3���B*�`�eȉ��5=�W9u�N�A�k~��P=�$�����X��Q�B�^����J%�$��3�hoǃ/�F�BR/�qc�SV��9�IQ��5��[���ob��7нw�0��������%��	��ϐ��5����_���/#��qo��<�ɩ=�%i]��y�.�W��\q���'-�(D������B1U�P�t8�n|���z�?Cx�&�f�<�%��v��#*�����t���[B69/M�������P*u�t=l�v�R�>��-Sx�p��#�$����4:�D>|ϓ� K\��� �D���ᡦhݸ��ｇ�������'�\ȥ�j�8���fj�Y~��G��"�3P5	�3����~3g�A\�Z��r�	�T���l]C��a�9��"t��Dg��b��i{2�(�}���Dv��PG!�w�n��:��.�ln���P�=��<fC&�R�,�w����ur��^�9���
P�������s�鞢i04U�݅�-���о�>�q�!�c��\.#���v:D)��_�{���/>A|�6�~G�F,�)��:�y�&)���,fYj�!C!\��c�_��sO�Z7��Ԁi�Q�m]ZK���D N�1X�h�P�	����d �Q�^@�P�`��р����%���n�Q4�� ���H��1 v�}���4�f,JS�ش��ÛC��q������;�М�0��|���ܔdYM��|��i���$VqyS%�$}A�������c��E$[�H�,���C��������q���S��,�x��9��Ͻ��S@q^l`�	��8(a�E;i
H;���01=�9�I��T����^+��
��}���;0�۰�m�t�	��5SD�Ӂf�b:�R8{b�����-�t0��*���C�'^x��<:i�N?�y�t-"�`6�et�1�6�76t��r�Z۫��HR�щ�\����B�6	M��&�P�1�m����?����'���/����=�Y�|�D"��C��g`p�v�2C6�9��;���H_��;� v}g�{GϞ�U�F�:�b�./q�#�u�{}1<0Y��Zg��U��0��z豨fc�騛6�,�k����9�/|�q���D��2��1�R¡�~�����IDJALJ�����߾���_�'���uS����/�p���D��@��X��p�Cg��^��Ag���= �;�RO\s�o��ȑ���:�s���8�g�|Y���g����� 5�@�h��D�()̱j�{e���e�#�G�h�dkTkc�9$�o�Ya�Y&�gW���J�|���h���֛o`����bߓO`��OA߻�u����4_s�������\����_�����n,�q�:�"n��3Tf��3� 49��B0��X�b��T8�!�*
ĭ�Tt������pÈtM�C< �0UU5M�%�,C��Ч-)��Mۜ��O�z�f�}�g�����.crv���5	Y��;�%�'�b�.\%NQ�k2�y,cC�Q*��v	�J
�&\��V>�[�~�tc?��VKFA�?����0�TG�Dݱ)苋��<#EUTǭ�-D��reL��z���5���(Gn���m�H�!|:����Uhj�b:�����O?��w��O?E����Oڢ�V����dJK�ݢf�BB��ચ��Z�~�4���;�<��0��'�A�\���p4n��U�<�eS,ͿW�&�$ؾ��g��IRF�a�u��u�s�x�xw� [_���P`�$�_��>�M,�.Ե��.�R��"�O?�/�
��Q��=<�jHd��²`plW����	DQ �6�R.�0�ғ��pf��- h���ZkR�l}��{�`6�(
��-���(��80��E��>BҘTR� �pz� ���_�����	�b�V��S�N����e�Lg��/ ��Kf"�2���8:�Jz���E��������?���?D!b����bR6�\P:Όr
�� ��\~�*�J	��$�N����^A��	�t=ز'�L�@2I���,b8m���q�R%	L%EQKPJ|ě��r�3���C�ܾ{k�lz��������n�v�I�.?_�{b��w*�W67���{�y`i	[
�M�v�[uD��'����4����d3W����g�@�H�r9��M��� EN��7�ݼ��>Fx�&ꡏ���"R	��P4�)r���}��w�`2I%�|�<�,�fq�{����oA�9��.��C�)�N��+�mݴ��%��dRH�~C�!��לDH�{p[W.�y�2|�	;8''�M,)s
� ���@��8�!h2r�㰃�����+�P��0s�I��y��N	݄"[U�a���1hg)M-'�l���v�� S�k�Uхhe�/]@��Ut�^E�ڀ�`RO�~��'�[�
%T
E����n�iXp��`�w��ē������>��s�8���.��a}?kNNn����M�hE�*z����47���6����Sт�D�\��i��9���:��U����+��&�|�.\�JЅ���4�g��lD�Xd�<fqO4���v�M�.U��4�~���A�9ew�t����>������3��֧��4��=��þ��'��h[�>d�dE�!Z	M�h1�UZ�jH�^��?�3l}�)�� 5�����&u��e����2�w�}�V��pcC����y?���([�+���_��'O��� 0щT�	��F�ъ$�zrJ��zj32��v�*9�H���t�13�ۍ���	<v�^��o�}�ỿĽ�WP=�m�q����'���{�B�M��Falq���ӓ0��S���[:Tג�@�@���L��<�S��+�c���isDl���/��օO`�=�4���4�w�o1=���i
�>V�_�Ϝek���������[跬lm��W.�#i�������2�1��x��j��G    IDAT6�� �82�9qF%M��x�BcXI"�b|2:�X(ɡ�+�h��\� K��"Ney��*Z�*��:����}�Ńf�;jUq��k�v���tI�9W�����1F�ۗP.~�Q"\���e����V��u�\�у��7�a3�ͼ	`o��
���e(��H3��T����Xgy�,�{}���.T���R�"�vo&����2ř@B�X�$
"?@�BYrƫ4RR"��`�;Bz������"�[�����ɩ3/r�Y� L%�r�#��"fa��s�AL?��^x��Ch�n>Z�׍Q+U1+��*�ckB7�	(����H�=���\�L=�!�����KX��	|�!��M�;}�~
W3g,l����r4Gɵ",�X��m����n!�M�z��=�
��9��ab��G�� <���8}���Cz��{�ns�ʦ �6��̃��6L-FEK5WѺs�?C��`m%?F��sHA|�r�X�	�c��a��W*��� ���Ӱ������b񹗀�C�
�l�`�����$j�Z�z����3���It��y#�h��hm7���l�E����]����Rd�X�C�	����Ma�%=�p��|^�,���B���,&N?���������"�z!:�����,)�iM�E�P%�'A�%�	��5�B�I���ؾu	�.b��5x+Q�P@��m�t!nf�fEۤ��	"�4�J&�AX�B��ӰOB�g^��5A"�����j�mG>;z��z'5�~��Ҟu]P�"2X=�݇�_����_ Y~�q%CY磔ȄT1��v<��ڈRfX��� �6�љIL�>����;����`��C��Ű-"AB��-�EM
�\w�I����{mt<B��Mto�B���l{����_6�t�k�|�̡M����c\6Lc��{a�g�`��Y�{�岸�>D��׎�2�YCD?s�N"�%�6�6�����C]{�`�1T�-@��@)-2#�^(K6�v-��8�����t�x������'p���������3�@�q�k�k� @������돰���߇���J�Ip����YLL�	_I5�+AV<Ͻ�&�}��[a$>
,2Sb.���Q�ܩ/�q
��n���8���y�_����(^�w�(�e����y�tKGNb��Jc�i�f#�fe�Лt6�H�)�0]�j��;�s9񈞅��.�S�`p�".��'h0c&
P�iH��ӡ���:�b^x	^�>��O ��Ȅ���|�~��A���R-�����	D�`#�����D�+�8-o��E��3��P������D��X�j�����t�vI����$�>"M������B����}�!b&�kԱ��X�'�aM�B+��*�IS0�<QQ��LW�4�fD':�o�RR��p��c����Hh�aw���G�7�um�{���;e�ޟc���}�S�5�_�M���Խ��q{M3^y��˗��o��V"�B�p�֒�]z����\ˢ��22��C�����K�$�3>�yaGh3w<�$�ۮ���'���(�H,]�9���Xn�����	�է��-b��^��W���Z���-�>�bI.��8J��W�e&��ì2Q�R}:(dR��(�����ښxT/MU��a��xt���G��e�3������v��ei�-�%�_հ�~с�8���O�ķ�cg�Oɂju�%��RA��|�R8eS@;AC����*��.92��,:=�0��~+��ǿ|��p��˓�)���"5�j�޸���H7D�%Ԗ}z�C���5E׈�E���X]k��Jp6
Q����5
#b�O�@�m����$0� N܃���=���-N//b��	R���7�ҧ�6����5�R�%�	$��~���K�:gn�G�c��S�z�%Ć�f���f�ѽ��X�"8��	/b�3l�m���ڝL��0]v����y��o\�΍+�ݻ��E�K�:�6D����3d�%$�L���,�i�Ve�XC��q̜}�g������ 7.��űZ���P�X�q�kZ�JB�I�8��HCI�����}��^@��}�C�t8����qYy9	�ot��<���SC�o8�	���:���v�����@i�~���
�	�|jG���I��Ƶ�IzK�ue>(�&�o]���OѼw�Շ�Z�N!e"�bW���(j6jN��1����V�q�[�	�*"��s�ƞ=�����^��^ ���T!���0��(
�I��0#�0����a��� x���[�o�E��
��A,��`!A� ?}N����0�$��B�ė�i�Fr�X+Ø�>=��'�a|�h3�2�%G=Pl�Cu�X蒢�i�4C,�i��G�^�����{Ѿu޽���p� �����,�(���:��(�
Q����`�Ed�?�ڀZ�j	��GP;z����cRx��S�/P��7 IqHA3����΃G�.���x���7h�І� ,���H���b�L�X(��ZG<VG�q`:�������o��{>����?��)	�0��>O ��������l@?�mt�M��&vZ����,��ZR��)�`;%�58&1N�b��� ��Mܺ��~fꋤIh�l��P�}I��(�Xh�?�\h.ÊEH�S��0����Y�P�rt�HL�`J���@w��[���^�n��i"څ�!�CdO\K��Du���JS�煟iԪYa�ֽ;����޿�2�	�ƁUʬ� ��`hXz���k��ne�؀66�]�'���Gw�p�6R�G��H-�U`�!����<�>O0��B[��5
�����M�JU։4<"+r�ӂϏ0l��YۄE(Q��ŋH�	P&C/���8����i(�����+����SD^(�g�����v�yY_��EQ��<�4�</�v��{�wpTL�m莆����>5�'F}�?W�՝�T�����7��_��Rh�v��?>��_��M3Zy�͋W��`�	���B8e�
�8ͩ(<�D��˅�);w�{i�t��0ϡ��W���KQ��p(W��Ê�I �,F��Rr���j��(�1,�v	��Ə����^�왳�X�� �D�2\�:�2��#/5-?H	�q:�6�o���2,�N\�����q�:z+�Ț-�q"�ԫ�'�g�8��w]�����#V����C����w	s��c����8t
�n��h�d-3�kخ#Ś8>0x���,C�Ֆ��R�E�Nq_����]t�}��O?@���k8��7�'U��RAăq����j9��zn��ɫa��Kai	��#��yϼ w�0���k�X~����n� Bi�t�b�Q�X��UeΜ�e>ҭG>����/0�wޣ�R����I�2�W$�%���~����;1��[� 6C`�Vk(�̣~��^�-�O](!�B���hwf�㓨�Ǆrâ�MH4�1�Bg�=K��ύC=4��D��M�n�@��n6�8|F񤄲��6�π�p�ͩ ��>r��n�}���GՀ�0k� �O���ӴL�hDa�no(��0N`rmmK�5G���#�����*���#�s��70�ZG�m���(�y`��g�����F���!����CW�y�W3���8����x��8���@���0à�#�S�>d�E �o���X���,�6v�H[�>@���ܾ�ޣ{𛛠��\��)=�%���b��0V���OvnqB'M�}�0pO[:��hn
��1y�$��i$����ͧADNE?�$��3��1L5�,����J~�����6Wocp����)���,{H�@h�!�G�8 r�BSx}���L%b��"�9w�G���)֩E�Bu�L.�Gqv��^�l��Y�1ZG\�N��p����as��{�70\�D��@��	��F!SQ�mA�X�r��.3#n;�@F��H�É6��D����z��ȵ�N�A���>?wq��f�N�@��ZB�}+��x����V���61\]E��H��G�}6���J�_-؆��)`�:�\L�9�=?�=�'�y��������T�q��a��T��Cl�(>����s�M�f�29��}	�J�է�=�d�\��3�g�%ղ�Nz��I7�dƃ�,4��dd�.R"���~e�$� ���<�l7�ܦ��� �?�{�_��$�õT���P+�X���]��b%�R`�V�SE�9ߋ+�צu��ؕl1��,.9��<	�M8(��Ѻ{��&����� �bң�`��bɻ��y���3O�$�D�%A��>kk�g�=ăUt��h	�`h�LG6M���Dl�$�]̘c�π�w��\[
pA�������Q�¤�a�y�n|�!+��C�M����H��Lq,�����$�G��!�T�@w�k0
i�y&�"�w��~v��w	��-(�Kr(Q� �m��a!�Rx�L���M��r�_���3E�~�%�/�MS�Z���u�lݸ�O�n��vo�
3��
��6� E<����<N5Ja�:,��3���R�Ģ��/�dH: �y��!�b(09����\qZ;N*��m��C��Eؓ��X�C��!G�"J��0v���>�����
���}x}^��KKКτ�o��)|���Nkz`j���t�����˗>~�ƃ�nm�����@!�Zh#�un(s��'=:�ȈxЍ�p������:q󧞆�g?-,$<�����)��r~�X�Lp�(B��@<�X00371���q�*�?A��%d��h�b��q�(|P6m��5D����1jfv�}x9Q��a'-g2g�MNA]Z¾翍�����0�n��v��f�#SC�P9a2E��!�ᷛ����*�K����Ml\��k��/? �[�Z2����E��,)ٹ��vD�&ICʺ�1эC�2	Z�5���x�N�C��a�Rc\-�0�f��ڗ �I�^3���;=�<u�	�5`�C��V�y� ��ct��F��B�4� �B�䷒v�+�MJT���t:Ml`9A$�4�ZT��tu�%%�^:���O�]8 �>{z&�s�M� }����:E��\�s����`u!'��kh޹�����b��!�4�,V�"`ϛ�L��s��<1z�*@Q_��6-��қ<d� o�z��}(�]Be�!�3�p&��0�2 >s��*L�&��\�h�G�i#�؆��!S���G��Vlo"�������<���(��2���¯5&��5 �$����[>��vtxEG����"ǅ�.��@��Y�R̓�v�7� ���� �p��Vz!iw���m!j�WVUT�F�C�|��֜D�2Da.���LRA2�`"�2Kf�����o_���#�Fwr
���g�@��Z�Z,�,V��IKF�	
sz]��x�kH:�666w$�b(�/�=�żҹr0N4�?�E�5�1%�d?�&O�%������>�BLG"�DHn�xz}��"��I��U8�)!ű�\8M��N;o�kHZ���`E�	���{D� �m��B�%Y1�$EW��34�;���p䤌h6����ۯ�P�,Π�wJR���/��Oș��&�jX����+��fȳ,}��"���k�MjuW�O�^kç�?@zPR�TAjwݜd�$���E��b��5	�{St`Lp&R���r�#5���CR��s��B��b�(��]�'N�Ic�MtXe$Q�W�F�+�ǜ��2�&����	V�x�fS>7=��ƴ�%ꁚ��?y�^}ι���>���J�</8L�9D!���m٧�U \`�/(2yU���!�1��f��!Ab]7B84��k�f���7���~�����S�$4�P����}�tSc�����8��ga��#%����D�������g=r��g.Ü`�4�K�.�I�8��T���s]p���W�?��_sy�k/�MS�\����ٸ��O��o�S��U�`��5i
t/E:eJV"�D"�-Z�p��Ć�*#�R&���˽P�[�#�0�S�� ��7C)R�D�zWˤ�P�ca�P.q��נi4��35��%���S�P{�4P+#�C�
/H����"$e����7MI�� I�z���
�I�7���O`�_G�����e�ݞ��LޡM��0��~�!n<P��1t�B�AB`�L@����w/J�`��Y�9ͮ��0�}�A T����ʜ\2��ǰ�D��`d(8���^���=to]��Oe�{ȴ�Q������hNf� ���*q�bQ��xN��Д-��={1~�j����Caj
���@B�ȓ''[�޲v�c:mئ[O�6�u[��W�s�&zw�#�܀9"����xi�	i�tlW���Gȝ�A�-B�r�I�� T�@i�A����}0�ǡ��C�������[X�<ȉqz�¯�F��Fw�1���۷n!llI ���/^Hi"E�L��μ-EؖA	�3����!�m�����?$�e���E��Gqn����P�5	�����8BDr�� *}�7��{��p����v<���+�c�D�,����hJ)^�,@������K29o{
�#l�P�6�a`��qӄ33%��E�,���56�"uۖg,�%M�GCD��$
d�5����������1=��3YN������,G,N�3h�� �;�)��^���)8���Z�cc��
cU���2;�ZE�1�Bj� �6����t�7��𶶥��:}�CA�H��#�����yB4}ˉ%#�5������"�m�>��fJ3��d��!"3�^.�����O��M ���496_#a4���!c�l��a���Մ����B�gK��H����g��\�����^��u��rO�2
��V��ݎB$Q(MW�w��DhH�H\
��lp�PzM1ot8B2�n�Sm���nO���=�����>\[8�,�ͦխ-���e]9��P��G�@�s����'0u�ʵq������\OQ��`�lI��f3(a�ܩ1Q�K)c#I�U.荅��i� �.v��\��.y����D=##��D1��-�$�JX�QZ$�0ҶFh;�����>�T�ܛ��A[W�
�!tC��X�+T��1��H� �Ah�}%�%�)�=�*M_�����^q��],�nnN��<�@u����zږ�.0�q@�������~�*��>�K�Xx�L�:��<�5hN�]s����(�����<%������y2:w]c��ò��c��aR�b��{�����q���5��'?F��MTiz��(���8�B���'��%�n}~�N���C
z�Gڶ��-ە��A4�w<q\�, :���-����/��A���R�@� �r19=/���0��{����kK{�yqj�o,�x�^}���7/�]���������kۑ�8�y��������C4���?័���?XO���%�m�"%�.�2����KfF�'rfI�H�`�b1��NwUTU�'N���ÿ�vg�����Cӓ��w(T���Y� %W4�bX]���n���m	�:+�c3��i�th��6��'�MBFf�f���s���h�Na5�H,���Y0xf;f�c�R��#:��cz�ޏ���@��#��ƴ�`�w����>���1���L!����sA��N?�=m?���G/�<����%L
m�++�fX���Qn�m����<��P�V�\���>	��߬MK�|�~�{t����i}�mjN��$�%J���
+�D$]�����4\��^_R���ϞP��S�<���9u��L�uőH ���[���3��؞P}���P�0ӘqtH��C:z�1?~���w��;ߡx��i��B�	-�K{�a��y��^���v/�Q>?�ݟ�������O�h1`c���w�؁��&���Sݮn���?�  �IDAT�7N�Λ)�h�ۇJ@F^<�K�wi��۴|t�"&�>zH��s-�B�I��8���%mO��4>yE��Wt���*���=�e��S�� �*X7 ����p��mu�Č��L�D?0H��Pq|B�w�"�V�>$wtH�''V5��5d�Y��Q�(�/���/Ϩ�� ��`��V}1U;WM8�cؔ�|�0��ϦEc��u;aܡ�U��lH������!��#M�ߥ�[���ה��������J�Z��ພF�k��4^"麶ʛ��������%�4R4_T$���&���M��N�C���v-X��g��ɦ>ct� �U�RLnE�c��	��9"ꖤ��4��O�+���O�hz}E�ۓG��dc��@%B�nV�X_���x?t�؆�&ɛL�=�o�Vې$.`J(�b�G�W�L-�և��m�̂��-��|1=�x}M���%0H��Ze� o1��7��]{�Ҁ3�W^��Z�c�@	�4�ۿ��	�K�$�� i0wE�ݸhmG�D�&}H��D��������M�E���G.��ʅaUE�U?�V�*)�6Ģ������A筇�6�l��8Z����%�ô���R+�h������s�^fU���5��[��tn��mr�Us�M�G�tT9�lӀ���{��9 a}zֿ��o��~�{ĻN�G��*uB����%����*Iue�QŶ
�MC.d,��"��4�F>�Z�#b_�r`;/�7�O�T���!>7�!�1i�9Z�H��`�{X��������{#�9>y�6�'F]�~mr)ۮ�Hh���a�\� c�FR$ |��È�����j�q�i����LP�cQ�b�wEeUeT������������r�i�[R$�RR�FR�[�J�)��Bz����ݳ�~�{�=��νwH��Ł�2�����pGV���r����=�x��3K��IQ����OA[$M��93:��!����C��[�W�l�k�ZWiQ]�|u���W"l,�}%��
�''&& D���G������F�V��<�!�ւ�l�"����;Aj$>��A����w��>���7M,c�vn-�o�b���٬���cDn�rGl�&sz�v�]q��B�;����ݻ�ؾ0�-�W�� q��A��m�
����ᇥ�>Ga=߾|=雱��}_��<�?�l;�*�ɿ=�U�⇅�=���TM���0毹��\/ʌ[�<O_|��~|=ݶ|�����f�lvF�L,�Y<��,��A�nC�/��vc��l���O�X�������������&'h�, ����Б����D+�[~�n��nl�l�V �+��!{t�Pɢ�Tf�v�u�wE+�Y���$���.�A{"����G�� 7�j~(��`���h��*�ׇ��}J/C�����ֵE�KFL/M�ƏfT��Z�(
����ZX>YR�j�)�ӐZ1y�9���	�`P*b�<mi�0�i4,떰�Vշ�;*�?�"
߄b.����eB9��+6&~o�-�;��%kS��;�_�㍝�E��~,-�/S�
g�������4���A�]�d/u�S;�F����Ý�6LPQ� �]���r+�w4�`�UZ���-ا��f��tc�T&�q"�/Y0'H����y��,F��C_DͲT;|��I�6j��o�F�����f�~&��Z�4�@�TP��r-�2�}�s�X���cN��3�7�����W;����a
*���R���3r�������i֓2��7��&�h�K/��)��ģX����Q9+��w��-E�{�`N�7�
U�w˨q_*:����(-cB��)��6�qO,�� �E'����,���$��'wW&�Cښẜb4�|�Y[��*p[G'�뭥Jû_���vCC�̪�ȩ-��D�b�Ѿ�s$ݻ�2�n�K�����OwG���q�:�pQr���w+3?ֲh�����J����g�r����{)ư2��[�L�n��<���E��#K��*�Q+f�k"���.ۣu���]�~%���f�5�F���E�~<��Z"��g���(�v�� �V��x�q��>d���S�w�%��*W�~��D�$yY|W����r1��X���3�5�d�o|
V�{ݔ\�`3�rI's%���<�|�KYf��lt�췰sl�)������O�8��Cc8Z}�' �ʉ��D��P�jӏ�l���dQ:�	b~�!�u�����z�1:c���,�]��b�.�]��?#q��&�-wla��Y�gܷ��BA|������Z��qr�;�w�Q��H�`{ej�$���tG��<�lC~E:n�P�C��m*��j&N|��\��������$�LZ�ŧc���Qx��ꆇl��9t�&Li"�$;���@�w��҄�%Z����y�����g�&~fې~�#O=��c�������Kǐ�����܎��A����Y�}��]���Z�uy��q䃧�Ocp���@`��PŔ�%_"��8�η�E�I�>a�u�B�>o#��!�����jU���5�%� T����~b1��b� 3V�u��^z$T���'��O­.T/)Y��sH�p(�S�֒\B���-�s���-�/8����pA�o�$X��Xq��>��bǞa�:���ZfI�8J��d!�W�U�AO�m+��^���������S�#>I$�qs���T��ei�X4�t�����W��o2l�(��̇���8��`U�� �@���{���{�VP��v�<��	O?��}��T�7G��͎�7��5��x�V^�ʴ��6�.J���Z���qVI�+���u	N1��ߛ��2��9<�7�ZgD�|i�s��#gӨL�O�-�*��j���w��oFˉ�c��޴2]c��O��2�/� �G`��"�9 K��?h�o��о_�:�K�A�f�)��x�7���z˶AMEX���ǒ�6�g���w��:��:�bF��?3}Bo �;�T���� ��z�7u�ب�9�b�2�'	���p<qNv�.RtG�Q��0�C��0����i҆�y�����MݯE�l�W�x�����#H�k�;��D�\�P��(m�ذ��X ���Eė�3��U34��v@4
SH��4xu��)��v 0=�e�(NVI�_|�p�$��wJ���7Í���M��٣��Cv��1��)xX�o�m�Ğ��Q�b���FNH����쀴��&V�T�*<���d�&Sy/��R���q�ڧ�s��*5,�p��1�a��P�h[�r�%خ����C���:]��LMWy
�mU4�,��|I�(�yK����P7�دK"b���z?2��۝݅'��]TEX�kc�2Ǝ�O�b���w�a|����,�3N�Q�}X&'��&k�h���F䨣,���e�,`p"�8�;�qW���Qa�����CS�|�d�7`8r52 ��K��i��b�p^3�ap
"!�I� �� }����vYK�Zl�P^��#{&�3�a��pE$-���$�-����i���.��!�|�~�.re@n��1�ė_/:lg Q���q�;�$���� )Ï�#?�)� :�yO�o�����F����$ۃ����p�����S�I����\}r��c#:�(��'w�����u�	�4��ȐL����z#|A[U[0�l��.K��g4�5��������w�S"��$�T��Mٳ�8i��k`�{:;����Vc��������Wfb���ǴĐ����Z�_Cuo�
8�s	:m�}��g���4S��^{��fZ
P�|S����n|�+���-"��e��ah�u��Z�!,$��7q�:���'���f�jl�����
Wݿ_� �}p`N�X}>E��ۙ��+�0��9�_��7�$�q ~�
��&W��.�o��?���/:ȕc�)����u%G5k���:��=�Xb'���hd�_�u�h���b׽L��Q�-�7Y�Zq%*�*��6���Hg��Wb�l[S��hҊ%6A#(��<P�j��
�5��:��5�}2!��؄�h�������K�tm�������df�p��%��I����yoڌ����U7�EnZ(��1I����,�;�w�
�!`����z��t	�4��PF!$����)出Q�k/�D��Z4��d	����siV-�A�8%�zňo{�b�j�3)�3���e���C�s��zσ"H��l!G?O�0 ��S�8#��2U{��������u�Ƈed���=� #��t��(V�~�THu��F�;�*���S25�H7>�R5�ө���#ġ�v������܎
��
�������<���mԦ�c��z�"o��@�CQ``Ш���n�����}WPJ�{��u���B-!/���Cn���R�ӕʩ��x.��U?6ވ]*������( �u,�[�A�"��9Y�(D����@����H��=)/X�;!�D�9T)������	�F�n�avnk.�$~*�5� .�[caM�ΐ4��%ޡSc�_ZL��kd*�78���4��@r7�(�c7�s�_�W��%Wr"e%���������I4Y`B���I�Tl�T�X���a9ށ"��B�_x���PGߎ��1�1�>�Z�mو���ܻ��D�=���3<��?>���Xf�!�������Y�V�©����ڵcke�]֞�U9�%�a�V�'���й^g+.�S�h?��i1
Ǡ$p>��	A��%}+��k���~E�,2�D��!G��r+���ʫ��JOe�R3S��� � �����(�L�(J��]�%�iK�e]C��P�Y�����$�
+�z�׆��Oβt*��ϫ
��+pMfȿS�����e���Gg�{�<ҤH�S���.�H�P���������6j�i8O�hOn�j�b�]�^�Cvh��8�������[�����(W$1x��OZ�}�Y���3�~���l����RYQ�������R���i4�&<�%On��@��?�K(߃U����yǽ�˺M���e�E�������]H��_�&��6LY�����}��$p�����JW���3��C{��r�J�l�m����u(�$������W�<��6X�L���{q�ӎ�T������"wEK�L��9�(���`^����/�QĹ�O�e�E@y&�[�FV��&�!R*��J ��vE\�r"0��P�!��<�1�]����H��C~e����1��ʶ�+��j�ѣ;7�9߹�D�a�)1Zs!������.�֌b�E����|G=�躃ʾ�wv�o���W-�Ә���k��v�{�)��$����m4��a�?l���O����%��G��c�]�����n��a�v��]�u3�������!��@���@�p[��R�S��|m�PK   ���X�V�4sE  iE  /   images/b14b5b74-4377-48a9-90a5-00abeaecdcc5.png *@տ�PNG

   IHDR   f   �   ,M�{   sRGB ���    IDATx^�}�]e��s��u��^2�tB�ЋA�eQ��*º�bQPi�uu]v���"��� !� !$!�L��~���~�9���3)#/�0�{����������r�7�U��<o���6�Sļ-1 �x1'�"$Y�),[f������T�x�'a�a�nԴs��*폤2�Dv<Y6��,ɧrqЁ�d���eeL���p�h���t"Z�D#����f�g����?����<!�s�ݞ��͏.ʌ�-�M�7�F��v��i�u#��ͼ�����DH.��Ù$�eEOI�:)iڐ	wF�{�p�����W)���7HoX`�vl��}��������UɁ�S�ɱz'5Q�O�8�lHp��J� � <� ��f�.<�V�`\�&)�顤��#ZQ�-\R�l���xIUWQ�~�l���?�70^�梁��ʁ]���t��3�նԘ�����:lU�\��Ep!�D�n�%h z.�y����\ׅ �E�$1�L׃�I�X>�1i�U��D���y�Yt����$@o`��zWwoc�Η�h�ybn��I�NT�='.�9v�gCU<h�Y B�k�`6�	���%� ��(�� �ua�6,�0\�Ux��Z�6a
�O�=)�{��n�3'~����yC ӽ������V�67�[���h{|�B5ґ�k &	�"Dׂed�
6��
Y��dO��I���E��T�'
���'��$r�<��\����฀#H�ۘϻÞkQJj�V�����5=Ǯ�<7� �C�!����k�<���:w���L.S�	��"!y�� �.�6\�ↄ$E���
�\Ra|��L����1�E@����>BG�s8� @�z�6ٮ��dlq2+h�99�)T�pky��|���s�?o�uO�3K_z����{[N6��B���%1�c����g���p/KT��Z�U]��tw h������[x�-��$@��҇��]�c�X�`�������I)tG�d�=����Zs�ϭ��?�΍+j�ut۳?jvo?&b��UE@H�J6Tх$Xp,�I�$�,C�����:��v_Tآ3�! |�&#��s�D8�W�I� �����J�ݓ������?5.�}��?�Lp�������m��S^���tW��J/���tM���bXD�g�q-�l�K̻q/ �
��A}��ux_|��H*�3��0��$J�C﻾c H�w�8��T�밿��\�P�1S����P�E��_Z��?4�zN�����'9�g���c�+bNN-�,���q`dlfOdY��(lW�M��L+A`�$E$�O�|ﭐ@�/Pg�3dg�i�����!���a��s�=+ϵ!�-)�9����;i)m)򓒕k���֟'���0=O�V�����k���|��Yw�4�""�=.lH���`�5�(����|Z4zI�E��W�֎Î��rI1UEƝ� i���`$K�$�x�����\�g�;Ǽ���,�!���s�C��i8�o�}�@�3'�t<~[e�KO]��ܦ����BQ'���0�K��T�(��TZ�kC�Tئ	�l�%Tʪ1Xg��cv���c�[d����$1~F�/2�Ì��c�$��-��x*Q�`�K.��D�'°���{~B����n�#����t`&w�W���M�m~��O�z�,+W�j���"��04=�5��eZ,�eB���E *\�1W��dL�r��Y�U��t�
}���n��ȼ0��ˤ�>kZr�OT�@@ư!k:<WD�4 	"�r���a���*�[z�߿���{��;_����Ζ�BvQ�A�*�PS��6h<��pY"�����A,��+��'I,�b���s��sS$p�/���s�)O- ���Ԛ H>I���� >=r����tN�n&��ޱ6���Gu+�{䴯��!Ю���A����9f�{�3��|��WT	axK"""�Fx��R#�c�n�zP΋�`;��+E�,e�UR��\*����������?#A )q\�/>��c�������s���D	H�	��� #)#�����Xџ�e��x����O\|)�߳��Ϸo����M�}=���{��~Ewm�e��@��L7m�Si�����6��)"�(��m#�e^	WF��{t:mo����>PZ{m?��sq`IJi"oo|C�����f�*�.r=9k�U�pSӱ'���K�׿?�zP$ft�S��w}hצ��
�ǫ5#.4~�B�R-*�'���#��W!�4)����|��)�x��%(�-,�I^�o��Br�J��گ�09e�I ���3s�ɶ	ț�l��.�m�3Zlk>Z��e��y��|a|_�9(���'G6o��{c�/Sa2��R�"e��]@�!(�-q� 00��T���[�Y�;�"����s��~n�I�(���)���,S/f[Xj���Wk,vb���c�
����0,OB&���pdc�<�5�<[����?�}/,[�~�J���-�U����e][7}LI�
�",��!���T�\D�?\H��<!I�{)ӃE�ߢ�h����-a��;DV ��9��%	rd�@ʸgGbx}�Gcꊤ��[Re\J(4m�-!�Kã��$"��ǭ�P��4u���p����P`(1��s�_׵u�7쁖#JDQ8P���J2{��It!���łE���-&_�@�O庸��#��Bs�#O.p�}�[Ej��cDr�|�G?��r;���mT aL*�~�甹��Q�d�cBV�-3�2�fM�p�X��'���5\12[p(0�]T=��]�lۺ>j$�J5��@�n\e�c���� 
ONR��mMj�2Я0��؞�#ENI�^P)a	~R;��L�-�EF���a��U���� ҵp�7�F�I��xlK@�v )�c[�s6$� �c�d&Z�T���Γ>�YX����0ޖ-J���#����~���U17��k!")P"%"%RK. 9�HF_�"�0�$lG�b11�c���W1���*$�D��腭;��X<Cq�M�7��d%��D
�+|����-��:���/��;�B��]�l�I�B֖1`I����=���a�9��;CL�)��|��8�lK��?;��ɋ���°��j[�h!%�&/�le�%�:��1��$��$,X���[@���
��"z�^�`8�T�z�
����X�����sK��f���H&IP����Uf`�(M$R�g��R�HB�qa�-�&��:��1G��)�-�G�v�)��<)�_�K3x0���������_d�d��{&$r���+$^!U�c7�bx��M�T�7�b`�}+�d��3��)��d�W�2�T�|�������A��T�ȓ����ç�0�5%Ẻv}g���լ	x	)O�e��t!Q��t��$�)ݩ������e74w��09p�oH�<����u�*�LUĜ�Ni{�hE|i`|�@]P:E���0{A��w*]I -S-�vw�4pC�})��	,��]�l�-~b��d�p�L[^V��!'�<��)�"ï�_mn�Xc{�JvR���5�/�Gޑ`DJ�톶��>v���|fۜ3��wM{�z�;�<|V����M&)`��b�pI!¢|�/�js�����N��$e���n!�%��=C�N��+KHf*�$(¦�X�ҁ��P!@�n,������d��AH``8R��1!w�ua樠ǁqE� �aAș�mi!�>[�������w�_����L��oUF��=w����͏|?ߵcI��D�ν*����s�"
.[��%A�W$����d�0ڶ���I��d��'F/f����2?	Y�\mn�8��( ﺰX�M�"лRCy�t�(�Z�n��ц�W&`�A.��A��c�,�F�iK�ej�T	H$$�Rr�/=�7M������^�57��<T���w^:���ψ#�E�0��(`
.\E�KYc�R���T�Q�90��E�B�c�6yP���'(��i�rȪ��
��t��M���
Y�)JLZ��i�dL$�,#��uH��lz��c&��)onZn��4�IJ���>e�e���X��b�O�3� 3/!�0P�`C���Z��럙`����=���������X�P��+$*~�2L2�䶲��À�IjHb(�� 
 %�
`�[�R��PcŘ̻͠g`��id@� �1�7��HP�ː%	�-a�p0�t0�ͣ�o�E�T��@M����(/� �H�B��^���\�����av���5���vf{̜�R0jx��v%[��]��[��c_���_���<q�����n޶*�Umh*��T�$��������������eȑY��ɛ�<jD��j����:��-�1�< �>�ꊀ#K��FGYT�#)�՟Ķ^O�A6�h�8&P�͋bՂ�k(�RP����B�Ar��@8��/O�E�[ǁC�'�$Ǥ��b_elY)<T���?�}���Y����<�0Ûb]�?��Ǯ�:ګ��@�(�7�&TN�B��(HU��������K*S1�g��Tlt�ضQ�n��@A����`x0���r�5	�YP��'��M;���C�8�(��"&'\�� �E�q�c8uU��I�N�]#�AQ��KLP�	�`�Tʛ�{�����h�u�T��p�w�dc�7�=�_�������Sg����*�=z���;���<��IdՀ(Y,�Dޒ"�S��2�����rC�j'�U JI�2��nWÃ�S��&c`^��#�T��� �Cx��!lip��*�_و�¯o�� a8�e	JD������<��7 �}[#V���Y�C�p�'e�h_�L�+d I@$��D�D09���#"e�ZQ�⢓�媆w�� �v�f���o�����F��w���B��`R�B���󪤳���t�1��Ea��G�eA&�N��,"���<ޒ�#� !X��k�FABG��86��ş� ���k"�8�~��C@E	��3+P[�"�F�����C�x��Հ��nr*eD4'�0�^�g���pwpX�K,������3⨉�,�#b�����V�Y��U���+a���I{�/`F���e����y���%QɅ#f�g�)9��aʻ0ϊ��(�'�@�~C������1��!`Ҵ�=�GK���PSQ����=�66��ݛF��=G�8zI	"����փ����5ub/���m� z�,,>pZ5��LĽ4��<֢�ƽ���A��3��s���LI����yi�0[��֣�xߗ^���0�O�x�3����H��R��3pe������+��)��Qv�%�x�]�`�����f"o�X�9?�AD
C�`3ƨ�Ʈ,6�؇^�Q�Y%��(�"�L�0$�uq�@���c����2x��,(�]� x�I���LD�+�_���wT�8��ӥ���r���WC� �S��J�6N.�R�B٢{�;��s~�kٙ}��n�z�9~����qx�wi�  �Pז�2�,%�yPe��I�HB���K�%\Q�-(�0�!�1��9�f
!�{D�!�j��h7tܽc��N$�,����8�)�"1�X�C�#��Etf<��b��hi6P�y��s��%��J��',o,�9�3��.5I��m%�d^�s����<�C
Q/����.�Tٱl98�to�ly�=m��#c=�E���/�h�ܳQu*�H�0�$3w��$(����H���gN�3�H8���p^��c9<ߗ�c�$3@� ��6��ư�T�2��q!�qL ��H)m�C����(��'���2�U�P�:;��|
+-x�������S7$� ��8��UM)�F6��@HjD�m�, c�H�Q�k��{�|�d�E�
0c��l����6�����p$bX�(Ѩ��T��L�ǣy��lr.)���j��Da���$C�b,���<\ׄ�J�"�h��tk�w��3T '.�[Z����́����H[��5<=l��ݽ�q�䀕�N\R���2
�$�(�Ep��
LVCu��3-;�WWN ��z�������=�b�Ԍ�q��|���g_���3>�� C˶�����'n�bq~<3]�dY�E#cϵ$��A� C�~0wY Ec����<T-Q�����Y��5g
�BU�1���$���A�P�]��e	�+��Z�+C�4`K*zRvy�kK� =,�NZZ��:ʣt/ǁ��o�R/��O��X� �͏���O��ԕ�}`,[�D�Ř��Mk�9��g}�L�凊w=u����r;�[9����b\Jz���Q3�˘�̬$���e���d�k1`!��A�E�����ї�pϓ�x�eCi �Y^���ceQ�yUv^@���Q�Y�v�q�(�z ]�7�X��k"����$ �$�|q���v�u��VR��J�Ⱥ`��Ĥ�u�d1�7"�Č0��#՛V�����A�/�;6����ﹼ�ͅ��R{��AP�t�#� j�:*�ĸD��4X��� k*L)�޴���<�u mC6
�/nĊ�
Th��c(���%7�<�3�G�Sش5ÊW�kKp����*�{e�D*0ϊ(�/���nZh^ƶ��4\b�6`�K����G�GGet��(�LJ�3j�N:Z�q�9~b�;�*����������g��|���%<���z&��D;��IKVǗ^���g^��j"��l��fY�`NƋ#
�z�;���,�/����T7��;
)3���T!#i�wK���&��+���
Dj>�I�*�\X�"���ڌ���Ęs""�5^#��	�@%<�$�;0t����T1`8"Se�v�J�?���}r�9��?����Go�x�{�+u2�Od�ߑ<8�3F�ͣX��ʙ�P�٧�r`�`�,��t�a�Z��k�Ľ/�q� �cI���p�ht6� )��X}X#&�>ԁ燩H���@D��XV����
Y�'o��|4F`�����U+�95�X1$M>O��/��j�*���0,�9������֜��Oמ��.��������O���b3YV�Q�D���^��,[���l�CD9���@%^�ĺ�H���2��a���ܷ���/�M�lA|�����Q�X.c٢L�Rx��Q��r<�۔�eE7JR�@B����aEe	ņ���F�n5�9Rm�i�:Lj�'��>s�d�nO�.�A��<�70��
rV���V�u���.:H�[�_z�잍��O";Zw��"APD^��j%݀M �]vTJ���L�O-RX�\���,p�Q��͑��j�5�Eޡ
��=#����,*��,�ԗ"��IN$1a��Z�IVYvA�T�r�5���QT����tPV܁"K�²��ض�v���9�Jc��g�L��Tee�`�򦀤) ���Ŋ�]}��W���5�L��{B�_�rr�#�!4ٽ(!�H�Tv�y�">"�(<+���&�����J��c�*H�)0=	�IeZ�Ia ���%#�R�Fq�M�X|C��,��)aV����ɖQ'��ɵ�����hR\��i��,<3��h��;�5�� !j�"��BQ�{f$y��DY�D�S��Đ��r�I��Z�[y����`�+F#���g|�k�#�|��}�vG���;j����i8ٱ�@0S(�^!���Bkpi�L.���ș�%�����"cÓF&dM*z����:��\@��3C4�gGY�P4jW`+�u`�)�Q�����@�l�<ZHr��Q1�K
�2��:����]��ef���Ez҃#��<`�R1~ÓG%p�m�t�XV���,^vҏ�r��˖�{͎��������돿��<-楥�h���4�%&`�E�%,�J��ψd�,V0�;i��+��n�"5�Rۤ��V=�$������my^�F�@$B� ��"��J"[G��<�~Ò���    IDATE�F�άD�!E!��XT_���ĩ�dщ��˔��K��%��$���D��$V
��T>GcԔ�p�KuG�~��� �6�o��}���������E�t�H~�w��L6q����r� #/I��J˒ˀdگ�i��Y��0����HaHJ���0�����;���E��D"F"Le2�f�l���s�=��,�@��D�#%"(��#�z�*
���U�v��':+�2��ef�>��d#03E�MM�H�sȉƝPV�]��·����w|�u�e�E�[o�������㥺�g!]1�(Q�d�:��%�<��\�������<�,�P�@����d��j�d���E�@��H�T�YU��:�H���e1W���U/hϠ�Ԝ�|��h��wĉ���:��Y�~�K��=�o�6���Jl���h�
9 Y�Ÿ+!��G
qǒ�/�r��n+�~��G���g$���/99�0��(7���(t�y]����b�ƒ����7"g��F�3��t��Y]��}@�ըO�"���<�f|�'+`�!.�ߘD;�u�Q���:�r�3�YC��yl�yi��D�NTYs�e{�a��n,=#yl��EUM���4�� ����!*�%�v��<�k+���ۅ�s^w��~C�������{���ڃ��^F����V1��0:� 2`hAh�S�%�R��3	�b����G�ar�H%	P��N)�K�"����˜�E��0F2�-�)F�m ��U,���|uƏ��d~�?��'�]']���\f���7`X�������0D� �nу�z����������o`F7��f�c�^���q~�K�t��%>)��0gK�G��f��q��&4�#~?#�?1��?���#l�h{�Ep`;7�
�g���^��fX����A�Lg�M�����>��rj��rYR�r_4W@R8ɂ�f
V%>����fy�K��{��XtH	*l1]|ďO:�j�}�gn�y��x���g|׳ת��z��!Vٮ��I!

���]e�F �r ϡ�Ae]]~;�	�t�D�]�<ک���{&Y|�:����*7�+Luq����Yd�x�|$#�z��@��ؙ���i��Q=?�P�܀�0�d����r<
dl�����5����\��mg�/,~WjN���ŭ�_=�m�1޵6��ňL�]dI�9o�R2�*3��~�9�� X9�;Ѝv)��t�m�l�Yfg
Z|��8C�+ ������
�" �I�?��@o�{saAcy���r�#'�3���qH�x�s0L��X���%b��P዇�yޥK�������x��������j�k�;%�@23Pe4�L&�7��L�u���t�#�}��3]Ϻ$?_��۴��H<���|�d�g��X�&�b�G���t�E��d9<_�ꋷZp�N����m8+	�aZ�ꚯ�H}�H�<��
F��`|�;;�ܯV�t��zc��Љ���e����?0����KU�A�%ɷb��U4Y�.�8�"y�ʸ��S��6N��J�9���"k�@��^���{CA۷eQ���T�0��Ž&��A����������Scs3�I~�!I7���cIa�24�1�Aa$²�Y��SF�N�J�/{�9W�Xw�c¼u������[���G�=u��	��U;�J���l@/%s��+��V^��$@��!W��Kr�(��u���8�%�~U1�َ&��~z&�`c��*��L�6����R=��N��,:m�W�����mR���'�L�t�μ3�t�謾��1D����ws��\}�̥倩2&5w}�z�#w~6��P��˞�5�2U�9W_QZ�%)����lv9`���%���9���R����(��l(�$
:>���=�k5��?��L�/�IVn��^P^��Al0�OT��t�E�m�����`�R�l����U']{�;�yh����İx񷑗��󉩎ߒ��i<	E�2h�"yO�-���ǻ�X��_k��s�+��K��4{�_2 �?�	���nq�>�6$���'����+�tC��@A�^3;5*pD�����6�E��"����vѭ���oן}鬇00`��[~wiS߳�|����=+)�&'���hG����)V�+Z���"ٔ>��1O�Ʀ��XA��T\2}���o���'�BM�A�X0�! ��L����71Ɔ�2��x�a�pe����[��y��3߽i��r@Uۑ�Y��Ο\bP�khD�&h�~NX�������ƣ�3WML��[%��d3x�HS�]��=m>L�Ŧ�y���C�!�|�Y�pU95%C ���^��W֒�O=gA0!�����	�C��7�M-?��u'��_�O�̌Z�^�P��1���������W8�+®���;�ԙD7l1�Jv�l�X�A��I��O��~��MSb]�~�ej�o��;	���(����k�z�z��x�_ʎRǧ-�Cl��g(�O�G*�d	جǈy�v��[��G�c׿n�����,0���o���V���"ٱcÎ���sah:,���|��@���T'2�L�ﭛ�b
$�/��N�� �_����D&�p>K0�cX��|;>]�}���H��0מ��&7�`��H�@J��󉚍�NY��s���L���Խ�֛�}�Ɩlx�+��=/]�M��g�(&\�CWv4���B�N��3'm��-Ϋ��X->�����z-`�c���H^��G�?�)P�0�~4m6s��7�P�q�yIE�O�\�����������<#�J��;b/���y�/���..���(Z�eF##Ȟ��X*D&1fc��/�p7�~���� [�t�t�^5�rz��t`��2�¡��ۮ��8�o/K3�w�\i*�Y��� È��sՙ����M�vs�i���{��
i��	�(��(���D�h3[C&E���/��H,)�:�h�������K���^|��s�M�z@��GIMGd !�.:7�SKbi��-~��h���xNĀۦ6��v����PŊ�h��A�1Cn��n��T���G͉5	�Ê�2�dx�/1��
=���V�4=7��LM��>{�'o�Q�S�| O�Y�g�������m>�wڋ������~�q�H.J���%��F�g�a�J\�y�9�^d�Ը�˫>���Jg�I>h�PS�_�_�����'{O+��x�N��"r�S�4
U*I�X�OJ�4�dn�QVXSR4}�<>��>�v�h��Rƥ��-�cK��� ����ħ�� ��n�. �d |�%e�=I#��0��!��1�;��nXz�ſ+;r���[����ؘ�ｾat��;#�k����"��$�LaM�J3�3y�46J��J:ˍe��}��"�6���,OE�ڴ���g���N� �$��+��`�m��_�$&�ό6>=]��X&K�R��DQ'#|H�d�Jn1g�rrD��2�
.L��	�q���Q3���=xع~q��W�	Eb&�����هϙhy�J-;�4�ea� g��6��n΁G(0�'!���)4�WB�v>1ȍQ͟X0�6(ͫQ��()��9ұ~[�χf���M�H�f�&IaDq�~c�R���.=d�$��$pM���0�L>$[�R5S���q�M��IY�e����q�h��S�s�N�o_�~�)�Q��v�Pw����Z���l9>!�"�|� �M���E�Bu;r���3E�uDQ
2a�:͂��_�%E�L��a�e�<S�m�l�����X�?~k:04��-���d4�y%���$��#b8���Y��eJH��T��g�eA�
"$
����W-F��D�èI��8�g�'����?��S0��>{[�K���Zk��\�,(� :ua�B�a���B��k��fMe m
=)��ϋ*ZB0�R�v�U�-�*u��ұ�Is�*��	c���!J�TF0��*O=G�\[Β��Z�oZ���hy#�<{fQ�d�I��Jɪ��$I�@�zȦ.J�h�y@F�u&���Yɤ����b���Ǟ����}z_6�>K�`�?����O��aalaa�Da��X��ő����=YCt'����k�)(��)LD�T�p<�N6���fgӇ�V�^r�B	VX�%��2{�K�S'�i2�r�q�B�a{gW�y5�I����-#yd�9�f�>��$���lb+y��IJƆ��a���Q-�j��+2J$;W��f"&�=^��9�� E`�9d�s�L�0���������g��Y8��Y��g`Z���a;7����Ӫ�VX&"!ˆh��(Cd�91ɜ���6K+�=R��w��V�s��j��oG�[��&F���񡣽|z>�t�k��'S"yVL��HH5�I��f��n'�#���1��K�}��k��9��0Ĝsr��%b`�լe#����#��Ñ�Z��S/�$J��1;=�$=��v13|d\p�� UVX�5�7z��y���ȦEd�qG�Y�p��|��_��q�?��}�"�=�m�������DCU��؁���;<HԨ:�i�qX��ԚQ�6D��i�cv/8�S��T	}�j��;���p,3�[ce'Vxfj��Y��P���8!Ѷu�FDT�yꞃ�K�3`h�����>�p<� Ĭy"����9R��*�Jq�%��Ɋ���>ů���U�Y<ֽ}y�����Co�VM\��xh\N>f�S,Xixy�d9��KY|�����7�Z7�G�0�ol��ؽ�|驳VV�jq܆�"�fY�]�4x�F&�f����ak���ӛ�e3���h����D�h,���'Ɩ{�T�h�㖫�X����!�L5uE�(����$�61k4-�y�e9N2g;�.�'�j��D�c5ڵX��+˙Ҽ��K.�?��G��ټm�x��K��к�m4K�� v� 13���";�a$ˍG��=z�G��=�=��5�̖�\y����*N�-[XE���A��#��5e�'<���HN,�k�µ7,]y�����~#����w^�Fs��s��95S��4c�eGmӈ���&5���QJ�+��(����*�0ji�tHIX�������y]?c�]Ϟ{���{l�n{�Q3yn�1�D�&QT��r�У�4�0:�`L(�Z�����<��Gg�:��oK��?��ݙ�'�sG�ʊ).�CVy[�,��LYw��P�|��՗W����cΓWw�r�Ǥ48^ �X�w��{qg���l��]��&����&����s����`��K�\C�=j8W� ��Ar12��p��W�}��ˏ~׌�ͳ�/<~ۍ�:��_Us"!��� KQT�j�0i�`�����'�wY���/?џ�c���fs������N)�HD��S�,�!����3�N�j\��K._�:}���a��>uG��������o*WEʰɜ�t=]�!KD�����E[��}ݒKJ7	���L��*��׷����x�k��q�;�D3�5�M�0�L������Ol�	6��Rf��3�T<����SGv^�X,��N�D�s�G'm���΂��?[p�y7�~l��f<.��������N�K��;��x��\�(@��|��+>���^s~�~I��){���p��^Z�"�(����tLL:�p&����;�+M��ug?��x�5��ۇ�~��o)��Sti@��E^�cȍb�)|�����h��n'�>�14��?�xq���/�����bz��I�ch�DN(z�l���i<����?3f�����|ߋ���U��A,\�"r#�˟=꽗|��m�����}��'�^,��֔�0�)�c ��V���EG�uM���y�;೹��[�v��և�˛�~LB2�
!�a!�jO/��>����<UF����Υ'��z��oIS%�LLf���ƣN�NӪ�~�8����f!�h�f��R���W�x��Q1&M:�l�^���{jŹ������gzݳ6�t⍿�fE���7xc{�ZZ�ɢg`8#c�o9���?S��k����U��H��_��o�߮-4��G�@.�b��&���/zׇ?[uĻ;gz��̋����oۣ_mR���\I+�r�Uw��^^��]�3��7�qO|�����/�o�񕶊t2�![�^{���x���KΛ�ò�	���͡�M��c�#ߌz#�4]��l��,���θU��٣8�L�>�k������w}��'/���0Ҷ7h�ϭ8���j�~߃�����ý�����u�������;�ye�*�?V�x����ѭ3����1��C�^�m�}ח���m�f^�]���}�|��3v�im����۞�:�� g���nlX��GM���qOo5p<o�ܹm׻�n~�1[*$r�^Tr˒��tEI�kO[:`���ݽ��|f���a奂��J�k6ΛE;�[���7����KX&�j�VR��%��?(T���o�%���Ծkl����EOP�/]*?�zx+�1�����l��Ap��U=�VP^�񲪵O��Q����e�rf�L6��z��+˗��C�����F~a�c4=�ZTR�����[f�!����v�0�ߓ����r9'�|�0>�������2�����r����͆�_��ZKYq�Euu������30��ñ��OF�l.oD±TWV���x�>3�g{�o�㻺^�?42z�i��t]o)-.����%���Z���������/��ɏ�|>*�Y]M�w��C*����޹`hd�V�0�u�����?jk�7���_m���r93������[�x͌���^�����݋�n1-s���]�%����Ztל�� �|>o��ߔ���2V��C8���?��ٿc�� Se�4M�-.-�Dm�Bf��Yޯ ����i�>��e�p(~sY}��ˣ�3&���Q?�5�󰑁�?0���}��f�_������f��\����[^Z����y���F]��\Ww��ÇG��`��R]�K��?Q]�D�̊����|�=14��t.���0�b4�sYi�5��u}����ڱ��{V���2�E��%J?U[��/�@�tg��g`FGG���e������ﮪ�����j������G0�#��7s	ILQ�����ŷ	�@O#��k���8f|r�l6y�a�C�p��ꪚ+
+_sf����Mz`G��#FGG~g\�%
�/k�]L�w����m�0���S��5�i�����U�՗��WS�(����I�� 344���0�%`�H$�@5�j���7�P��ew���zdx�w��T�Pa�����E��)0����S�ɫM3&UVYQyyqq�������߽vxh跦i,fƿ���aV��}Ve$1���E����h��޲���JKKi�����CCC�	�I��z������řLꋆ�E���J�//++;�㘁棆~c2w94�((�|C��?�-0��K�'��7�zA�ஒ��+�ȿg`������v]w��j0�S3���Lf�������;j��>�U�5���f(QXD�����8f`` �L��[6��B.��ⱂ��UW!v�'1������c;�5M,L��f�-s�0���E���������P[�x�j��m�����[��w��v�%���&J/k�]Hq����<�;�ښ��dz�L6�D��k���LOO�ʾ���ڶM�_����yu�(�U��>�˞׮����7��Z:�
0�_�:�%f����n氐�+��Lâ�g*q�q�����7���z:�E��[6�]}�W0����t���ƶ���),*���n�s���N�ƾ�JO0nj������-���z��׾����7�c�i��D��3����z�{���)1��;69�u�1�H�-���^�O`�wt��Z���vz�\�1<�We��_c���j����Pgɐ�t���H+T5�UXX�����ΩĴv�z����W`���]�O�i_���~a��h�Eş�_���9�]ok3�O�\�OU�w�{{�u�t�: &QX􉦆ŏ�50�'?��G(�	���4�]w�{eLgO�M� �P�Jd  IDAT������M��@bB�h�֦y�������.��%`���0`Z;��r&���b�U44\}���C-M]�]7��t�(,�DSC�\�2Okk�u�xr���X,Vpgռ�/T����=�{:�oi��*�E�%��s���s��ã�e��H4~Oue啇:�op������W�����M$�?��4��r��Ԏ��3G��m��H8z_Mu��JK�r#�fc�_���_6��{fs:v"�����������"b��V�~����w��V:~p�k~k��_2���>�9Mɨm]{N�n���#��k�(.��ѳ��J`L���������_���$J/_и����~ILg�S�G�k���H$�pYM�g���i���P낖��_����S���s�]V;;��><2�=&�o(�+�lUa�!M�n]����S��ʮhjZt�5.y��tt��}d��{��+�Dc�U�V^^Y9��.��?/�b��%�\U0=���e�����#[���,������}����t|�pۢ�ֶ�3�	���0s�QF�ֶ礱��2`��U�U������)�oQ`��(Q�����s�Q�y����r��hߏ3_�Ğ����Lyy]�[i�g{/��m�Z���8,H�\�4��1�%�I���G����0r5�h|SMe��ee�-������CC��:��8�1���|��q1����G#��ێ�������Fc�5�uW��Nt��ji��e;'��:���\3>cb�M����lY50��+���Ƣ�ǫ*�>w�������ͭ�7ؖ}����D����-�Y�Y�rٟ S��kY9���K���E#�G��j�<ԍ?����G�圤(�D����M��$���rf����Ζ�Cý����h4�pUE�uwyh��������,������ll,�� T�ռ2O��lY98L���F�U�U~�P0`L�&�I�|{����%0RWW�����_Z�Q�F�,���?��n�hn����')��,L}g��ҟ
BYz&*�@Pd����U�����|U${�����C�Ɛ�t������)��L�|����s	���׺������eTFñ��j�9Խ2r�;[Z�g��:EQ&���75��v.�Q��������i��c����U���|��aO[�wl�>�SX���yK~?����׺v��秦�/�E�)/��֡nc����[Z��bZ�9��N&J�<�2�(��8��TWW�����o�V�2��\UQqcyy�!=k 5Pֽ���M��UU'���45Fe��.�?<T��E�H�    IEND�B`�PK   ĺ�Xm.���  ?�  /   images/b2b92e47-5c05-492f-ba01-c47f59068786.png q@���PNG

   IHDR  
   �   Ks3�   sRGB ���    IDATx^�i�d�uvޖ{fU���t�Lς!A���hRR���e���-�vPG��I)¦�e��EKa��-��	P�pؒi9H�d�� ���p�Y���R�T�^k�/�{��;����]���%wFtWU������|g��<|=���3�p>`��3�p�����x4C?8g@��E�p����C���)zx��x8���x8g�g�!P|�=<��<���@�p<���3��3�(>p��p��C��YEQAx�(�H��!��{|_DB����q��vcc#8|8+D��w�w��a;�}�֭�(
{O�(
#��<WQ9>��x�0�z�^�h�H���>�*�a��z���{"{�Z��·߳,�j�Zj����<�y`0=��؅��	��y�&�#��˙w߶��'�c�����wܘ�y�q6������-��(
,h'��H5��V�sr��(����jL��aV	�,.�8�,��:��0��<� �yNᎢ(�?��d�,��q<��N��QQ�y�$�<S��0���,�"�x�$�2@���y����eE�E�e
PI��</B�5���E�a����4M� Ȣ(�E>��"AD��E�GE!�8��AM�	q����"�� "�$	Q�0�<O1�Y�i�<c#�7Y'q�e��<�L&��,��H*A��8�p/"�L&��8��<�'Y���Fc�X] tpLZ�ׁ]�~����@��>O����8����1�� EQ�����^�E��x<�FQ\�4
�0�̂�VH\�YQ�����V��l/N
��L�EQT�8�I^�&y��g�V���0�</�X�y^ < �d��A ��&/ĭ���!�V$��<�"�3hj��(˲��18�'I�i:��Ss�iJ6�L&z�XǑ�y!Y6��$���0��5�d� �G�8�̄AH�!��q�q��(�R��@*��gyF�d��ؓ~�($�T*�c�f�d�U�$��"�nR�V�,�ܒ� ��(����g�#�9���d�v+�dP�L�(���aQ�0�q� i��a��$�GQ��1�@⢣j���ߋ� � 5�8�1q�"���Hݽ�E����E��q��X ��$IҬ����5����lY���Ȫ���lH����%��^ь�J=��V���,�VF���<���lE$O�<���OӴ�eYUr���)��$���72a�I��q\����,�dYAP ���I�;�������Q�ӂ� ��I3��Z��wը!�c  x�����?/��k�8���?�H�$�9m�8/~�q�o��,;����#=�������j5�m4�x<�wn��$ɾ{�{����1\��C�%�tAEdgʔ�b<�&����D�DqZ�E.Q@T�"0�0��x�� �ʋ �e�� ����B�<!��w�8�.�b��DqЏ�x7�q�$J��0LSe7E��0�ð^�Y6�V� �q�e�t.�,���`��';�W��� (���N'ҕ�2K��SAQ)��d��+ �4M��tT/&YuRL�4E��d2T�>Is
b�V�(J�Z�K�ѐj���A���n�e���-~r�0��m@��h!d�)p� ,�&�a�î�\<��������PA��̀�d�a f׶�!;I� �;,�6����}p���y�q�w	D�γ\�þ������(���{<>���k�߱1H��v�9V���I�3���n2s�$�T*�3�2`�`�'�Q��8��A;�t���v'��(�F�V�=�Z�ZR��Q��y��a8
�`��R� Xƣv{����`�;z� �(n޼	&��5�:����{�|�p8<1��tԚ���H����d�1�k��%�D�8)ta��
\I\���EI��4�-i�ZR�5x�=^��F�0�m���R��cNk��}�	�����	$>3���� ��	�1�ϘM^�|�a��b r���^E�������@��@��ӿ/���@��������׶95���v~G��(`b���@����gN�\���r�|������>�3\www���~�U�O$����I��A�nRM֢0�Eю�͢w� ؉��T*��Zms���	�@'���G��766�<?�K{Om�l��[��g{g�ذ?��1�����; 	#I�P�@�N:)%��ք1��V���URo�dyiU��"�f[Z� @�b�Ŧ	�Lpn,j=�δ҄ ݗ",��A�csf�-0\�^>P(h)�����Υ ����R��9� |��� ����Rg2_#����#_��0 �� րǄ�L����(j���vov�f��0V���s��
f���k%x��qL�3�p3�l|>��������]�7���5���K�$Y�$�8�YQ���H� U�x�R�_k��_K*��U��|�^��n�7�(M�?t��s������G��v�k�������;��mmm5���z}���jFP�ҪU	p&QHM0��K!aJ�¨7Ro��
���ȡ�G���G�ӞW{���MS��$Qe���f�iV[&J}Acuq�@��_� ��b碶ϕ]�w��o3%|��kU ŬoC��~ӈ
BЪ���O�fL��o:������ݻ��|�7k"ع�^!��L�{w��	�{�}:�4S)�Y�>�0�{)��)c>�: ��l�{!*h�����I!��P�N9�y
�!w�ܑ�~���1@�ұ�yM�X2�XB�U�D�8**q���o�k�sqR�b%I^J��ۇۇo�Q��?4����ܹsGww�>�����;��ߵ�����M��ٔa ��m���I (�[M��k�\�!1�D�K>�$�\�$�\T�c��;iw:Rm4%�Td~aYN=��9|��
�&P�Y��3uV�V�
�e�*���4�>�T{N��% ��Ms�v�[!�@��0Ơ�Q��i�7�0𳅦c �PǦo6� B@J-�9z}!���m��1c,������ϙ]���U)�3�d{4-���gK���uD����_\ާ��.�S���玿gR�a��<���E�דq65C�u���>'����Ql�b��qT�J�h�o�Z�8���f�s��C�X�?�@X����|c�������^o����vcwoOv�{���-{�ۜ���lmnʠ�G�XY���\G:m��� jW�]T+���$��~�@���I{�#�FS*ժ4����#����N��Ҳ�q�@Q�J*��K�f�ʀc
"&����[����Ej����.ܐc���`c���6\ �Y����q��h)�aA���^���΋Qj�,�Dar�Z��Q���,�>��(����7��̬�Ҟe��8��>�of��ó3s����|:6�,MKAg2GQ�x���H���pn��������e4�l<�x��ԫ5 ����/.-v��V�������m� ��{�=�����w������L
�^�'{���`#AB�d4�[7����&}`�jUZ��Ԫ�41a�`�+u�C�c��|��VGZs�QTk�]\���Uy������cR���P{��@a�ΔjO���f�S2@�ى/��
�/_8L��(��0=f}:>���@���<WV1;V΋�V�5?�A/f��Y�)� >ڽ��=�8�}����珟���58?5\ ��`��YX@��y�ݦ/�4��HF����ڒ��-I��
u�IP�wl� $��w1`�k0����ޖ��M2�F��7���j����j=w���;`�2
�<Ϟ=�m�/_�Ϯl����px$MG���o<�0Id��:͆d���]8/�.�Ѫפ���T�XZ��ԓXb87��dAH�d�V[Z��4:s�h�dq���u���G����RotJ�0A��O �v0ScV�����;׬?{8}����׼��]�g>�{_h ,��А�/3I�1��p���5�f�,H�ޗ	�]��W(k�P� s��M�:�I�����= �����j@-��p��ADm��:0i�sۮ5��ڵk���.�t,sss���"�nWj��
��l�9-��Ϝ��1N��$.]�$���4�MYZZR�?[�6��t^�����幅/,,,l�`�"gϞ}���������W�\'aww[�w�@Ɠ�Tk�̵[�8ߕ�/o�����֛2���B�-$I!I RO*�ۤըq�yQ2�4Ϥ�lIg~A���0/��%YY]�'�C�I��r�A#�&>�
�����������و/���s
<��� ԃ�����UhF��/�����e/�;(�1��s2k� `@1{o&���YFQ��9/����,S2�2�W���e�K��m��g��8�t Bp��2�	����v�
�F��3�Ao(W7�	X�G���B�c 4K�s��;����,�������[oqlG����^�ٸ�l���������x:8�vʇ��Ѐ��8�ȍ�?t�ʕ�Gq���	CA.�J,i�J�Y#P̵ڲ�yG^y�����oH6I��R�@J4��q"�J,m B�#�I&��H�z�T�-��ve~iI��ќ�գG�ȱGP�$��R�\�Ʃ��ܼF �i@��z��q��?�8�;>e>�NK��:0� �j_��3u���ՙfd������
_�M���0Ytܦ�}�?��ٵ���iEa/���@��Y����v]�/;��*��`-߃��3ӲL�7g+�/�·p7��~�ˍ���������dn��N�(*}�K/�ec�q��������^z�%y�7h� ��|�I*;������o,t���ӏ=�އ��v>���={�s���?s�ʥ����=	g�zv��,X�@,�B�J,�z�~�J��[7��/UΟ}O*Q(�JUBh�I*IJ��Ea�&~0��^�яz�#��9EgqQͶ,>"��+���"���p�����2�}�g?��D�&H)�n���Χ�4=�~M���jz;�&(X��]��o2�s0`M�(xM�{��,x)�R�c(}���wV�}�ʀٿoc�&��^?tm�dsa>�A��}g(���	���<���<	��� 	z&�8ll���U~oyuE�S� �Tk��)�u�E��_��A���W�&^~�e��׿������G>�2��Y�qT�څ����Y92�k��><ŇgΜ}f���߼v�����US�I�У�̵ZE���S�+��(��~U�|��~i��Y��l"A"U̐����6����A_ñd�H�ޔVW��5ߕF�C���!Y=|T:s��A�V�B�R����f̀�4�-t_��
�F���L����s|�9"�'L���Q��U�,d���{��e�}��g�����v~��,��	
�n��}Vu��s|�&�?~?PXF�3a���G�?�3�Ef/X�����ۣ����䥕e��	�y��a��K��Tvn���`28�?��x�"}��G�X�g��
,դ6i4��?v��_{��co~��CagϞ�ll���W�������#���lԴcX�@��Zo`�䨀�J�5�_�"o����XߐXri�
 |�(*��L�j�!͹9�[T��������
��t�鐢Ať��@��G���%��~Sd��5�`g������^}�=�� �guP��2�+)���t~�����5�����<�	�?'�,�X��,�*� U6+�Q	^��A�����XnJ�j�/����ܸuG.\� W�\��+�V�G�CGK�Vg-��d��1��5߈]߷p:��ښ|�_���yꩧdqe�̽��"�j������X����S�Nm}`q��׾v��+��[����'�:��A��B��ZM�&*1j�IGٸrE��ƛrs㚄�DZ��Ă�@jq"�XCE�fSCFA���p��$($�֤�nKgaQ�s�Ҟ�'P DZE�1i�6�2����?f�w����^w{�mVs�><^#��	������a��>����㧩7�ie����>��@���Z��Y��K�2g�]`�V�,��Y�c/3�!�D�;�oe
�����(,L\�ÅELx�n�(p.8��)��}�ڼ���B�z�}	G��2,k]
�6��d��q��a��6�pM��/}�?af?�����X|��7��]�*��:����>�я�����_|��?�~u���v�@�73r�Z��
%�:D�K$ÏF:�ɍ�y����ڕ�2�e�=G���T����F�Ƈf���P��c��KҜ�Hwa���G��(�3�( H�9�@R�ݴ]i�,P�jǃ@�#.�i��A@1���k�7�4ZS~N�ֲv=n6/�nh�@:禍o
���t���ܻ؆39|��ǳ�y�sɀ����nsF`wEu�)��� 
���.�h}�+P2��3�(�26���)'^w2m9`�Y:v�@vvv��ٳ�/(j͆�>}Z#w�jYO��+/�љ���B��³�>{�+P�+�x㍵����ҵ��cw�ߵ"��d�)ցE���E�/�f- �<˝�7����ʕ�d�ە��<� $q��Q�J��t)��&��"�vS:�e�G�P�ʡ#���Ą,ƴce���1Ӽt�9!�Ot4�OԞ���DBu_�t������j֩�4{�t�iV/oB��Y�9}�1��?��k4g��,�Ͳ]�z��3@Qv�������s�M ,�9r	4S�(>ϼ��Y���a:��2
M�6�����\�z��Z��Q������vL5�R��xf�Y��9�nMb�H�����^#%��<��h�H&s���L�V��k��_���_�0̏�
gΜ;q����������`8F�"���~�'#�'�( �.Z{<��'ٺ}�@qu�"��U�d@����F�.���r��#d��c��W�t5���\
�����>"���jiҌ=CsAὃ�b��8����_`������w�E��h����w�Tm
�
|����7P�4���3>����E9g( �� ��k=���g����^��dl����AJ�!SӒ� ��̴�ŝ;�e"��P�D@t�OTӊe�y0CC�mD1��ѐN��^����ԩS
�id��,����$��͵������o<�̵{=�?���(���W�]�x�����w"��IP0M6G��D���c��P�Y&wnߔs�-�/I:�K%���iz4Ҭ7�дf��e8N%-�I���):��Stey��L�qV�h%���hm��J��Ͱ�(f�bV��R���"�S�Ժc��AO�	��9 
&�>���n\� 1kJT=�ߣ�*��rZ���\n�}�j3�g��)�z��}�l8&��Q���B���HC�8�H���rog���k7��>83��W��p�;�2� =0�oǣ����X}=X��OR:H_|�%y�wH�{�1FTMq�S:�$�0(�N������_��O|��)�P\�p���g��;ۿP�	tN���Y�2P�1�p�D!�L�L�F�����ݷ�bx�H-�=e�" �D�7" $la����ǒ"Y`�l(��l�$��������Lsh��В�P��pF�ʰ��|����J��l��1��X�/ld>hZ��s��,Lt}��-X�0��,`�}96.�Wc����� ���d��g12 �?���?���x���%�M���^@���y8�@�5��em�t��Q\�v�aL3��8�,�wU�H�Q_�R�a���ٮ��9�&`]��&/����u����������
*�BWaoo�Z��V��啅�����o�A�ý�w߀�7��wy���nm����x�<�h*b�F0 , ���+�h�˗l"7�m��������L�F���Wh0������*
�S���d�,�(&c@����ai/�K�=G��.,1��h�V@Y��`jІw�Z�N\���'1c#[���@�ʉ��0f�paz�A|`� ���N��Mp�������i�F����qn�I�F�� ������A�m�������~7'�1�YF�o��E��    IDAT�%��}���i���t��16cxϜ����Q�0F��ˍ7iv�t�b~n�IQ`0U���ĭ/3ApnF/�=�e�n͑P�  }����� {~�'e��j��ث$���P���V�W~�{?�X�x���W޿|�/߼��_���6J�y�5y5� S@�D !̣(�Tnn\���g���u�@���'����	S�^H|�]WI�L��/�.k5���t�e~iA��p|��n,q�7��d>
K��|��LW�y�V���k�w���ʹ�A@q� ;���AAw7K� ���f��`᳀���A���A�K�&�3�?f���̨��1k��ٴ91ǆf��]��=� ���N4����.�ꃓ� �����' ���tf޸q��[Z\��Ph�
�MPp�����;ח�
�(��E9���<��'��'�"$ �[��עQ���������O|�~�r��K��~���+?}����d<W!�� �U����Q�q&�
�-c�ґ�X�&�.�c�`o�@Qeg#g����V�I$���n��I8�F�I� Pt��(�K2���X����|�U�����ȱ�0y�K_��<ܯ��WC�\~�Wgژ��_�i���wf���k���ɽ^ը��c����Y����Aa�,jtO��d��N�i��>�R�o���(����.D
n�2��p-x]�{=��s�d�?�|���[��ׯ_��9�z�>
 ���6>P{��P��˰lM���_y�%���g��/XY1{�*�5�wWV�Y_��!��_}��S.\�{7o���I���f�e�SD���&�Y,si�E:��k�r��E����EL?7@���(
�3�FP��"@�̀ٱ��fW������JM��&����pe��&Ȁb�&�@���n�0��@�:�1k,>(���˗뱡@�?Wï�8��(5�)г@��h�A � �,H�;�3g�RQ(�!��z>����V�B�x�((�Τ�yP���6�Ɖ���>P�<y�E\zܔQ���o�m݀V��٩V���x��V�Q ���l��T1�Z�vnu��_Ym�?����&�o@��+�<u�¥O޹��=�@�X3��^
D�5��S�Ҭ��K����U����dGM4�u���ǯT��n(������^�BW�5��j�|wQ�an L� �pnvK� ���8�QX��,P�Ty�Ga>��?��4�~A��T� p/@8HC�;���o��,ׯp-)���q�i���>��3g�i`c0�}�������~p޼�L����z��\�#6~מ�L���Yc�'���]6N(��`0*� ���@���ͨL|͜O�8A��Mc�'�}���0!l�=�
®/���|���x��'hր���>�؊H�Z�xx��O<v��g�9����������w�]��+�;{�FpݑY�A�I�&�.��K�c�Uc6��b��-I�=���L&,(d�@�d�m��qqU�5�4벰�,K�W��MF�������k%�0�ia6
c����{..�sA�,(L+�������|a�e��f/��cQ���l�;L�	�����դ� Ϛ#�B]��T3)�>��w���$8>/�j(�1	��et��pXgs��ǰ�����y�<� ���|��L���:P � 		W �[�n�<�ˬ5�(��@�3��L6�Ȋ��m�cNz8H_z�ey��O}�i:��X�+��J'h�R�������;�ϞZ^޽O���7���W���/�]���n���
�Q<��1�"A+��v���oc����;'[�nK1И�Rcc�jU:͖�0�#�2��D�FR�23�Q�Ç�57�Tn�*������CQ����k�I�@ �������&���Q!�N���b�����Ĭ`u��#qM�{���[&NͶ��V������c��Y����{~���g���f:f����-�}G�}��3�1�e�l͙i�`*�S�6�C.�E=`vP������L
�G͙�·���5�m�V��^HM�}�������/=�jR���0=aq�q�n��%�ί�,.����+����μ/@��Ͽ��r��?���=q7P �a"Y���Z=�V��$� G�rD3B���Kr����u� �)f��2	�@�V+��Z"�H��g_�{x�whI6��$�v�я�y�w�5����msg��5.0�o�}V�/~��-�w���B�5�b3-�(��I��g����Z��SD�͝���\�G�M��\��}�b���g:�Ε>�]yи�P�]�}0��
ʟ��Y��Ӏ���{B��{~߈�h\�(p�z�QP�Es�����)�q��H(Y�r_&�\_�����/Y�ߺI�x��g	V0�y?��ͅ��$�������N�?�>v���(Ξ=[��q��._�����NiHKf�@6 &b��x�d+�p�q{ajN���W�����Q�G�E	æp9!+��L����CP��( @�N[���e�    �ݙ�O�;85�X�ա*`�?Q���lڀ��i�?�pSF��k@|��e��� n������4@7_�����.pj��G�ìF>�f��,��e�INe��1�+���_�a�c}�cU���vO'C�������<�'�/�Q���3�h�`/gV������+����.�X�Ǐ=¨�Ǯ���"0�aR/�{|n �5���G���_�^x�`�Z�O���E�f#~��W'�Q�V�,w�?w�����������}a�_�ּ��{����q�?f����U4Y�hR���*r!b�� ���XꕪLґ��ؐ�ߗ���$�K�!R4�a��PY£q%a��>�X�&�pj�;-&]�'�ΑՉM��y������im�m�k�Y��ll��W�^@1>����m} �c�Ţ�1J�m�(]ޕ����S�{�Q�@p/�*�Q������Z�k]g״�l��<���ij ����S��Y|�[9D�L����Z�2��C�
4�°ޱzqQ��`;K
�����&.{>1��	�����ߒ�|�+��N��?�q��G:�~���v@�����'VN������1�s��ͽs��������tՀy����u�lĄ �� P �d��@�M���s�3�j��� �\
�)
��?��ժ�`z�z��bau����f�M_Eg{~�k����@�3
<0[`���2!M0�2bG����b��&v> �i�{�0&�����Y��O�s�  lK ��p��gE���M/��25�]�3՟�]�;˹�oL�� ���/|;!q�-G�|&��$�	�P'��g�)2۩��Z4G����V�� 	��g��&2o(p<�(P���-|n��LZc6~ ~��'��:q���[4= F��|��;��X�n����9��������;v��/?~��3�//\|띿t�����'KF�-^���^� �[�"I*���Q�4=PÑ��(��҅�r��Mɐiɢ�@B��� @��M�8�H'n 4@��8"�讬Hwy�m��C�=ߕ���u�(�D�J�@�G?��p��W��������05,�o`�@).��
Ӏ~
�	�	�><?6��Vr��ךK��/3�,����o��{�6/��mn7O&�>P�{%s���mn|BE�� e�m(J�����~�T�[( 8�ݬ���i�����B��x������G��X�� P �� <
���BM�x�5k�ͳ1FM����(��_S>���(�?r�	Wh���cN�ũ�jۋ݅��Щ_|�����x����ο�Wׯ]���(���U��E�L����v��6��Ѭ�`�X�\P�X�*�/��;�(jIE�x�D�t̽'��� 33�f@IE��h�7K�T��mW��G��.H���G1��j�usd�v� )eW�l�(l���΄�Eg����iӒ���[�>Pئ�& >���`��Y��G��oދ�(��L��cKF�f�7f����Q� 2 �����7�J��� {�7O�́g�S��ހ��qn�h B���<W��C0g�m�c��#�4�ND
��ٌf�p�ZD98"Ph`$\3���(�ӕ�[	����}�7�s�����P�;��l����˨�j���������S��k��}�Q��ڻGϝ{���]����9[�X�;���HG�N�2)�F�!{P���	؜	W��_�[�|_@��T�<g^ �f�x&�*D��h�(:��p	W��,,,�Q������a(�(e���@���>:g�5��;�|Va	�n�
��nZ��4�7ma�7A6�`�L3`|�H�$�>��@�rO\��,����4�o:��鵢�ǜ���^��9�3� �@��f��7��??6����yl�F >�軻eJ����V�dz�H���f�U�Z�1�
�a ��NW��i}#����^�/��^O�LK0�(@AF��[�/|�@q��#�uA�B��k�g�
�j���|�W9y��:qb��c��r��ŋg���[����(�r�B��P�~0=2�)r�
��Y� ��x�ܺ�@Q�©�����Il�jR�ץ�����5�c��.���d	W 
�(��6��8�-��<
�UT��hǬ�4&�kU��'��]��{ڟLW�$�������0�ڧ�v�;&w��8t�Ge�5L�NK�E2�'�E"�Ŭ�A�v����?��@�t���مL6��bs��LF?�	�2�l�ג�A���( � 

>M���2?�
���yp�n���
(��1 ��Pw��i �	W�G��䪛1K��%�Y��u��n>u�h"�3o���?/.��*�۾��diy���� ^c����§�����=���(~���x��������o<���zQR c��x�M (@��D[�իh��h�(�>���7$ذ&O'/��1���Aa¦��r5B�'lL�AP���n�A��t��nIl$�C�r PP ,,:Ӽ�
�����0�5o<������5�i�l��]5��hm1�Sf`���y�)<��c&	~��(�V���3c�Պh"��m�j(|����/�@�����B�-i\�	F~c\c,�f��E�ٵ!�"5����`��
3�A�޴mׁ�K��GYPmK�S�S��g��ҍ��}�X�N ��f��[�´{c��l'Tp�so����17�y�ݳ���/�-�����}��a&�/�.
*����:v|��<� �s/�z����~ikk��t�V���6��[��~��G���?ӕ����'6��d���d0b�U�iw <8�rBkv�bG-,9��r��E:3�\�cяN[�5��&��Դ���'���[4�_�|�����\8SM3�6vȯ�Y��&�^�}Ŵh�p�v�e�=���\�m�T�@ �hڸ͇�Vc�	j� ���\�L/���fw� 5W61�H�L���Hs�u���o@s�j/C�郠￱jfY���12��L�谖�u� �c��1�����#o�8r���[�>v~A���7)�K�L�Fx�6%��k�@�"4(o�ml@!�����K_������
 ٙ #����k�Dqoqa�W�:�sO>�����_�s����?�iL� @��(�� �]��U5!�;3r{}]�^8'��]��ףɁ��2��6$w��V$��e"����{?��ԫ�^\��e
�O4[mv瞛_ �лm�:X6���\Zl�]�񧦄���wY�P�.u�7M�&1�A�^s�y���C0.pv�*PX~*\N�	�
0��9�aSܲ�G"
����0�^�̀B�jb ��}�i&)^6�~�l	�n�%Q+�v�fzhB�4a̮G���Uf�����
d�ZH����k���<�ObU,�Z������y�I1���#f�;�k�3��a�0M�M��X������Cs�{���Ñ�h0֕��
5�-/-���N��w�>��ܧ�}qf���מ~��s�����nh(�pE��Q��q	a�K�Z�j-f�Q Ũ�'P\a�պvwDF��1�.�I��N6�\��F�>r)0����t�����$��y�U��
��,P��XF���rN��Y�Uj�S��~���6�]�ϡ��@�2��e
����rMrՙ��C����Qc3}
�D3 ��VS�P64��G�I.���f�>Gs`��	;�-�7�8�HA�:�Y⓵~PH�޾�Ƣ|0���-�@Yդjf�_��z�Ib�( �pe�E�=f�|��,\߀��VQ�bc0ӵ�1k�F������c����9gse���f�).�̢E�-yo�y�����1o쓁bl<|*��ߝ_��G����(�{�o�������.h([�LT����E�淮�#BO�D*�D��`?���p(��m��������ܒ	���_��"��W��`2K%�0��	��Md�_�H{qI�WѬfI؂գ����9k@����t.���tӀ�Y���)�����Pp� ��G��:1�C�(10��s(>NC3ʺ����X�9�"�ͤ3Mu��d(��` ��D��Y��;��:��70�	P(��­��Pf`��O�O�@�s��b@��G�+��J�`nm3c��X�ۢlFk�1('�V��"t���F!�Vu�Q��������( H�����U�l��Nn3;p^��Źٱͅr�r4���ƛg�P�GƂǱ��+Y�:�??7��G���o�����L�<܏�}��>v���O�l�|��SP�v1G�4c3�G��l�H�V�F%���nܐ����q��l޺%��]�H��c�Q����E�:�g)���B���,��23��Ҭ�]?�
4����$� ��&J��X���}2T+����*P(t�>9��0u��be�T۬�Mn~���n�S�u�8�ٹX��z��4��[�pZR�mG�H�U�z[��^�&O�tW+*��.�!��D���4�LstRHf�� 
����x�w��3��˜4Mml�s��1�`pf�}WD��� n��h���������O'�>z�\�&��780�Ga�kJ�"n}9 ����݉Χd��k�c���]��|���Q8K�8����IR��p�iw��cG~������Ϯ]��ɝݝ�(J���G�E!�̱�05h_�ِF�&�J�\��;w��ښ\>��vw��G�&	��'�5�1
 Ec�+��E�B�9���ך��,�5���K�ݛ�؅H�sf;�! �4�	�l�~hPx����)��2�H=��zXw�J	 ���Z�9�������>�ͦ$�����W��,O@Ao<�"�]�5j���(,��"��@��A�FdpT���f�z�v��=Q���^�6P��P��7P5�)�*���,O�ܘ�s�v7?������U�Sߐ�$���|�*��]?��|I�јU� 
n)���Z ��-��:�c P0�9Q6���K�a��s�α(vq]T���P|��Xn�b��vڭ����#?��c�]�$��q_�g>��w]\��ɝ�ݏB@TcdJ�4ڑ��a�2�*	��(D]E���m�y�\|�=��c{[��X�4��a�wE�����:GG���BC%��έ��Q4Z`�S�	��\�ihS�汙ˌ�-߰��EM��q2��zU�&��Z�[��n1P#0�[O��3U�vB��DhV��49�O��N�@H��V*��Yܾ��6N"�߰�?�훆��40�G������6�qє2����I1N��S��4Tk��B�iKc`Z�8�4L����vt-��F6�����۹0�`�(8��}�9+}�ޫ$jf�AXnRlQ|�滈z ,��@�Q��gGf���G�l���m�i�#���a;�/~����}���駟f;�V�-s�]$#���v��.=�ן}��7��?q���O���>�����£Ԛ qz|�    IDAT�܄!8:�*�4Z�R4*UV��vw�����K���b� 1@ο�4r*���D��s{t ���`Wb��E{i�졎M��qP�C�f��`�U��Q�m�⨦��=<5tC>�1|�w�s�iUDS�=z���� �7��(�!��i_4�1?�<k��.}��:r^s���P�jB|:d>�U��4�5����&���74��)�	fa���K���Pr�Kq��L �67�0PE�9`�e��O��A�����((�eW��΄4vb ��d+
3W���=+�>}U����΍=+��`��Q��9��\��|��2J;?~�[N�sǵ���]wy�5���g�+/��y�3@��5�l1�PPP�����o=u�'���G�8F���[���+���' l�X��-����~-� �Σ�H�U�j%�N��vx��m�zᢜ�&_��v����?a$�*���	����X4lUI�%0�XY�a!���	w��n1�BY��T 5��v�N8ԕ�I�Ӵ� ���٘�(�~j�'\��C�+Rox��QС��l�k�3��u��i!����s&`Q�).mס����ǫ&�C�w
������s�?�:4��!ޯ�aU�؃�1L��UFa~��ZRل��+�A:���������zߵ��d����GC��X��h0d%��l\G�	k�΍g�� �>�0����2�4�Pf�HO;u�~ `fJ ���J��N���sԜ���ŋ��ӟ����Wyn���]\�����9p��w:����C?񱧟������ۿ�o�]��ˣ��1d:�t��bf6���H�գ
�^�Hju,�:v9b;<0lP��7ަ�1��1�[���
DKH�Q\�Q�0)�l�4��X=:�]�J9�Vh�04��VzU0�;�D��c��3�`D��Nd>�Rܓ-R�H�XG�ѥ˙�31���R8 �V�7j�:e�r���/���h ��i��J@^���j�Y�� � ��O�����(��=�1@�P(�М��$P`[ Fd ���|5��4�F{,�K}����J�]	xS)�P(�Q4����2�&��s�0�p@���ܹS�QAT��8��MRe!G�_�?�)�e$e8���� �dT^����P�5%8N��k4�ݐȅ�����
�7"*�|`�;<8S�v��q���͓G��{�ԃEQ���O���_���pxR�qa��>�
�S�� 
Gs]xt�ݐ�N�����]nP��7�!W���/�y�Z�1
�'�gL���I�-�C����������5�?����D��:�2���FELs�e�i��ZG�[Nj�v�½���"\�v�[8p��v��q��:5��)TkM7sf�ŭ=$\�G�()������}��%�KB�(�T�5���q@a���(`VN#A�� P�=֨N�۰�~Bs"ⳁ3錉���aĽS���v������9+`��M�XwS��o��@�|��ԎUf�Y���ဉ�C�L�v�Տ � T����s\����6f2�:s�*�E.qU����������c�N��XXZ�P���G�i���ͣ�N�����Jrn����]�����B4�A\h��r&1)��� Z�n֥�jJ5a,�~On�o(.^8'�.I�4�\A�Z�x6Mdʹ�iȤ� �H�ZY\^����8:1����0a����ڎ.
��@�u��\�.�Yh����P�ؾ)��[];r!�^�� �׎.ת@,R�h�셚�L�r���vۿ5�ۺ�4Ì��I�&Ȯn�P�3�k�W�ԞW�`��������B�x�T������	Ts�v���	R����P����ޟx�6/���44�j5n� `{ 0���M�W�a��AY8�"z���=Fq���]F����v�NYr@⟏�]��[:Puջe$�
|@q��:^(�(�2�
��-�p&�z�7��.�W����+�4�]���/]^����! �4I� a�á�V���_hXc1$��h5�҅�{��c�u���3r���r��j��@�7:[���dQ��d�H� �-�"1��bO�#�Npsb
PiM�҅�l��0a>
\�Zх-�Wl�B���	���>�n��=���� 4|Z����4&�..��I��v��^U�.��qޝ�Ø����.e~�$.	3�>�'`粄&�
6CߘQ�ъm��/��4�E��7�L���B���J��a~
033el��\�P�LV�G�/�`Á���m�=�	��!Ϣh�'`�o��y1v�ޘ`��qi�R��y=��������L��o��2\��[�DAٺF���n޼-��������ٜ8~R�qVBc��o�YV�Tgu���w<u��Q<��;��_}��.]��[��h15t��,3�nD+�P9�b�Pci��iԫ�E"T��&57���ٷ�!Ͻ���&Za�lUI�)��җ�6�U�-V�v��+�����5�JY�c��edZ�	��O�t�N7ۓt%-M)�]�Ù*K��4m5�g���=��u1�q`_F��9�q�_�F	L#�v�P��\5$mǤ�L.P׊�L��6����Zp���9, 
uRQ�0���1��L�5�5Ѓ���4 .��ܦi�^�
IS��4���,��rp��>C�8'���~�%���q�=��)�XK�?��Z������ ������Hm��9S�&g����&�������+���_{��y��)&t��|X�`�)8��ǎ���(ξ�Ə^<��l2'��2v�±��&��i�sIlTKbi5��\UL&�Eq��YٸrYv6���眛kjw�<�� �<�U:��m���V����V�d (3��ů�>��]9���2	�3���=l�rL�]�氳Jɒj��+ن����'ʆ\�������f�*M&9y��T�n�r:�9�b#�PؽhX�$�]&(���79���sE���|�l�;e����۬Q!�a)��&*8������V��Tv�Q�k��DhG75�����t����%Ѽ�-(���*3u���Z�8*{S�]M�SƬټ(dļ���֯������(L���uy(�m�:�y]��K�o��.�����D�h�k���N�i����9q���=p��o����7���s���'Yс��R��ׇ̐%ʍv,��F�	��|i�݈t��x,7�_��Kkr�"�Q��07ߦ�!D-�u 1�BKR���\W�]�t��6��{crA���ӈit/�B�� TUb�>/��@���Pk2A$���N��yǦWQJAp���<�8H�/0�]�e�ގ��<��2���`J��C	0�/�{��i�G5�����x4����^���5J��A�E��#�<��Wn& ��T�c\��u97���g"2,3u�"o�P;K�����P��WWMk�jv`�� ��.23��U�b��Cj�/R��C�47�Y�*v)�0��ɛ�40�֜TQ�&�j7Ċ$�`��_�I��cO�"�r|���|�>��֮Й�0)|k(X@�����֓Y�uZs�9u������W��r��ş��q�G�I�\Aq���E�4_Pz�3ʟ��v�Tc�Z�H�vv���lm˭[7d{�C�Ӥ�ެQÇ 
<dך�����&K>Bc�.44ԅJQu��� ����Mq\ڮ�Y�q���̵)���:�Tk�w���1Õ8�3��v�v�଺�L��I�({2/ĺ�	4�X��W��B3��@����iT [�2g,R�k�.�S�i�If9��.69�h��o�(��)�`|�FCF�@��>� �ɜ�?7��``��=��|��1�xee�=8�g�\�XXƙ�<a����*\�U#u\�ˁA�L��ؚ� a�`�"���{<�ם
��w�|<�V�	r򨢬����jR�EtRk��fW*   �ߵ6�<�UbM1iP�(�дwkg��8ϯ]�˗�r�!Z>��
Y�x����ϝ8v�G8F�/�p�����������h<��&7�hB�W�Td '�	aף�EH!6Y��������Ζ�>XK�nv
����$�B&�9�,E����H�B0L�ij�UC�����ۘI�lu<P,f,ƽ�niWk~Ø>ێ���:�����Qn1��f����!�x�����2�
6��	6�e�\�6 u��	�;1V0>���φ`�����Z2� 5���[K̵FDM4\���!^{(P�I�7�� �hu.���Ew��d�eڨu A-���n@C�D�f�����{a�����5�g�*D�,�kQ2QY�X���z������3^�_��k�{�Y81�C+p���6j2��+1 W��E�,oaO�����X�ze��>:�2$�6	�򦻠e�f��9���AK����쉵���������4��@Q�k�+'�/Co	��4�'��y*{;�2j�9�9f9+K�m�9T�֬J���+e�i�j,\fN( 4�����H'hC�"�0% %�Mqf�$Bs�'  �Tq<<�q�������PC�"���櫀&`��-\����m��AC!�ʯ��4�g%R��b�X�$F��X�� ,z���z�s�4*�7s(�.�,Z�����Ҕ�m�DqE���h�3jyL����a�\tA9Fhp�  ��'�>��K�29'��턅/�D��L9X3�1(����p����f*��Ӑ+�����_������9RQ����ڏug�~��7s����ș�\l�vD�p�;[[�ǉ��V�"K%P������j���Gy��o|�O��s���vw�L:�Ѐ0=�na
$oؤ�p�9z�8�v7e<P�0<Ӏv�D���p�š���Df�eW�xF�5<�
�����J�(LG
���kB �{c8�Qja�N�р��(�-L
�h�'>�ɴ9��/��@)�@��k*2#k�o��f�C�UX�2�ҋ2mm��N}��1��/J�����r�!��+�a/�P�l���F�&5���,f,p�9�ر��\5<���[��Q��T�P���qD�>j#(�(�
��/	���_����X� d�>X�	�n��ﳚ�s>���A�������� tD�Թ�ͭa�`�DM�i�IjL�%��g�m �u�BSa�ɐ�2A��~4�й󄕌�
��̱P�
ߛ�N���ܹ~�&MDV [X���qZ4
1˲I������������sϝz����᭭�g�e!NEPi��Ja�@���fC;2�A.�ޮ��>x�fihK�]!M�D�Y� ��=d�M�ZBG(��MD���k)(@�2�9R:�ߍ)`�Ц�j֞�?�a��/�p3d�CT������Q���l����'0����X�h�
�0'jR�5
\����Ԇ5M��lQ;z�����>N�R�paN�oĞ��sAq���x�d��48f��q�(�%��֍B�M��z/D�!�p}P��&�a�? ڸ�' f4�b�'-��:E��D@����>��ld�� =�> -���U"'�����u]{y��{:L5J����f&�1Y�9i�,��`����ZV�	f�MQG1�O�f���5.���,DG��
cksGnݹ�Κ�z��|F.�O�&�j��KG����x��=��-��-��(�|�_����}A�;'P8�C�N����A�PCpTƅ�v7Iu����v�$���`�� �)��5��ٝp�`BU�k�nب�,\�f�#��Ij�̍v��4����F鸢��c��)X��EI5�l�����**mA�Ԏ�ڛ�3vA�%GF�P�%���ԫ45j`I49����`shj�$]�Le. �
��aD�R&db�o�z��#�G/�����&��@璟�>��ό�c��9]��Fʻ����,�l�P}��:E+��@�Gl�Ϻ�1S�1cL�f��Fe��t]�pfZ�sׇ"��a�df*�:��e�Ztǒ�pP
J� ~}
����v8'2L88�%V1��=W���U��.e��mxl@`:%��t� @1��ޞlo�1�\	L��z�ˡ��jRiiy�ǿ�c{�[F��2P��o��cg�~�S�{�?�q����T��E�K�#��D�p ���m��we{sSz��Dj�]93���D:�/��)�7�`�?L#��FM˺M Y߁�7d����b�ZקFqU�(�P��w�!��l�٤S��Jj&o�M��'�I�1�}q��waY�Iu0��ΰm�Q�f��l����$�����^�a*��nK�ӕa:d'���6�H�#��0���r��,�b/�A�ХaL	�[6#���ѡ�v�2�%|)�k�H \pm�~DTj4��p�5.��j��Z ���DpV�s���r�i�aI3?�ܛ��1i:7�r�\J8MI�$ԁ�ϟ5�^9j����t�{� �����	�/���}0j�J��٪91��3�Qx���D�<4�]sc��!�@��4=8K]q�:h�L�ZS��O�7����w����u�����2P����'�9{�WF��ߪT*:����6d�ud��q,{��Jl��]3y�uw10m���0Pƍ>�.����54�I�$��.�EA`�0�|J:��#��T��4�~𶵃w�����3Ԛ ގ��8���]�������c�uںZ��Dm��Ԅ�I;�����.hל��@c�rX���{<��;���p�����L#0�����g.,#wab,ȭ;[���yз�H���f�s��M��N2�]w:s_����x&0,<�2��P�����R���0����9�]}��h�,���`�xj����±�}�}�sP�� fU�(L�g?C�&Y�قp7�
��,z��F�M���,4�y����8ƃ9�u�ɀ�/s2����S���<�A�ڗ�;�����A�Z���:ݕ��h���ةS[�,�P��W7�rs{�{� �aXX!#�s��D��} hf�._Yc��֝M
 ���%^�j�Ea�o@x�
�;�u� 4tZ%5��hO6ͭ��X�
Y�$-44^@t����p��8f@�BY�љ����E�k��8?ƄE��%�c��� �u�KX����+�h�:(a��*v7C���M�q]|w���L&���ޗӝ�pO,C�p���P������b2؄��}Z�d�d�i����v�=�E��}�� ��ݜ�Ϙ�̦�3�قs`� ���;G��=���а����p|S��M��V���n���0,��/� _I�@�|��p.�LX�-�'�J�5H�4L)�dzhe��s��w�VÈ��g�0�֜�� �CX��a|`�ŉ2
n�P�^�Gņ|�������sm6�����?Y�t^\��_?~���v���o(��o���k����[�n��\�HM�
5�!#b�lC�ﰇ�����?P��ՙ}�1�c�4�u.u@AP�a�D�vu�&t�H�c1�5�^q~,V,HDG��+�:<���Ts��~����F?���9�I]�8G1�ZB�1�{Cz�Q��s�{tb��F�}�� ��{��;�9�۷7y�j�^� �jRU��@Ӑ��&Ǎ�U�����K7h9"�p9
��qN�����!c� 54G���ɢ
�< J�B����3�I33R���p���_�йp!y�x�	�Ox�P �<����[��݈����q>�fp.2�r&�n�̛O����a�i=�!��PG�%�1���F1�h�V�j��%zA�R��螧���
~h����m����|~�fK��nv̼�\�:0^M��0�Be��*��:���j&/t����P����ɍ? N|�]����?��������[��7˲�H�m:�����MF7���Z�񳡌G
t�:p2M
����fC&Bi�
��8yYz-����|� ���Ή�(��"Д[�Er�������i    IDATƻk.Cą�m��r�L���e����2���-e\Z��K[�Y�+E>�'4��)�)�$��5��p���Q�9������[i����q6O�X�s�E��/��ugy+�À�����;��s��/��1	hn���i�=��1s�j�����`L����q~2/Σ�k��#���x�gf�����!j煂Cۘ���uq�J��`d�27�bc�|Oh���������<Me��E��G�������O�F~�+*���"�2L^G��@��`
y��(�j®o\c�̗��ó���ӂB�b.Q�vn�+��۵j�������u���fs����hV��z}K����l���7n�����c�#L��U�Ɂe�"G�,9p�0� ���A3 U�@�`a����eP'��ϡkW����G�v��NX��E���
�&�` <X,Ko�CC:5�`cQ��
�"8�2*�(�Ę� �kF�5�,^��nqr&dԦ0�\�I�V��6)lF��M��N��������e�sԶ;M������S��V	�����d@gJs�@Y?r���E8?����o&����cse�RgFZZ��	�ӓ�æG�������4��U,�9��.��r��g
��iL$s9.��9$p�P ���m`d̏�m��* ��^]^��md���S����P��Մ	�{�Z�* �{=m��&W�i�2��d��.��4�۰�)�Y%W�(y�լ�o'V�|��g��� �(���#�/_��+׮����ݏ��0!p#Vd��᠐�Zo@_ �=f3�j*��r�r����lgؤ���� �dΡ`\0��:� �==L\�%��k��D�q�6���58���D�	��P�T���A�z{{�dŢ �MPS�=��> �5�����V�@a�������hd} X��� he�lw�<�L?��Vo>ܿ��C28X��;�}8[.�����ۡ@���9�?����S����L�͘g����Q�	�������1&�&[���kA)�Z�LƌJp0���N,	�S��\��w��Ӂ�/��󛠣���g�f���<th��2�1��D��߄�{ah�uJ-5+���<�����,�F�c���;�2��D�����μvq��8�>�e��`E�nf�����-&��;=#n�!��dZw�I��|w����=����`���3gδnݺu��ի?p��忸��s�?V01�T���j���k���^NM����w�y�X X��-l��ʠ5NM��+�2�!�}>�F\��i;��F��4|L*��|��@a&�i�Z�m�F �
���F=(�e��ڷ��֨ �կ�f�ua��,�y�ʦ������mx�����NƔ����#�����	�x��V�F-d�b	D��[BFڎ/A���
4��oQ_͉\[ �9��S�Fg��q>�
BC��� �����gL 	��R�m�AT�Ri��Q�.��`����*��ni�D���M!�rs�����(�,hԨ���cA\�ń s<��M߂K�um�5�#ڂ���Lt����!�������k�M��<�s��}4Ҍ�}_lI�e[�e'v$�!�8?��Z %��@m�аJYH=,�á�
I 	�8���ڭ}_F�F3�}�{?��̌s�zG���M._��O���w��r?�c���f�ǽ�s��8G^>�"�⌈�/�Q 
���bO.��#ZJIJ\��\�h��{K�J>׶��Ƀ
���g[@q�������k���n[^^n�x<%��zqp�R��Q�\��>z Ȋ��-M_ �@������0���DS$Ɵ�Q#P��"0�<b���e!�����fzq�4&�����գ"%+Z襄Y�&�Ɍ�1���RӋ�k��&�0U#J4�v 
�����dT>��#�K����H���f2�pNA�LFX/�%@'�0*`�K��.�"�L���$bPPG��$RoR_�N­A�b8� b)����Z��^XTJJU+��A����:%��-���b�($�KpVDXa�pKlЄȢ�B���t$vr��7�@&�V��{�����$�&QE�d*�Z4>8.,Z8�wD�	�'7���t���B> �h�#g�-tPu:
P����9���*V�$�Y7��A "�� (8L�$�}�X2~��;SUVr�[����/�
er����t8眯r.;�ZZZ:��x����/0���|����h���p�]X"V&�h۲�<Yإ��H$�@��$�H$�M9]�s��Ƈ�d��ﱳ�./�~H�k�"-u�����
i.(A���E��d�`���T���N�����{�	�(pY7v-�B)������	�b�D#e|h���ƂL[dE�f��E,$�Q�@5"����k�K _J�@"%�I,,~!( ���d��t$ԭE`�3�J�#uA��s�4�u	+"�	+�RȒ��n[2�I�'�(�&�B��m�Y�P/�p�ŇJ�+X����s<J	H�KnP���ի��������&ˎٙ�Em�@�1@iM�)��T�D�z<���O�fI�k^�[%5����:��[ Լ��F15�� �-R٠`|!@$U�Y߄\��W��D�2XΜa�E���ܼ�j�*>�ӧ/�؝1P<����ǧ����z���5���[a�%�GRy^�[(,���BH6���J�HY[�|w�BT ��IB}�D�r\E�� ��ԑȔu�����C���r���9|\,X���nX��&L`��,%ב���	�Ȟ�"�"�pJ%RGwXK���e�,��e#J-J�ޥhq!>���[Wt�ta���R�՘��`��KHcA��$�s 𘐽c�4�r>����Iiq�O�B���O�3�g�����@I���̐�4�Ő�ܫ���/�& ]*�,R�󉠺�?jq�
^$�#�����HN�]K�.ŮP��0�n�oh#��D�wi�EK�+b��a�:�<�x1�	�	��1�BkF��w�A/�1�M��*!a]���B`c(�3�� @"w�H�5eg+�Y����c��0R\Xrg[c����;�K|2����⾾��LOO߱���� Y\#�@D�1h��'�0>3)Q�X���/�I~�$����+K����6O
ق�l�+�Y2�Y*�(v�WS�	�V%8�^%X������-Y������B��<��;xv\��#`0F��E�ui�P�J2��eC*�^"șQIxZ{Bb�a�V	)9���,'�J��G��
�d@(_�t,�H�>�z�|(&��@�慌Ν�zE����!�#�3��H��_��)Bgp,�ǁh)�G��܍�������{����S�BK���Kp��;r�H�KX0DȳZ(��in�m(�Y�	�P�9��T��z�@V�ۄަN'��9O��".�Ѐ �6' ��O�-R�����l��5IA���U��P[�+I�s���$�F��cF�7?����Ϟjow��@��#��mm����Rm���u LE�H�K��I��0���@�RO�%�@M@![ı�4,
����.��h�L�߬j,+-e1��ҟ��`
5h��T��~2�W �x��R������P
�дP�U|H_r�C,,�S��BJԉY�@b�cE��I�����M�,�jP��n�D4��濘j�r�	^4�4(��́D<��4:��}̄O��J�@X�l���dB�P�.��M�K�>Ǳ���Ȩp�*��FA�I�$#C'�Zg$#��X���H.@t�I��6�%-
.�:7���'�cH֭�҄+"�/���b��s#sA�I���I N��)� ���}TЎ2�(�$	�'�.�0���b3#��J��(�h��Y�%�!��K�"�^��9ϕW������^@9��щ[&&ƿ����x1�^P��)I5��#�. H'`bmX K�S��n$�����e'aj���O,.�Q��^	����I P���v��>���.`�"-^x`�Ү�=*��,@�� 
,8���&��������{b,� ,iJ���e��TZ9�G��~�k�1¯MP��Y<�pRގIih�� ��;�wq%�Ol�q�;74�]Z
�0��KOz8� J��C}	тPX|)*vʢD�/����R�N$#A�-
�E�w�A�CE�-�p �Os�%��D�7Y��T�<����t2*���k%}~��c����G�Z͂���/�W�����ڱe�`�$<�� �Kmx��%5Wa�Pߕd�V�xp�G�x\���*���D�B$>�I
���^�y�y�mo�{�t]�����e]d:��;99ug0 Z �`�+��$v��n�(ǎ#��9Df<h������K%%Ǥ=J.;g��$�c�� wdL8��]�9���<�;�_�E��H\U,p:����h���9�a�u	T��ŕe��3[
2���� b��S֘��A�|vi��T2h)�BZ"H��ye�aA  ���;�1 ���"aVIT�u�-]\�KA����Eʹa޾(h��q��Jն"9�\C"�,�e�%���5��2����QQ��;�����kCϋ�@4DV�׻E�2�����!��@�D�����3	R2�@@�4� �)���S�.X�Hc���P��/�pƽ��)�iI0�Z�襘�Yi#���E9�!I�NSq~Q�-�R�HN�mӞ����O=��;�c�=[<>�w����;�Ѩ�'�t ��`��?��b�$��}���RgP�Tز@��w!zI���J�'���_ è���>�
<�|��� ��/����C	k�d�I�O����pXԷ2$(�d�Z����u��
�AJP6�<zj�X�ٯ��F'g)z.�#���n)��>"z�>�#�D.6a�� �K��I@(mצ!���؁�J�҇��t�	-,�0�� �������!��L{
\�G�e�X��,;Jh�)�{��j�q��ủ���t99�o� R�X�8:^�Gv1��%��V���A& �u'�Wj�HKcO�%́l8E�@�G?�d�h��QXVP9�X Ԥ����N4ub���%�����Ú�?��a��Iw��Vj��Ǥx���G�95��������V~�S�^2NqY��g?�u��D��KKK��0e�NRl[��Iu��n��~,�y�LN6�|R���wlQ�X���1T���j�ll#t�O&@��DP�w_
&!� �^&�Zs_������d��ԑ�z ]A�R>��R���T�� Ar�Ʌ��ˋl^^�p�I����v=8�C&+/�m㒱��/+uD��rRM+���^�����,
�=�]�3�)�;$�m(&�s���ba���F@#-;�bR؜�h���:ᵘ|v
������QZ`A)��`cQ���(R�X��(dL��}��aJh��m�T:#�oq}*�B�E�\l BdA�
'��Q�@A���v�	(��1P�W.�o���J:9g����C�d'�/ទ�z,XZV���j�?zө�h^(Μ9�300�ƙ����
.~��QM�7@^�C��˄�2�� �"�E��|�Ң/���s �G�@�AMPPЇ�c�o��9��d��ًd!�%%��@#&�^M��F;pA��G�R�l`�lJ�2P���ϔ�K7�c�WN�t)()���n�
�D͋��8#�4	�wځif��#t<REk´�}9(�(,
���y|�܏BlcT{$wxQ��`�����_lj�i���&,�9M��k����� �뉭*���l1���^��N�VP,F%�(D��s�D��`A�$�u����h��,��wp��n��H�,i&������,��S���Q���V%�iӼ�*O"�+���b�9���k?)�H�����	�%w3⫬������p������,P$	�w��k&&���x�XЅ|��ͤ�#���Z)ӛ&��)7�o�'Rj7�`�V�sV�a �AAz,�T"U�~�?��~2��1&�X����왉4΃.��nb��L����ْM�*�"���A�A�7�[��Ơ��b��Y��%�K��A�]��b��N%�H,Pv�dI���\<<dp°#q�#Z�rg��B��`%����q*`�Yn-(D�Im[�]2�(�7|��]��x�Mo,��h�8�����҆"J	P�A��ԡD�X�Hm�lH��4����	@Z��hA�y⿔���(�Y�IR�E#&��u�AJljd�������ng��ɪ"D�wB*
j$I(�-A�heV��HKb���;�GW�**���l�7O�>��"7�
\���������/��o�.
#�D?77���7�hϓN)Fh)˞�HI/�w~�y!C���;�8�@�5�/a*�@�,�}ZX Z�"�	 @P@A���Ҫ ĕ1 ��_�1�@a���솝�-$�Is�������B[
ٟ�	��"ԝt	@B��\3Z4�%�~0,L��\p�f�0�I���\�s`w������ɪ��@!���)�֤h~ڽR�	�I@��Ѹ��h��7� "���3ɹs-�(a��Y7�z�դ	�l��@�p���G,F�;PH�].hVv��-G�9#%�v]�Q�rD�9�wT�I͓ ���n�����":!#�k,}���F�9�fB ��j�q����=eyyϞ>}Z,����(����ه�G����@��d���&��"˂�$=���R��|	l6qT��/f��v�a
��)+��E�Ԗ���B��M' �Gf��I/,��º����{v��tOrASg4�dz��j�o��A^/�*��2t$^��� �s�F��(bE�� �IK�_`�&�9/�W�Ks�!�'T�i�w��ݏ'�{�����c��I�B!��;	�,�|����Ks8�+B���V2�ʩ�����'�\�˂5����%�,J�^��E!F�nc�E�ݺ8²  ��㹸����BJ��c�cGŚ�ƭ���=�Zҋ�j��@1@S���$�/eA��(j��@pҪ��B��l;������w�	���� �)���b��¼�V�T~���|��K��������{�g�ΙOz����|�&7L?6��T�_x�0`e��,,a2r�o'/�~�Xp2�λM�e����E!N!�ՉX<n�@ດ��.��$s,�<7,$���eZ���&��Қ��AG�l���'��5�%��J����".�3�z\�!�"v�na��#~�j��y���(�AZj�=u4�.0��Et�U� ����t�;�d����I@��3��;
rɪ�_�s`Nh�e�W>�� 4+Ȣ��Q�+$MYiͥ�Tx���EU)7��e����z P��x|E��J��a�%�X���Z�ؘ��i�%�4T����bVɞ!"8����Pp&�7�z����c�%���>}Z)��'c�x����'��V>���aQ�e�'&SwɝY�0P	35+N�F�|�R������E;���4}���/	�WI� ���c��]��a����Y{�ep�vE�҈;��H��Dz�fN�%_��R�LѼP�(]z饢4$��G�[�̩4X�y9-&Әp�,���D�_<��KW-��@��lH f���c��4�����k�0�/2E��	�Kr=R.H*�"�����"x�n/jW�
~ �W�R% ��h�˙_.�4To��}T��r���,s��{v)�/<�㸑Ȁ��)E��t#A�&7K�Wy��¤1�Jc!�������4K.m��A���PF�g�����sPŌ��(��Xg�9�J�˾{�+^�����H����������[�~߇��h���7�d����`'>����ş:VT~e��'�Y�\p    IDATO�$������#Us��X:P�#S��--0 ���@�["������럊eu-ҨT��d$vM�eT]��� ��5����mpwww	n!���������0@�;�ν���=�]���ݫW7��Ҹ������):\�vԓQsL��&���4�e\l�4�9�T�-H�on'7q�͚�=��mi�z�ip�A�(S�\�2�����2��R2�ԁPS�:f�s:ZA&�a�h��S�ҮBuK�Q��*!�
�	d377G���_�)ܡ]�/�f���j޸Kǃ�;��������	O��4)P,X�qd�%��	4�l��Q9#��ZI%���-b�.�N,�%�p�q���e�5@��6��\�D�+o,�b$̉��p��|��=l��jr{᯺7wGF�8���[^|���r�����Y��8����CFrrNx5i��)��G�4=�#���l��ۍ��R��J�_�aN�
Ϯ�盍v~��'�N�y@E�8ߧ�u���]q�A�ś�U(����H�����
1	I�j��݊��L��D6H���~��ba%S���J���ߺJ����}>��A�¹BS�4�4��e�!r�/$㎰DhW\j}G�J��
t�r2q��ٹ��ߕR0(z�ư�Mٺj%f.���ZBVډ��!Zd=K��e�"���w��拏�cj.
�!o՚E����I-Wj���y�y�P:�+�ZS�[^��FE�l�y����j|K� ��������t)��G������N�x���&��-�+&u_�uO���ڪ���Ы�&A����2��c��[)#��pe6�+����������@^X(Dz"�4�F�y��:Wȟ�D8�x!��cV�RX��R���s_~�Da��3A!�a�o�ӯ�J�Z(�1��ƻ3�҆^���L��^��T�RR��@��������tz��.C9q]��K���5�/ :$UA�d��t��Yp%���y L���������<�I7�a�T�x=rb_9�5^�]��"�����7�qLh�S�i��5
�i���/u�K���!�|���p����j0VB�r�����5�NND��C�S�@�|%�F>�����k,������f�q�t1Q����z'�;�7�a���Lp\7��^�I~]6!�z(�?�~xe՛��U����W��i��m��ի�6>��p[�&y���k�$
�1�c����;p�4hU� �>+-_�����,��/O�M��Pj�ps����k$��H8��X��O"%C��X�$�̬wd0��,�����zȨ��f��p��\�'�JQ��>=�P����'�Z8T�^�Z� T}��7��l;�!�/f��G� i٬�`W8 ;0�<B��&RLDz��;-�Z��X�[yׅ�5t������J��b9%J�HyQ!��0�T�� ]�u����ʴ2�s�b(Սe�]bB�H�`�"�4S�*�P�r2%��H|��s�s��5l�Al[�7�Z��[�jP�_��
0F#֩)<�����j�_d�G�^2M-oKW�e�ް E4[��g���>+��ؾ�_4�g��Њ�a?������Xz"y���F3S���ʕ��Z<���yzR~/U��o=l��W�/U�b�&�m�W�-��nf-��IQ�.�e��W3EV?lȑ�S�*.�Yv�g�`Ri�5]��l���e�YZ-LB�17���w�K5?�|�.]����쪢������9
�O�`x����� �I%ѸIB��}��+U��Я
L���M���̯��@Ah�t}�fFH�C�ｾu�p���94��y &~�g�_�S�&��l�dU�oZA��Q�ݥ���E��~_�%^$�*G���tNe�F1�s��Y2����B#�WE��`e�Dx�� ѹs��~ /)��L�Q��	F�T�
��{&]�8Ƃ����L�����̢;%���{%x[<�&sryz��6z���A+/Ρwo���@%5���%;�b��<hU����Z,**ꜘ��`�����/�U5�جD����D�x�._��aG��Ϙ���7jce�4v?�p�
�-F�Hx%3)|ͤ��ܽ�U0�璀��ږ��jg׭��Q��,��Y.�Y�LS�2]�A׵�������]���������"0�
r6��);х�7��P�/^�8
��h�Ù:&("�=B{��N���_)�7#����^�N��wXxT����r�O�kk�r�M��cΗ
<9*�5=�?G�Ӝ1�Br�F�W·"~ڥ�K&��k��y$��1)�$V%3�t�U5�����^�[�vf	�e<�7��q�YFȤ��Ck'���\%���+,|��?�u�#.~ҳ�D?wOEu�s��zשּՃ�A0c1��ʪ�����ӱ��!V>���E45hԬAo3��DI��MG���g�Z����L�b9P�\w��}K+��d�$���'E��"w��T�&�-@<0~���]k�}t�;��@7-��s>���G
�bmt�ny�^����$JK�2�F�P�q6���\`Ь��M&Ճ	��S���R����~TΟA�����S!v۷�Q|�hjq�AE�a�љ��p����k@�گ��-��>���!!k���	���3���%��:������8��&�z�"�ԓ���*+WOm��h�	��h�?ٮ:�#<�j�}��e)u]50���
��)�yEzp��'�04�� Ț��z-I�ƜYBQG{��i�FcyqI��B���b��ԑ�cQ�Z1�ssssyKs3�y|������T��AM⏯��r�	,1��x� 2�وzi���l�t�v��:4�ࢗ��mO�^M� 7�;!�	�+� �� Lj^���i����q��.&@Nc����b��l�x&�I�h��I��/�$��I���4�L��(��Y�I8_c��c~c�t�~ru��TM$F)#t��'s���WDm���)KN��]��v n�Q$=¨W�  �U��S�W(�����;l ,T2l^Kdr����/B���:TLSy\�w�tG�����<y �x)���+�s^�-mĶ�cI�?�R���Z�@7�����@K��$=�A�}Ԙ#��5h>}�Q��b�-���V>Fo�~叜ęS��ט�����U$./S�WIz�������k�Bkk�K.�	ul^���?FJ�c��ʿ/�D�i��J�Jt�Tɩ�0�#��m�֌TC^����f�ASL�b�~qHJkby��|Y�S_�mll�9��k��TalX�P���^7��*�-V7b��{�30H�6���Ӆ�ey��R����˖��s�f��|7�{:��cd`�;�O�I$��]q%RM�������ĈK��"Uʾx;�g����:��i���H���^_(�kaGܐ���[Ĥ_�ȩZ�@�!�����qC8}�9�,�����Pr!�K��7�Y=�n�,�`��b� 9�?���$��?+�ࢦ�P����eD�Q'8�6bw7_�P��6�ar�g/�{����W�sZ�οŗ]�zѬx28=[�6��ݥLk]uJ-���"�V	#q��䗊@_y>�)�0�f).�@*�H�ob|yQ4�^@ ��ߐ|=��hPJ��0��X4�l;��������M�򡉉��n��{�_����u�qyy��M���]Y��b�T)l�o�p�v�����Q��C=��i��H�����S�"#SQ:��%�U��?;�NaP����G ��#����m�M��L�w;���NB��u�<���\�*�ۉ�703��(&�Q�Q��,��cą����+���<�������K\-� "b�v7ŰSb2 bK~�rb����g$�Ě���Z��	&EEu��3���ՏA�>����J|.&+�򔠨k�+A%�͝� ��ऌ�|#�+�'���`L�M.#�^�r�K�Q�y��}�Vߛ�u��������{��@%9Ɣ1�ϟ�gJ7��$�-�Ʈ�9=��"5走㆜w#��}U(q�_*��mx��2���*�uR��1���H��zҭ\F����s��	�$1v���"*+��jvѯ�Q��gD����?�NI�sx�>�����0#{��Y�S�iwc��ϝ��h`U�.e�#�Ӡ�A|F�ճ���J���g�Z�A��(������r#EY	�V�|$a!����HFtx���c�ۣ �Ns���~�g�O./�JA�PS$
��x��R�F��#\�x�?�v�ԡ
�(���)ic�~䠈��1�U�����+�K���?�l�#�ND����@ٓ*%�4��Z1��B!�`�ܓ�b=5S��o/�/+�Q�����֖�32Rk����P����1<���G�	\0ц�G!HJ����;����g�9H�ndLX+:���^{�z�.�62����l�-��,��&�Q[t �07T~�OK�#Ϙ;����Sc���^�}6Ϯ/� ����Cg1����;���<����T�:1r;%�$������5K� 	+�4]�.����?fOQ?�z}��`�x�t�]�њ.��y����g�N�	��T~?�6���ڞTBV�1t+x`�L��Ĉɶ75���	���m��\�{�jkkӺ	��(��"� Eb,�=3�Q�F���\�=˵��#�}JHL^��A���ؠ�U�q]E.]� �?E��b#��H�����i��0�����LǚD�����$J�o����)0܈�ƦI"�˚Y0�	3~O�L�݋�9��g����3p��\Ds��aMø� r�2)��?1 ޽�$#�}T��Y�A�
�,@qj���$�G[��|0�BD�"w���Plem����2�/�'(#3S���:1��}zߠ��S�2���0���� <G^y{i9�P��lɜ�э%N�W]!{f�{����Z�*�d���F�(I~�.ǼZf{fAN��d�Ahi.;`��A5,�m�654���) <V�ަ�U��K����x����`�VA��/Y頥R�+Ml�v��0B��'�8�3���zsm�������a�=unjZ�pf?PM�9����Cl��XߓG��>ro��a�r��0`����ub&��2qV�I��?��C���fLb"����,���"�+���
)�d|��H$~��.mB4߻i9����I��R)Q@U�vJ� WÏu2��-�V�&�g>v�Y7V�$�M=8���S��rh@fPo*<
��1�`�d�
#�SPԎ���#���h!����A���!N�Ur�K��a��*���J�-�r)SWw �,N������|	H�c�Q���J՞��f�)�i�{����R�3d���F��Q�t��\`
���*��><�|�0
�y�P�M�݉��qݟY�n#pg/���$����-���}x�+K���M���BѮ� �yuk+.����Ep�a Y���,�{����'����0�yd�%}Mʹ���p~�����<�>� ]��:*��~Y����J�,�;wj��4�@�%�-�;\o}�İ�r�������{�����	k���n������v_���|2+'gAt\4Hj��e?���a�8��kO�=Z��[e�R�����s�����3c'�ȡHO��~���}͑���%96.fo_c��x�S2��j��A$<VTDU�ܬ�v�0B����aA_O�(�F������^:m[p��4#9�5ſ4���r�$nΦ�q,3��D7TÝ��BJ�|7�J��-�B��rE�pը�D~���p5LB��GD������n���.����4Z�TL��B�Z:���h<����6Ҿ���E�֖�k�/�����1�iBe/+�K�HP�vHp��bHE3T̅�h�mY#����ljjr=Dh��;�a�mw����FFE�:��٬kl4!!"*�V���mZҫ ���o0��C[A���,3FGK{X]��ݝv������q{c�CBџ<"r�;�@�$���]�E/�b�ս���@��D]��uA06�������uw�?����̓>- %&%}�VZ} -����%~����g��5mg5�J�����m7B�����g*-QTV��seL����I�%=f�-���o�s~�u���"X�φ>�{�顑�kSeM���dHQ��������
sCg���]Ɩ����*�^�g�����w]dd�7�I�í��_��e�0I	�RU`"���s�#av�1:���K����bM�@���{�~&`��j�����Ch�<E]��d;�?�Tͮ�����Uge��+Zp�����������Ù��[��v��hG������S�fo���za��G���_��߻�I]IW�6m|}I�4�:����g��ó��U���&�?�m-W*2y\����
��@B�f�/�ͫ>�75Ř�D�,\�Ҡ�������O���������d�)ǒ
�+��������k��. �����9���b�h�'$$P��ݑjh�w�::����H��\\4;x>�/�_��(&Z�cD�)��N\,,�O����qt�����{O�9?�M�?�j`�����g*�«��6Պ��ؼ7�������������ƈ�"8�g7\�a�%�i��ӧ�V����F��gE�rc�4L�����>՗>$�����!�m��#��~o%$�Ow5����w�b�"^XB���MM�NVZ�!A{I�M---͂�喑�h�|�cU�mmm�EIO\���݇B^.VV�eUUjzO������d�����p 9HK�,=����Q9���H��A;�|������^�Ge���v>t#� ZZ%}�P������5�FYh�����Y�+��S4�CW�<�=�4J�*k�}�"G�"'B���k��op	m�S�Ϸ�H�+/��f�
�Kԗ��J_+++U7�%9����p�~Xu$s�8���6}'lՁ�T/��z}4�:qc�����l]�>d�6��d1!r�����g~<��|b���i��J7�Cx�����;�hr|
w��?����:�����ӭ8j<��HW���q��-�y�.m=���j�//�[}-�h�W`�b�|��c���&Q�i+�4�Jr�P���������i��/mJ��.�:�W\2l���?����c�_�^xfm]q�8YZ~m#60WS_�I��m���!ed�zN������w�	SK3t���ѱ+&f�����]������lA�x�;jB��1]E��z��^��n|;o[j�ogw7݇y�)��;�#mCb��b	n���Դ�6"��%LϞ`�sJik�Ք��հ�5�ҘN���rH</��A�����`�V�F��%.���1P���~r[�A��F(�������q3��~�2��2n�(_�?;�J��"4�@hY��ST|-[=]�����p����f��4e��*��[�67+�p�kSD���@@�K"�kJ��.��^���\�d��-jE���x'2E�sP�?�۴��ԉ0��+>���l�eBz8�d���_���N��陡�Z��?9$7<��}��C��w��r�6�48$ע��1����e�+�A����M����Iu������og�o�y��666���=���i�q$��sKj[������x�]�hE��۪m1�<R�c�	��*���{�h�K�F����Kk��OІ��` �N����
�,���E��񾍍���ɬ�&��Q:::����`bAǠz�{WW��(�{p�$o����|8pU�qd��O�kb�G�m<ƀ+E_OG�*��[�,���Եm:�+���P��.;�e�\��>w2���=\F���s'�!6����l��\y�HB;.<�+jg�ҧ������-�:"БH�V&��e;�y/8��k��?���
%xcu�m������Wfg���8��o �x˺\�s\�wL�/���>�Z�y�"������]������Nw�&�¦�[V���gum��|��M{?]$��ڣ,�\Ώ�OmPR~_�MA @^sSg��K�k�]�����[���椙���p���*���0��MJ^��$2c��}�{��gQU��yݷݪWU�p�aU8YX\|�n�����b�l=�a���,��WVV4����P��'@wȄ�#S������IY���((�8�q�h���^׿g���0UG�3��ſ������kg�9����blxy�����^�
�>rt�`�������K����S���v����6A��0y��璐����3�k��a���o-hRnf�$q�Z��٣��OYW����}�Ȩ���$��`�eJ��Q%��q��v��Z�~5�P�U�/���q�}�"8p�H���F�8�-xKG[{n��&�B�}�ut����65++fh�.'%E}��������v���?�gd�44�C�.�0�7IÛ>�1Q����Z�ٹ�s�h�_KAq�'��c�k��ogS�����/�P]�[^�5N��������(v}�<�?l�{xxH{xH-�������O��Ίȭ�������G��u��)��P|_������6g�wK0��h`��oB߹�+�* ���@D��r��^Y��m�u�2@�����3�Dˍo
p�<��}���r�ȢE��:�FNp����4a�S7	�+.��i�P�dN�u����h<�k�d�5@^��׏0�����|���vgC^����MdO",�������+�"A%�}rbB�'�x$�x�o�gv�����q���G\,�W:�1����ٞ��%%/��G�h�?^ 	8Q����?M����eM0{e��v�x��������I���J�N�<��͇
\�J{ylRbFb�,**��8���r��Sje�2�~�Qv�����n?!XU��f�j<����%�N��Ɗ��#�E��ZY��ʴ�u$�	�\ ,�`}s�s�S�&"X6淽j�YeddT"��1�\�3���*eee-L	��ߍ���}��Ny��o~}5g?�&��h�G_Y�9����b���Sc;��C?"�`W}�+��'B��Ƨ��`۰9����[Rk�h-T9i�ຍ��,^��םͤ�"A�~� �uqv{^�pz�m/���������&jy˄�����\�dgw�
����󐅖��8�4�N6W���Ֆ�f`�u��6Xi���;ᖡ��80P� A�].�o���N]��\m�� ���Z�s���X{�������\!f$2�PR�`@���������V��\��+!����.��Fj��n��V��#P~Á��
 Tx��Ӆ���à��9���� �(+��kb�O����Ĭ�P=��H�嬮��GSU�ARE�`X����8� d���fn�����W2&���1���w+*oO�b�4 �N�8k����1m �jdɗ48���.��ݠ� #�LL�*^�q�H^I���! �-ϳ����fs��k��#B�����b�.�L�@�E)J�ˑ�)o�9�G{�1�Y+Μ���LO���7a��y�����->m���M�F������%�/��e�"@5��k:��	�i�Ě&�2�zz򼪮��m�_�]|�^�����\�O!�����iʅ�:�`<<=W,�R5TU�1c��+pcc��n�����Ա��{8a]�BA�Rݲ�*�ݙO0l�T3g�]U��j�F������v_/�]9߷����+���`-T ���-��t�ь	�oc~�.�V�����P"�+��o����f���Y|���m�ӆ�]L�49A�V�;��X���f袾5�JC>.*�cy��6\�΢|}}���S pk�t�C5J��� �o`l�m�ho֏�������5���6�ͷ|Poh�9>~��5b�G�.a_�,e�ot�T��Wl�M�k]-7�ܧh	iAG�2(4b���#f�_\�����L$�J���U
D�-����޹:=;�qM_]D�:�ST�?])�;��x�wv4D��B��zV))�G��(;㷭O�����_�A�:��G�S�KQ"��B�tt�_�ݧ��W�'��<����F	v`�������=%���Q�������VC�l��g���cE��aT����͂�~�+C�*M�5�|��9Ͻ��>&T$$v�h(dy�_:���w$C���Z���e�`'K��z��|���fK}��7AAI��e՚FR���@#[W�I�u]��*�:X�ߧ���<v�����փI�j��.��ɓ�Ԍ�:��Z��f3%�p��m�����t�{W�*�ߴ��`��QȤ��G�� ��O�Q����Y	�U���<fc�2��/om���8���H*}��Һ�����x�Q��,/o�WY#�'��r������o�؅�dt��
���H��חǫ�9��b�䬷�������[ۛ;k�V�5� �����չ9Q^��ԟg��YFX̦����<Y�mS�YŬD��t~�R��~�=qs���P����'t4��N��7h����&?N��,1nlb��#��䏌��nn�tttXJ�X�����r�"#X�'�@p����I{{{�Bq3"3��ӥ��[��$a�SS[���:���X���LÉ�	�3.n򖺦&<l��8X%R������)�������Q[�4�=��QQ�,�.)��޴��/�hm��ơ������CWK�'d���S{�����ΗrSf��Zn��)��j�{�ա�B�;��(�x��/���Æ �`5.;׀gkt4�	'η���U�����|�`���5X3�4޵ytW/�����U `b*AP~,��dbh��S�V��$_�N)x:�F+Ȣ)�����\�����uv����P���hX5b��sb����]����n���I("{e��g[�R��&���v�
��#�{���^����yzD]�%gCh��3H3���iGK�����9��e*!�./���_5�`�jhh8��=���'��غj�L� _[[�A��n6յ-�u+�h����U�nkS�.ƿt��Wmd�><��@�aj��V���J�u���{.���Uȼ��������[sva��q{���ͯ�����j-k0|��}��AOx���*��	 �aa�+�x��l����>Ͽ?4E���$q� �:�����N^��d���K�o߾��3O?r��=o�u\�Ki(�Ў܋|6��JX;��m4suăp5�.�h���z�tힾ�6�'v���W��!!����J��3��(vuu��V_�%��00--���/P����ն���k�^�jA�v�u�i9�?A���>��)>����$�$�8�YX�ٹx^����-?/,���s���UV�-*u�6�Ѡ��{�����nq��Q`RR��N�������J[[ڬe�ql�#�������#�i�)-���P�
l-������볏���A��*����\2vu�@���S�Y9���a`g7�����o?�kfn^�mF��B{͆��
"��w�(t]��7����Q�� hna=:�yp��X�Xxc-��J�4�G��2c�����;��*v���{	��ń�{^i�9�:{]_�E��k���sH����o* ���Ѣ���вm[��l�뫯>��d`��TϺ��2�҄�-�O��
�[S�
2Q�^�	*^
4���h�Q��Oݐ�{ͳy�N7��?X����J�Rh9��g��+�@��]���GG^�\]����?xt���������e�@��5��%-�-.?.��Ɗ�:����7�j�pģ��|��������ʱE������2�%in�������􄷇����֖���#36ր��ե���/� !jl\�o�	k�S����l��wdu���y������Rqq�P� I�/�p�A�}�˦��a���j�9Ϊoܶf�� ������p������|�+^je�?���l���"�¿���Z�љ��ۋ���x3l�d�B���,/��5~e��˙0�J��f�÷s����Q_g��
]<wPyrv����pL$A��N"걠@r�����U��j��>���h��o�������|M��S�>y{Y5i���o: t������,QbcM
^ǁ#�QhC{�]�44tMVf��n���=Y�{W<}��Ǘ���������F�b��eg�z{:���Xd�N����;�<E��'�{����v*;0�O>�hgT���9O�|\���Eꙓ}<h)!�H��9EDG���XY�o3��[��q;��z�5�JMK�LFTlc%����T^E%��5�:�1�y�~�y=ǒx�}�X��y�EK��tS�w�ᎄ�ZA]������M�F2>9���O+��B�C����w��ÿ��s\ޠ:שh�$\���u<e9#^Lq���G�WG���#7�����k�Q��V��F$�3�o_se��H&���Wg�o�s�;�(���;ݝL@�!�!)}�m�e�#P��.�L����+EJ��)���)��2�QT*!��i�Ό��ˇ��~N9�����)V�m�+2:8mev���[kw�����\6��N�����y���C�F8앫�b������-��r�}%����o�\��Q~%6��~w�}	���̘3N�U"ll��[�dh����G�ݾǺe��-���ׯ�>������6���4���d%���4�J_z;�ll詰6h���l/�uu�͗�I�'�N*I�{<��՗��BC�fg�3y\��H~*G�Lᦎ7�n6(��D��%C/�����4>ϻ���0F'3�eR��6̪
�OM���8o�Vq����n"h&>s������zy�h*�󰊂�"� �`��x(��P-2[&7u���nmi����|I�濱�ϯ����o��`QK�Ι�q�X��t	���y��a�W׻�`����-�CX
�?�����ڽ�>�ۜ�?��T	��!�_�U@DB�ۮ�\ml�8�i�¼N%�N��&^��`i�:��OI�M�����)����"��t�C�s&��-��Ј�}�N]�1�@�O��S1�p��)�{_�P�$3^������&J��w��mն�j�p?/!"N>��0��R�y��~IĤ���kǅTS[ԉ�:���ꗕ;ٜ�W�ޤL���+�b�B�ϩ���,,����7�%�tQ+��5K���\��k�e�f^��x��;3;���o��V}���Q�]��{C5Tz��մ22t�U[�����=��-n����tK,<=�L��^���6�NOOYE�~�L�y=P5C����K�2q�H�Hx��'߭.`�:JLL�6wR6�}��YRB�WS���|�E���F�3q��$�1/(((�
�����$���e�����km)9��e�a.��O��@�V�326v��O��l{A}/�B�g����J��np�����)000$M��~�쉣�Ĥ���;�
{���?��yAG��./ή��Ҧ�e�v݉邃�B ��v�ѥ�����N4�F�tS���4��"�Ēv����qr�I���/-.҂k&Qn)tv~>���	L	3���P�!8��� �稹�n!C� ��M?Un�m��,Ĩ�Ԏz�f��E��x�h�g���d�����ܙ�u�cq����s(��v2qL�+8qa7�Mՠt�*ד��#;߼�WIo/��N=&�?�B�~I��w8�<(��/	����k���Zd}sX���D��������������֤�����+�g��j5�d����<dN��S0����n����ŀ� ���外�>���b$?���y�M]}��e�ܪ��r��+Ѻ.}���P�B\t�'���$d��WF��slA^^���|��Ä������4��.�g�%�/U5�K�����㮠��v���+Tfm<���uwr:��¡��T�o���#37�pZ�^��wjU(h^���f�wa���Z�˭|R�"����/�
e56�r�
�liY:t�(ӧ��2x8��
wh:�y�m>�JI1�R��:��_����Y���$�#!����3$^�� ���������$�_oZ^.�gl�� }��D]���^�̖��"ڹ{��T;�Yɡg��Y�C�(�n�I�Z"6&.v�������b���O�j�^r���u��l6������S��ɺ�$O��ǅ�ɬ���Ħ���ee����ʅ���Fu�d�c����{�չ�]s���yxYޚn""��U�~�Z\	�����M�N�:I@����6�v��E>�����慂
ZN� ���ˋU��PK   ĺ�Xq#Q��  Ț  /   images/bb187b5d-1fc4-4a4e-a882-8dc83b4f659e.png�zW%�u�[S��d۶9q�mc�o�m7�M�&�fs�]�߳ޯ��9��v���42""����
��p7�QΕ���p��v��@��C�ң�C@dy�J��y�w��ُ{k��	�n�ct�c��^�%�k��¡U���)%2Sࡥ�h����"�c�D�@$�)cR�lYؒa�CT�6�MW=ߟ��*}{+�ms�.�+�Tk4L��}�Z���U������+]�ע���f��a������J�q[*��N����8:�����Boq��_=y=_�_��ݟ�g/7�s�Ұ�B���ؔ������6��{�?��_��`�Q^<���4�6�(������7(��N���v�[�M�,��9��-y��}�|��I_��S�:�7�c�{�;>��rFV���g߾J

"�5H��]|�ɡ�gtQ���z8pG�����~Z�^�%��y�
}P%��9i����q�k��]s�|,�${����u?��%+Ξ�_sp�ޮ������mfp;;��!`�Ä��N���m�ʊ�<!��N�=H���^o�q��h���hm6��"�U����ãgY0{(�:��><:+��yq �	�_Tc��H��j��WQ�
�q�/���e�T��bf�7�����[����6�?O����P��:���w�O=؟v���p�%75���h�
�E(�?!`�բ�"}��S]w
9`��a0aL��ה?��0�w�����'� =�����(�1ꟜѬ��2�������xI	�J\'e$�"��#�C{�KJ[Cv
�=p�?�<E�)�`M���I��lʞ���zA������ߧ���Pg��ߨx�����׍���J`����� m!��O�e���� $������4V�pF���͇�zI~���b��<UU���G쾽���BT��}8$�~�{se�%�ۯK�T}�81�B�s;{�ݚ��#	Z��'����J�X�U>���pU���qd��`a���׶›��iw\;<j�j}}����Q��������M�#�������U�G-��|WC��%=�y|�#��g^��p ~*�.o^�jnЋ��"�|`p�ˉ?�	�0��jO�q��23		��?�sx:���I�Vϊr�_Ð��R���ؘ��+�V�T�`f��B�=J��l�.$u�&O�ё`�t��?��ɰ�zLYѴ������+�d���hn�f襣#fH�ZvL�����VN}yPnĊ/˅vx����a���v՞�o�O�<��� ��a�
ۥ����^p����x�=����d���ۗ����ba
�g?0`'ᳱ��I����2|�F9���1�䵣Z=�?U��+ݙ�\ 7�3���݇���߶
���Is�kS[���s-����ޫ�[��/����|��BRW4(]�t�,y]�e�rw�cɅ�;sq�hw�$��3�u&� �@PXX�����G�UoǪC�����J�c����uM�o'n�͝���^8����P
=ƍ{ۄ���k�&����w�*8?r�a{����t�Zi\E����Yy�]��z��7h](׌寃����1����G'r�!��-cXm�QAo�{��֭oM�Xsиx��O,�]{fd\�qSW>�79n�n$)��}�s:�2:�n�?�o�,�4�i�ٯ�-�퍍��;:P��ٱÚ�z���[��Ao̝�-1��ds�c�ұ�Ҭo�){ȡ�mw2���|c��̎�"�4�%��]��n��Ydp!/��J�Κi77�X� Y�KKw��6��7��"!6��|.<}�ӟ=��=Φ����W�)`P���)� �����$�yT��&��Kk��%KK98��3�6^'(���Q��]��KHjesv��x�,��͍�o��G�-"N���
b/�L&�V�P}����r~bM��V���N�$�[p�u�W�_T��:�ww��f6cS�G���������ݝ����?ꓟ�J�*3��|;'I��b�c���v��]��m��H"|���~K���8S�Q0��ɱ����~���8]�u������Ϥ����;���xkA:���:B�����K��O1X�÷��^	�a�t%����sn"a����i��f}�K8t�o��S��XhB�d�
Y5*����BB$�":��<8w��D�=O�2�yx\��G�I$����x�/ہD��I�7Z�Z��H��>�E�O[$-���3Na$�C���8����#(df��f�Y>�-`. 5���b�0�s���6o5~m��,\ay���2`�Bk��d��y4W��AܙX~�S��?[�2�{�tH}�e�l��Y�j1�`�������:��c��eh��R!iV��rB������MH����)}�ygo���~5}�0>>..�S2�I�M��`<9�i��s&/���������=w����>sN^^mkg˺^�~�z�w T����pN(L��DV�m+m���W&���_F�����VA>>���Ws�_�J���˭�'�}����������,*�����P�gؕxۄ��q���|]��i��j����w}�v���"�%'}�s�p��J~�||-r�?�1N�������q���I�%"	覸��}���뇦�B������-�3q=!5����/��_;�]�G!���v[���d��_����7�m��.V�H)A^����9'И)4�x��n���~5�u�a�ھO5�ݲ�i<�z��qix�vSRdf������8y�d.�X��E%~߁7���&�\^u�5������/�����u17W�-�jc�%���ˌR��8A�<��RYTΈս�͊�S�ݷk�,�ux��_�nH�'kVD{�̅��p/��8�.����+b�R|q��(ߋ�ȓ��8J�Y�ܰ�?κ���_|0��o}�h���7���ŕ����{�of��'�)�\5�\轸�dU�.�zǫ���ՍKK�Ԁ��Q���V0�xl�9�<�
aZh��!�Q`�G�P�@"6k�,��>� 
g�*�k��@�rm���7�֤��{z�O������~�2����͌|`�+I*�BL�|}\}��	�[�����,������&9���ه�5L��%����\���o"Mq�=�<U<�!�s�)�G�w�5
vX��ڵ�v#���M��#x	-�Dw�?'��D�(�8�C~+|���`n�ni�}����Ԙ��Q����p���n�D���V�p�
��xE���G��Tkk(�c�x�P5(���D����Wqt=.��������)th��8U�d�E-���a�'��l��-f�յ�F�)B~WJ��!B
��埥9ct :۝آh�e�nû[�
�b*M�\�a��P���n����������Zl�T{����f�DCB���}�����sՖ'�����l�H�����Tj�A%㱗H��f),k��))7[�Ҩǈ4Hz��>��a=,d<-TJ��ċ���/,�qli����� �+�պ̗M{���]���e`��K�Q�S��wY�Fܙ�W,��ʠ/�K�B�m;x:��+�?#N���i�\`6)5�~�����t��ě�n{��h"4kd���7���ɸ�)�������n�
:�T�2����^Q������8͎U�{H�մeifb��|��Tc�j������W�c��Ɠ�U��-��\���`��Ϗx�W��4�b{�A}�Zk���!
��g#�G|Qά.�?���;�:x}r	⺍�85�I�?Y�EN
�W��g!������WE��Y�1^3F�2�(/�(ф�,�w��7����SO?~��JFG�ڍR�@�����O�>p3��m�VO�}�x,@"�eT�e�H��s��+?E�Vo��u9��5�� LT^1
?3@���k�x���i��uj&�6_�x����$���NŬi���d���wO`���r"�v�(�p���H�����^QQqÎV̸A��8���q�9|	�]��>1���z��<���ub�}g�:r�s[�<Sh����j�������w�w~����l�&�Y��yz��{%v�m��,�pgZ���l�:(�|���yM���7t*%���0X�xE-�8^�� ��fc�z{��rIf���IrQ�xʶF)���ȣJS���9.2l���hߞ�?N��mo�D>
�t�����?��h�����A1�ZWg�M���BA,gps��DY%iȮk����GLCD���=.YY�
%޾E�N�3��a0Na]cjݳDcxe9��/��S��\��Ŵ���x����0�{P��XL_}9<���~�������u���<�v���pK}�99���M,��Nl�v^��2W[����D����q�
�E�2eC�~cR@/S�!���r5� K�!�toB�5�3��"G�h5�M�0eϛMK��+�G��<�l �g�ws�� �ꇶ�m���w�m1xw��W6��ezq6�-��0�sȳ�����'�ji�h��J�����J���ZA�N���>�%��E@�g�c��a��9��7���y�>=Vc6�����{{vE� �<�~G�>J�v�HOLLH�t�)-|�T���Ĺl�5��1��lgL���=�>O����|SO�+B�7������	���u�W�y'��إ�k�Zg:D�
�d�Df���B���Y��vM :0<B�4+�:�?�yZ�C�H���&ɀ*���?XU�\38t$�Y,���������և�-��4���Eu�����A�*���=�6|��sCD��%6�&��g���!�$��2*xEЎ�J���
������F��Q��������)m�X��*�e�?�s%!�טM��9e�jN��z��њ��hz"���]��ʏ,�ʢv�3��:r��7�f�##���g�N`���ý������A�T5�1�����+y~G��q�I������9y�\��"���purE��~��5F�l����o�r4�S9�u��p�^z/>ykM�.����snp�L�r�n���B��9�{yBR��c]���/��LF��	��~c����5�,F�y_H{m~dc1Ź�!�|Ԫ$�aW2��N�e/x�����MPx���)�>����U�c�ؘF�����ro��|�Gb)/�IT�mG�F;
y��sz���� ��zl��|�0���~)�u�&��}+D��ه�	pm��=3LlM|����ymF�+8/#�z����|��)��J~L,�@p�h���I̳-��`wQ�BT�*�[{����ڍ:���~�_v�av+?��53�-��\T����Ͳ|�<�*�~c�^��PxL��d'���o|s�a�H��0�*2���_��� �#�58
�{����a����S��R]^�L�fG�������M��W��5�*���z.�$r�޳�ì���bsoB�ہ2�E�v�(Rp�u�7��ǌ��?슇+e�
1Ow=��LA�����RGb�F"��Wq=�P��.��#���WCR�������e0��a�UƊ��i^����o�
[UŽC��H;���x_�&�*}��[ն��)���{]#�1S|�f[<�h"���S�.�F4怄���n0O�� T��L\��v���W��"{�Ա�I$����R�{�c�9�����N��x��)B�����}��b(@p�5Lװ���=����6�NƟ�38)q�� =W�煀iEhp���t�y�_�bLA�����~��ś%�Upm�o~kv���d�S ������
$���u��'?�����,2+h��o�a����j�M�O�B�e3=�_w\�C�l�s�����9�.9p���d����$x�eM90/&=:7{��oo�ڶ��>��.l�򂼫@{�۟s7����o��t�5��Y&	c;�Z�8&t)��W&[����&@�QI��?����;ƖR,�த���� q���q'}S9���ƂF����O!���͞�n�??[x�6�Xo��d�}���C�0<?z���S�|���6�q����`�:�w�UY���L_����I�&n�C����&Sp���|OG/�M�v��my<��#E����l��ڎ��׮�ĳv��&�|@��7Rg�i�}���N�3���r�B�j�U�"��b��7u�.���8��E?�h�x�.�E����l�f�y���q�����@: $�}-����М����B���:���C@�kd���˃QQW/����*כZ�@U��� 6�r��|YٰP��e �����U4�w�����m��c=W/z?~dѻ���L���We���6h��y ������ς��F\$�m�b��ġ*:�4�j�_�o��j�����u꾲�}�s���0���#'�Ӣ�1'���x�c�T�/��ń��x�@��� .a\Թ���)�G���@�Qg�����J��I]��*l��ezQ�8&�x4��<(����d�Ǹ#T��3_�V@և��8�♅n�ú�;��
Β�@�� ����?G���L,��T�ڜ�h�Y9\h��X�ѻv�w���v�"R�I��7__'d��A*i0�S���]����6}������P(����鱭�>��sǞ�pd^Ŵfa�8)�j@D?7�ey"��t(r�0P ��$��|�}�A:�ϡ	9����H�Z�B��n��j-���z����Ֆ`���0|#��*�)�������+|���A(U6~�-���h�~�����myP�םL0<mf�͹sF ��g���c@3�����J ݋H�����^ �x$�^6V�l��0g����<a�Yv��U�DN�a���9<��;����-e�j��g
82�f�������8��:��4Dm%�Y�wZv�>��y@?vNNzE��b�`��(rOwC����J����	9p$�io����}P�HK&�*l���<�����L=��Y)��� �d#/�����T S�3/�� ^�����߸��W3��Îf%oT!W���l	E��r�&Gh���9�f�ȟ6C�pg�
�v9��jn�x_��Q�������O�W�-�?�����Z�_bJ���*��+`d���7��H��I��;��,��*x=�w�%ԣ��<�<���f��=�������;��%y�[CU���{�R1���fy�j'N)B|"�]M���U\�+�dw��,x�;�5~�8����4
:)���2"o��H�po?qR�-5�f0fX�|���z�W�QD7B�`E����o�T�mux��H�bG��|Z�d�;����N�u��oawO�/,���Sƍ�%!�L
��0�%���n�8����i�Py���8Y���D�(ρ��	m�v\�1�|hM��U�Y+	F%�^��F�S/��)c�Sy�C��3�ix��eH&20i2 �Ę���h�`f5@�=�����BOd?Lm8��܃ml��G����-�܌�˸<A�>k���r�t�9���ʭ[P��=~�_e3�gBr�Ǜ�jNd=>#�e7��N
$�,B�n>S�-]���23k�OY;��X,�l�h�_�DB��������4d&j��&���^������j:d�g/�%K?�]�V���C&i;"�E"j3��X�AsPDʓK THtv���ձcf8�./�ٌ��)Qz^݋hVD�,Y������#m����5����7�5_)����vǃٞ�B�)g~�T>����w��e�fH����ĀbK7)��F�*M�B`R��x���Jթ����SK~^9	��,���>��h��FL�W�v�CaߦBл)�6g���3��Q[�QѼ��.(����V�BXe£��kt�Ϟ�g��ܷ�<&��h�c�&45�u�,8ʻ��p��9��GK����a�(��"M���{w�Qc��$��W�8u�HR�ʻ�r1fkTib��Fvm��k��G�z7;� F�x��D�=�V$R���zMx�&~��ՇU�q��,����l/�'sG���8۷[�w.�t"iԸ�Kn���rhѢ2�������ѹk�Ԓ�F
5����\��_d�wڬ_���+��� ��`�j	9o,TC��B�)�����x�XJ#N�["��l�|����d�f��1�5&��W�o7=n�ݒ�zdŷ��G���ء��ڐ��|��s�Ǩ��tܛ��mo��x�S�+oyg�30Y\�F^�wbRB:�w��o�D?����'��*O'��T(c\u�Ʋ^�Hz좐O4�f^���ڛ*g��Ӛ�<ug3u�q�MA��Y��
BR?��6�3o�W�c��e�K���d��p�|��<�Z
�B�9Ӎ�zuI)�[V0b+��b.8l�Z�������/��n;�u���*�$�	�q�ב*�ܿ��-{ׇ��v��+�l��-FXs�i���|_$w=���{7ʻ� �p��}������ǎ������qfY��L��UM˭�8������j�]}�Q;���Pޢ��W/
�y�>��Q�f��0�@�~*"8	5*~9<<VU��M�_}�Q2��-	]�;k0A�Bۢ�*W�p�Oy��(4գ��~m��ٵn�F��hp���N��D20����d1�h
]�hCB�k[J�l��]���k
G#B���tc����e�6=/���&�x��U���wV�Ǵ* ӭ�5�����ּ%y�C�`�������e'�g$�����HՆ���D!9g�?Q���D�o�	�3i��V]��fD���F�f��~�����kZ��*߂o4x¡�l?�U�l� uބZ��V<��	�^6BDq�����ُ3��GY���� Ee�6�mi��pP���.�
�6�0Cy0��LO�Iu��~%��R�&�f5�@e(�fc1��8#�7ɱ�~S��%�&� @�+���%��.�F��;�_�qC�_��g\a"�E&�È������2����S��x�k!�ݮ�����[w�x�ۈI듲���i֕3�_����-�r8��T>��AA���N�(���#H�F���:a��/4>�0�s���¶3&d蠽o��`���5,�F[>��$Z����Pt�3	�D�W���J�����F���_��e��P4�в��7���r��n�������و�;�ꝸr��b�d�t�3"ң�y4\�5����/���NN�R8��Xqm���LN�f^�rIʵ�5̸���"� H�gC�lwٿ�^��Al��N�z�D���9eM4�6lR�D*���ʝ>�](�8H*��� �~�����q^�9֜S�����*սC���$���7�%y���̼T�.�6�A<n�GR��w�ڙ7)�AA��ȳ��`L��S�J����������%��5d��֥��R3� �ML�#�ZG�a�7��vp���6�y]� ��!���9+�k.~���G��ˎ[B��£�43W�,����F��9Ԝ�ɭ7��1��Ɇ���OG��]��";���9�3B%g�m�q�-�Ϛ�o�ݱ�'r��v���ͨ��i��M��`���FVV�;aR���`?3e�
�#X

:G�B�����,|�QAO���{g��F[����Ҩ���Tf�0.Jn�B�M��E^�-��Ԅ�>"+/���?o��t3���]�3=�9����7�Z��}����k����
��ޝ���Y
\8v��%;�f�;���^�?�}�?��(Zβ�����q���Rl?c ��s�&h��N����%�aು�_]�h�u���l-K��F	���A�`�4u�����5N�4��b�����f�I���Wc���>��uQ��.`h!Q6��>��q���\��h�Mۤʛ�5A̄�*��s�k��ew^?���ө�Z��l8�R�C���e����g����4�s�q��j��2�V��"�iQH�(E�����Cl�c`��R���id�(ċ5ʩí$>�1j�R��z�QAmu^Vd�%�����F�8A<�$�zĝ{�����1s�~CR��-7g3�$0ʉ�<~�������0Ow��H�p	��b���!��V�P�q����\���ł��Ĉ�;9L[U	zg�jm ӱC��Un����mUחa�Z~?v�F�q
λ��������c?q��N�O<Ύ�����ޮ���t����`$?��R�_�	<M��=d�H��]S	n��V;D�bIH�|�&^Iܨ_��R�����k}Fbު�h����f�k58�h�\�Cz���ͨ����`�[n_����2f��?&o�z�Q���� o�����Q�qQ��Y�F��[n��# ��;�Gݔ�ɫ݃e�8���UZ�3ג��g/H�!�qTe��
��~4r�9���r�v�M�������y|����8�,pQ�_8����\�Ep$2���&v+��V٤!!�P��j�]E[
��
�����*I����,��ʪ����@q�|�H�b2f��+h0�lpE�q�̵����K�(�N< L��Y�C��]y46)�v�1]}�R�z*�)�2k���]�'=�w�T��c����_��-N�l��a�;[�+0L0�˞����	(�����L��rjZ%ksյ�PӛU�7_�m#���`�z{�~2�|�~0�߯����	�<<���T�#���qFX:JreU9}�h�~�}!pb@���G��g����
N�×�f��p��A�8yy��+l���ue��[w��[�2�rm�:�>Ɠ��9h.3qBo�%�В!��h7�/B�ػ��\���_���ݲ�p�U�kDՊR�^V����C�y��?d0�`9��Q�P�sH��� �4���H?����?�q��}-T4N�G�����}��ᛛ$�e�9���#���S<�f$)]�Z�� Œˇ�F�-�py%t�b���������p_+�L��L9^ܙ��!�岟ɹ���m�����5D�*�9i�š"���~��V���j���"��5f���hd���v�������@��9Y_�-�V��ů_�E)�4���uelc��q��Jw�x�r�� �0������C��� r�yt��C���x��Aζ����._.�� D5�w�[�Q�$X���`G�����yղ׺�p�U��d�P9Üąv4�v�)��4;���-*'?�r�n�Qf�ߥG���!^0�'�d5f. +"�h�+��ʊGj�bC��Y��Υ��Ի�fxs��Q�6�Zet ��(/���]|�#�c�"����z�F��4�-�4�~�_�"l; ��D��m�5�S$M��2Br�)�yk8&!e:�5���j7F�3C`�`�z���j�D�t{�#�h��Z�ۂ����?��,E�Ҧ��JlU������R�O��<��"'e՞t��h����'�5�ʻ'�Qw�ӜU0��=���6�m/��A��x�@B�/��䒶��)L�o����
T�jY���GV����w:�=]�`)�jy�*��ID���B1g�cS��!�72eO����<��v���X��P�&l�L�iݳO�����>/�P
r�+j)fܪ&����|�Y�:���"ߙ�]����g0BC�v����"��D���FVP�g$g�7z�� �Qͷ�30T&�9�495�K����ҫ�16y>�;�s�Q�l˨��HҎ��K�]����և6��>��g�&����a�B! %�y�]���B.�.����H�D���>������Cq0�M1�B�i�3a�a��?���'�^_��`�M���&�r�M�8)��')�P���E�/$�"����=���+�hB<躄5ξ��4�r����ow&��n�=��tEj/#*��e\J���/�M�LB����������Y&�������<��q=A�B��&��E���ي��8�@p�ZR��ˆ����3��'=�C^\[��0�U��ke�������2�=R���k݆i5��L7�lL��	��M�`����p04�Tf.\}�{:��7{L ��b���u3���IP��z����%�łɵ2������+����RH�Ӈ��KB7��Y"�L��.�.i�N�u��+��r3|�-5�Ȥ�$�½�^��#�p�r�k�~'}'j`ei\�4�O,�r� �d)��#ץ��	^1���F�?C��ͫq��������t�D���^wA�/ʙ91Y��{o�S��57��'V.�����.�n���$��Hu�%���V�8��o�|�;�ET����̪����x<Kuw��n�%&	�W�,��]��%��!���Kw���׺b���Q��Jx�D�'��%
}v�a���C��FP}6r2�L?F�u?��戂|�B�I��k�X24�)�`��D�[F=����vT{�'m��īU���)���#]�/�&��y]")d��M(������5�ٜe��[����~߸���'�q���d׋�&g�������J�v^�zD5�*|tV�Q̚sq���'U
�`���񘧲w�ͻU�T�4����]4�	�l���@�9-���/����2��r�*˾"*0ھq8�-f�8��Ϋ1�#����U|x�HY	����Ԭ�z�N/�8�1gd���Ŏ��=T�<:^�\���t��n$&jdD�r�@�[ҐG�}x=�'8�<,���~���"EPk`����<�R_�mF�������������d���Ժt��b��������nb���:?	@n.>O<{	T0�4e�ll�Bӏ>���GEq�Ė�z�̙-�xv���v�����&G9���`��8��=��bygd�?6��'�TMٝr �U��bv�z���}6��2e��|G��H�'�Y�i���Ȧ'���H�]gO
Ц.5Z��ӧ������L�؍z�������7F���:�����##(fk���8nl�c)��,[.�:�O�똋z!����P��dI�����~`��l����N��"��A`��'�d>�>���Ĭ¸�۷�g��{~�d����/MR�;�z��i ;Z�d^Z]����?���F��d#M���߀��iG`W}��@6�\�{�2����k�F�%/Kۯ�_g�{(Rt8� EUP_�x��0g�J��n��&�8�O)+��&Q@TRpH�����}�KbN]Vnq�e=��F"1�1�:�V~���6}Vέ]����٫EP:���c�$�/�E�)��:Q2�0M�V��`�qEn����3P�;j�
'�Ak��M��p���uYu3q�����D cN��N[�]�f\ a�ʊI�h��O��@k2��J/�����c��F�qLb?a��X>������-�
���Ն�<J��e����8#�q�X�Y~<���A2J�z/��f�U��b~�M/&�s�����}?�q���][;J+@��x���4ԛ�&�3����	:��(��W��*s���y���s�B%�8h�k2���b��~sL�~�Ɂ�-(�'��ң�?bw�}�'�p�m-_9N!�Vw,z9������bg��dQz�AZ��L�~�;�jQ��̬ʀ�]wG��O���+�y��{},LIR�d�M���콂���L���;b0�NAVNr����R�J�:-ֳF��]�9��)�;5��ކ*UH�1uڽfݭ~9d�D"�Z�'5��Y�&�63c�I#�"6&&%���L�"_߬��j�)�
��P<`�-pb���C,p6u���������i��):����eǗ�k���|���5S��A��{o2P�<_�q��ve�k`��?�����&^�sQ�<�����t`��m�r�2�剂�6g��#7[)�>b��k6�W��F��m5+*�؝s��s����s��)��$2"�K��a4�R�>��c�u��95&j�}�9����ju9H�kܘt��o{fci	�vN����Z����S��y�ҁ�NV��VY������$�DN�T��k��:5�`r���?�� �0A8�z���NF���͎[�ř�x��%�!ʜ��<k�S4�.$4]F����y��?�%3b��*�|� ��q[V"Z�.�^!�R~?��WN��Q��,B��c��b�t�7[�~i�������iN��L�l\���?��iD]�]��Tk8D����0�����=����/��4��r���d ����1:�X�[�������xm�C
8���PEB��o3�ͭ�Z�윘�7�+�api\�����+�f^�=+��HD:+$U�	J�GkI��H�P�'��=���S��ϣ����D5�w��!m�u��5c7O� ��z�9(�9��}Y:�t>���%:k.lE*�xY�8�y3��*�oz���S����4c��B�-��6(�t}�V<��Y/��9��9i�T��s���FB8L�V�8Ep���;E��{V��=��	��%��_:�tʺD�#Ky������.X4��p�xΨ��FX.�a��c+SW�
��#
�I�4�xlA��a��\[o	�S�s�X�����������u�"70�?�a�I�d;�g	� Vk"Wh�_�����B�>[%�{a۴�9$mM�"���7����v��̽�:��u^_�z�}s4ou��t$�]ʢ��^Fc�s$@aw�s���J����ΆrSߘx^�M�s+ݪ��j��1a��
�j�p��v�9���àt�j(H3��y��'��Y���,b+z���~�&ˎ7nfo��hz�%�#�xay]�6Ƨhz��Te}O"��(�<!?����H���n
�ɩ��|e�slz\ƍB/U�c�,(�
�C��/�?�}jLt2���i`��GE�Rڟ��0t�WD�ښ�wx#�Z]RVv��ߜ�����G�2����q��>5�(��&���A���N�#Ƿ���al��� �Z���)T�<9���PF��S��i�~CF��>̝ɝ��u�����K�+��r���x����T��
)�w�j`o��`9��
��f��h.�b���+��6��/.9 De!C7=����I���< �X��Ts�@�T؀ZI�)	VlaL_��s#R6�}�E`�0�XȔ�uۓ��h?���$�%��?�di�`���2\� �9<�	+%v7Dj5<GB�d�U���PN
��?zv�>W�\�FK)O�ac=+�?h���\6�qO[�1�
�������-:P��a1ޫ�ݿ�	�#����� {p���'�B��-�-Z�SG� 	55��Ԥ�+�q�2�	��N�d?�ei�������f�z~qcr�#�07���� �60a��s��`��l�VȀD���L��oV��X�.�rl#���۠�4,<q�NNr��|����aL��2�!C���/��ś��z~u���k5���KF�N���ِ��d^�Z����þG]g;,}�M�Ղ3i�D1����<��f��\� �_�l!�ș 8-���I���?�r��y=�W��%�,)�NY���?��@`�<w�������e�W�-k�����Z�gJ���3�b���x��/ѾA�4{vi�m�B-<x9���N�f�;��Q��8S��H,I�!�<b�awD� ���$9d��x.�w�o[@i���n������G8p�f��A�@�G<�\�;l-�Y=�y���T�BS�ĕ�u��L�tQ�4�x�Ŗ@�<VR��=r�m������'���ȃ�G#s/�l�W��W&OV]5�j�>�B(7)<ِ>�դ����L������ˀ�SO=�s��x�tQ`f�N�Y.j��J����X�q\tA�.��U,��G�h�H@Z�Gw8��'l���6�Z4�?0�M��gF�.����E!s��&�?���Qj�?�u�T9�{)m�q7�/Y2鱎RKYǙ�%�ė��6�[d1(��JP��WA$d��1�QFl�m/��f��xzõ^������i�y
���+]T@Ir��b�� %�<�U$����|!7|t��rK�@���H��N�z`��T&���/�Iw���NY1�����`NH�y�T}��v�*Zk�=�a?�|@}�c�+��1�=h|��6�X�e�gP���xni){�����~�*�7o�hQ�@Xd�K�հ(d������ @�H%�J�v�s�(��]�ĕ��v.d��r�ꪶro��[�]�s���,������p�K�跡�U�Ja�ϲ��_1$�4��TS�e� ���+��X���5⽩�t,��%���--K5ċ�������]�1RZ�`%�J�����%2���k+�-!��s� DS��m��?�g(��%�!�c�����-��]K���{wx�V� �>"��P+G���ו��z���s��}h�L������E1�c�~�q:3|#(�K�j!���!%�pI�����62��+1�Pj��L�l�ϤX%խ�u_<Tb>�Aι�N ;P�J ޶l>�1	��sc2�c���3@Ap[��;��ۮL~�+�!��!���<TT�Ѓ]�W���Sj���i���ɾ'�X4�8HX24'bv��+�:���e;JW�@�-HV��sSI�y3Q�%�J�7p"���i�5K�������� q'�e��j̪S��|�Ƅ�5� ���-p4l��R�h�<�3�����!��9�{�"�Q�I�ʽ:�D�����Z�-e,,���Q�"���M@�b�I� ����4��I-���T)���(�,nE0�]�)*B�p�4�O��=>qW�6��9VA��u2C$%�/n_L܂��Ń݉N�����]-Ռ1_�Y��?ĉ s���ٮy �W6��eEK���3&�=츸�
�(	U�DC��5	�-H��A�]�%��)w"�g`Vh��qi5엉=҆[�AC`{	��~�*�	?�&d�VH��՚�	�iܖ]Le����Q�|B�+��@'�0�&A�ry~�<B�J6"Ʋ�n�D�
��%����9!G�Ҋ���#9���a�D57��x� &W������o���F3މQh�s�J���7D���a7/B�sT�Rr�r�/�9p��������@_�P�%���#E�>JF7}	�7zq��a�!㹐��R�'��$��v,x������i�4���-Ϗ��5����6���V�SLdV�pf��7<nAP�U�b�s��BE�PW5b`��-��(ݴG�5�<��m<c��X�fCCpR4?W@
n��d�DV-һ�������M�5��i"�$��,�5�1e�F#a.AnAϘl��u��Ȳ ��K��!g��-��f�ڹ����~ �a3��,$��I�~/��,�&	�NK�G�ȍ
fޞ�^���d#{��a�G���|*��a1��d��W7����)�	E��ءTa)%��'ȩg�>CN��	w�eKH�_"��ۺ�߲{�k2 ݺ���$A'�@~��5���`�X���&H,M�y.�W����;q^��Y ������� 0�!�6M��@�+��r70%蘃�V%+�?�p����Vp�9�_���p�@}+��k��1������K�&��P&��DU�:����ŪXylPD7�M �?ۨ�.�gA��0J��DB*���!��r.f"I*w�Hi� �_���JZ���?/Vn9��Ĥl^��[�T6���I�d��eu��(� d�Pߎ�+�?`r��-�䈰��<����*WG��ebr�W��`R��ٚ����:�9�R�B<:X����՘�<f��RJJƈK��=�~C.�/�K�=v,�V���-E����
���lb9����*�Ƕ���nW�y�^p�j����3,�B��@]���IE���X�bE(��i�|�Q�%��B�0%�b�Y��,��.��L�=	�sI�m����М�(�+��G)L��TT, �
�B��g�	����I�� ��n��q��m�^<A|<��Fꮑ����0)�^���y��"s���pD�@a�==g���R�Ǐ=Ij*aaY]A�V��y�����)���"���-ܰY�9-�7
̅E�MV]]\�����Ǡ���1�ԛ��=�W���"X��
BO=��߻#�hV��r.��L\ii��C5��t����k����aR��1eB���M���vY�63k`^������lEsYʦ9���ca��
SEX�I���QT�|�������}u�&��99�F?���D�y�]P�
ώ� ���d������&>G�BkR����(E������fB��|!ދ1B���p]\J���k�>}��8����F^  �C�ˍ�춌L[�Z��E���� �:��e��N]�VV?w�㚶/�|^�2c3�`����ք�w�h��b1�!��[
:�|��*�?��?�Ms�
~jA���-�ў�����xI#��l:H -�̌.nn�3z�WLbZHvW�`�]����u%!(.NϒF�����i�6}uN|����ov�բE-�����ݻ��Νc6qV����S&%�,U+v�d�ȃ�n�k�l,J
��h(�.�w+Z�@�՜5�e�O
!Ø$��X��1�
�m�������]2��*�	aѢ��f�gh����e³*^����3�1��`� >9,�̴�����#�"u8fZ����n� �j�"A���\[C|�<�&g=�~���<;;K���\�"¸2rQ!aq.1B`���}\�-�� F��H���ɵ&x�H� �/L++h���iaSlb���jc��kt%GZ�$w�9�^�I �^9� �1����w{M�՝��I���}���w�y�o��ֹ�����n�-ip+��]?l���)�X�ЎNj��.��L��a?x�����#E�y�c$"Lzd�Ѐ%�'����A���n�|�2I�Q��#�0�mx�"W�
t�ك��?��df�{�]���_s�m�Z���K�#�ƸwA��� f���p����\�_hCxiE��%��	D��ta%/�@����Xۏ�i���}��۬�I"0!�n�ҍ�K��/�>}rʹ1x���q8ǂ�$;g���8??�>�H�6�i���x&�!�ِ�%!���z���Ǐ�Iŋ��[ T9sA�|���g�gݓ'O���A���)]��ӼW�$�d^�~8KTwC�u��܂�&8'�>�GNǊǯ�@7�o ����������R�?�����1�81�����<��%�嵫����|�����~��_=u��n��ع�ãН������n�R�;@ �շ��ۑ������=wzzJ�l��4&�,x���w=3ۖ�M~{v�$+�����%�z�dV`���k��0蘨�XX+F�4ځ��̈́���\�}�YP�,Z������=��w<�������	�/���K���x	���d@x�+����D��kY���"��C��s_�k�b�����TGZԮ=8�����	"��U��%A-cs ��H*H��kԟB���b��CG� �32������[̗��1~M!��_�g<;���������?F�X�'_9ڹT��<�R�׌���|��78���{w���l.�J���B��Bc^N�F�K� ��'�Jq7�����Q���ǡ��	f~�y����\��礜:+�A��?d!���Hؼ�$������t��Z]'"<��)�����!�������^�s��7�|�S��Ԃ�����*W�Tmi�@�]�5��d�ҡr4i�5��������9J��1_�z5	~�拽�������=z�wDj�%k�K_�?�/��|~LVLHxG0�g���ɬ-B�wb�wlvi��1�Ek�Z4q��F#K�W[f�_z�%>�	�X�*Xs�}��@��-��O��x��i�s@����Լ��%0�з���s?�s�*0�q�y�H-y>����K�M���cWL�����I¨� ����j�4)r" x*_J�]Q��1θ65�2恹m��o��j
$�K���*3��X��16����#E��8q���V�q$ ���=�,�z��T����@3�gװy3$W��զ��3a�vu~�&�ӧg|op�3G��|��o��Ί���ߊ=6��q;�J ��ݬ%��g5:A
��]�¿��6o�//�|}����?��/��W��y�����l9�רه��!��)9s��ɨ!���VXx'�.	�<�̄�\����R�2��sQJ6��D(5X����kK�rA����s����ֿ�c�x�|	.��Nb�.�Õ��Ъ��/\��X����½X��R��yѢ�^��@Vѩ�jy�<z�N��|ȓ���0+��ѓq�� s�ms���@(��?z�򕯸w�C|��ߗ�=�J��&�=�����/��3�S�7)����Ã���{J���Ï�o���م�Nȵ+�Ű�7mH��c�f�ީ��0�	Ǣ�W�|=z��h�N�V�Q�eJ���,v�&��!���%#i\��#�SӬ��m���\����s1	U�F�kv��_y�e�3�#�仄B��'�q$%	}����3g4N"�#)�Zb"C��_��	Q�l�IA�MM����[���{�٭*$��rj�`	�%�����W�T���z�?������������z��OUP����ޫ�~p�o���d�-H2�V4�����%-��n�"�O ���'�5c϶������D6U�B�[�-�d���`��g�M2������=�� ��~6��ÿUb�Hx����1� *1� ���v�����JK�᷸&�T��acBk�I�z���C�o5������1�%cpA]lU�㱀��űc,&+�Y���S��Gt;vu!U���\@�m�E�𛝚K@F���GZ?b�@�"�!p]�2����o�����.�����_%w({*��3&s��Eh����r�:���i�����~��iH��s4�P=9R��S���E���������?���ޭ�y����S4�.e���B��gx$�/U1lt���q�^�c��b�iO&�	]�Ww��+O=������o���_��ϝ�T��������o���ߧ��EN�%! ��4���j����=�
 ������.�V�C��(�Q ��{ɵ�yW�u*T��\�����"Z��p�H���?f����ثZ���s�[���j�*���N"��]Zt@;������r=*ފ�;_XnA�u4 8�kX�;�J:��	p]L��'ց�9��({@��'�?�14�"?�5Y��l�ތ��ia�������9�n�nX�K���u-����\3/�)�:����P��BX�m#�1Έ	@��%��?���k��0�f3�Ğ�:/�+X�zv�q?�*�ǈ�Ģ�Bqq���*	bo�1"���q�"���_F���������*���cx�v=�h�Z��=��#[��D`����J���&����~!t�;�^fD�q�$�����+�J6?d���t��N����^@l;D#�$��$������'��_:_�����~������}ba���|�;��JB��{��������o�wۙm`�("�M\@3
Q\¯E����	D	�9!Q��q�����n��� �a^ԕ��v�n�H��J��<�9G�-W��==;�H<f�!���Ic V�mZ�.�[amSI�OU��� �*�.�o޲�b��`0�Vc_y)(��}>���G���Waѻ�N5�P�'���q�"r<6��?���,��T������}�;,\�5�EF�ޤ�q���+�&h~ˀ��ؚ�❡���;'��UZA�t��l�B��~,��z���U�H4�"l!h�G\�b�/N%i@�V+�k:x�D�2~@l��g���/��!��Ya���㣻yY s!ݰk�����!����W�ʮ�$G�+��dCW$4ꕃ9�s��;�{O�*�<1x��0@�4���l@�QKBP�y�Q��H�~��G/�$��������_��_��uA���/���;����G��$e_��Z��\���z�q��X8t�� �H��n/\{�wX����`���[ ʌ,��H	K��:M��`)8�s�h��9n�w�� ����G��V������0T��Ru���@Ֆ5("V����sp/n�vŻSϘs��y�������ѩ�t��K�T��8].��EA)��=�ਞ,0�x�^@q=s�6�>�����Fb
Ȝ��"i�֠0�r���\��:qyy��\){e�(��v����]+���i`�T%�/Ũ��:νn����S)H��	�q�8zA�r��8��#@9[��-
�H&���2/�]�h�d��Rh=�Q0��x��f��`�����6�xW=�!ǣ�8��Q)eOO���f�AD �-���'�؍��L��BB��S3����X"ke��@<����Ǐ��Z����

�*'�������~��Ĝ_���� K��3�۪`c 1��ઌt��B�
`qyc@?+DSVi��;��.@����5 By�#���7g�7��;�& �T+���ث�C�t1$�s�eǨf�[З�.���f��p.Ȕ���C�(��%���M��Ԋ�b�lv2�,j�& �d��_���uL�Z��&��_�٢�]=���h�'q�I�LhQ�p�6=���Bȝp;���\���q��X��=J�l�ZY� ��ˢ��}�WU �r�&oӀ��Zܶ�Œc������GqAb���^�W����+jd��V��^^��킆���a�yd���Jρ�.u��x��%!�vHׁ���E	�%	&��HC�� �J\��ìW.��|B3�8�	F��4ϙ�%+PTlC���C�;�
+����/6*�4����Y��w��âH	e4 +�?���/���������������ӧO���W�=���fW������Mvv$  �x1�"���D�1��$!(7C��a��\aP�э��u1��J ��9�� Đ:�F��n8k���y�@�u�l�Hظ��Q_��x|�f��ژ�	\��J��$��&qrg���r
F�c)��_�R$��@�Zc��Y�H����Rk\Z�@������/��<��D�Xձ��Ӣ�q��!h���Ǩ��H�͕���]��21��r:#��X��T ��J$�lZ/�.�h�tC]͙qVq���!���R��/@y�^ꊦ0t(�ݿ�՞�����:AQ�\4=��e/H)���u����ߠqH<b'��B=x�jĢD)��i�}L�N�ŋ1NF`�K�G�c��/sy��]HG����m��¸�I&�P�gI�Ì�����Rvsm�{w�Xʴ��'�f~������w���/��/5�ZP�-�귾�����=��(T�oRS��B'Qy��u#���U�M>h�5��b&���v�������pYZ��U���3��^�g�y7h���
H�˷�2��rR`֙[�q�' ��"�&�;�3<�
M���5"Pσ���g�@�ެ�#(YkI���\���v��˷'���|�XX�m-Q�z��}�y�"�}A�<���(D�k:tZr��j�\.]��\�*����%����t�i��	���Э$-�b�ut|�J�Yy>#�g:��l���!&�>.䤂�!e��,�~���0��WmȲ�`��P�&%���fڍ =�*(*)��:!��R���a
�ʯU�~�i!ĳ��������w�u�&�y]�ۢ��`R�Q���Z"���K�@tKxɦIYI�^�Ŝ�2��i|�V�-�/�9�o?����>��S�>����?~�o�-uW`[��L�xR|U�,���%��ʾ1��%*,x���ZAZe�v� m��%0Y!�l�QLv�R2���-w��N���6��)	W,hj�oh	�N�ClZ���j�<Lv���1�.��2��� T��ki7���X�s� g="��۸�o,]KL~.��O���|1T��}J�o�
Vs��q���x��|���`��a�Z��5�1�y1�84�>�B]�����̄+�9U�(��
�����L7n�y;6_@*Kq�˓�1�;]̗4��Y�T���>��������u��4{'�P�F����ܞ��B�1Ac
=��R��`tÂ��B:؎2K��tW\�$U��+9�Rj����+�.�����*p�(���7R�G�*�Y��}�S���~{����௮�W?�?�*:3�����ф��=4Z�:�=���K"�،�!1��o��Ɗ)�u��6ь�1������')/�Ȼ��rա�L)�B�/i�����p)??l�+��e�Ba�5��܇�{��)�Υ��S��}2��*F��] � �k[捅'[��K*;�B 8�� ��QJ�I��O��`�a�������]!�pQjlJ�m٫^�x����Z��_���cuHQ�T'3�0�>$de^�r_�-,�z�켦:��~��}A��~�]�/�<`�x����P�9.sI+�sT�����kzT�c"�I)�"V�\Q'�yYy�PUA�?���6��V���}�x|��A<T\�(F�z��]�]�z�ir\�}������՗��w��o��7�z����Z�vۿ�4�QZ��BMP�d5��:��:?�s���(ۥI����"�e��Ί߈6��uV��Ќ<�4y�+�e���b��W�'IQX,�ƙ��� �EʅM!��.U�<l����.�9���'TAW�@*��DMKF�L�����
-�*U�^o��P�-�(��U�3����	�^��@P�֜S��b��u�D��9�ꂔ���S0�s\ժjJf�;}	�y��\��$��ݶHE�Y��R�'���I���������f�
jC�_y�Nv?�聢�e;��F����a�ЗJ�RE��"��躀:)��!�;7�<�E`�k\�\={x8Ƅ�gTT%a���9�X�W�o)��3a�A�NÐ�<�hˡ������Led�`��ܩ��_>~����3vz��8=�J29^nۦJZ��g4ᛐ2'9��`$���Tr�|m5�<O~>l�{A����Q�`�d�e�R3۟�X7h
ל�v��\i�Ka�᳝��t��CWo�jT�g�w%k�vt�xC��Sa�8j��pl�Fy��E1��)��i�ȓ.�Q�����
b�#�P3����&x[XbE�^EۿK�Sa�,�B�fG6�z�n;�ۘ+Zq��l�ll$���9}44$�7�/��~TTf��J�n�����E
^��Yu����5�͙aZ��3d��A@(���E�I0_��I`�����A�B^2J��=��pQ�3#�S�����.t�\�V�4�	�_l7THg��v�"5��\sR7��>+�c�dr��n�3���\AA�?��xB�l���i��Darރz=�*5�ڮQI�%;X n�y�c��-��T ƍ%�W_���	.-��lw�T�,����ITlV��TP8�O�6E�g�ڢb@�U5Ho۠�& ���B�&�ǂ@�P�,L9��YNA)d�����~C$��w����X����tk ������6�ObɇJuj��Q����8CN�T(��A�;��mMc�ַ�HD�L��G9SAaCr#�"jQ��;z��E�[��n�,�Zd�Ҽ�
Q�n�H��DI()�!�Y���;�RW~[K��V���L�ɥ�O��}b�;��Bv�������ṙ���� +�qx|�qG^�P!�T_u�&�B�, �IH��)�+(�ޭw���t�Z0�)��K]��Ն��ه�U��m<�J!I<� �ԭ̥_�.&�b�%~&(��)	�-(80>�4�1�N��M8(��V=��;"(�D��H-R"��gh��uIPX����������q�r��g��
�ڞ���n�� C��֕������m����<��*<S����^F,m��G�R/��PC�i�H���I�BP��WXА����������Y����D'2;$~)�}��X��Zj^p�`�5�G�,��B�cO�f���Ժ��� ,1Y!�!���Fd�ܔ�=L%o�@�����hj~)����Ȇ�"���^E�<����y�FM�aB���q.�{tpTvϒ����~����UU?�q�Esa��3a��2@����H�妃8�b)�ދ>myg����&�j�:ۖα;���3��P��'����s�Tp�^�X9���	֋�@+RqTa�-��I������A0� ������jz3g=�l%o��F�<?��I�=���k�5H��ݘ�b4��p�0�J1�<u	щ=��k�I�B'��d�&
��l�����UGJa8F�:��7j�E��j�� �&B��%/�])�j�%����f�n����P���mR2��9�ʉF��i�K�E�sݏI�Kf�3��	
_J�>�d\^q9���h��(D��n_A̰�IJ���;P�=�W�@J�����dV�M�Y<@�
ɚ�y�J���� �aym9q���)�5	�͓���(�B����!i�wh��
��2�"U�쾱�kؖ]��iհR^\j����#����`ȵ��G���ԌI�x�����U
~���R�{`�nߊ*D��&�ݰ%��@J"4��e�V�C�L�7'��	���xa/�f4���-�������^�-C�3a��L�a<��w.�߉_ᔛ�֞�֍����c2�M���|y�M�Lѥ�\��RT��C
{�|鳒g-������>E������鞫��a���e����GΝY���;<:J�&�X8x�:q5H�M�KZ �ْZ^(I�Ej����^N�qb@H���QLV��i��<K$'%��y�B�j�\><\̾���{F�DqE�<�n�6�	�
=�7YZk��fn�.�pXG�7K���i�T����~t�F`�潉H��b�>��iew&N��¦�*Z�q���%�L�
Q�� �zK��0�_��`~X( ���K��Ω��CA���p9��� ���?^#զ�
3?��6r�4��QCN􅡟�ס0B���Cz:�&���}M�d�u^�������rf$��lI��y�8������BYD�d!	���*I� A�bx! ��I�0�![�Вi$Qəyo���?U��s��:�CIV۩�h�y?�}�V�W�:�;.��#|e��ؒ����#�������|���y1B:a�XO"fZn{��ɬ�� �mf�K��[+J��Z#mci�]c�6z��s+��P�����$�P�<,�PC��S�wp�G��#[H���\aM�s#I�[�>����čr�}�!��$�}B�?P~�����a9��~ml-4�OmwNP�=��q5�'rtt����?��|��?{����t��D7���F�q��J��N-��T��.{*��]>,p�]�g�c������~?LR�~��&�?�!�Y�(4�	�P�q����]��)�������`��$�u���B�r�"��ċ#N��l=�ǰ�E"S��xkYaJ���kI�_p7��;�[�{9&�m�a�ud7׃�}c��q��V�0�/4&
���\�!F*�<"��:gS
Q�XJ��4��D�(_Ij���`-�\�4(xK�̏C��������q#DT�D q�6��2�}����Vju$�&tw�Ӎd0�w>�w�����u-D2Y=N�ӏ���v��k ���_�P�ߩ�ӗ�i��z����u��w���_�������Ct[���s�����Wy�wwb��=F��=c|�1~��y�����y5�v���jC:G��$���%����o J�R�|����s��$jK��O~p�`fs!�d�7]�mx�9��/ J�|�Q�?jLF���L��O���E���[��iD���WI�Vt�<���٠��N�tl;�4=��|�X�Z�1�$3�	'�!���v3\�X}�}�ِ�织{���Ҥ�ۆ�$t�7���bEb%�{�ti�^��9Rl�g�C�ȧ�ngh�Rs�7�޺��z���֦�>v����p��������֙��_Gc��lY�+��U���&_��=�O���+D����� �&�O|�ݗ��������W��?���~"�<����^n�?-�=ypv�U�<��,����(;r4����_����x|���3�we�>���t03l�nOo��!��C&�-�R;��'����3��-\�H�ס�3՚b�oͶ��{���m0x�'>��*1��8�K�ܮ�!1%�J�x����K�V�--~.���(���$�kiC��u��K�l����-%�����m;O�R �U+���|�llɈ(d�`A�ck;sEl��@��/�r�̋�B���ej��P�0ڧ��8i����<�m�2��F��~�:r�-��ykX��O���2'���]OV�w���7�W�~�o��/�@�'ң��'?���_�����w������By?Q�u$�A;.�w�?��DZ���t��I�D4N�L�ᦸ���� {)s��.Q��]�NƷ߃ږi�c��ALſ ���k� �H�B�ԫ�z��i��(�����b	����R��c�n�W���B�mс@���ud�I��%���`������fX�I����i�Y&p��Ќ�c��Ё�������/���Wƅ*�d���gŭܦ�6�.(a75B)!�J�t>e�Q��([r�%�w���ؠ�bE��2�L�XI�����'�o"�%�rs4��R�r�fǾv��y�B1�vs-ǟ�Z`G����sG���9*J�q!I��#�s��}U���J�e>M��vQ�u�ֵ����k���'V�"�x�3��̿�:��D�>�)G֘a�ې���H�Z��l/���)��,|�q��&�Ns[�`�E���";C���s]0����Yd�ꐃXF�D�)��*�u"&h;�&�!���tȂM��Ӻ�6}E����IO�7�X�O��Vð�[rH����[O~���o3vc��޳���v��O*�?avcC>�5\�
�:tu3�	Uۓ��)�.��!F#V$�f�VJ �ZA5���,�#�I�<��Lf�K4��gO�� f�烖�����9`��j!�#z`�CR���6�rJb�b0!_�� *�����߃���AG�y(GO��3�6tG�������EH�|^d�kU���I]�4��������WO�w�������O�ӿC�-z�}��B���]O�K`�0l9��\Vǵ����_C�B�ܞ����ِM�v�E&�|/ݟ���n�h���)�48[.�qj�ؿ�J^*\����A�Ai"+�d���2�j:S�	��,J�	"��)�'�-���i:�4��c���|(�I��ٕ��imp���B�u�qa��(�,�Ɩ�U�m�@�>�Y��� ����v��n�*�R8�~X����K�����{��`��kě�6������w�l԰9�}�"\6�V3��|+�Y��{�uk�4�cj:B-���K[v]�X�!{�P�4�,�FR�|�ւ|��k��y��r�U����{`C]R��3��ƶ�1[��N"S���\�'M��G+�m9ݖ�c.s��i\���y�8��8���s\e_�{�������wO��߱�����{����w�~��o���%"�ҍ�I�_��<����%�T,���*��Q�#��W�5�[m�^bc����m��q� Q[�ٖ.�o+�B�6�_T�Z!�����8LzP�2\b+��-*��i��L�5�n���5<����H\��e��'D�H�$�H,a'6��w�k���rpcwG�w��p:e�e���$�t?_�D�f�l!"W$DG���k6�v�`���$���`!�E`|;N@�� �
U�t� j�&�&R��d������X�D'��?Cc#Q�O%�'���}������)�� ֪��
Z_q��%���!���D��9\4V�p��#rŌ3�*�W�:����?]��B��ݏ~��O,�/�������/A���/~�?x�7~���7i����z����<K1�;�G�=��A���vk|QA�O�m�`�\�G�/�x2���h��Jb!S�+;'ş�CòM{�=�Tt�]��Ƀ�����LL��%/>�G��W���<�����ՙ��j���N^c����]���q���.��w���|��������$�ɽ����(1>M�?}e���	�x��>�Ey:Ty"V�$���y�@��Z���V�!�k�5=��*d��sY�?E%0*�V�	��H(y"~���9���C�ҝ�9�bX�n��Ɵv�!�s��a"E(>c55�c9�Q�zغ(�D0�M�ީ��+7o���鼺�37n�'�E�X���S�a��:��+4�����Ƴw�����|�Z,ϒYx�h�4�R�JY%8�jA�FIu���6,�����_�����q����b����)���bX��
c�q��轉�=���V*���}��Ҁy��58�r�
qU��EKb�t������b���;6��xQf��+;�`+]�=!�'!
�I�k��J���F^3$)5����d�|��6:�\�q0�N�_/�+���.����������ˋߩ!~!�E��ߧ��D��������y�)ǘ��/܃-��2m�JS�x�A"�ȵk�;��w2z�wqx��,,��zQ��ݪ,��f��G��W�}��w�ί��]=��Q�1"�7>��Ͻ�����Fs�ߟ��_��� M�w��rk�^_�戦BA�6�4�����C�E�q1��Gw�G]	�3!l��k�Cx]I���yٶ��_��%�`Ą�L�E��LO���SjL�k�_���hB� ��^;���B�PˤH�x0$j��4�XZr�>�.����u�u��ϕ���U[�I������80����i�)��3Ix>�)����얠w&?o���>�v���d2�s���Vp}Fȕ�D#N)&��Х�5��d0�3qy�ȸd|l-ៈ�����|�w'ճ���_���%�O�R�"uۣmv!�o�����")C/_��~����Γ�eV�ɲ�ϒK��'��E^�9K�O_x��9�?v�㳟��9}�=�I��Gt�*"��W��Ξ=�w�w}�m�+4�pS.�cg���pr��C=/�v��d��B0Ԙ��(Ϲ��.�b'���>��Kw//\�ٷ=�t����][R��Hwd�.\�,A�킒�	%�r}�]v�}��}���0�~��I9��.޷�1!Ջ�du�ǐx��o��͸���\�]��u|,hy/G����>�NH��߃�[fd���v���G�/�8���X��x�ؕ����+.R�;���mr��C��;IZ���G���+�K\ڸԭ�,9#��^Y�w�"�F��_��ߙO��:*�k,��þ���E���ދ/��5������]�X?X��~9{xr�����}M�=K7�܀c�8Ǵ+���m�i�H�N>(w�%�;�AR���_�@W����;��W��.:���'�?))���f폾�Dî�lRߛsb��Oi��˥�l��t��3�t����C�&����kz~nӔ5]G*f��>�C����8W��/1Op�<o��_LCm������s;�u(Ix�;@d�l
n�&��j��8{��+ǽ� ��F:��=X�a+r+��K{�|$/ �#��)'������A�	�5��L*W����X�cL����x�C�<��׳�|C�ΐ1��Y�7y�.�<?-���<+�$�|uRU_/��������r�.?����JT?)���EQ`���c ����o�������$����Nm_���d�X��b�y7Y����ih�׾�L?�IR��N�е�,:�Lg��%n����:��Fk����h�v|�@��m����T���Ś��󃕽�kw�굯]�z�ߑ�������;;_�ȲrI���5=�;O��֛q����r��b�����43d����f�z�z�)iR:r�,�0�]N�V�5�m��'����������&%�\;��p=�-�j2r�Ak��>z�$E���w���1�kL*�$B4�����8@'	t!aK"��"�|\��h33K�Z��m-Ww<�������V�j�#"�P{���J�E�Yj�V{�Qj+j׮U{S�������}����h6�\�˒�`5)�L`�T�{6�'��S�D^�Z��Bߐ�e*#�^���J�u�xdc�d��O����o��\߲?}Ru�Xm{\:��(������LNj2	�<�{ǮLeI��s����&���"k�?(J���]#�1y�Qb7bT/u��9��贁�������T(�^r��d�D@�$�.ۭXb�RL�K)\���#��$�4nX�z_�ݤ�]bٖ��\}���dAY1�AS����l��¯�����E+������?X���1����:n�'�Q�;����R�P��?�������`-'8�8<I` �|~g��~!��͕[E���K���P"O�������*���ƫD�gʷ�G57���m�?���mR����R�ws��<��Υ�TNά��/Vq�v�����Z��y*�t����&m���0	?k7���ǆzr���#��e��2w�☪�{��n�h��Mr�xM	�\����&4�k��,ϾW��dG��Ĥ�O��m[`V{���"N.�)��
�AE�Y�2=&�����Z(�B|I?����<)A҈$:���N�G�\�u�Iچa4�W��D�.�L������}���X+�(їՇ��@w_^�ʀY��r�-�\F��-+H(�-ToQ�a=j��*	>�����ӼK:�����8����[��>���4�;{��ΰ�|��OJ?�X��x��bD��-&�&/���W1A<�`��X/��7������6���n5R6�.��&y�g+�Y��ؖ*�h�y�v�ف�����u���~�2ށJ��j[�G/qk��m����ղ��(�X��_^�<i�#lZ�I��P�(w
�����F4}Ub�b}���F�x}*yc������H�;�q�Bс��R�>�$�*�K��.�ƫF�}��,g�0�<9#�|��q����0���ưąٺ�u����v��M2鰍K�Xu�����N�O(�c[/}�inth�e;�Z}�3��ۯ��xFZo.w�b-�<�.�M�y�ʹ�S��3䤆F��%����̯��v�~�}幕��{oNom��E
ր����e
C������I9������d�l��[��:��w��N<�zRJ�]���v�����[��.���Z�p��Z�2-�����o?���9���F}��c�r�`��D�~���q��heu��n��,7��"D;S6��Y�뤘n����l�~�$\~�k�}bt����v�.+�bɰM=�j��cy]ܪ�ԝ��~]-y}��]^�LZL�W��/���˧w^���Cd\�mJ�c��Es+�.����������ʒ�!5�J�/Y_W�W+_�]'��U3%Rσ
��4'�J���/6����R@B��r���fp����ʱ�kX�&W���!U�T�H�^��������y��?�0Sp�D4���gK�k��^P�_��t:K4>C$O�"/Ш��I�]�e�S�-ה.��Ɔ�����u�=c-RL���?��0 �A\-����y��X�`pr2�E	��ާ�I�
��;Z�4q�*F���"Q�����|�[�M/4Ʌ��	FBI�۵��x�_F���JjS�"$t�r]+.���;�J����B>�+Q/�ѧ��t����$S13�=�rӚЫ��*^�=y��=��t�6�рM�G>7�d�����Å3v�$mЈ�B@M#k�ȅV��i�c�������	���,�uǹ�_R��vk叿DRh�'�jeR�g&B��?���gT������F� G��H���H�J�K�n�?����
駽I�v���s�4vﾲ>;�.��9צ�KS�\�:]tG-�C�[�ck��!�Q��<<��6�fw�i�z��U���[���ٍ�d�,��?�4���F��mT5���א��\��l���k8�c(^��&XX,8��������n��Ti�3�>����K�J#��ݧ�m��Y^+�l�-6�,�/>_�m%x㘎W%v�P(n%��~J���b
2~��_g�H,$˲��8-��X5-쓘$,�e*���a������~����꧜�,� kA��R�%:4U_��/Ȥ��hH�S��{2�c><؎\!�7Q����eq�-8�,��$��1�F�>�sx��dN>J!����ڬ��N�[��[�"ʸ��p����a�����n��i�����\��`;�G5�]N���^߀- il�$^�Jm��"�I��?3�*�m��dfR5��|7�d�xmjJbm& ��Ӈ?!r�\�B�	���;9�|߅2FB���I���za*y�� ڋ9��͟�e�#	���b~S�q�a?��a�+u�Sj��b%*'�{�	���}���t! -�R.
"�ź�}~ndw ��������LJ� ��j���u�tYP�Fy�ھ�ە+7sBCH��|�蛊P�эƔ��򚪙\#�ȁn�����_�m�it���D� <�B_��؏�<�)��6f%�~����/+�I��]o��o὎t����0�Z�������|��0�m��f������(�����n,Lsn�Y`E�q�'�U&�:�'<�_�#�s��]�Q��z�El�m�Lmf
n����k+�݁�Y�D��;�%�������E�j�+��˝r7�v�?���;��^��,3���Z|��r�o��:����4��z��5G�f�N"0��.놘�fQ�����A=c�Q�p�'W�iT�X�uzt��Ը��I���o�N�s�r,%Ն6t1�������7���5����𲳮���[M�c�:�1�2�D/���ߺ��ZI��CymEMb�i�4��ݫ?)ݦ��~MB�:��霅W���E>$��`���j`�Võ�e�V��2Ne9gMz�S�!v�+��NlZ��>K��OK���U	�Eg[�����������!&ۃ�0��Z�S�mk6w�T��D����[�lU#5.���2���(�˫{��d�[RǬ���}�<��'k�H����#�|V��Ypu�Gz�_���W���)��x��+jg�`�|�0I��ok|�WhF�\?�����q�a���0�1�d%����5:�$K���A��?Qȃ���xZ�=�C/�[E}�AU��nP]Y ����8����QU@�o�~>4bԴd��H_����t��'�۸�+ǫ���,w!�L_�|Gko }Wx�	�j��ʊ�T)�e3�;����m��h�����Α����v�j�1Y�_+�~oWA���2�+�X�,K��.���b�l?Ǯa�q���Qx.z���������A܌]Q��~��6+U��j�&A���QI�ì���k����s��S.�]�*��������\��ٌ�AD������?e@�ik��܈�T��3�n��N�k�/���}s��;��?��{.2>lg�/W8i����vmt��EF��Sʨ��W��-V��H<6�l�$�b�
�d�/-R4A�l�O���������^�5��\��߲�_�o`�j�Y{�G�})+n���]�<ߩm
�����l���{Q�j�1I���wK� y�g\l1d��ͩn��>��AZ���'B��o����ɃR~�-������[���L��ļr4����ư�{��DpѺrA����}Մ��'e�'���c���r�"i.��D�@[V0�M�x8���q;��e6�9��#o�8�U�k�����:��F�.
�,��QW0ii4�O��5����|��Vz���t�+��V Q����Y,힟H��U?��n.�Uy�*ݣ��&���)�I���܁h���[�A��%���1��
�S�c	L&��B��st�@�͢	;�J�_�"}d���\Y��o���a.�Y�:���PϒHM���?�з��7d�hU��̇f��$Z9���w�Otc<�)�W̬�.}ՈF<��I)��@�����5���Q=Ca>�#�F�;-ڼ��$I�B3)_B?НFjV�\*4;[єvR㪓,�RY��r���e�z�ż��$�!L�	0u����<�p>dO�����y�W!d�oa6{�-H���4�B�x��8@ ɸ�^�X��������`2c��ܷf�i�XS����b���}�#c,�����ׂ�ak1\�)�N�%�zV��q���d�e���$�%�f�K$2�2)>�K\�(���2wB�#1���I���vU\�v/��~������>ar2h�L�c����;�nS�u]t��h��%�O��$'Ë�
����Լ��4b�a��3Azq��o�d,��,w��gk����l4!C���5X��Oq�l��K��\��Ԟ�L�4��z\�������ae���d�T������
]!W�x�,\Y�j��*�������L0v�S�=���|�1�E&!eNm�;	T؈���Х_�!���m���$�}����iԥ7��yީ��j^�� ��Te7k�w�l�A�wU��$�>bF���$7���z��'W�Z����A��	�3P��jV�P(BREGF>p�����RC��I_���4y�'�+�-hM��vi�tf]����&�	Z���jꆄ���{MSٍרܓD������Cq�ƞ�fN�o2�|z�J/�:戣���	�,��v��@���vw���dr����b9�Ъ�Q�u�Y�P�tU�?w&#��#eG&�����~q��YUJ�'�L�č[ی�T��:-(8�Y�0k�:S(���M�x�d�|�LlP�P?v�h�~MSl��tY�Tּ5z�[��(�
\%{��)����(VҰ-I}8*0�3��,�=��{���t�=-#����Nk��
�8�F}�a����d�>�9u��zz�=�g4�����N��}GAs�ڱ�T!��;�Nj��2o�_��*��Y<g�nx���<o���@����WRt�������r�� pL[w�Am ���tS�?ȯ�ȇ���7� h�&�����tc̃F·>�T@X��R R�meNz���z6r�v*��'�FV�1���K������֢��m�d#EB��>�'ț�Ҽ|�.�����W1b~
�B<�?����#�����y�&�����R����L��q㼅%
�ʝ��ڋI�?DH�LZȝI�N`ڒ5x�2
:.U�M���d"ߘJ���I�F�	�p����JD��X�� 2Yط<j@'���*�yv��6�_��r��}
}o�@����و��J����z�-��`v���)j����ԕ�LN
���[�Pݥ�ec�ɨ\��8��3��7\2�������|d�ܜ��he�U.�}�����HY�T2j�/��OD¿�
�7������K�t�;�N�˂�����cj��L���i=W�W���V�w��Jo�ye�RN����W0���x�@�����QȒ�>�n���Z�+�}	�{|�_�!�`�"o��1�������v��S#���:=Y�Ԝ��O?�`��2 �M�X	3�Y�n��7�G�)����g�A�#���0l;l�YɞH)*=ؤ�G[W{�=&U����ҥ�~�c���[�*���l���"���u�P��>Z&�����Ǻ���97�M�4�������!�b���D���A��yKH{� ]1�N�5b^�����w��א�#@�j���u'gF�q���"]���<Z� ����o���3x��!p碤����-肹Z
��<[�n����f�i� d1�<�?-��>�1����EE�}�A׹O���+@F-=Y�Ǉ��c�(��gQ\D�~<��E����j�H�)��(Kh��'}�-��N��;�e��TG�i���Be\��qi�2�"��A�<���WXOQ4[�a���q�����D�K����+E�_4D(�1n�V�og���̛�����ٿ��3�ݕ��n�*ӊ��]���Pg|���ǃl^kW��U������<�7Yn��D�+%���i� �8�*&n�$Ψ4�m����Of`��VM<���J_���e���+�`����~�;��I�|��M��t�5�V�\W��+W."qt�0Kf�e��4ӸrMx���m�/�+o�碸���H�	���0�F%��c�H��%�����:,Q)R�Tsq���W<�G��l�Ğ^5f^t;D�L*�Q'����i#�R�A�yk�3���Anqk�I:>� ���,�^&��V��������4�?��O�R$�V�w?t$E�;�Q.����]X_������"hץS�`__�:`�j��?a�����s��s}��>��''�W�4OĆ�x��ozj���-��H)�!\z9"��̌I���O��� _��HW���ʸշ�(-�e�؉:���g/�����ϹV��K`�ڨ�~jZʁ;�������=�J_g�G��Ǽ�HRy�l)�^�b%Z��u���^��3��ޙ��F9���_&���<��JF)�H���6o�1�����F��>J���\f�=:ǒ��H��5��ID6��@XY��,*;�����"��6.h���>K��p�T<���h*��M<��h��)��PK   F�X�x�</�  �G /   images/d8843636-1db9-4a03-89e7-cf770aced3d6.png컉?�{�?>ս�-ۭ.�IYSƮ�����}-�J�6����n�d�4)��l3KQaD1���%�,c�=��������{<~������5�z��s���|�׌���$���;�9�c7�Y�w#���g�>��~�GN��O(�h��&�?l�0�j�g]�����6��g�q�|�08N��?�S>n�޾�),mQ�W���O�~�_���c,0&FXe������#��g��Fv�]j�j�pI����[��5��	�{�X�}\�����$�j�z��ɤ��z�-��_�>r?�Z|L^���M�u��0�.�az��]zǴ���`ܼ��9�/��,)�JN�6�jm|bG����Xb��	0���Uɹ�.6e��k�=�����sQ�IG*�%����D���*Bجb���)��x��y>KKq� w�v�L��c���I�a�~%7���H��T���!���R��ݎ��IAIi�#f*~��ލ�8��8�.��!��H����R�B�]n�]��7�
hL��rm�d���dͷ��v��a~	muUU�i[W-4��9�U��3t��C��2��l9߱ܒՏ�5<�84��@�J%�ˋ��+��JH�y<p�G,�����Z�:�r����#M�7��<�u��s�!2�2s����^����<�o�2/���t�^�XÑ䋬�+�ض�[���k��r�,�Lo���_��b�#i6�=�����6���_'�jC�7�����؀�_�&��y3*�}�
T���>��k�Z�-����q�R5��%���^��ZN%t>��k���c�� �̓q.�"�%)��ް��`���(M�B1w�w5ޑ1f�[9�{J���]�n	ⰲ��@DҬ�[�8^�����gtim���*�:�޿�����rUɀw�JGoc�_Zɧc�N��zoݷo_�Zݼ�'kźy�����������f�9��Y�&Z�%�1+��&���(�0��7�:�����z{�8)\x��ʂ��\��Z�})͔)���~̼�%���W/�x�����諍�P�·=̻�P_Ǚ!o�M�|�^1{M��V�[y8l�3),0pnD���̞���h�<��Wt�{�f����j���H���ب��w�#bK�r��}z#�7����Uy��^��wL�R]#]'d���K�-5f���m�u�6??�ŉ��1��A���Y&���%����m���LFƿ�'6�<��1��}fv� n�uݑd�3�N�}���=~�:�!&S/�|u��C:n��7$�6y�nO��������W�+�1t��y�������x�3'yO�T����^�	����?� ����"��_�)���"i�>>t/vF�e%s�GmjZ�g�:eT���)���wnEb��[YY����)b������k-��B�q��� fʗ�X�` �33ۭ�eVj� �8�xqe�y��8�Lh�+,,����=��^�V�ޱ2tA� ���|�\4&�k<9ů���@ѫ�����:g/�	�ٜ�O!_[����-���Q*��{L�N�82* .�~Q�Zڇu��MT�3#.Hb��͆���ڶf�B�s��[ƁH��[�o�M���i�|��	1���0ѵAJ����*�h��^Ɂٍ�⚯\/]�4�S��#���Hk�K΍���R	�<!���k�'��*q0������Wɚ	��w�-Q���8�� ���6͓#R^3��*o��������8WdG�Yߦ��e�_�6Qc+z���C-��%��na}^(M����,��c2�n�=J��r�����;tE�Č��w��^�v���Z��)�<3�Ϻ}�O�u�R�����3K+�w4�*P���C���� ��2��r"Z��'G�0跛C~�mc��&r �����rחv�!��8hm���:H>u@t�Wjr��_�v����t̅X�����
�M�m�/���}{���> �vF�+��!Vj~��S�``r��61�\IW�s)�׽�G�vNSވ�%���pw&��OKKVL|�����s}�w���^�9)�?���P��) M���'��S��ɽ��}S��#�X#��gx��i�n��Nٞ�Y�%̯ó���U~���x�^FF����։��H˞Ku���/&_7��V�ج�b���N��T�sl:;](���)�_�.m�srZ�R���S� \�D��3���T���1�[�}.ԕ:q��v�D�W� G=!�{M�/*+u7I6r h���I$��ԝ:�-�E��t���<<�A{u��) L¹�R��nCKˇ�	���5}
X�$���߾���r����IR�Z��H�7>Aת]߿l�s� |�ۣa��Y�[=Q��|_�Ǆ���6���Iz�t���^�__)���S��UQ �kvR�n�S���ۅ��Ru���<��u(�ψME.�۩䳻n���ui��?q�pqw�.�sR����^�����k�U6��Zd�}��&I'$�x�dv����ʅ���F���r�a����\�"�3�M���G���~�ܳ=7^��v��V'bai��
�%�����R�,%Т�f*UW\�T�ݸ��/�e�;Ǉ����Z��ؼM���^�T�#���uf�����Nu����tD�Ǐ��}���>�O\8��R�0?����Z����q�S�5b���N��K����L�:J��ӷ`^Qq�� 3�Y���Y-ݱ����՜(U�? ���3��lc��h�tK�ߩ^E��=�Ҕ�����26����8�"U���7MOO��R�R�Ȭ
v�t�A���[��(�����y���O�x����K_]�<����?&����9����/lnb+v:&C3t~ҹY�ŏr~� �������q�ƙfmd}���2��19z	���_��/�>}dv��-�ݾ�9�^�Jj�Pv�O+x=\ݱ���@rZ�c���ӏ#��
�W��c��߹�rw�ƫG���\c��q��N�Pփ���Y�/��U�d�j&�v+�D�Z�i�V��cc';\�鶴Y��4-��+TS�Ï��7��qph�,�Z�8h<7�X��5؝*��\ߒil���s�
���|ڕz�T���� �e@������8�t��dc���d'g>M�,-�Tu}�i����x$�V���7}�5�3�O^6$8ҸR���m�����2�p��S��I:%|m-E��_;��߀�����աTq�Y1J��E555���낺�����v��ݟ��f��Z(PW��W�&v����ENNq�S��^��������tL���U����w}��AW��i�n��� ����"~z���"8�<��(S(11��k��>���?PE�������?�!�͛7@�o;[&ص.�o�cd��S^^������T��w���������ѫ�eǖ���wx�-~,��}�Z'� | ��SQ���AG�O�B��>&����C�����3=9���>��hl~��v�@ʹ#�^�8xs ����^@��H'GZFG�7��/j�@�YiI�x�Q�T@6��
g���4,u����V�O��LZK}���Z(X��Pߪ�	�l��VKkɢL������L�����K)��sj��tb.�����Vf���b,�m�=���������
b_���.��+��l�B]g�s���[Y<�;�W��"װ��{ mb�2�w�B�_��}�*I�5��TVtmO���T� Gr��<����s�(�}b�d_�Q��u�H�$�u{A�/Iə?��y����Դ��G�0~p�v�1qP�3�Ұ�Ż'g}@@���k�}d_�Z9j���)<^W�@ʛ@�tvK���k��1�t̔*:�&�]Nq�(Ke�\� ���͇���F��V��_ݡ��Ƹ����G��w���ę؎]]�䟠/�=|B$�Bo��՟��~�8���~�?��s)1O{�>�xƟ���2֯����)�����R�q��,-W<y��4�޿�r��Wn�����4��3�u:fͺ=���"ڽ$��2�]�7�ى�񁣹Ȁ�H�ʹPOo�� PX��Dɂ�f���?����{q��U���Q_���,���t���'{�A���$�d��p������Ka;4ǵQ����D_�+����m�Վ�D	r����j/� t�����-��u%T�fۛ�A�?����7�x��l�+�����&>6�ۜ���	��]��[<߇�q1���������-�n�����S��C/��w�r�� ��Z��=��㖖ayP�~Q1��"�l}I@�7�m矴"2@��4 _;�(3N$J!�|��K�s�:[g����7pCΞ�>�|���Q��ʰ%�w�:�3��oe�?�/�ܮ_��n�OK����<S��_�v�-�L��Ž-��*놮	�7"��������o����|?c�x�R%tU X�q��'��\�T�@})e���>^����߲n�uV؀�PC���0�w�����5�E�d�含��\������p�zLq�i*[��J�^�Ϋ��b�4m͍����1[u]�÷ϡ?��	�}����K�߿ψUY}���b����8~U���va��L^kbY��o���#�8����V���iV�,t;�����}+~����"�T3�?r{吝�v!��H��}�6�x�:,,l�s%�y� �n�q \�I���p?k!��}*SW�8�-��nq �{�')�!,��J����n��뷆ծu^lM2���v�yq$S��!�p߲Q2t���̍��֥�9jc�>h�@�Wc�ی2O��Gي��x{A��]�z���'�Q�MV���Ӈc��Ҁƃ�+Kk�υ�]���kCSO��m�ZQ�fgg���< ��+VL�|C���;3	��7���wpҁ��i!���\��Hz�\ѽ";�6��Z�e�_&��޾]7����Nl���%�%�Ճg�߼!���MG�qX+�����O� =�BN����i�R�
�����f-�4ӹ	*�*����-�/͍/�g��=���i�վ ��EY�,�+��5��T���2�{��+��W�E�!����*-�ބ�Ȉ���@<Ō�=�~#pϊ�>o�&4��~ֵ�m��6�+�����4"�ݔo	�兌���ܩq^%b���'T��t�υk�ץ�_g��^��Gc��^͘�������<��u+9W.����̧�� ���Ʈeg�aq��9��k*L%�BG��R.��q�����{m���&��:��Z�I�@�A�e�̬AB���At�V�XD�B��D�v������{ق�>���4M0����i \�3kW��{z����~�h^���@��ho%8W6�lw#;�H�3��A(ȝ�RgV�#����L���"��?�zڀ�����lNn=/���+(�]�VI�Z�MV��e�o՞(r�����R宪=E�ae�-��������T�b�:���W،�/F����ͼ5�D"7.[�6^�3ѭ�:�Gp[i
���NJJZK��f_�����򎺜���W��(o�(|(�&qy�,��E����;�YwWȜ� ���N��o�<W��+5���85����Q ��5>�Ӷ������p��r���w ��-���f7����3
��)<�����#��žaB+Y+������ �CW�3e��R�O����Dژ�)�<�T㼁SH��<b�
�tɾ�}�9����8=䠚�<�{�?77�θ�f�����q��ǃ� ����U�4A�����~��*����9�U�.>~�`��#�4+��ȴ�;��5M��ή#�			Q���_쥊��������{׾sip:���B�ˈ��xL�b8l{�Q*��~*��g^;�=M^�����XX�T�ݝа��asN��)�~�k7Ȑ^�9���)?�����M>; ���f�W�U�טĀ%yKyL��W��Eh|��^w�G��^ ��΃ܞL�%�H�K,�DR�����M�z����<p!�'�S��� �ER��Yw�M,mQ��]jm9��ϋsː�z)�?�S��?���h�I[d�C�,\1r�>�x�q��_Uj��:�ޟ�[�d���mo�JE>�	��3G,0�NMgU��BeZ�Hv�7�;6e����Ih�ou]��܅�o����1�&��BY��xb}���۠���.�f�۹kg3'�.�Pʜ�<vSs��@��}�j���s9?��\���î�!n�]�3	�%��(mͧ<�ؚ䕑���3}0)����D���L_�ޡ�UKFJm�=s�{>r����@W��a,���'�%�x y��y���%���3a�2�����!x�Q�D1S�>ZE���w�Δ#bX�����];�r����I��H�%�r����W�K�=���w�{�씏ݤ����CF���\m�O4{�ѤSl�6L�3t����DW�/���$W�T��J/��'n�����|�f�I3C�P��C���u�5��T.�s���8�R�;*��=���L�g�T�d�.(�8������T�?�,2@����UBq[XK���~{�V2f�঱i��3�ޟ[�}��Չ�u6���7��$7I-O>����Nf7�"�fA��WzQ�5��:��4�k��g�m��xI�-glq��Q�P�{i����s<�jg~��E�r{���^^��T�u�s�S��_3-��N��)=����P�<�w3^g�ƒ0U�LQ17������tϿSV��ب4�C�fbg�����%���	�5����1�M!~��a?W�s�y���#�bdl���J�Ւr��Y��nam���g��*�*+�a>J���𜏮0O^�(��z-.y���/]�s_5�+J�,���W�};����*���.�yq�����~ϸ/�.�	���q�R��g����˦A;C*���g26r5ĒÔ�<�{��j=|~��(%{@4��G��������|�=�IˢS��SWC�>vR�9�It���4����u��c���~~~.2rb�[^f�(�� ����#��tԾ�7��c�ø=]���?ѽp��5 ��	��,2�@�[Zla���n@=��N��r��R���M�4��E8FQZ�̘D7���h����{L��~��ف�qG����is_���і5K��g��u$���t��U��̽���q���^H��%�-�-��{�p+�ι]��^��c�{?SUL��"nm�i~dn:�o̇�5�g��|���fG�s�(Hp�a��Οu�����z�쉷:2oa�-כ��[�7���M���ꁱ؇�>KO�g�����ĉ��E+�uJtAr��7"׃D�i�s��{�61�I�k�f��Ⱥ .���5�tmdW�e�\7�l��j�N����C�;s�������Q{���F6-x����˙N����i��gA���هy��D|�\�^�͗�Զ��=eLDAܧދ�r�0�(*8�����{��
 C�$y�'.���r#s��{���^�\�.>��(�r�!"�͍�-܏��7n�~8+������{��U�+Ǯ�������M�x)eii�Hŷ��|L���5��%�1���y�^�����0����uA����-���%RU�^�x|sSd�����Xlݱ�NO��ZJ�^�;)	,�i�6Sj�f[�,�v�Oa {?�oH~)�dn����_J����o�sC�cB�����H^�O�N������G{�a�����9m{Ϻ�3�r۩�O{x9%o��:�Y�R��[?��,��b/�����f���҅\���9ʪS��l�����i�^ؓ��_"�ok����������x<|p�hl]lJ����t��(���x��X8��ƫ�Tp�N�&+C����f�4Bk�T�XT�)�(з6^�.(��#�.��b����c�8�Qw�$]��î����IF�MabӒ�4�X#o>�r�H�8W��*G�����:Ԕ�����8	�";w�Аѭ[��0geΞ�ie!��c�}>A�������1�{��ur�Yn��MBk� ��G���Ϧ�5S��v�q_;.-��Ӥ"G�_ ������c.��)��
��^�w��Ӳh�Dr��Tq��$�D;��
�lQ/+(�@�Z��d2⮩M�0��qU�m������E��$E��WS��k��3��ф�\7�Rq�vؘ~�1���S��ވkv�z�j&]P_'�����mٷ{�i%���h)p�0��_������qll���MH,��� ��+��-���p�jri��gu������c���^�ƓМ&�-�ikkc���Љ� �d�R���H;	�3↚hlz��aJ%��i�bn�~��~L�i�G�y��sڂ�3�i��4-�G�=�dL��i���[�wNLX�)U��K�B)�i [����)`0��S˧�����xT�`������Pvv�T+�(?�����~)���.3;��\��P��Z�=�?�B̻|j��ݷ��1�r�����ɀ|�ZZ:������ϝ�hE~xO]��PKq&OՉEi�X�9-���a]D>��M��V�-"�>gg��z��eaUU��R�+ˊ^��7�}�V�LU���ӱm��썟N���;ĀW���A*r��g~���)HUTT\m�-�Y̳�	0f)�v�<��&(��Y���*��Y���J��v������4e�,azf�`�ԉ�B �F���W�!����@F���Z�GN$�0�3��'kʠ�a�&ڳ�:/ۣ%wg����C��)tꍬ��5�$m����k��g�i ,Mj���n�
�X�-����j�f�����k��+����xك�+|��h��,L3�&�˦_+�t{(����-���;��2 Ԇ���?yO�X[�%��AS��RRR�|�.�T����ɛ1�)�הwÁ=�+�&��=��ȖJlPĆ����'��"蒢��� �|CT4kׄ���-�������7�,];�~Ӑ��oQ�Ǥ�ĭ��*�r�/G<�����:::�eabdt�|�bzU�8N*w�����.~�'�ξ�%L�V�Y��7�8K���܄�7���guy�Q�0�B����k㶂U�E�k@� ���L%�}G0���6��:?��,d�>hgg���J-LP�7I�?�]�9�QK|��I˶��V�����<Ƕ��VzY
�O�(B���Aך6�Sf�=�Ҭ�v ��U*x'�dd�����`;�D J ���#��@�e�a
L����_R�� �ڈl-��Y��k�ܲ1ĳ[G�����b�]Y�DO�T/>q�S��1����@�;v8�S5
}���!�s��������-,=�rP��´����WHY�,����E�AY�2���0���j�3��u�#Y�kǋ�(���щ/>���,&����k��r�#��uB�Ҡ*�F纼X,;��8�2Ht�����2Uw����,�T�H�'�!�i��gd�}k/��e=�8 G�]HR�%vO���S�G�V����MT[����)����N���\1� �t`��݋+��zK_�i�W�j?���IK���IT��i��iG*�4�^��$G�X�&f�Hy��d�7[�����ޚ!s_Mx����LG��WV�13��rāg��փ餙2�P� �d�&L����*����+��ʰ�|f(2M�� Et([����
F��؀��Ut$���iV8y�&ט.��4Ө�P:��m�*p�q��=��3#):������A�)�e����ۭz�K��1���^}3�[/��s��%%E������\�1_���)`���E`�*O<��7��ޯYg��WܭSu�\�,5�΍�|1��s�O����Ǭ� ǉw���r�.\�6Ă1%Θj?[X�'[�D�8�����3����z�kD�3 @��^ ��}���f��e��L���-�d�۽�o��t�N׾���\(�*��~O�4��
�'��v+T�����a+/�1&�β��!ƾ� �H(toƫG���D\BL��G?=å녯���<ai�S'B�8�u*��blT])���`�:L�
V���
C;�MIvvl����Hw�]P�N�=��%�^��E��/�����M7�nF��Nr
��P�Xьw(����	eI��������fg���m��ށC	Y���wA/��8=i�KU���)��#�������C��7��{��?���e�C�<�EBe��VȮt���gh�����J0��V- ��.�y���7ѹ�d�4�����	�A��}h�n�g_�,,� �6�Z�C&�&U��ͳ>vޅuE��M�-���=��w��҈LF�W��N~�;0, Io֞nT�",����G�ዪ� �Rlh���r�)p���R��At��ȴ�)�Z1�5M�9&W���\�X[�*k� ��< ��wEE��⊉�*=�.2`���މ���@Ia\�Q��>��Z��bW������g��V�PX���|��@g�f0)R�W�% ��4_+
K���Nwk0�s���>��Ws->��k��q��3�	��';�j)7�BՔ�A�����_������2M�����r"��k�,tO���9>�T��3E	����޾+d�q�iƢ@��#�,���C�е�z�=2�*dBq���A8)�Ca�R��Ћ7ʜh��W~���e�'��0�@}c��R�x=����Շ�YV8��"B_!w�S�{��fg�ކH���Ů�y=�9+�)�?�잾 ݣ$�����Yݥ��?b��D'��;�㭲jd��2h�x0Ug�$�9��3#�;��2ފ�/��;b�\�����d����?�id=OU�����%�)����f�T;}�U�5�ia�����C!�F��\q�	�&��8����bO�8�˦ܧ������{�PU��eu����3b�`
|J����A~( ^�Kvnn��e�IK�8̱;�L�Y *̢셆��0�b!��� &���Y��"�F�L�GD���`��R@ iD܃����G刦,AL�%�������o`h�Q�*�a9��Y#V�߈�]s����E�\7��5'���׌��v����{G�ϳ~������S�Or.�l�ؕ����n�m���G�|����6&��,��m⭂_o���nW���ܜ	� |��=w˚�i�F�u�^���&����)_�gn��>u�
�:og���#�tv�7����� ޠ�-�������\�pU07�d���$$-����
�����$N�¨Z]Yr~��JQ����셔rF_��f>���1L�	(.�Ϗ�"BA�"�g3�$+�2��@�QT��Ÿh�r���Yu�#�l���h}��@i+�׺�sw8��������GsS��@>؃��
��US����iL~��NH\���碱�0�5��K��A�	���B(���;V�YYY:�~y��<Y�����j�"��Y%����,<������r�'*�ڡ�A���B���˵r��PH���L�E`���h�@��v��ԁ4-^�zbD��,��4��4���qE�i��*�T_SSs�(S0��>���#����+�ȵgϞ)�T���c�EW/�ӳ�Y�L�(��J�x�dϾ�~���ed �6��_L�E0裾��մH�""��;��!��Rq�%��c2�:�S���D��W�B �IɆLU�#��7��567�����,��H0����#&ba�G����M���s�{L�/K�rYi��X�E���ڡE���ر'O�d�znC?_dڬ��ke�K��Ցn�ޛP���C�6��`�znI�=%�>�$���.1-s�t2Ѧ�G������E}gcc�x��K3)�P2$�%=uzE��&G\�>mm��u��%&*�9���z\�;����x_�U������_а�a9��T����%V2�|EZ���<ձ�W$��+�s���1�,�V��kaB����V�L�j0ɐ�$���h}����X>S33��NO]Y��4s��Lj���t�R���>������(��:#�<��+UW6�+ҫ_��"��<�J!�/2>|��|y0��G���Wi��i?js����t��P���i�Ӈ;�'&�R!p�tR ���+��3����!b5����Z��_T���	���;v�嶞jh�"����<��A9�=b�|o��@�����ᒍ7R��{��݇2&Kz�t	'z=���77�K��3z�]z�Z^�BM4�Y�5.�Epʏ��#��6lؐQ9���N)|`�(�����EL�*�_h*%�z���c�8����Zb��.�ۧva<p�mJ�)G���[�?��~٪����>���9͙����f��,�S�}je��5&������ޗ���N_r/b��i�.��&�~jV���ȉ�ZdhTW��y�)��~�K�4J�>T��Iu�����ҽ�?��n�ݿ.�戳"�_v�.�
M}���&�`M��W�֜Qn���EY[�B�y�g����x`�i���0��xu��2��r�t��%Bk�	�D{�{�
;+-�3���;8�Eggg>�J{����űbB�`�E��.}� ^��_��8�k�,)Đ\�])��Y<��s�5��ɽc�a��z4��V9W�?�J/��g'G�4k�-|���!�Ǆ�%!Pv(�9�o`X�(��۲Jjq�n���?�hR�LE�K�\X'�\�騽�`��ֳ�+[�W�'���&�o5(�ڡ���i�f{���#�C�2/�NT�Y��B��V��&#L6 �2��B�mz�Ɍ��=v9��^-���/�&9&�HHZ�s�ӅMg?�o44��z�Rg۬֚�WWfiz���'��f�׶�������3`+�ap���3�� �W��	a��kg@�2�g����&/�ȓ�w�ޅ���W?O�>Z��[�C�U�ϋ� �f��+���]�d~��(���k�lk2��@≫�b��M�Mxo�E��H+*�k�=;�w�թ����W1��&�ѝ��Xbv�xɟG��^�r���YRܕ�55�l�6���4~��ƣ�K�T��fi���}�C�p��9��ݠ\�B/�o��z%u��}�v�Z�wؘ��E���c^�yt����i�
����VI v�XhKpA����|{�x����/rำ#ή.r�s�Y�Y.'�nA��u u5k0S�Ae��sh�}�C8��[�J�tuA SKt}�ї:�8���"������&;��[|f6ZY]]=��@;4��DDG���]���9d�|�dD�<*��y\����|�SW�|����?|�9h�f�A93���u�(���WN��aW���1>�l�XKh-���1�?�]�`,U��եN'����JP^U�s�X�~!b��6���9�ef�xt����SP�O���u�K0�R)`��}ro��T�U��� ����1��g� ���Kl:�!���������%��¶�+��4�B����G螸��>s�ï�C汨�5�[��F�M^��)�7���9�!$4�b2B
$�YT8e���P=Ks729��\��|~�5�{�O��r�/�0��	��������^�����P@���r0A��2uB�hl�q����#�x�o-���y��q60pn�R��K�_��7\>G]���.@�$={��i0�oEc��Iv�a	X�q"��{��d��Q���А^-�{Q�>>9�K�������jg�+
�N�$�30��U:Ag!�(��hdsL�IQ l�t�Ď�F�B�[�f�Hh�Q�B���a�Ԝ��E ��o��]�CBړ�db���̄�Vddd��Q��4�n� oz�B���l�bF��8Z���|2TI��H��K%i#-cc��k��ﺘU�]n��������:+�2���:�->nU��@=�8{V��-�| ?|�p<��e�Q%��! �Qkǀ6V�J��P�].�1���T�VG�����5����G���V��i���;w�P���O-�#�D�WLtV����E��+W���θ�i��Xg�j���j��k�X��7u��a��a�Z<�e��)B*�$��ӽWV)�Bp�(�y��wﮱ�ZK���O���̳qc^`�y��7>�pO]8H�O|�|V���N����5��Z�9m��F��<�MF��΍M�0G�A@Z�N�� ���Vϊ;�T�NS�pg?츱�1���r�װ�B[�e�j���Ӷ��""A^��G�/��������az'��������U��c|O�~D�AjS
����J8�qk��GSr�����$-��9zR}r�3�d:��\�=�_�}����Ev���;���Z�\����nn����8DE�^ɮ����e��&�oO������tw8e>h�	�T�7--��6Á�������6�U�}���.pF�5|i<uzRSV���xaaA��ub�B�/JR���C
g��x$C'�6��Wt�	�a�����*uh����4xS����dOC�.��f�1������#^�'��4�7�+��Tu�>�˝cj0�Ư�L��(����M�G�6�묉1��/��6999�v��ˈ�l��,�c���c�[�����Щ�_��Acу>�Kl��������b7sy|�K�.�}�
O��---g+�$�L�f)�?����䕵-u)�9v�x�,�B�����E�#O���Zk�`���KU�m���3�@J�gپ�� ��󓅜R*��{��V�ᘕ�RU��L�q�%�_Iw*��,ƣ�ˣ�nD���G����Ƞ<���σqL~!>I0�D�%�'�-�E�AE�d�b|���U�B��
�g"n %\Er�+�~&�x�ZX���ru��J��%�TU��@�q�9�[^��0f�װ/h��Q攁֫�Zs��A�~��t,/��.P��V>x��:t�O��,�L3Yç�_u�����D �]P�PSJ�^i��@��ĳ \�`L�;0�X�AG�K\�����\��U��E�l��-�/�V��m=!zΚ�1�x����T�F*��1�Dn�s��	{v��3��05�ʃҺV$��xg!�9�#��BQƭ�D-�1S��0_�oYQQQ�&���M�� �C��D"v�fh��$�����@/&/�f��C&���-և�E����3*V�ּ��>-Z���X���B7� d�z�f����34CF���vvp�##��]nDO�R����K���G]@����(��-�/] z�@k��s�B��d�����7�!�<hv?T����0��2��0i~ Ly,�:�Y~3X$���nB}�B�sWsB��������(���uA����0�`��^�����K�����!!�}t�� ���r�+9!�<�9�S�{��3=~|�k������\�,X�3��^�=��������u���h��zt�8��G�G�am�cPߵ�ï3�����`1:�I�R�;�Z?�R^ϓ_�A.�1�6�*�BN_�T��Z��3�%h�,����?`����^�r�̙��<��o�rj�sx�z�7�R)!�!Ń�P?�����.4�mS�.�R�|��|�r��d�"8��1��ȅ��Ѫ&8��"�>���C������j������:=+���q m��{����]%�$��q��[��?<H����J��Z��&z����Ї��r@���1���M����,�)1�g�UOHh3�5XueÅ�(voP��}(�fؐ2����bbbBI����9�1��!#���Λ[��/!,�b����ծ��2��'���b�1�������1�R�Y���Q��I�erpŪ �6����p��p%Lg5����[�
&Q/����f��$��̙W�@$�1��?qa���~�(���L;VW�(N�SrD�?j>��J@�!%8�����/Bs�� Tq����r��-+�$�0�����D����܄��a^q$�ۙ�3̏������ �;V����uۭs���F�>�7ONM��ȡ8��&��9��#��5)� ��`'�mbB)Gq��@sR��?�Q���ƻ���kG+�֜ሉ�v�V�Ѹ$������Cq"�L�Yn�O[�T$2&#e���)���|z��Qt��{|�a�B/��K/�A�d5���jP��>l�X�1}	��OK�6�W`��PWS?�G}��*��}� H�v ��EK�D��l�5�~̡!r�d������X˂�c~B�����}@�/~�Ki���ʏu��&*5p��9�*|x4'?]ʹ9�l�~4��B*�$7P_�,�0,�;��r���˟Z�o���{u8Fc]��g4h���,��)�c�o�6G{�|+G\S�-��?_N	���.��Y$��M�$��ܘ�e���6�l��f�wJ�Ƣ�ⓐ~o&��R?��ţ��hO=gO###�bS)����'����VU2Bf&�&�^'�\ι���bf%����)*��L0W__u'6.�ʿe˲��9��Ļ�X���y��}?'GR�.���򤌵��A�AL�xvN�gq�5]iQ���Ď����|�B�T9nj:7�����3|m8háx0�@V��N��7a���@.����ѩx�_{���)?�!�O��̙3�I�g����P\�Ǧq�f��#׷&�/f@%�Q�.��BW��R?����U{���M�234p$n��t�d律�85h�Ĥ�\iU�=}�T�_��;Б��={V��kz:���q}�3�hvN 3u����ђԈi�"��0�\���tQ����&� k��z�E���|��ڹ4�&���q�+�Ce�S>�As}�db�	���X�ٳ����Bx�`JS�z�3�8�e~�O>�`�wr����Δ��ID��3	�.������A�����k]�Ĥ>�ònEgDG_kU�o�T3S�P�s��̑&�2�&�n��X���PMi���[���
��>�E'���{H�r�^t$
��1��2�i0N��Eک��kd��9{*,,o����iU��b�/zF�!�Ɛ'�pD��BMMM:�kO )	�m�6�`ztv�.GtV�_è��	!�rc�*�ܕg�5+P/K҆_�nd�/�&������DuG٩�f#6Z=˿^hy��4�A9t��O[�����ب� V地`����߽-�����6�K*gs�R��}G�42$����0.B��ٓ�|�M�;�k�T�ǃ�E�_m�z��S��}�ca�#������M셸��iP~�^�
���0MN��������7�M��w����iY�_n���c��A�;���ߘ	6�0u�۫�t�
c�	�a">���>��d�	 �ܨ6��fy��q]��44�ak��訣��g�x�a�?���W�_��
ş�Lr��S��,0��H\=�ﲄ���ӓ}v�H�<������G��Cj9_DE������QL"�9�2���x��#1	�`+�w�W�f����j	?'�~�if!��1�2�/����ӣ��'�� Ă�#���n��!/K{Pn"&�9�u/%���m
[��k_B��~B�w)�����.d��o޼ق-�OQj)W������7F^ ��\t���뀤��i<����A!2_H�x\��ȵI?�pj:��DR�2A���e�
'v{f��\+2�x�kRY��B���߁k0�J&��(ZgSgnB3z�3<�>an�O�F�W��mv��U��v�z�<��c�1i�k3�P�sƆ7J*�N���_[�AV"L��bZ�W_�gL?*+�sЗ��H�%bB��5�,"4��x1*������L�f>��*�p���iӕ
o{wa(��Vt����{�N~�oW�2/�F�o:$	���]h:���Cg���gҼ\Ah��0�}���)A���8�G�Ѽ��y�����_{Y�`~���%0���Ev+����L_˳�0�������h���Z�xLtt4L�{�|���Y�9�����ӞE�V,2[���0�)�{.Ȝ6��K�s~��x�J�ẁGǨ
���i�)�����.9�q��;1�P������'�ra f�'ںW����K����] �0�E�����|a^eW��=�/�(>)�L��S�o@�M%.2��?o;/i����R������Ar�-}Qo�\�u 5i�y5u����^aQ%]��FT"
"Ia�l �	
B+9�����GGA����TD$'��I�� ���&���<��}G��{0\s0v׮Z�^�Z�v��3������Aݤ�ݛ�~'�;��v�	
��j1�c�7Q�P�F�ƢR>|(���� W�Y��&�6{3��.��a(�d86�$ɌL�8�W*s��d(������,XY��
*�r�2Ms�[��C�.,�(�E�9.��T����n����y2�bb+fʳ�ͫ)Y�@��mPQg9��Ku��[�DK�l/Qv��m����Q��F̸dgz�MړTX��R$/uS8~a:9���NȘW�ߐ�)~����Ÿ��ƈ�� �����߀e7�+w��8��J��䎯,*�x�m�(#08A!�h ��)]�i���I�Zl[�S#�Ӳ�[��6�H��E ~��t���u�YEE����h?��<���0���Wl�_$�����h�V�*�����^Ηs0�a�x&�Y�A�DԻ=n�.���Ҍ�?,��3�OW���^&�`�߷�Y�0��0�4��&J�d�9�Q���������|�q^�:� ��д3�%,�RS��C;$x�����u6Zu}�GCz_�%Z�y&�:�j��?@�K�o���9}�zYMiF*���ƙ���ۛ6Oԋ(��C.�ȷ+�Kn�7>�1�u�Ƙݚ��Cs��e�/l���H�{�rr�7KJ�R���ك��Ʀ9+(���p�Fo@+�{*~!��zۊR|��5S�'�&>FT4o����7D��bo��u���>V�����$:�_��
�n�%�(��۝��X�m9������f��j�m՗{H�t	�b��.���Q�ƙ�ē�(��'8����>��j4�X\e� }/�HbK��������г�l�]�{]GMK��#�K���n**��$����A�xzq���a6*�O���NKM}>"i��PRRr�j#7���z{�܀�2����ݲs319�w��*��<����-�2ب# .�.så��Ν;&{�iq�|�X�(ecŧ�Eiih��j��/R8�*� �1X�\R�N����%?�4ΎG��|��d#��y��1={I�{�(j�󮃃�����C���P��GH��F��*�h���I�m:]�Nbm����DV�(���a�8����W/g��M,
8��Xo���Ǎ�w��5��ް`��#�uY�
��vq�GJ|p���ݑ�P^��j�(�܉Z{�d�������!�\,�5�%�5���#Ԟ���y��AP�������s� 
~h߶��eDEE���(t�D�yDM�j�虛��C�J�p/�3�ؼE[�nK(�=X;�E�6!du�=��=��I�Gл�e�Ѽu��3M-���(V�I.--U?F���o�N������P\ ��P`k8Gg��������p�r���ІF�~�22��?)^��N,&�-Wmy��<��B�.5l���W� o���]y�P����a&�x�}�V�d^Y�v;~L�3��Y�]{��9���{Ӧ��d�-�X��{�X��J���h�ek��C-�U��o׿Z�_/��1,�*q'������/V�wv�>����Ct[n�kC�vB����8ScN\]�����N���W�L����6΀��Vf��\lll5�+��w��q�[-�M�;0�Lǉ����f��W,����ө��_*ʬ�y����FƉ�uZ::�J���헆E{��ƨo�5���˂���#<Z���}[���ܗ�Pt���ڪ��w|B�&��s�h*�1q�Ӷ�ݕs1�\f�ѿ�+�螢��x|fD2�kc�6|�1��f�)�"�A�"�T;T1������tccuq�������9Z�m�S�OwlZ+V"92ɫ��>��.^���G��Y�9QS���xN�u7��؂R��zfC-f�m�C�Y��Rl�1X�܋y���,�Γ�M��s��\�P��;���bϵ�sPh��BO&@�հۧ�'6��HDX0�c5�|Ý)rq��r���%��t~Ь�N]8_2��I$(^�=v�kK�o�N
�=\���?_~����"@	1�W:+��"C�^jXYS����̉mo�M((*nPS`!��ٷ��\��ܒ[:�1�oLnM��h��uJ�lo>ʭ�,��=�M��L�u"���_��5����E{HQ�ֽ�ϕ@���Z�t�9�����j>h%��������y��jQ��1���� �P�p�Y��ϱLD P˹��tMN2�"��"n�����3�B=�4��F��ɖ�ٙ�g'M�t�F�$�z�ף�P:�� ֈj�s�8*�.�f�:�Q�F�w|�k~N�Ѡ���ά[��ڊ��s��8��M�/��1�h��r� \��V��]]�}����	W�Z���{���^��=K������n�\�����HZ�p=�0N��j�E��n��({%n�(�8�0_9g�T���Q�p�>�fw�׀l�x�q������ɑ(�K�n�/�A_t7���}oDJ]ys {����ӡҙA3^m��� ���<��ʴ��IG������\]�$��6��55��� �r�����n�)so�A�CmjjJ��	��0�h�}����x�hSb��x��.�ì�f��i{��.�0W. �UѺ�=vu���8[R`ոBaD��:��Қ$�3���5��bv=6ײ�@B����r�\-:��n�(�����	����OCG!@'}$�Z�p�:Z̈}��*�)|������#o��KL�9X KϽ��,��h��D�Bt즜
�������߅zţ"щ.����� t]&���{��9~�LmJ��D_E�׊����D���jJ2BBB��!�E�=~�������qC?����7�3�]�o�C@�FU���v"κ��KG�������Ў#�/5S�>��Tםk]�"y�u����Uƿ��j5'�w��Á���}���CB���jG�|ʢ�s����ڊ���-��k��P{6���	�effvW��V��E!��!�#���nmNF}-=�֙��t�L#Z�� ���6Fb�HAb##a��V���z$ lT@�סŤaEٷ�����u��{��`��j���y����a�/�J��PSz�S��xP���P���J����c���F�)󯼄�y����K���Ey	H��{kKS���^�:��`?c�[c�ۨ^sb�p�0���q�p��L<B��2�(�jn�@BWd�ޛ��rВ��L@���J��J�+M����yKeި�OVS"��0�Ļд�[��$뉶T3�\ _l㨂�N�ݰ ��5r�j�
���7~�;~a	�6�񵰪�ʈ�N�Q,�<��(B�XI��.�ͣ��}x���Ld�	�m����ܺ���.@w���	h'ӹYJ��?}���
6�pa� 8#L)�N��5���X���g���f�t���U�Y���G�er�ԓ�`�m�֞J |~�����৯�W�?U~g�|���g����߅!k�Z#�#��ns�~1�"6��62e���x��|��FУ�����1� �j��Dąu���'�-�{�:@�ZDӮ�;�qB��܎�L�<�D8��A��G�šq�l�ڢ��El�\
o�l�(�;�ARZz�=ں�����Ϩ�y/�s��>!a�@�ܡ�,_�`9낖nO�̽QΧ�H��Xȱ�uӒ[�+�Da!�����f�b4��ѮA#pN��}�3����l�e�7����F<&z%1u%od��h�e����Ŋn$K�J�s�șnTo4��xc��I�QJ���f���IF���O����(�D�S����Or4�����l�X�T{*`zQǑ����W.�P����6V���\DHh�9��Fѧ���P�o�_��֏ʃx��G`�ï��t;{��[h(�����ZP�n�"--�G{�	��8:z'��jK�aeY�?=� ���Z ���4t�/a���Fk�Dkx=�lDVD�Z��]�b#��ю�k�+�A�n���oN�:e��ʎ�PE���"��vu�{�;�m֣_UOF���	�2J(��g��y��V�r�
��8>�9�ޟ�4�A�Y��'�zdcTz�ؐ��U�=�_h[�{��0^�x�܁yB�=Bԛa��̧��a���Dׯ��d�A�YpK-FQE�[.C�@�n��9j�4���2L�̐u��~�L�o/�'jn�P0�&��5;d�-��.t�2*Ff��H"P���:!Pi+b��؁Յ��aǈ�����i#w��+W��(Ц��$D-)X��n�Y(��*2��I:Ա�D?M+kP���i�e>v�gx J����f������~a��fG�����G.�W�����τM�������A�� ��/�a�[�1�*��Qq�wc�c�S�d� a-h&���맶���h�#
=��%hy\=�|���s�����C)��~<~͙�΍�Eg#hu��9���ó��LW�9 �?a&+��
{�99@���P�Rٝ�^�`��<t􁉝��r��E��Ѳ��1JQQ/h��=P�5��G�99��*>qcX%�H�j�J���(|�z�G)6BV��G�v@�i)���X�(�����C��O?]��k}�5վU����$~�G�3��JԼ�(*܎�h�D�v�\��@�U �h0�R2w�]+�qv+�9W(<Ƒ�z������.59Ab�)��eo���`��W�B��Mre�eT��>�����r�Vݹ���e������;���o�3�2|͹^�#ao\l�X�)|)׽�|�y�U�ۿ�]D��r��5�vk�Z�3}�(���������T�Hh�3�U�74�2��y/tУ3Ӵ�!Xj��[��F]zkI�ᙠ����I��uD����޽�,���/��y�ǣO�Pb����yg\���g�tu��'O`!�U��3wS=[; N;�L��$�s/�����/v���h�熪c��ֲۺ"I/	���Ӥ�1q��K}�a�1A����E��
ʹ^���s6����F{����K8���>��;-V�ڢ������aK�������*���6�U�Z����DDD��4��/1`>ѵ{�1���K�$�����2}uߎ���-c�0n+��	�Q�����(�;��[[[;$Pj��$sG�Ū�����qd�I��P
�bz�q����w�u�� ���D�;��'����X���hN���;���].eR��K�aaaɧ�װk��W�a�yj�19�b�`��[ï`�rq��ٗE�H.Q�{aB̕S�BѪ%�'J�����2Ѫz\I����(��|4���H��.���RKMȢ��VVV�VS��K�}��2HE��~���Z8���ljkk[CK�7"{M%j��[YZ���4�p�!�u�""ޤ�b�4�����VON���-r��v�*m�*(X%FFF�Ft�`6�E����-r���{26<\K7�\�x:vCv��ҳ��X���wx�{��[�h����I�C� Yn�[���ݩ\ŶÒ]YY�ykk+3̍�<�������UG�.�Q�q�g�JB��Ƕ>�� �s��L�&%i[[ZY���Z������gk^��-�S�<Mg(��n���TR��;z$�=8�.�?���i*Q=��:����^%���k�Sy�*�tq�ف��d̵��.DWG��Qs�FLr����|7���O ))����cw����X���) ;�a9|�6�o���ɛي�,+�>����g_���l|E��bsT�v, o��N�hX: ��_Q�ш^Ǥ���9�B��߉u��z��[A�>@�����e|||*Ȳ?���L��5c�5#�������l;֭�kd-�5� ���w:�s)�M�U_O��cf���C`�$--��WWN�'&1��}�O�#��H[�/ϙ����-�v�����Z��χi.��9Rc�i���9k�Z����mJ��y�m����9�T��V+c�
�aAO/IJ
�h@��	�m��"zFF}��R�����#ȩ�	 �@�������U�I�ǩ�ڭ���a�����@)���:���l�Z��'����w$��1 و��a�8��L&`���鳥n1�Q.��i��x+��9h� /X4f�Yqq�U�jx����A�C��P�!Fr%ܴ:8�՝�R���b-7'��D�<���m{<�ɛ�D	��.-��֢n�$ә��������]^0��b/Ȇ��;����d1A����	5hQ�JdOL��j�D�0� �`��S����0�}��҇���i�I�>�I�h�O$��Ƕ�w ��^��T����w]]]��������q]|Z�C��Kk�URjjj?�V���2��1=WL��詹H�\�������h1�
8�V8�'�4�љIUv13''gk�3��p�9��L���I`j$7�'`	�J�Ұ�/,[W[[�6UN�J�ŅA��{�K�m�:&66�M�e�Kǃ�n��x�E�T"��hi�)��p�d�6=�����}�7�u����f�׊�ɛo���4!���|z�D���KH
�m�s���FƮ_��o7�8�gy[h�/��Ɏ�2�s:I�	f?a��*��A��_�~�@�BU�qI�P�@]p/��d6�q/��+���W�x� ���W���Յ�Ku�};�Ҿ�1R�QV���NGFF�iX��AzwQ�� =��Idkn�,���>zpÕJ������(;gJ;��E��Ȣ�57�$'{ �_=����i�s���>O]��.�pє�#�ܧ%:�p�hZr�D�xWR��/^[6�	-�S\a�xzҸa*��Q<��D��H�CS���J �Ă�yM;��V��1�����#��f�
H����7W���ƚ���GD�g[��|l���HOMz��L���(#gӳ`OIr>Pn�v��J$$D�ٕF�ͱL�)'��7�h��t�\�@]�q��mh1�m:��ى��p7���}k"i��bj�m��m@@���u�ݶ��B������X����ٗ���ͅ�ƨ�L2Ȱ���tk�A�3#i���`BB���藗網p��ʁtc��0�E[>���K���e�����I]"K� ���%'i<.��=M��#.5%�%Mw Ŏ�����6��\#ϔ��Z{zz455{ݽ�f6.�y�;b؇3�b	!��P/��ȅz��$�"��\RA.���b�/� !i���J�_�����������_��:L"��[�H�]��٘�2�����::�2�DF�Ƕ�����$�f�˾5.}����޾�wIl��c򚎗-�����4�Ҵ��xv�7EO��ԟ�x��6��Hl�^#�Γ�Z�������/b���o?�q��3<���FY��t��w������>r*/d*��(U��.�`��aRmO��G��; �w��$������n?.}�m����)�;vn?�y���G6���0��;�� ��[��9�A��;����w��`�����K3�i[[kKN䂥P��*͡�Uv<�k�����5��YyFPKL4�ǦJ�M���h׹��`U�?i��N��~�'<������D*�{5���&�7zG����,�5�d{�tO��gCOuN���P�m7�1YX~W�O(e��2������]/��G�ߕ��(��$�N��$�N��$�N��:��^���\�R���cn]��;Y�~~V�̺���F�tta��f��O�)]�h/9p��|�A�R���/^K�z�_���.k�A�i��m��|B�c��dd��~k�l��L��߼um�S.����_8�DMK��|!���m�U�����^+r�̒��5�����2%�n���&���	�j`��V�q������Lv{����d���tJ�o߼yS�Ӷi�����Z���l�K={����#�$%Y����ŏۉ����t]���&s�ۦ;r	-�sn�����2�v�%ʑ�B�H���/4�O�Z
S)��iwR껗'''�tѭ�\�BN>hO��:�yS�2�w%�3�v6S@@�D{÷��o���E�riik�޺u���j\��5����:l��h��'R��
��9����$t�졡�!P&���G�
3�����5M,�5�[z���L�mm�s���������"/><M6��xx���c��"k
G���h�G�f�
�j�kj.����x[�P�9Q�P#����+Մl�>�S��j%����,uu��10lmm��n��Y�G�w���w��+x���_!���-ujK�s �����D�/���%��5�薙�w����aq܆�n�<E�ף��!sss ��\rKfP�$	,����{��2�M3��X��酄������=|�L��`��]O���Ell�B��WL��*_����C:�r*�Ύd;�����Ɨ�|�t�b}}=G�uS�{ɏ�u�\rr2z��Q66U)��ׯ��G�~���OnU�:�h7N��(�"::�����6��/4D�eO�����wO)@��q���Mݜ���;z���I�o�2���g�rS:�	1�m��7����dD���\;�������^�륆��o͓56��q&��H`�Z��b[�-ݜ������k�j�g�jWs!6a�ل
��!!��W�������7��{Q�C����xv��O��fT㏈SK������V$����]���{G���w'<P~�~��6�C�k�Ch"`�b2�.0Ḏ��}tYu�v�p��ϗ~[�2`J�y��c��7u�D���V2��#�6|7�Lo��P�z}�;���K���\�� Ο?
Oi�������ұ��$����;�̉�G����n���Y����!�߿���9E!�.H!κ�z4r`SÜ��d����.C�L�ƥ?oݍ��O�GD�\_yNZ#�6=z�"���͛o�o�R����R��,����-�B/����8.(8q�4�ޘ���v�pg� ������o��ۯ�-m�����Zi�?�������<e0���,��h
�eJ��}�g��.=1R̩Z<c���t����xL�㟔y� 8�H��~�[g�}�B'y��ʯU|E���IK�����H���t���;I/�x�Z�F�:QOO�? �E�ٟ���c`d\�Y��|A�̳q��KW�^�9����tKD����U����O�f�`���y΂�/�W�K�|P��j����!a�5Du6[܄E�bh����Bff&�G�o2���l��D�=��<uY��?� ��\I0ⓢ"�Q�.�[����O�u�Hŷ�EΝ�,��4K6]7���Ko�~֮|W'�d�������Y���A�� �6wr~U��}�*0+�����]��nR@�"�^B��x���[�v&��������>�_:�\߸���|��2**���I�3$�4���¼���x�7@]HF����Y�8��^�@�{���?~�7�8+$D�4�
�mDK��w�K���>�9S�=��c�Lj��e�
2M��t!))V�޽iit+�R��vG�����/yxQm'9��Ka/��/_���j6Lq�Er������="�^988�������i�	��4U�HnUY�(t��[�%�^����Р���ec(�{�Edd�j��j��e�J�jWTT���y��`���[�pAF��;�Q[K"�zK�n�!<�����|ڸh�O�����.���<b؉j�?��Q�v��*�7{�4�-@G<�d+��sGV� �0�*�x��_������ύ�#��8� �"i��#��-��SN�!bv��Wm�&;�I����+�}����
���KKI���6�?����M�k ++~�� �❸!?�Ú�Wz�����],��lSrr_��Ea�s<�$��e0k���� :�4D�]�f��vDGW�f�f	 �E,7EN2 8G{ö�g\���K�y�o�vK(@�ۤ�_r�v���a��$\������Qj���V�J`~Zj"N�6'�z�
���H��K�eQZ���4�s��%�s����������J�+���S7S��;�/�iPx����!�,�+�&爔IqY4m�;p�e�����/v����������ɟ3�h�x���rA�o��=�U��,W���1�Z�G�*�I�^ę+x$< '��{O�Y:�7w�U�Z
�������A�7�n4!$���<@+9l��m�t�MG�Ť�[zzz���#�l��22ޚ�1�="M��j)))M�S�n���/	�@�P��{M�.(	+���Ԟ���
�2������"I3��Ak�e�@�.�Vgy�Z}�dR�$^e�v+ �ZU�����|�����n���jrzJJ^^�����6�HF3��Dl�9�UG���k�&����F*��O�4;W:ۯ�T��O;#  �N��9�<c�� ��0r�Yg����oŰ� �ֈkʛTG�RQQ�值�eR����G����T3q/�i���	�=�ș��ub�M����"?�A3�*N9�e�?�FY���]�����❸�9uR��?��[�g'���m˘�ru��0��=�K��wO�$'���Ѓ�Y�ᶵ�Er|�b=`|��d����ӏ��Su��۝�%m�������[���~�Y+�z��_���\נ���z'��y5�8�ff�g��8���ِ��T�vbf�8"�mf��oۗs�G��|4c��oG�l���5{�E8v�Oك�ِȃ�NK��}�V�g^Js摟��~'��w�(t�޸��Sc��r�=V�ז�S�	8m�Rz&��\,��w'Y�cFF����x����W	����B�z���DŅ3ie�S�	p[hW\H|��a��<�a�M��ߡ�Lj3�����Nn{�A`���iy�/���'����.��3�~PlW�[Pf2nl�����ٜ����]͞�㭮�Q~Ǽ���M�<r>�6��;���z �N��Ӻ�YG���D�Q��m7'r�e��ڪ�����xci���Cx$���w�.,���F�ǩг�W"A/NJS�R��

I�w���uH�@X�5�v�B..��/ ��A1�7��WV���1&֠M��cI�I5|��t��qp��3�+����,ٴ�n��o"��H}�S���z��Q��ch(5C6�,�������T%�@s,�I��o�a0���M>�O��z��G�pc]児.2����d�d�ׇ}��НW�t�~yǄ��6��k�m"j�R��{,H���2�H�JȆa�N<��kݑ��}�B�������uޞl��L�l#�aސ��M�э���Zy��;@X�~����9\w.2f⦿��@�<��d�����c�W�[�A߳?��r�s��oY��RZ��?s�o#�*u��d�U.�>�2�@�Jp���x�I�`# ���m�%ﻗ�ݾ�
��&M=Qoo�*�6�7 �+l��-Iȑ���3M9����-ߞ��6�4�6hb�vU�̣�b�9%U�h��<1���E*^���n|��������{��׌H*;�G�'6t[(|w�q���	�j��.x��Ag��x���ϕ~+����l��wi�� ��	j84��[,��vt���}�k�Ǖ⟵LQ*ذ���7||�8!Ҳ�A{:�f`�Ej�?�h�@RS:���P�	��6����~�S�9�y���׫�8.Kw���rΣ=Z�鳽#u���ŋOo�3��d�.8�e�Kyz����VAռk6���9�uèc2{�	�h�9��� 4��aH=`�;My��Eԍd��e��)//�}I``��g<6˅߂����n�C=T~���B2j�K��̣=��:���\@��:nCEEu�q��kXb�y�6�E����{����)�qh�ݨ�׺
S~����ʮ�0.����{lߍ���.ڰdKۦO03M��l`PP|���=k���Νυ&�LWw��ǩ@�N	Rx-��O5�v7�췙-�����>یuZ8�p�K�L�[��߽��Ch����v�������md m��Ǐ���SR�W����[�&vvgw�=0��ދS������}��@'���,�]n�AK6S�y�g��1�����9`dȥm�??0������O������gƙN��^C�B�ƽ����3�:���
u�3���K���)4τ�x��Ҷ;�_��4���!���eZ�)�۷o����i��P���ROn�ai���������f6Pݷ-�N�T| ��u1W�˖
%� �&�"]��ɎLN\z�G���r!Jv@�N߻�i�� y�Ǐ��*#v���Z-��d�d��`�����X�]&� � ���T%��2�.F���n��N
��:�Qȉ"����+��ꧺ�<�|}�
���\�NGl�E�/u�:v����۫d��������o�ޡ�t�E{�QVV� �b�#��4��o�f�o�������_~��ٯ�ϱ	���	�ӞWlfԩhXl�m��
��?/I=�㿂���]���U©�Ǐ��LQ�PPаI�p�#�k5���@�?��/{�IF�m玚B��\�8�j�=��y����}6���8�Hʟ\�6�ai?�J��XF�R|�jtjO�ĘB�[o�<}��V�L�3�3*��--��MwR�f~�����b}��Kcc5�2�e�ݲ�N���Ċ�)��*�]�z�R�ͅv��ӽ�Y���R��xC�S���u�ܝ'�H |C��2p���9��Y_��j6w^����>r1#�g���X+i.�:�"�$�9�=m�\cĞFA޽˽x�/���)�,b�m�U���Ǧ�����Ճ��!$w�)O��˫���G�K����}�H[II+y�F��gN�rJY�4�R���\V��j{I�$񺄄ǲ��|d�G���g��������␚��	3pb�s��D�����$r����M�ǡEŶEED^NZPk�	}�ƃs��%��>W�����t��4�1�-�z�`CH���#��7b���Wä/�v|#�I.���j�G/=�|�gDZĪx�'��~�5I+�vuaL�sաhL�ڿ��[��WXzED����B��z#%�S�"�������J�;��o����u߳�����lN�Ġ%�7z�+e6�d��	&��#��E��#���5cS����h��K��}�Ԓ�������\�q�Ç��@�H%V�͔����k�J����$dc_�|�X�h�>���۸X�do�����U�T�2؟-v�gd0���M�p�c��^*@>dƋ�����s�52�y� ��v riM6:���7�Syw)�LD��؛\���������q�$+/��� ��n�9�q]M�������gG��H�gLx`���\[n�\��V��O�o���� �y~�kp�vM9�swĔ>�T|���}��*�*��G������II����&x�'�lm����8�B5�W{\�K[�|"qB��B��,���D�6�����y��˗
���Ǳˏ�;���W��;0�w�߿G7��}�8�Jަ�/d'�>�S�R�Z�B�@�H�������|}�z˩ǾQj��{���(tc��l�M]]��5�C=��ggmX�ܾ�]�:~B<.u[��s���9���]�VOP�䒞{�7�t3�M�X��O��NK _�:mM�����DoJ,'[ߚt�k��E��GN���%���;�!��*�$�l�|�]ֻv��)����\]�z�m_�;X@jƵ1 N1�*v�3�2�dc�=�:�m�^��+�T��9U�$F����Ӌ�4�3��3�S��೾�>r����:��EA囋��.�y�o-��O-Mv>�y�y�����0㕰�LL@�.�^�t[�Ѱ�v��̕��:��f�X�8c\S�>P|�z*Z�+��^k���0",��n�MH\�Z/�ς(��k��
��Pfw8������>>���콧N�m�Yi/�.u�}���{'*��������WX���c�9�Mx�`z|�33��7c��=d�	�����&��gp�ۍc�=�D(�ۍ�=CBb��h|gA��\�0�s���a�$@3��"��ѵ�^���,�s��m֕��	j
̇���;��M)o�X3:z�E�K�̑�A�R�s��,%+�%L��W��\M�2�q�F��n����IM�
���r�-=�c<��tI�6z��,JԖc�p�_E�y������r+��aA�zje���A�c��;�6�e	OD��֚%
���Xg\�\�֡�j~�J�(3��T��Nr�����M	����k>r(\��2��H��~&܍�
9� �I�-j��e�TTU��cyi/��7��q�h}X� �@�jz���0ٓn{QZ�訨+R�,��;
����5�`�K?j����l�'�Y�2JgD��?�~�ԏ�S��x��A�.ѭ�!���a��G��zg�ɤ�&Ka�F�l�^vH�h\�!g��{D9Şkj�v��v�m5�5~ƭ���IF[k�!Tl.&"-������n̫G!��D�j*o��bH��Mk�;7}�;
�����݃���u2,���Zi�����y~1�/�h(*�==�
�����yC��M0����\��.>d�y�/{�B��&����	t��x1պ��x���߇Vs�^����؍I���X��˞}�1���j��t@��2�A|�v/�����*|ɦ�a%�5`nn�:�� �����A�wSi����0��� �P����l��[��K~����@���{�+���22̃�^�Ճ�\�D/jY�[L����-�������]m�5 p{�j�s7�~��7�4(_�]at�Ƞ2��[R��=��I6��=�<�r�u�U�s�v��Ҽ�͵!��e�"�����[BBBO-[�OʗrK�����2���j��E���D�\L%����j�hO3��"�3ln^�:΄H���q��<4}�a�6�����1�|��_WYo�Zo��]�RWW7G�5K;G�Z �N��V!2�ˠ�y/�p��
o�²r�?mdB�\|iXx���������VUg�ދ���'$�7�kmm]��%��5�C9�b�gs�x�d1�������*e���b�6��"�|�=��}����O*��5���P�:VH)�!k�����	*�;'T�(dKttt�h=(332��)M�˰�]�����<sOC<�ٔ�VVV�{C�yZzk��Z������{�2�b@�r zw���|�/_�\A<��C���b��%!t�2Q��U1W:ayԠ�t�|���\�:��"C�4���vj���!�vC�#�92��2,޳T��Vӷ��`nT_��x>�G\�Q~R�K�b���lB� Њ�,����wmmm��_���F�r?�14V���G�r��ϖQ�:x��}}s1���k\��1��oqAk'�h�Π�^6��Z����]I(�o-�l��x�H ��U�ж'@��H+uަq���Ɯ��^���n�-�}ǀ�ϟ?��7mƙ����dv���L
oݠ��� s���8w䍛7�0Z�jc�'��ٸǱ�1���D�c���$o'J�Q��΄�[{ٯg�|#�C��8��5T�l���7U��%����c(�'�
Ӭ?������Kw��Qk�!���"(��d�����}&QoMw���^.���ii<* �
yqjl�l�[����5�[�
�߿�f��3�����S���\�HM�%�%�nU��s��3��*��HwkMV�ռ7G��g�%�	�H+''��ѐ������&r���\�7��,��U��f����
��`�C��qU͐�?��SP=B�5��ˊ ���e:Q�9*d�H��+++!����疹�#5���tm�J\�x�v���r��Jv��PI��.Q/-����P`�:2�J]��ZE朽������vN@ʣ��=���!v�����a�2쨡��[ӽ���vc��mI���*Q������s@�v�H �Pd� 3ây�@�}�����c??�BV��jo{{{X:I�*�$��j�.����팶иkx���� X��z2}��R6�b�:�X����j���{�6���1�S�b�!����E!�*|d��j��G�+�M��%�uj�W�7����7�?�K��L�9�h�qnBK:y���Ꭸ˴�/^,oB�@�T�l�<���CG|i����^w@��^��pD�W�3�Z4��� 5�F��w�6H�*�=uS�wY��;Ǿqg��`��<���]�S^^n�<�tY�}D�{�4J��=L	���H(�}x�~��Y~���۹6��d� �ׯ��c��9p����oh+Q����jÈ���rsD1 �e�[Fþδ}Z�y�e:�MI߷���n�n�3�ńb�T$U-EiX�B{�+}C�]a�1W�x�]��LB%�q�	���J��H7���Y_����R���j�݁�9���Z����d?��t<�� JIESa3%�0�$�;�'L�א�gUU�������ȉ+��ËeN�W��=~p�_��K�Y��\��V
	AxG��ϧc�������E(}�v��O�y9w�:U,�B���o,u�~/O4KYC���sI�[Ux���Hu�9�{-WHD$���Q"I�oT�:����y�A�/�3T�$wr����痗/"#y�h�=mҵ�3�$���u�v��PtD1�6<Y�4�-�=�`����T�&�b��QE�c����F�i{T��d��� <�M���B�������{�lC��d�:P�II��w��BHk���$�7#��']�����M7�.(h<(�{a�ǉQ�(�AKK��˝A!�\���U��5g��S��O\�;��L��(\��˗1/�GX�2i�<w�M��N؆�S2�҆��?�R�;2�?px�N�۲�����L�O��s���G9�:��B7�q����IpII�;́�r߶O�K胂暆�?o�r���=��-�)o�A|'U��I��rr1����B�vF�	����/CS���_�ڱ%V���]K���7>?9��.�0T���<��JJ��G�����RR����O��k��i�UZ__?x���5��'0^�Vr�[�����:s"_=����X��8����:�c�� -��l�:�-�W�|w������ '/_v��[�bO�<yZ@�q�n���D��������g�>��Ç�螆�U��ϵjf�ιWƣ����2W�ͳߡifⷀ��D��M��/&%��m����*��`���L`��<<]]��Kd�;*�����ٳGVV[��3���X���й%zM���~	��І�t��0���rg�EyDD��{�\[��� �;���dL�U�x�2�5��G��C��p�5#�`�}�qYY��Db���O/L@@��ݽ��=�A���oi��N���B�㝧g��*p���K-���U�V�@�l�sczUgl:5�i9���u}��[NRb⟷n�<��s���k��_�zu�v0V܆���}Մ��孥��G��"SS��p}��;O���<98v8����.�_�6���jhT!�l�W�^�yL=A��V򑩫�4t�O�wH�9��o|�{�ꘆ�v����/\� Y�!5�a�e���ǲ"~~~�Զ��#""ʷbOpp�� rT00�rxT���H�i���ӧO��.���^�А (VA�<r�dכO����_���p��)ٽ�Z��9�r��B��&UTT$j	��{�b��Yyp%xk�-�y����*�c;
�T���ݼu�2����KKK73���3dd܍��<!��Cx\<J��ݻw��m�-�Mk��|y��{���m�5�v��n�:������W�� 2�S��R~�	tw{��ސ�[�%� W�����*f��~����gå����2r�3+�anӽ(8?��.M��`�e��(o6�M�5\���b�}wM��>|�̤dhc~�;~�����������:�b�H+YS\~/��y�纺�6+++�{���ؾg��Ӈ��q[4W2;]��o,������˳o�y�<ƙ�U������G'��U��� {tx��q4��̕�zd�ts����2L,y�ttb��!�X@> ��\U�b�	{?����pg&m����Ɨ;�r����O��R*�-��g�^�v�D�[��} v���O3�������B�C�f#����d0
m��l�s�M��/���5>��퀪��Mũ.by��лs����˸^�{������e.���\�%-M͓ѥ2ڸB���;��rɭ7��揄�$��^"�?�'�28�?�����2\������Yh�&;�jnomn|����WXL"���{��1��-,��q�_¶��Z�hq���ˀiv`ư��1�.^#	D8Q�~��ʩ���>���Ǉ�*������N�q����O��̠�4tZ�>�1���I�}5�Bʣ�s�ū�<$7M��l�q�?�!^6�A����c�s ������S�����ZZ�'ځ3����v~4oU�����)��.++;*j�ڡJ����g�6s[�:���c�M�j���SI����F��s*�̳��옧�"�8�!2K2%!��L�L����׵����=�������t���Z�;�k]��n�[A�Oe�����W�#��4ٖ}<�7~�I��zw�q���w�9�O��f��D�~�<֚Z���Ƥ�m����z��'O�:�����y�]R�H� ��Qhd�B�f���� ��y�<��L�ůki�k���L�G��+�b��V������{��Cn;z��-��`Dq�?M[Z�#��\�,���诮��Xw�D4�V�Ѹ��K��Ɋ���P�N�a�E�
�,ɮ�ظuWW0�_�|Q"���>�N@rW�����Vc]���E���`R΍����_e��xbX�!,$����I��x����.gqS5�v�`!���8e%��11g	���G��NgEt&�w�ᮧ����K_#h�"�.�*�< ���,.�翀O}{~êQ���4�444J�{����
7!U�}�ol@-��y����t�HmБv���L����Sl�:�[���R���ï-,,.���4IVFAM�˪h�i)�T��Ԭ2�yｚ���S��Vɺ<R����OH!�|݌�L?��G�
����L�<tԱ�2��Cr\^r2�$�E�;9p�J\���'���9�c&�r	)*��'��̒�Қ�1N�{SR2��\f��?�	�v��|��+�%.	��9::B2�s���.D�s�L[j���d��nd�<�Na���J�Ǵi#��&_��"#�U��h/=�X�ىk�F�}�c��FĲ����xz
)��#��/�X��w��o���.v�j�!�I'�MM��x�$Ĉ|���9M��p\��6S5{��L�Q`1W��|
� ^����a��/=��~�̵���^Z��� �b?>C|��2���C%�N$���>[��WU%���EAӊ�d�C�N�WK�G3�@B��Q��^�����@	

�C�!!��Π��N|7j(��"�������u�Wq��7uϵ,��VP�8�ǵx�t�0��}��$v��Y�"�@��TK�}�〴Q�K�`a��֫�C�q��kk
i.'RK����%��hf=w��֯@O�T{��V�C�x�4�E+>.�����j�������!�������?���7��٩m%�p}k�rw{�\n�9~~����v�UQײ��6rr�Z&��﫫c�=��u9RV���7�;K����MăBC�����2�C�{�RT�x�(aP�������,��,��w*3���w:r{�7ϸJ��{u*�S��\Z)o�J�y^���ӎ�FNPN��\�����#Xt�3�k��8�[��r4���m� r�=R�o�撺�*�t���Q`e�K����~9�D�|��7��X��;gϜ�"~��#�U��������r�R�\��L�mNw�Lv��"�$-u����qKvVNαp��/����9���
�pc�5'�" Jxx@�CP�.��.2��s��_��s�7e��nDDY\\�kI3�3wZSx/!b�ٮdu(fu��s��j>'#c:���`v�ɾ�u/�D]����T׶IDhhJ�!�s�Ҭm�r��#�/���������@�`�G�8	�,�>�N8�u���_M�OH����J�����!�j��'���[�y{�<A#�XU~nnn���93>U֭)��6��!o�,#���'#��޾sG	AD�!��W�C�� 5�N�0��e;	�~�O�}�;ȼ��n�XU�����o�e<��\@��=E�
n�Qtt(X��e�ߓD�]�U'#�����;d�u���{����)鹀��3/�p�aU��*ݴ��>E@)�3�Ғ,v��77�@�nx���Uc��w6ϲ�ʋ��.���az�A�/�k;�#c���"ػ�)ծ�.�J�kͪ�2ǁ���K��
�n0�?.\�(��s���rb��/��ut� 0C����_�8
�)�q�MVL:���hk���Fƚ׸�iz���Eۣ��ƧT���b�>}�)8��N��$V$/����⨈����:K@�������Cy���A} k��Jʌ4������O�r���Euk�������A!]r�Yz�;a�T��p��4���XV��7n��qg�RB%ŷؼ�����"��fs)`�*p��9]>Rsi�ڝ;�Q,2���� <����j"��">��7"�В*}���3�ԛ�#���8��Z�!
���...8I×�yX546r�^����)�˃���c���qZడ\ȁ2��d�;�W{����}�w����>����3���>�R��p��$=�e@���*����k���c���έ����"��̄K��G!�C�"��wZ�de��Hq�EN�~���%��v5A�u�O��J֡?&��k�X&6�W�
K�ah�	сǿ>�_�)p��66.�#_�ݮSSS�s����U�f9����ge��1��}�kY`o�fQ�Ј�����Jn��w���`e3�����������K��u���ii��!��芧3���7k?�5�k������j|�S%(����!.����ģJ��GZ�o���ӛ2��r�J,�Q�h�x��n��1�oO��f[t��h���s����������C�%�:_�M�N �:��C� �H�C�Ƕd7Q{�2}�v���˿�ݜn�S���D���RT(>&dvG��|�^��d�R>��S$�H��d{[�B��QrIz���q���#S*�. (|��g���.�L�ӳV�-�ÇC
��A]kQ9u���y����g6�ڎ����f�S�Z��8�,	��}�8���A���P(�_GJ���9ȷ�ٖ>w������v��&��{���I�P�yg�����qj���=G��K#��ds��{{�#�$���~��a���%%�9^�ܮ0 oL`�-����|B�m�-�`aa�'�H#{/0�䆲�5s��c�7�]&���6���w�M�ORm�TN�u�'#�AB.��q�ZSS`�|����/46X��)�'5�b��{R�<$oLL��C2�j$��))�q-�ְ:��;�x�߭�2���[?~��1^B�G �*�+����{��L�5S��sv.~Sϣs Y�2��ǽ�G�ɟ�:�AP���Vw�uD�v��)ϭ���pS��Cr�F�D;^�@R�o�N7��0�Rl6E��l�+�I<ʛq0z�.��
�R��S� �F���P������v���˧�����:�����G����ȍ��_o��!��	���bb�Uτ�����b�[��wYeTw�<�w���"}nrt�\\�ZS�ݥ�&&&�'�_�6'�ƕ�_Z]!�{��4���m��c2��uyLU�xЇ��1���O������G���K�/c@���y3�  ��J��ם����C�v�߲���.8���x�e� ���0j ��3� �40s#&�fl�>=� =���ͯ�����;!�e�o�PT"�GٓL���TN�����d�����Kr�@0�X5ёu��g^ʪ�ݮ��V(���ď�VjP���F�NAC�����:�������?�ɩ$^�[����O��+��D�0V�Խ~��&��Q�߶ �x�Hyn���wJ�G���Δ�DOY!^)�011�2ۃ'�����A2�Ә��%��Z$�[ZrC��]�dk������G�~��s�y�LD���c�>�<~��2����s�~{�~����� �t�z'���C����Adz[���K�@C�.�%9�Ԭ��c#t��ñ���[�.\�pc\��X�ߗ��x���K7�1�&����K %T^��<~�,��U�BU���V�������b�����L��l�6n��9��0_H�(��(hگMM;;n� )�W�M�1A�����k�X\\���Ql�v.��<�%		�����!M��������@�
:-.����z-�~�h-�� ֙��њ���8!��0H�P�"�!�b<d��./KF/x�1�ok��r��(�v��}>�zw9��HW%k�C��@�<m�d��Bs��k����L��9J�dS�4�&q����L&Fȟ�]J��������˓k� ���EW%���n}&l�* "�\���\��hn�$
����[�� ,@8��.�v��� r�.�L �k�F���b��6�^_�|��K,[�@6E�Iu؋g<C���iM|�Șĩ�K��r�*���^:�����^8���*9V���@t�B�#ff�&�.&~�����V��xY}]������ wq�����ir��q�s5�j2;T�����V������^a�%''�wsr�-?Kh?c�D��a��E�����Y��u�2�XA�g�$�xM?D$�8�UKS�v�O�h��+H3E�@��՛7��]��o��V{��� �>�L| -�K���F��?��-�;�nU�3�m�}���ӧ3 #*g�i#�}����
t>q��Ƀ�4%��Ǫ���Ev%Q�L+e�T���`�;%t�O������X�^n��̪��A�u�j�p�
��a��	�����f!s �K����5L��Ra�,ɸ�����F�A�?ږZ��c��茗8����_fsm���636�#@����G�;f&H�������m]ݺ�n����ӫ�h���ÊC�#��<&($^����!�m uYU�(|��b�#���Z�Y���ӈb�cդcT�^���F��_��:�=<�W�N��o~ �(<`�Ī7$��Z�f��~y �J}����,�tĔ8ր���ձ��QT$���#�~�1o:�<�w��x�"^\��}Ц7�B�~��j<����$U�bJJ�Z��Z��,����&ޓ����G �c��2z����8G@O��N���~��p��z�G*
�N�f��lMu它[�D��E�X��Tw!˟2G>�y�}�pt��@_���)����~55��^��ݵ��jfi�P�{?�k�}K����-�^���=.^��0j����#��44�������������GH���n(���cP�k�*�"��6�Q�g��;���Y��g�Wz{�Z����x0��b3���5{[2��J��y�e96v��֚z+\|��-�0��ד���[q(P����=}|P˦�p�E��B�l= u�Dr��M�3D_r�{�p;�g[^������|&H���贋u� ?�;Rw�m�S�*���}��q��0�by�vý:Lg�*�sbQS]����)O�~5r���gm�=SS�g�[(&�d�[DΟn�HxGX|�M��Z�L�}iY|�p�Gѽ��-ID��*0
8��T�~�}���B��k���Jz(lY{�|�w�]A=ⷆ<���f�h���L0�-��j���״m�����;42>><-�V�3�uB�Y����b�~�-��u��\z�W&>~����!�E:S^�>������Y��H�MI�~3����/^TG��sK�f�rB���2r�G02�}����2C�niii�J��q,���7���-^��?�c�\ ��PAJo����v?���.�\5�
h_Ԡ��	v�#pg�ɞ"*��/}?�����}�����V=I��Н2��7�6��i1ҿ�B$ 6������J��rrr.l���(��W�O�L�^����@�� }�[+�<855��T�ҥ�����R]ZS�D=��|y{CEE�ͭ����A��U\�M�m$�.T�y-��$�R�1����e�
i�6?0>�~BO_?��[Aߕ6Q��|D�5X��}�/'�u��sqŪ.����t�J���E�K�T+��l�.ئ--X�t����W�����m�t��G?K츍K��U3W222�����Q�fa�=
�?�S�|[���
�1'JY����R7�|��2�Q�?aw��-����������hE�
���o��}E��G�v�����6xs�K�I�ژ�
N�f ��B�;����}�">�J?��$��K��e�-N�C+`.&n����!3��f�1� �w����W�+��۷o���1�2l�}:#++=-�xfT[��8�ޔ�Ra�ne�iV��˗�{*!������IG�j�.t�?�3d�?P���[塆��3�۷G
3ϣ-�|���.�L;�AhW�LSP�p��y�Uw�.�A+b�D�3�ϕ���D5m��<ŏ0q��;;/�l�|�J�I�wv�E�6a�
�Cp�^BBB�����ٝ���jq���F�=��_v�"��R%I��'�ߦ��C/;�Ï�GII)}v ��6��ϝ�$AQUFQ��v�#+S��a�J��#� �O�Ǐ�0!��oؖ,� �J�͒ �K�TD ӿE����C��W�au@�g
�6�~Mp[�9��#13�$q�3�ֺ������2�ω�2+�?ئ�3�5e�� �O4eX���^)4�^�#�{�H��mň���F<%j|O�xOt8ߠ����_Iʨ�<��Ĳ�p�* e�g>H����FwJ���@DO�)��l�l�-�/2;��3�g�ⶶ6��gf裧�#�s��c-��\&��/�M�p cEޫ������'Cș���6C>��Z����j��(&	�����	�Ϗcc!���3Nr�Ȃ���z��ƍ��_�:���)##�=c-TXX�'�J
��ix�`�%��Dz�\�z𭡛�9��jo��0����w�$u�,00�}�ٿ"({�+_�3�v��2a���k�C��c[�~Wy��y��+��+��=̓ 0�����%������қG!�zS�����w�?l/)Ú�R%�=~|���=h�󢢿XZ�US��G�(=У��E�+4
�6��}��J}L��R�Ф��,��ǚ�H%=yr�J��.T{�-]a���̧h���+s}&&&��==�rb�� �t�f%\ǡ�:�ɛN�tN/�=H����Tc��Ne�����J+�Rc���	UJ�ks�/�=���_IY9p����T���':r$�q��2�ܰ8�	��'������b2	�q�Jy��a#�o�uݞ���B{��������r���#�FG;�{!)(H��N+�O���+��R��JIa���B���l:z�X�����m�����w�F,&L���}��Y!������@x?seER�f�(�1P\9��(��,3�$��߽q�2`OZzo�V�Nk��=֝2�6 ��lS�6�n�cN//���].�p�\��-�x##�G����]rd�55uEsbpL*--��7��W5���� �?X�3��o�ɾ��~��Mke��t�z��ɓ'q�� 놆���܈6�k�l:6E2<����*�1��s�ˉ����{K}4��#�D3K�uJ� �pFb84%t�.��tǨ��ܮ����R�>��u���%�|]4�3(R�q���]SS���t6�Sb��pX��T�9�SrN[��wOK���N���V�h���Id��.�d,�U1%@������c���ذM{��9�� s���rzq��Z[OȬמXh���6�:�vww�>}��8B�q�84�_&��]�:.�)���u���2^���~n����R�>&%���p�Aɝڞ�*����3�kk��p�����V����:��^8��� Y'���Ж������Y٪�� ����ճ���Xe!A��v��M	6�t��iK��˗O�_R
�}@B���X��P.�����d�;�n3}Uz��Q�*"D
dk�W&�B��ܝ4��E�o��p�������_����'{��U��n��s��g϶��V �����tȜeg�!�di��耗����g��|��u[m[K��ņѳJH0`6/~�� �O+p��l��)%E �����...E}∁�����h.^�Ϫ԰�g�a�̥ha�i{J��.��C���<�j���k\y#��[4�P�p�#K-`j��{:u������������ݻӐpAh㴸m��{?'!!����P(��0v+j�@���{�0�r?^.��̑�?�\��2��P��c������o��.��W�8�t�!0���2��iϾ9��U�����J���~�;�����������HfU^�w �g����ɖ��r�z��j;�u`�2(?�n���кlXA�mi�r���W������Ե�����B�6����v_�����8� �\����Kw��_k�-}&�'�_�2�4�|��}���z�9����\���s�S��Q�� ��N;�+e��<����L�8�V�(˞�i�A�%���ʊ�i9DA�VRުv��BF��M)��_�Fp �Z�n���r,h>����.�A�i�'��������66����}J��а0�Rj��E��<��w�F4��w��뛚ď|L҄�9�a}�w��슅E�e� ����|j�����{�[G�}�r`a�oݽ��;~��D��y�����w�,jRPC�t#O����$����x ���}$������g�eh=�f'<�$�6EU`Z54d��CJ��,������]\t�(:�N���>���5ٸ�0`1�$T�� �.��%#�t�PL��e���(�TAQ�@�+��?�?�ȅ+U��9w���C������VD��������!蔧���P3�*$��5m���}���sr4��:}�a�d�Lթ^K�~ǨO"�>�ܪ���3h�?8�7����ܟ����H���t
�ԅ�eʻ�9��!� ڜzkg����T�z���]������֜�{%���`Y3�Q{�)ϭ4��8f&3��w<H�9^���Iq{��J/h�x"���0��E����lH5\�D��ڱ��t#��;h�
L�y}�b� ������m_�q�mm}�*I��*H~�@��?:⹵u��� 6;R�MLx!� ���bCs(Y8���0Cn略��Z�#�P;蠓��A�W�T�+7o��/Ŧ����ݸ�m]�v^��f� 1�
qAy���q��$)�,��6�������� ������]c K>�O�{�־�E��|ͻ�I-`S��_DUzX�1n��hd����[O��UF&�*��u{GG��oV�O�۷T`�vvQ>c��.�ƑGJË���n+@фiz�K*�����*�θr�藖���LeTd�3�K�Ŏ���.�g@�{)�k��Ж��P<\�����F����\C&��	iPfX?��cv.�gm����j����`��j!"4��ў��Y�ڞ���squ�tM��R�و���+C4�������`j�u;��=lV�{�U�8D̾���"6�4sAR��]9;�m@ǋ�2{th	mwG�U�F��g����/;�~�fX��᫝�y!!j��&G�k?+͜:���\�[�|#BTd¥i�����{���Z��CH'����J��Ul��P�+�����o �_���vZT���o���o�:���\V��"7���m���Ǻ��q�Ǎ@G��u�Է���aXd6�g�������c��|�rrs3]��j�������!�&��yx������?f?=
�[U����o�KC�}{��U��Q#CJ���UV&;�:B�� �(��<�*����"�YC��ɬfi��������a��`#�
rr����s���C�98bZN:�/�c�M������N �N�t^!��c&"bb����R�ܖ�T��������.��}xBf��	�8U�40�,2&����44�ϟ�&^?�0��{�O����'''���Q���5P�þ�&��Y��r�>��7���('�]��k�$��.bx�\���oqå>!7�[�'>���C4�DV�l]9\o#h�8� �s����?P�J֢���P�y5��d�L�E����Q�W_<p�E���DGV4��؄, <���pq�i���n%=�}d>�ǰڻ�i�Ǥ���cǐ��ʞ�Y�ٚ��K>��M{f�G�=�v�$ņd������>��m@�Ť}i�t��7XĨj� ���l�43͵4␎����7V5�h���DP��pR��ԧG��[{�GNbRy����(X+�m_,=�����`;���n�>W��}�l�T�MV$��9V#�$N���2���"5�]Ƈԣf���v�A�o�׏��[v��` @��p�e�]���<x��%�^Q�h��;;��{��A�X5��ٞ�L����g����!��Œ\���	'!�Z��l7�_]��C�Ň&�9��2���6�"������M�پzD�V�@:=
@o�CMf��򻺎N0����������v
�<���u�j1��;������>��T���&�8V|1��]�O����j�^[�a�����û��5�}�rW��~���ԀF$���<bg�a��ǭK999l�)���'�Ͽl��E�����~Z4�	OuMC��k�� ���(Pi/^\���vNJ���Ö�O��HKC����*6�s�^�K8Jd
<��� J�#x���Q,+� ���8��(�rr�����gzH�T�!C���!�fq4�l"?6�X���}7\�1�,A�|���~j�>�����Nh�����Y��͏!��k�J&xV�q��ddd M`��Lk<�y<�W`�RH}�?y�0�����h�h֠o�@Q�/�2�%g�su��S��A��T�fF�vs�n���]C�-Eņ�7TT��1q�����!�3[���a�H�/�ӝ˄�ZE|�������BFmzlճ�W�3K���ݞmx>�`e%οU�/��89�[q�0��A���x. �:��P9�;���tK��%=�D���i]�F�ւ��l�>�l�D�N���bN^l�>���ta�@v���́+^^bؐ� ?諴o��D����j����׸u���d�?��kv�V8�^���m���ڊ55\ı��� B֥ѯ��E���Vf{��������~ܲ@���;�`T���>h�@ DB�*[KvW��<��
�A��q�g���˿�7�؊��Lw�@ei��>Id�
�;��7~ ���8��U�)�3gp��вpp�0�K��-��������GL¦L���uָk�����,����2@�N��^P��:�j�;�r���<	Bsa8�����v����G�99Z)�r᧛%s�w�6�������JX����������}�V ���ǿ|�J^<�lz��B�uuW��ݔ��-�>�tmR��q{��J-�ap�96�8����\�<,�����7��6�'l�Fir�����ml���w*j��X��>��zU�J��1+5�0�D��7�=��us;�yDn>	n��x��c��ZX�9��rW���)b�
��`�aN�CN�͛7�-,-3)q8�t�D��n>>�ć렐�<,7틚ַf�����tb.K�Aτ�Ʀ����ek������ 2���Bќ��߾�DS��'�g��9�U<~V�Z����|1�ɓ�32.��OR�P 4�������ҙ�����D1��H���L��D�8p����;����{�~�dBB��}���A"�UkG����dtߤ�)M.�L�}p�`QҪh�x	L���X�xdtT�Z]�m���(;'g 8��rm�/���'�4����O"&�$�u��icS�=F.0b�)�������Ĳ�)���.'�Ȇé�fr�����C��������� �PTtN��:��D/d����u�����A���P�8��o��/������ ��ϳQ���b��F��l�����N/�򱥎�hآ��፭-˶4�f��N}4�P���l��+�R��/��W@�cm>�켼O��&H��O�bd$���e��㸸���&���I�s����~4����K�����/�f=6�=��]}�*�B�Q
r��فr���Tn�� �N��8�6::��f���"1��oP�q۽�`8���3���x�;��h�wI֩eD���J߻�X)_T%�tSL�q�	F���c�*,����*(�<���s�L���]��8'H���1�X�a������L���,�Ĥj�ꋬK�7˽�_�CN�FT��Q�uOgj�����O�$�hY������.A�+l?��]Az���pjeU���z�uS�����\����`UME#֢���\O22rd��SW�~�O�=D�ಱ�d�U穮Le+f����-us;@ �D&�0�����$Q�i�pltP4��F�Il�ˮ�&a���׎�>6���]hdp����2�vs���(���]�"�uO�{��!���#��x�.�`jjz��Ŋ�K�`۰,&����ozB��Po�i��s;} ��P��d��K�M�U�h��d�188�H�;�8}��#��Fm`����Q��u������H��^_�t �.�o��?�|�
�o}�TG8�W'��B�Ԇ�jet��\�G�AA�jf��kf�9��1h�}��hc���b#�%Z2,��1�x�(<<H>=��#xQF7 �v���s��;��s���N�w��4D�����n&�#ȒS
��ܾ�A��,v����?��U��%<T����z��&=�I�zc9��<y��/:9y�b�sLs����[Ef�M&��oܸ�K���d����w�;���#	�������������Kd��?�O���zL8Nw�<�Ӗ�B���&��l�aS2�&:_Ǟb�o��������yv����Ԕ�$����2[���У���5#'�"��Ngkss�gb�P(��^�JL�Td0�e����kT�o�@�g����H���⨉�8{c^�W�D������Q�h�m�'сU�����ch ��� k�`1��P���4)JM\��˹-��mY� N�&�E��33X���;��n�����" �F,�\�����s�턇����s�{t��#���i��lZ�@��%Z�i��{I�?�IRX��9>�e�[
C}�F��҈���H5%��6��\��c�A�.`a�O�Ǜڴ�Eu����f������	���7ɰ�OY����aU�Jl����j��H�lуX�Eb�����x �w�t��f\�-��7��N��A{t�[k�M�{�zu)�����cǃ����`��]��/xo#uOm7�}�*|��m-��E9"flg���4O;�.���"�G����E�Xh .���=:�|��u�1��D��`���,,�g���{���C��||M!�2\�P���b��X�K��؝��;�� #8�\�G/%�\���	H����9$Ǐ7`Ho�}��)ϭH[�Ǘ�:����㓔d���¡v3��Q��y�����r��4��=F�1ױ����N"�����y�5t��2��v9eࡵJA��h�;͢�����w{=�f ؕ���!Pa�? g�0�^��.��* @9�B�]��|��M���P8�[)E�2FK���w����tބ5ޡ��ͳ��osH]#�G/ƨ����;��k��5���TR���i��F9��'�8!�I~�h��PS�7F�SA�hn=�����$�Ua��t��@H�# ��9�-x�������^\��r��+����r6&�:EA8ّ�lݹاsy�c�3E����U9�ݷ�Q�BCo�m����u`���Uy-����ڶ�ʉ��������	��;;	��T����Cn�_|�k�>�I� ��3�?<<AE�F|d-/�<�{�z�x�G��� ?���1����ZDw�cZ8\��h���>��>����r�E���^����x���'X�}�8�|�x���g��hͮ�w�$�Rhhh@8.^���p0��=�ξg>�$�|}D��7�T��.R%��~�&\!�E�>�#T-O�����3L�9������ң)�����nN:�td�؀C�C��3���@��mQs�o�e�la�yГ�UD��יh�p#�Z��a�82J��J�0�^X�)���<����n��@��A�L�/'�n�����R�R%\B�����p���=�Q��A����r"�~�(�
�m��GY
f�(�e'F�=5���Vɧ�χi�}��5%�\D�܏HY��|�O&�8:�x�y➲�r*k���N�|�%YL�7�+/#���ϼ�+	II�Sb/�'�!�A�-E��6U��ǽ��1[�KCIc �"LhN�����24::�����vO�[��� ܕܮsbbtH�7��^�a��t~ȱ�p��Ng�:� f=z���6���уc�_���ԑ��m+%ef��c\VW�cw]�OO*(�{�ե0�������7����	�-��x��V3��k���@��oO����˞����|v�(4l����3JW�+6���V�;l�[f��k�:V��[�K�|Z�R���V�H��*|�!y$��xT[�PC��ݸo��9�ѓ��f�Ih��5NH��/��ӣ�1�4�����bO�-}����N�����3��d8�A�+�x��-v��s5���6�����5�9Z翁GNۺ��S���J��00�s���)vd�g~�-�j��������,���i�(��g�3�����;PT��4qZ���zF|7��Co��������~�y����X��&�X	b�ۗNG^�l�LR��W{��.6s�D]9�Y�<(�IeaG2�:�#B��\B��I�X���d����x�b�ϟ?�7�r�_����܇�P�05M���@oi��ZkeJ��t�J��C���m�M[Z�Œj�"V�B|Tlo{�tQ�'���D>��)>~c��;;�����\�#Q���MѭL�L�wn�ug����@�~� .�!���7P���իW�5{O�L��m��L�>=�6�I��E|:���z����ԛ�|����*w�޽7�Z]]]��~r�㎝�:p%A�A�q

��mt'���{<]w��hX��=����{/����L��t���.&i�&��9����I]K�Ny�^3��<������s�IB'��g֪+3�<�3ѽ��B2�Z�q0.g���M62H�$�<"����꯰���=�5�#���mp��d�/߼��虄<���'ۢ�߶����kMM��tE�,�U�li��㡒*-%A7��U�/���c BsCL�OY���A��F�`z��W�2a]�rrr,jv�}e����`��)O���й��N|g
T�q0���s,J�1-�(�)O�`H��r��ʭ��T�x�tt�K�|�o�ը�pnl aK~,!π^��)
�qp��R����\i�w7��!��{�=7��i�����tT���#1
�yn�y��?w����%>;77<���2�Y�EMjU[rw}ت��`�w\��:�Y~���*@�%�z0}�v*��̄���9����H��S|�hqx׆mܕA^�si[�F��}�
ף��O�]�xȵ�tr�v�?�G��ݻߎ�t������᪰��Z;�ky,������f���<-U���]� +���69==HR� �ϥ�]���Ĉ�Ľ��/��Y���)�P�?;��{2W7��)���o����#U����'&j�q_�Λ�̖�88�@�&{=���^��^_N��}��HOO/~�a� ;//��u����5k�N����,)hm�7m$wV:��Qi=�	�7�͋\�s\Z�����UrK�tl�r��M��\B�I�%�_��\������L����ל��Xd�3�Ud���VK�"����g⟪�������♵AG���49~��s�q�����d���ۊM�J �@�D�:C��$?����m��k���Z�6P2�#��M?�Jh����b�׵u4J�]GG�r��ct4~`�أύIx�Қ�k$&�V�1��!/���/L��Q�P�I�?MSG��������g�������@���<n��^sGo���K!�/��7S�5�*)�wA�����r�D�e\@��\�#Pv�Q���2#H~��!��<��#�B/�}�����=I�	4�㽎���՗DLHS���gk��(����A��_rGż�����3 �9ھ��#,�����Ρ׍�R4�A6��;8�^��KmN���Z���A�v*>��.O�|d�@��yX�0��˭2,_M]�l��
M�=�z' �s�8�yi���r�"v�N����������ϵ9��N�G(*[U��1Ϭ��ZϤ|�_6�h��Zom��S�}D.�}ɚ�J�Ф�DK0�c��w�`:�	l|�-
��ڄ{��ђe��L>����L��Sn�o����c��cQm�7/_��%���=Ŷ]9���Su�|ܽ�O�i����$K46MMO�JrhfJ'�J
�&�L6���g���7<>$�s7HXa�~F��o���ZY��$P�S��.4���������xP�g������I�eH Rqu67>d�f�x�f�=��)�/�<�b��6�G��Sn�S���#���H	�Z�N��r�|8�+SzdHH��[�9�Y��o���� '�rrr��rrs]�`P/?�~ZN��yq�V3�]�� �M�ں�]C��쮃C����7t�NfF���d�x��`:H����&���� 9����Di��������H���m�a,(,<U|�ޮ� Q��3�xj�?�C�<p�i�U����`J��
K_���1��f�F�e29�>D#S9�q�{�k{xss3ʕ��>	�8af�l�ڥi]{uu�y��<w�#��#Lx�9Zt8";?�9����dhcc�Ղ2c�,-�3+,q?������ ���{HkC���u{R-  -�ؘ���ݯ����x��l���������3�z����?f����>�l�~��;�s�J�Q�(� �5��̓��Q	��SY̜�'�ta�{y�K� B�u���7��C`[�bc��n�RKҌ�|&��`.��x}(��e����#X�h�6'��X���܏~��Ί�ٕo�by!dt�:��@��IiN�C��5�/o�d�1zWI(�����XG��7���
_�<��@8��x��k��h�����'��[��Zi ��7��`�:!M��a�b�V�D��X��ء���f��h9����C�뭇�1Yf		�L#f;�RM�$s%���zJ}���.�Rkו��!��.�ςT��/�x3I�'JzspR��|H�d�"�z��p��|&�h�*�ȩ�0�͏���o�vX �Bl"#D�8�h��Aw7��
�I8�!��!��7
�.��?���#q��[P� F�h��ߪ9���K,[��5!��L�*���+8��TlV�_]��o�}uƢ��R��VCK�,ϧȕ�� m����fwD<��+K�a��`���ڑ�-j \��y:������r�����oP�3GA����/�
K�`�Z)��eP��0��w�#n�Ps��s����U�`�3�ٷ`!N
		-��!�������7��95�m^B=Gv'.���<x�нcn�����,��,�M6�鉵
�����	̀X�0��������;�@�g�-�>����L���n@���_�5;.M�U@�|��(�xr=��;�!� JɾK_�s�:p��ę
���#Qfn�Ga@j\���L��k!041�ބ{��Q`�K0���W��跆<�#E\�n�M�GG�O8B?2�����go�[���i���Z�d$JS���t=�#�e1(^HA$�P���D�X|��d�Y0�<���V&ˇ����c�ݦ:����>�R�����Ny�	

Hc����A����~�L�w����	�g��N0�B�'���"�{0����B�kss�*�������tR��? ���T#uu��� 䔹�=m�O��S�P"�L�&srqo/�F���e�\@Gi�]�P*��'{+\�++���I�>tT���)���.-�����k�3^���=s��F>\�"���M�c��Q�C�ث���Gw��Z��]�6�f�%\W4��'
��UN�����#�o'9=h]z��v5��(�J�iHV(�H��C�����@b���>9 �ʼl��sUP��S��)M.��7�*�i��P���u��?"��Lq#�=�E�P�:U�͵i�&�E[e�Z�F��t�;�l�0?U��挍�=q4�S���xB/d���7�c��z�ǵ�ve��(aT�g�"1;󻄴����u�e֐��z��k5�%����?_+?0aZ���9a�P�[�F�d�\ ��zk��S]�z��^ο�� ��D��?8�d��o����qmڸ	JW/ϤZ�#"��0�Oo�v�i���
�Ё,�����aK0 �31�-W�fm��<I��N����F�+�Q�aq:��[e�[nþ���j�id�c������Ca\C��a��{s/���P�:7sdQ�7B}������\�D��^%
͌��u���E���[*�S��|��7����c(ZL�h��ԋk� ������4޻E�czA I�,�|y�)�IE�/N�Q�uAAh�&��Z�D�-�'��=��ϼ�:��;�z̕v����]Y5v����%iEXE6��W�թ.�q��777�^YZ��\S�cl)��:�_�[���л�m��9��	��{��!�5�P����=���'J��/�o/}F�J�x�b��ƭ[֩~���Ȅb�T�~�[��V������B�H���'��J^bk�����V�S���E����hKb��a�<��"�N��3
-&	�4%1�`��.��V��x1�[��)�]���"����4��s[�ң�ED P*��8!�I�Rme(B��)A�&B��ZQ0PED�R����<�� �	���C�{���u�?��s��Y����w���ϳ�/�o]��l�
o��k��3m�7���lu�P�d�V�0=���Κى��A�}��-ݟ>}�0?���-_c�8@�Mؑ�w�:��/�*�h����S��G���fl�@� y���{���� �I��1e��߄|Wo4ձ8H.k�_<�V,���t�[a}e~���` ॎ�m��IyO�`?/���Uf��/PY�6�P�`R<�z�|�O����1�m]Q�?�������xu%��
 |�E�݀��*[W���α$����L�hNTA\����e�~��Tu2����M���GW�aVth["9��*t��g��+��[+�_�^��r�t���M�ni�<��)�zL?��D�[���25f��
Ô�6�)��&�n�`srh�h�{e��TDh�UUp��c�Id��=�+���.]�����,'�vr�f?i�{���ASk ����~��0���q0� R�M��o'$�� Vb����w
E�,��y�C�WQQQ�B�Q�l	���_�Aj��E�����Tq[f$J��?�G/��Ta�RP��(M�CW��A��5��� �v�o4n�l�&� "RM˒��w���m������%�F�0cPRv��0�m�����$쿕\�j?SN��4T5�+M>K3]C�UD'��эM�W��%$���� ��ڂ Ѯ�+�Mǚ�=�D�G�jjrj�F3���	։x�`��&X�}������8|ŭ?~����ו�8��P2�ܾcG�y�l�֌?u���ґU'�@�a5BVh��b
�1��/�wf���ڷ���p�p@�p�6�OБ�%�G�?Yylyr��я�O/�}'����D�ʾ�=�:��_�l�ʮ-�eT� w���ԩk˔w�����tC2v{��2��A��3�[�ђL&g6���pT0X��Y�ku�{��?w
���#,~qt��&��a�i��I�tU��S9�Z� �4}�[�|d:	"���o0���o��@��2&yxO~y ��.��	�7��1 Bב�o���΅�~��ڊ���_�:u�yh��(�D˚l�B�4�	�Rz�����f���V��̞(Wq+��.vhhW����8˸��98��sU��W� h���ʠl�C�9B�W$�e�x���"��=2�f�p�����Z���������n1)O�OMj	�2'����_��d?g8��C��P��������z���,X�3s�v���8�LⰄ���yF�m��=z�3!1�Hw#���WW׹ш�s�mY��]�b�����pl�A�~N��QBy�cN�'R��r�Y�6?Y��iyۺ�N4�TZ}<����Ic�[��������qYYz�3�B!9��`�[��ĸM腝��U��A�m޼Yǣ-���[��ѩ����/"�y�(ګ�.5���m�@b2��`��Yla�c�AQ�����=��Ev�@Sε�����*+�⧻�̘���G�̻��+`����2�����h��+�ϔ�5x�2Y a��%�Q�F�]*0F��HJ�C���F-*L�� �[�/�2�5��r�G[4i1�|��؎νEZ���Q��|�m�/��}!J���*cJ���3� C��OL ���}��i�:��-S�!f��x5i@��y�C�Po~G���i� ����ӝ��oG^��o�lt�t�ҖA����uV�>)v�����ĸ{$�KLjԛ���XD����ڝ�7��{U/N��rM�
!�ͬ3�%p��^V��21 �{����4D&G���ZvJ��3����/�S���c����]���qw��$��ny��@/��O(ݺuK쏏o<Gc�V��W�������������Un@��.h�y��LK�i�?�jꠛ��V|]��e3mS�wO����W@�''�b	uX�`��dH!čS�&���>7�q�R��υ��;ؽ��G����e��Q�=��cH�AX���k=F�K��=���=ML��� "f��$�ब��=��|.	ĭ��eq���zs�������҈��hn.�?*c|�QS+o��QBB9��"��ؠ�H�[��cϬ� �T ��W�6S֧��C�����)+6�k����4��Hq��& �J����H:[(!]��}c\�x#�1��븷����,���8���@�Ӱ��W�YBMʵ��ʁf,�p��]��q�2w��[ϒ����2��
"^1�.�I��y�����Wů���2q3�t��Z���Oջ;O�b���o�@�ah�՛�P�X#�	|�\i�ޟ��ȗC��#����%TU�as!ͤ���A�p,�+5U�aRR��<73F�y�ѳ�p���+��K���ݱh��L����* H���.�U3�c%�&=���4/eu�ͫ�V�U�|ŭ!	��y����������Jw9�����(���P�!9��_�}X��<\Kl��rA����(��!f� n�)m�l8�p�3q��?���U%h.�MO�6W���΃1*���'�@3M�"F�&]SSS|Z��3{ �c-��r��͹�$kUj嘿I;iut%��wF�?���B�o��2�Z�d�a%�g������/����\39����0wУ��a�P�.�ӻ�;��k�0���x���5l��o8$֩ѵp���zL�5�l�P:��:}�ޫ������{%1���ݝ	x�",�i�5��bB7��и;d�����/�f���� �-��U��J"�b����3E�U��bu
=��r�y����.eQAm�)�����+� Sm��2z�Y1Ll�Eq�{S������n��eo)o�n���d���t�X*����9�:8n�c�}�+*^A�=��o#^ʲAl[䔈q�jQ�X[�(�{F�u-� ���^E_�[�L�����ِ� }u�ņ�=�C�H-
I���wE��R�}4����;[�|F��N�]Yi��^�7������T���y�I4�&��s!���`1�)U�UE�y����� ��Ws񓥹��π��^a,�� Gk'	��) yÁ{s�`;���%��5�N���ɥ:^⹏�ؙ�qj��	#-� �m$�Es�"<���޳-��s9�V��]���*չ�&Nʒ�w�d���`#|�l��>=�Ν)l�
;��u�j+팀�3O�ǟ;�p��^���C�L ��U����4p�S�PU�h	]:��[�s�3��f����UU`�-fO�y��y�\Q��h���7�.��	0�/ыr�N�/�/�h�WÝ�l���,^���L��0��_5O�,el9M�u���4I�5w>I�������}��+D�J?2ᬒX��1Q��Q#<Y� �,}�6 ��C��E̥N���Vh��Ն+͍�i�M/�|eq��rՑ�}|Žŏ,cY��B�w,������|EVM��f�H}z4}��Ͷ�I�G:j����.��a�[N��&�����p����$ܫ	���K�t�9�(�Ǉۍ鿯��\[1��5�%+noF��B h׊��KQD����U)���r(��#���Ց,/'d�#����Xm͢H<��&+[Z�	x���տ,SV����p:��vSSJ@
�|5Q���07��@�*y��@�� *�&P�o���,89������rΎ;���J'&�QyL�P e�0dL�Q-�����������З��R`�...�����`��>8��i�8!Pj#U�!0ɤCF��?@���/%`f�X��7��#,��)��&� ���͂�#F��F8J�q��=HM��O#<�5N��	.Y0�`���ȅ�e��;�^5֪e�����­��_��=�OU�>��_�޸�L���uv,���suuݾs�mu9���|���^�͊��{"���R���A���"T���ښ�*�ǘb&$�%��]�]�ֵ�Z�-�?�wuq	��y;G�e8U(��ɉ��ՋeUs߆Zg�񂗌�Ļw�����v�O��>�-�����p�e������y䈃qGrh�W}^KV��С�Z�U�<
	��]��@�?�
�5��}�+�˔w����ف��VeQLX�����7��~���6#	��Y[���b���;}#YҜ�\��IƋ��9��eA�Ko>�3�9/D�/+�o�)y︓S��_$�6�t��6���������O�>=q��{bB��8�Uu&��H��nL��ن��%����o��F�^F��It���M�ô�.��g�}:�ӖK�~�/��~.�Xܶ�aχ�gϟ����B���F}�S��K����_R�y�=IhC��1�[]�6m�;�w&��Ǐ�����]���RR���G�|��C������9���^�0u�W.z��F�M�*2�Á�f�N��#*<Bt�wLɴGns�W�<�i�P{�r�&��UUUc:�Yt�/�+d����`���ݻ^JHLU��N�I^�Z����!���9��*Y�bA$C���,�j0��'~xhW�/,R�2��>���4O�1��_us�?9�
�Rgj(a�U�P���F��}�����y�F�.{\��[��������֧�s�fO4r�OX��>�k�}�5i*��T���P^C�m���j���9���@��L�2��E�뻺zS�[f�zE$Nc��z����``�������	�)B�ͣ�T(s]����}g�����l�%���Ւf��Q��`�@�O{��ΌxV�Dቐ�ĩ-W7�����xz��n���i#���l��(�9�&��S���r���������y/^�v�)�z�*K�S��ѡ�z�!ͪ+H:�5:�eZ�s��A�Q�� ���Mb�T�]���[�/�N��̻T2*�\�>N (~�`���u',X0�`�(��K�ޣ��'|�� ����-
�j���C7s��Ϗlj�z��0И8��\�i�Ml�H^$=K�R�"Q���ՙ6i�p�;���>��2�K,��ު{T����K���o��.'�"�� ��K�``�������K_$9����<��loҞ�PK   ﴣX��\�  � /   images/d9fdc4f3-0336-4129-9adf-d1b56d6d3ad1.png��Sp%���V�c�;�mt��m�Ɗm۶m�c۶:�������S5fͪ�>G}�j�+ȉ#���  DI	QE    ��@��X����`�%4�  ���w��4Hx �������{�e�x��Z2�k�o_�ؘ]%u�B<._�o��K��CV�q�o`��n ;MM���H<�����3[ps�1)����Z��f�X�N����[;�7N=7et��?�o������U�BSg��V�C��A<&�VQ�4�ny
5S�N�w�vE�(�j�[[S�a�+Q-N��X�Q�����c+�f���+X�?9w�P���
�s�ް^-�s��C�5�
���	�� ��i�n��c!8L�������R�-��w��oH�#�}�3}�Sh���pS���f�tﷀ;i�}��d�g�H�4�x%`��W�����&�D��؎��yc���T�Q_u�*��a�����@CQ��I�z�@K�Y���Ms>QYQe����K�!�˃�K�<p�d[{���K��=X�Vk���|��Z(�kԫZ����zأ�&@�����G�;�6��h���	6���}���A�SZi�۪���_X������u�n��MTI�\����;?�pQ�E!�Ӹ."�Ъir��s2*4��c�������0�y5���j�dtg�K8�Y<YNU�<Q��w�+�\73r$��}��ԛ��{�@�\�wq��/�^A1dd���H/���lg�����y�
���7���4�ʢ�V#B��
������ۆY�K��q�����m�1�a��wGy'}/U�}(Apa�@*]��B]����|,Jʴ:ny-�~~�/�4lJyT��t�~���J�
H��wVnЗ&{���0�n��wN��M��q��|��W&�Wg�������Ln��o�z�8EZW� ؃U���h�G�jk�-Rì���@H�說��k��ajs���(U�m= !����<o��]�R6d����1�G��/�k�Ξ��_+�RL�)���o����HPcv�+ܗ���n+EK�B��ڢp���{�e��ӜH3t�5�@bm�!+7�w���@��F��ظ���q�)�V��i^Zk����l���'���g�����?-����e��vx)�-�ԇ�L�����y�C�����O���ԩ���P�"��x�a!�Z��ߐئ �P��gT9K�ZZ���uj�PbjwPÐ4�Ttp��2J ��+�U7%��[����hMb��j������RS��.��d��S����
NMͮf���8���-��"R0�Z�)_!x?I�������D���GLU�Cc�k�5Sb�������$�|<��.�l�/�]� V������Mu��g f?���w'P���T�֌j��Hˑ����K�'^����$��(̞�����]��v?����}��}z�K`�F�Ճ��9@'}gr��E��ezjt�����p��e�Ixp������/�>��hZ�x��s��r���w�u�K�}i?4K�	���鋵Q|�bY`HQ2	�L�F�Q{��ޅ�W��ʜ�-@6�T@���:S1�z�v�G�K5���k�;ʘyB{�yGՏ��
 ���u�vNI�&�w���rX*�Vj�ZJ�"�z�F+0O�f ��^Yś���yS�\B�'\��T�.�:���H�21}�>6~����z�M�S>Y q�w]W�rV:tj�����7���JU�@o �T�t��Wj���	!�5����#��<o�<��TL����U\M9i��X���c��Y��ߔh �2y�Å��2-�g�OaG&����g*��2z�`7 �98ȿL�Mu�7��b�
������6��6�x�T���_�?�A���cߵ����:5�����7�a�j��/�?3�]���Y߲ܲ�&�*��c���Ŭ�B�"jv���� Ewׅ�x*���c��l�����d���+f�f,y�D�M<��=�� sx�k}3*@��չ��o�ł`u�������ml������B�6�-.�J�nY��*���~�k�aF�s���ڋ�E�@'�c�×�Z��N7�V��G���C��R����Χ*��jA��p+����ք�r��W8���k���Z�Ձ0����Y]K=�-���jR����K�@�k	b;N>���g�i�Se�7D�<8R�������n5'K���������L:��x��a7����h#�5ٰ�0�4�l`��20�^�n$/Z�{�\��3��<u��������-�8�2�"����/uM4��{:���g�%��{|= �{X��M����}8�(��B}�²�i����h�5�����m�#�أ2����kh-��]+��#��wQHv���7Ġ:SQK+
���\S�����&�C�稏a!Y$qq�t��/�%B�鶻�5��ڄ�(bI��^qԲ����)�v%�Bc0�P���W��P���Iph���< ����$�[�p�@�DďUW{�a��?h<�`� H}k�dV�{f�c����,K����@�eRn��ԑ�}Q˜�/5'Gг�q^k}(a ��鲦����B"�dh��y�Y�^�1�c�E���"��Ur�v*�_j�R�/�F�	8?����y�v��(r���IV�9�0��lk���*G5p^�s��o�G��V��:N�K�m�r�|�<��M���� ��SuW����?�~՛oe\�R��"��F���Sc�����mH�d����I�;8!|�\�����7 �R���-�Չ9:p��'�C�N�B�Я�m�1�`w�`�.��'�pQ8<�aO��"��=�(�[�e�`j{ )��ܝlc�G	n�Zo<=��[rs��@��)!Q��P{*<�������Uf���4��,�$�������7N>����GIN��l��Q�D5��g��s[
��]!�����i�����E�y�J:R�B��mG�╼d�%������vH��j@餆�A~��P�B��%�-i��SY ���ҏt�1���������K0�
�X�@�(�XxH$BH/pҲ৕'�SA�}����0 *�Z����q���?Y�'�x��J��OT"�># ՟c�bڇֽ�%�K+:#��K2��Z��%�h`���B�_�	J>�����"���4���>OAX$>�(l6�i�@Q���SWhuz� �5�hv_D<z:�n"ai���G�v�N��P�$�9�.���t�	m�ǻ9�7��c���7��Idt���,��M0wթ�"���k�έ-&�'�^0�aGg�;7�ƇP!����Bʻy���1(A�J����u�`A��t1�4`V⏦w��[�(�x.�#qp��.���bU�u�},���޷#˯G*�,�A)�W�n)
�?�`)�o������՟�%�^���f@<i5ɝ
a��`t�v����x��7�Y�6�*����E�����,����C�����5?�ځ�6S��Vۖ+6�[�������ɢ��������_Fb	��x��(�QG�7�$�m9C��zFۑ�RTÞ���T��_�d��.�w%���2�f�@_��>|�g���7��6��k'�P3����{�MэF��'�}!���p���Bu~'�D" x��fz"Ms��P����>������,͜�/0Շ����M��!ٿC�Rn�� AM�&��~N��OF�~½������<ּ��3�%�|x���u�w^7��b)+Ж�mb�[�Y���×�����ڴ�~�򫾆z��J0�D�|�+�B�a*�B�P�^��.J��C�R�b�d1�%-cP�E������
B�[�Z�����NN6p��	�ژ��O1=T��UQ�EY�t��I�t@o�N�|��J�yP�5I�\���Vl�u����	
C�=,��ͳ\�ZD�<%��t�dlobbf���\��V� �O�ܛ)�i��V=#o*��|L�9��,Y������i�TJ��h�!��� �{\a�g)����kV�c#j5����諜S:���Pӄ՚xߚr���PCx�� 6�˜A���{�r�t��j>��
�l�@iyx�����\�Jyb�*ѳ�P�4|��XL����S�G��W#+t�sm��+A�
b�=��M�����1R
T~~�Ef4���y���i�1g���X@Z���e��6MRI:K�VLi���G�v Ą:K�o1/s�8`���Kf�Y1lz3�̽O�S)D��`�8��$ |-ƪc?עZj˲�g�Wf�ZH����Añ���ޛ6�J���ГX_�ӌ���kd�/$k	��q��ïSlO)�У=���]?ݨ(��\t�K�g�h�v����&��X;^}�M�P6F-��L
H� �� �����b(h�JC���pP4.��m�f�)�V�M��k7Q��P$pi�ڋ���D%MM>c��o�G��my�����/!���.�]�R��t�E��EYƦ�%�Q"���1�:�f����D��+���\�g��
_��`����j�}N�M���6��`-����RoyU�B�,�lիԪ�%�N^���Lx���f��q�t$)$j;H Õ-��U���R�sgi�P��V�6�w����uɉ�[�!�ẹD?����/��N���<�����|,,m\$��	� ��;;�Ʌ{��T>X
����Ј���fQ�m�VF�k6 I �� y�����O�i���U�\As�����3a�]U�fc�ˌ�X�z��C*�_�;���.��s튊�Y���w`���.�`��1��}�vF���	�\)�V!��G������E�����D�r%JUh�<S���t�冕�R�k�ߗZB0�7��^mOT&�1d˖��T0�8@�+,�84_
ȕ'Έq+YM�ģ�����ԟ�z̒s�c����%����9I~&��z�2�3�?���s#1��a�s�<#���#�[�*i*���sf8Ӝ����-�EMj�zɱ��
�i�����?Wf�Rq�F�bM���`��sq�� ��{�6���z{�w'ƞ̼ v���Wxd�թ	�4�7����i$���@�h�;��N�hW�[JV�x:��X��1u��_d�rl꼚�Z/`O����$�rZl��q�&��뱗���������%���'G9sC�$�3���v������f"#R1�Lq�$����x
LO��fB;3O��2V���{h���;~4�X+U�T��MI�F�ב�*��<�FW�R���ᳳ��w��k�v���fM��|�b�nHV���u]|��9B��}�� ����f�e�1�DRB��9y�%u�+HZ&XXL6���a�%e�w�k��n���N�s�:6p��YD�|��N�hff�����Ra��O��Mf�쩫���s���`l#l̏�v?���ώ�jvq7�I��8��'.W�1�
�� nC+TS�w�|U"��6�#�-ԥB��ہ�<PПD���G_��VH�d�Epr�6�t��SAe'��F-F���)ne��G�&R,N�Q$�pjR����h�@u�1<��ʫYL��a���ͧFhr�0`�J���Q�7xڱ���.���^�rj^��*�*�lt}�Mi�Dh����8s�cF�X���c�:ҝ�4U�^s%�4B!�/�,r�{3z��"!�5�s�<�+��<E��R�Nb:�_����Q��0'�M��	�h<�� ."h�K�I�u��LE�(� Wu-bM��,c** =���!йb�mO�(�]�'�>Ǐ��\�$6�r��4�EZ�YA�O�c�S��IwkI���@��{s����*�za�b<�?�q�ԟ�o�E�/*1�A�I�9	-yގ��+l�9NB�{~����a�i,���}�ֳ1`7� �}�?�v�I_��⥡��gO��ƥ h �X�D���-�0�+�#���<�����S�F
����pʕ!&"��7�ξZ	��f�V�˂]�*˭��!p��F�c�s��Q3����33��� A-�q8՛��Q]4!�3r�&8��8Z6dmd�C�~׵(��].�&��=_W�Q�����&��J��I��r������7�\�[pF��H��}.i>�l�X�l�,��92�jI��k�z��Ţl܊W�%�V��/y��F�=l�~��Z�~��%#�SE�#4�N׆�����L�)�9��	�aΟ&���q�Cyc����;�P'=�F�;�l�*Y&%ttV-�'��sI�~�1C�rA��IR]��ޫ~�h̾b�y{5P��q����/Y���<4q~~�����$�⑏DF���eޚ�S����`�R�Q���&fS��6zl��Z��H)��m��v���OR���<��c�7!��]����$9B�t�8pA�l,�HtL	#!r��ȳz�>�5c��I��j��픱$-�9St9��Jt����l�(����a��=����1�*8�\��L�a�HeB�����y	oW�H��$/@$ �ڝ�O����XH0�*E�˝NS�r����I?!�F��9lY��<↽�HКv�j�U�ц\^MoQ�;� ����I}G8�Ikcȧ6���Qu�ǔ Q#
�[ހ)���j�KMR��v�]���3L5ұ&��)�ۥ�u%� �\��R��*:�,T�s��P2���C�d7�b$i�6�f���e{�nn@����7�JҒ��ޥx�R23%�9��G�v
�C����'��ٷ����4��0��4�T� �.�"�/�0J6�)E6�);��,�9n��3�\b��#E%d���tV'��;�8E*��羹��Os��%l�����5��'3i�M},沞9��A��(��\ٷ�B?M�����(���f��K����Dk� �F�i?R�+a��@'�\![�49.�u?��� ��]������� e�6�����
"TKF7w�
60-(�6I0�t��;��ڻWHy���~��CLLDK��7��[d�y'hj�6�㥠 @�1-������sn[���0r��@��+	~�1�ٔ�����ib�}ؾ�A��� ���j�yJ@h��|�M�e�s����{�,'�G�x�{OY���[��YB��W.O�t�+j�SńZ��a=�A;q�� ���k��cHoafnd5]J{��K���U��m/F���kR����
�/���G�;���Կ��}�G9�I�h��B�QDF���Ga,(Vv����ĴS}K�`ӊ��8�a2�E�D�';�၍؛H��>��;|�Z��H�8�E�y�&�}��{?�_���g]�ų��P@�����Z�B��ϛ�7h�,��N.թ�# ��&� ��I>�=�60(��C{\#=`U@ݡ�Z��nR$ǍD[��HG�nL�
K��Sc9>�Gɧ��EB��w��v
 D����(�Aw�s2n�P{�EKS�����A�a���q��������_uZ� ����n�lm�^�"�񮊎�
���
)�˘���3�?�I�HL7��J��ZW �$X���]��a�ޠSB#�#��f��ޟ�v��JY(5�!���{e�������,ݲ�o+���Ҡ��_k�\�o!SɑV	�7&wM<<)/�K*��2ҡD�?J'yW�Q��$]{W�������!�7%��<�L�T�(*O�>�V1���/��\����Hx.����5}F4�y0�]QFfaC��L�A_6~7�i��cQ�{�A�`�2��f=��cDoK�J���S���V������Cz�Ԭ�|���1�}hgmx�_x‘�v\_�LnD�J	Q�3C�ǎ�����Δ"S�2�*N���Ћ�LX�j8j�"gK�T���Z��jK��WK$��a#I�їt���E�~�?*Mc�wTԅU��-�͵*�=�%JAy�V��rKRZ�R)a;�O���u��4,)fs�|��[� �<:MJ�k��/`�a-٥4�_Pb�[�Jկ��Fz�r���3�<�,+�@� �ֶzj���作��[h)6[ִ�3���~w��P����e8���l,��v�m��P�4�|;{RAy)�1������de�2��,�g�6=��iO���&Y Q��+��ʈc� C`��=��6%_�W$��L����g-�yB�b��ꫮ�H�-���J�P�(
���ۊ���V�g��D�+���P�d�"�䊱���9�?*�}g��R&���&�!�L�n��b��ŝue��'-W�$�I���^�0C�O�9��4�a�N�����R��N��%�JΧ�o#�ߤ�d�A���8����$�@&{�C�h�C��|�Â�F{t(wWC�e��c��W��HJQ�t����&�k��L�04�=XD)���6��J[���x����q�hu���;i�`��$�&��Oyt����$�&H.m������)W-���#�aHD~4o�K�4�l�Nl��c�+���7������g�	U�p3,����Q��A�M�ّ��耸/$]�7(��u�KQ���s&��u�a(K	�úbj��?܀�n���\/I��&W��.�o�ЌERe��o���8�W�MpnZ�u=�n��k�	�&��<��Q�(����;�V����=������/.N.T}�3���֫̐~.]u�=sOv]��+�<����1��-�
��d�ß��ي��I�XU_{p�+���Ž�4xjvֶ`Ů�:n�?����a���ktk�=S9|�⹓��Ȥk�s���;\�8���V8��l<�#4��<�s6Q���	���*�h��JF5m���ܴ5U�m�h���;�*Wn�v�������ms�ѓ��R�\M�d�{d��������2x��1��~�����]�c#�zZ%߮�lH˛�p�,��/$u���G�`���QI{�B�"Y�/Wu�Po�9;o���A��%�B|)���~T-?��2/�I�f�*�T�) �g�V��(���V<�1�&l���z;^�M�&O�U�������P��XB�W(3���`T<e��#�K!f��W����}��n�O�{��q���Ѡ�q��Vǽ�>�xT�9S��&�n;��q�`Fc��/Ӓ�H?t�R��Z���������}}C��Ez�+ҽTW�]�B�J�1=_����!/��@�M��{I��?��ZB�&�b����N��%�C�A��i��WhT5��}}��z����'ė��1�s�f�Λ�Z*��,��l�/G��"	�t��W�ltZ-hJ�m8�\��G�y!��Y�K3A�\A}'Lw ��P^Π4R��Q���ss��������*�����ք`�5��[��:ȫ�n��Pǘ�L����'�U�O3]RIn�����t���9��Ռ�Zn��k��^b���9C
�7�����0D�5M�e��Ly�5s��G����X�K�+�	�2��Y28W���-{�(��+���I��0�_!��0���P���ej��Vh�A���{��� �Ȇ��j�S/c��+������N8���{�ό#��,��QS��^E�g.`�7� "�p\��9T�{�<~����X#s/C�^]��T�v����|ށ�̾�;��ю@nA7���O�t�xf�������������)�t!�/",�X7�=×�k ��8ђ����:D�`�*'9��.Y fU��Z��S����������v(6{�l-��ew�t�� �pz�������hO��ƓL.�O�2�)����m��f4�(n%��9D*��9�^~ �ckE��N.Q�k����n7~ı��M�.��;ü�(v@X��U�t����\!C��o%#�G���pWe�Ŕ\ ���:�$i�����8���k�T�l�c$�3c(¬ZS�I�;�ؘ����y��N\�kUeGP��:��]�C�U�[��z�\������/%
��_p�K�f�&��������S�|�I��)����*R�+�ې��Z����l�]��%�t3�'��v���o����!�Wy <J��~�>6��z:�v�۾9<�t#��#�ì�*Q���_�T����dT�'�2�*�����P���*�a���O����8ݽbB�y��+�M/W*yI��ʔN�
Rݵ�lh!��\)b�TZ���.%�|���1y;�~�lYi44���+�O�,a���h���{ձP��W11�08�����_)����K���������C�gZ���I���7�
�p��l�}��.�]j$��]�'�*x_��/Ǎئ���4�NT̆��X��F=2��_Bb-꥖~���\F��"�T�#K	
IX��0��N�c4`��_BޱJqf�
#��=�z	Jp��aH�b�_X���	�ƨ��γ.!t��h���Ŀ	�v9.��:	�R��}�������l��o"F��W���(�Ț�8��d���D%
�9KV�u3&-�I�����*Y+?�X�S^f�D�z���֓�B?��B-�[��Ф�/Xv��C7�� ^7��6-$�.����w�}.cщ=B@���O��&N�����6��	�t@~3���N0�����GB��:J�qr�A'�H�q�r��(�_�fa�|�S�0j>�)qH��d�4��K�I�ZN3�I8��0���o�}��(xV>�d4�ǗE%b�c��S�1VPI��='w{,Ioב����O��h�<L'���5_����i�*��Wj�S�j1�m��TpZ���%�eٟ�݆b���/K	�aMGC�b�v�m֜M:򟂴'/c�ǹ���{7h#�v��+��� ������i�;@Ǚ��}f'�x�T[Ы��m� ��03��r���36� �K�g����#��J��\��g�Es=3M?�M�����a�"�mm�}"�*�O��x�v{$�j��ƭ��`��K�p��T%�5���܋�#�>�>�Ձ!u��Pݳ������hwA�4�"az�2���8��Q�@ؼq�k^)���k=�Pe���`n1P�-�R�˛��:�s1����p;�[���S'^Wo�1F1ڪ�.�qh68��O&]����ɫ�a�~m�[7g����FJ�5�x]f,�����G/���a=��;E��	j�[��x�jNH�1�,��R�M�����N�,�o	��,�Y��ݘ�z$Hʿ~��mvpn���*{#�v�.�f|;��{�}�L`[<�W��f��fO�r����:�,#.��U�J*,��<� ��Kq��O����
k ������VW��3Z�Y����v�f����'f���g��ͺ��G~�?-��L���Wx�a��O���0�dT��*>oq���h25p������ߔz<I?h~#�:�i�j�+� �.�I"���P0�൴����7���]F�"�<�wTm��/I�!m�������a]����c�IO@H��cT*bת-�bi��a�Ne�@�/�"I�O2=��W�8�0�RN�| �Mv�c���Wbك�I����.?�T��]�c�� ��=^BG�ހ<�{矕�I���2�tVp*;��Ƙ��*2d�kNrTDEa���6�CH�oƞܶ��vޝ��tI�H!�ݥ+017�\&O��{��1�!2���6�}�SZZ��و>��"ŹK�'��{[n9��&�$/c��t�9'8���e)*NKYv���1��U�}0kx��#mh.��3*�[��N}��;�+�j5�g�b>2kR�oҋ��h�f���ү�&#�ɵH���C�J�Q4�\�my��',m�Wj<ϼe3��a=G�ŧ�������b�,�؊�ߓ�<�(E���Rԫ�DE�ft���V�J3�	f���)�S4^%]=&�]�� ��d	fO�4���0SǾ2�W�w-.�}Y_���Ap�H��N;��/;�q��7J�-�A���C�ۢ�G�	Lw��i+(V���9�N�`U�G���%�\$K�kL�Z�3���ܘ,�\7�U�db�6&�u���&x�('"V!��xP��p�t8�������b�۽	�י��u=���wa�}�}�ߣB�j9+��[�P���p��Uq�s����
���3BXҟ��6D�e�]�@�y�i9���Q���a��)����"�':`��T{D�s.��F��p��2���&g���W���R�)�G��]���=�D&E>�q��)��|��Qt�ֈ���B�2����h�pD�g����ɑ.���'c�LF�B�6^�C�Ϫ)~ڠYd�+��79�&�iv֞G�-,��q>����N�DK��k秵���\�t��Q�����glj�b>\�\|Ŀ��HY �x质B5|vߌݪ���|u~+͏"���%B�n���ǫ��h�����)�Z�X���۲{���!֕�5�|��uE�u�����q!�::��5-k�����R�_�<���۽`"z��	L<��笊~|����v3n���j��S�
�}aLk�Β�w��:�U��Fΰ��1w?��5�ؾ���-�-Ϡ� �}�m~��l渞�n�N���8A9����	l�q��[���L\��F�K�ix66�{��lr��x|M�J?��;:>j����j��OYe�����(�%T�,}T����M��'X�����EJ��z~��:ӛx��*�)����m�0�ºPT
�h�~{�f��9xM]�q��Ix�69��������pS�v��K(�PzN"�>��|��T�ݰ>D�&�-��h\9��:#�(3{F���t�x��P���8���<"*�;���W�Y��n���-�/�77�
��/��XdeHw-�����D���*|B���"��h����\��k���-�\���^U���k���D��$[��!�[��{�(B�sj`c�>{�rD7�U4*Y��R��ˀՓ��ʊ?�TEHPэ}����V`�y�Gq���r�&�{�p�
�z���5^�	g=��k�2��J~�S���$5�r���5~>������=p�/&���+���<dJb��ˈnM����-\��+������r�!�5��������2�mP��U_�nC�&=5oCjr8UׂW���\*s`�_dӺ��<Ӯ��g�����R#�N���igZ�5�sF�fcx��q�I���"�>S*�щ�Vr6чB֒���C���{o�5oB�4�d�/7|�ϼ���h�q7�Dg=r����;�pZh�H�c�~O�V�mw���ބ��ǽ�k����Б�l҆��as|$p%��5P�8
���j�p���y��N��}��&s�<2&J�c]J<�����Ly�B���><�}{\�RO%��y#W�J�Sk�ǐ�q��H�ŧ���f-ԇ�3%͂�ou���ƒe�HC�t:��\v���B<�X2i�Y�5*�Ty�>9�z��C{9F�J�Ѹ��Z�rA�nĥ�Q@3g.֎�XL7�����^�p�mchw\\{�o��%Am�2��������4���LΞ\�����Oe���p&1옿BlR���j�ŵ�y�EK���}��������@�a��Y%�~#����D��ǻr%!U�	àt�ć �O�I.3TI|4����e"�i��nn���J�Y0YyA�[M9~$�SR�xFL��8��L�Gv(���2I���
A%����H,I����b���� ��!�A�����1�O#��������&��;I5�<.Y!�<�E�׵����¼Ůߖ��<M�l���v�9?]g��ט˟tiМEn�GةG���ju�'�OK-���W+*��������	I�o�p��L�"����H@��}P��!�K^��H5[tHn�Ĕ�I�pYR���m�y쮏��&�B)+\�&�Vʊ#.����cA �+d�ψ�"����W6M'`����0t�+O��:��A�C.�3��� OR��D��[���d�$�x�5M�'���Ֆ�X�V'��ˠ�N�7v�����PcuS��f����Y�)��] �_~��n;�ɣ��n�?G�TJv��w{&����˗ۑ����`1�(c+���;�x�W�;ߢ���u��䬤]%Y���hN:�B�+�?�i2��J�#C0QNO���
y��<�|�k�n�j �O̥ː`S(0SAnI�����+�<7(r�a4E����$��(��|�jl�ƅ�-$|�0�x��ڞ�p�)�����~���n^]��G��j���������V������`7�*�g�~%����Wf�6:���Dy�E�appM� i���"k�E�`�xY:4c�yN�����T��-������-~���i�}3����d��t���Ҥ��f5��Z��>\����Օ4c��o�\�?TGOj�~o�ʚ2&b���A��d,�щ{I�p�s4�N�5~"Қ�q�B�zYĥW���?L�iy�p��h����B��[��/�G|�bD���FKH9JpO��M�ǡ���%�-�G��Ȓ��:�]ۑ�H�`�k�?)��qb�St�M��Xo�MA7 ��4�{���J����9�Q4�f4��J�\���P�7�s�j������!pH��Pp�#[��Vz��J)��a�>�'JZ�Bp���@'�E.S����hE#�N��4X�#�=tj���뭅�p�~Y�4�T���!�7ˊ��ɸ����ȅ�f��!Iv����j��hŉG��y�2-�eb��ӘEa����칺Q�����3�Vz�j;_�u_/4�e駠��	�9ug�DN�|X�
)��d=�_j1����3�0�'z�q�7_����`Q��?I��x�R���i����%�����0����x���$\q�%��a\�L]�"3��b�?R_�x�~#_#�,�_>=Ogh�N��N�a{���D��&�r��������Ҏ����_>Sp�R8Z���Մ<I6bw����!��-���屜�~�����$��%���^XNu��%m�cI�03{&�g{h����h9i鍺3��g��N�򂇚�3?oB�]J&���8|-����=�R���P#TժƁ����	�3"(�Ep���j%+�$�� Qݬ����y���:�Qҏ��bi�jw�9�C\�vqxȳ�!T����=t�#��tp#��}�}�6gOܧ��M��լU�R־��D��v��{�ٗ�-Es$c�ѯτ|)��*O�z���M9�e�b'"��ś�7�%O�1-��V�Ee��a!X������{]�IZ$�Ez��H��B��|�v?n�G��>z��cE���3o�hw��?������|k� ���>.j]Ł�P 
�����<5���+2Q�UbLUˇ���N��ܛZ1��XV�W�3�	ym�$ ̅��C��Ϊ6�ك6��^�w�b�J"M���������
�'��H�w�eL�B$�$�F5�2��pܶ+���N�e���ڼ���Ƀ�!xe�sσq~����C�n� �,	�3��53VU�1���0�u{��{��ګ|�/P�kx���X�QU٨�%YZL�HZc��qƔ�K����M�D-5]4�����QRw<E*��D�ɣRM�i^l��3L�,k~jkX���bo�/)�� 1;,�/l��|,�'���ŕ������.��ݳU�-��J�\CVd4��*ev����df�(���n�$����2�)��`���!gxCț�շ�%*��B�B\��f�)�uڟ����V��s���h���fR��-|��lJw0P()�-�g��}
��^#�=�z���IEGS��Td~Z���g�d���'�"H+�B$�X��]'ȷ�xKo�1|9��4��9WLHLj2��[m�y ����^Ą�QrQ[>y[T�5Q�e��o%_g_���8T��L�ޕ�L>fv��/N�Û�qV����Y��f5)� Y&�k�Z����I���f���D5��S�&�s@�"\��F�[/1�#�_#מŗQ���T�H��N�r�����|6�w���ki:.�/-us�|�:���H��2+y��Ӆ�eڣ����/?����d�sg-��W�BB��E1�̠��̗�Mr~B���a��"|^�L4F��&B���b]P�Uw��yj��Q�S����ُ@6���Bh;Jc�͕+�Ov��<nOƋ�K�2ì&�k�㛔F�˼u�3b��|��eQ/3��qP!���މ#��(��{]�HŌ�	��E9��|��/�9� ��[=��s�{���
��9������!t�iƱWv��X�IF�
�ҳv1�)� �I����� (@׿�7�����L� �Ki9ʋ����i^�`�v���1���R��yJ&�	��s[X�U��,��糓pŴ�x���6�G>��hr&�E��e�~ �:��jO��I�qMX��'�0~�Xe�� �'+��B5�T����k��4���:��i.�z���YUF4:�e���O�O2E�$)Xj��]���|&�F�Ĕ���sxqwKn��p���轙c9;�����L��n,�����R��-� Mx"��#���x���T+j3�?�)�,�Z*�q���P�}O�)��>�7�DO=�J=qx��x�E���Z�0~i��fl��ı�X�zvă�jރ�h�}�s�]��j�:p/?�e"��T&=�3|~{Е
ccC&�7ev>��=�����R�a��j/=�V�=[�������=SASFn���A�Y�Ya\���̬l1��I�<3)�Z��I�. 9,��3'��S���e�|�ڂ|EZ�U ���Ms�ـZ��9#�fB&V23!��D&��-clU]7��&�ʻq�jk�]Y6TӞ~��mbj��`k�QF(���o�c�̀4R ���`m�Ϋb�lI
�����ջ����}	�X7.����0�PzZ����/	��t4��s~��c�/����W�ۺ �۸�ʲd��Ut��X�,�P&�y ��%��!1*4�X��T=���{�CT���z����H'��^<�p�T�b�2\Y���8��� �U	���Z
cqU1�g��Qf3���M�Z�x�4��xt�@��U|L�F
(U�V��U፜a�y21hm[�|�r�Ͽ/D���P,�hx�� ���T��M��1�M�!A(]�@ ��ϥ���\��_{C�,�Ƀ\��HZM�Ѧ�O0�Pra�kM^�)���־�0�t�*7��]�I���� ��J1��MO
Ofm7���0XdY��h�'Z�/�1I�$���&��֫X ����ixO��5�\�ʥ��T[�"X%�Ѽ@5U
��d�:���.ƶ�{P]�M# ��9���T�S�$O-�Z~��P��(	�s0��ˈ���Pvn_���Hf��ԞK�ua[���ʔ�������k����L�z�M���x�廷����#�;���''�R���MI[kA-.�JV6<� �Ic�q��rm���IK{uY7�w�����@`
-�5|4�eK5>�}�_�9+�$7�xO��C�|���'o��,ɘ��0�<xJ��KSΘ��!�4��H�?e���/�4�B�T��퉷�.�&O�'��{Bi�5�c��R�2YUS���aM>Hampqdl���s���w��199�(�Ӳ�Dm=��u�������g(L���r�pW�+ٹO����g�g�� 	��nJS�3.�%�d�7�:7��+�w�<'|��; �ۋ;j�>i�!�-1&N�Sn7g��:�w�6�M����6^����e��c��Z@�RC�~�9�ZcIG�
���B����L	�G4�2P�$�R�4��e�9�����a��Z�)��V�������#9z�P^<y�R�i��B��-�,�a�c���107GC�&#��0!�|�L��R2�׉-�7F7�@
����� �K]3ޣ�#�
��Փ�$i���G$��g~�	k�k���c�Q!��Y_��݋K�!��:or��4��(;0־�uOs+���JKE78��j�>����8�Fb@rd��%)#�{ ��~<Ý-	��(&���1�:rp���J���:�IS��k�������F �4�t@H)b|?ًAy��$��Ҋd,��<��<��1K��moH6��<�5>Soa�o����ҙEگc��O%�,�*{��a:wܔ��9B��� �fY�����FVS�����S��{]i�a�B�Ғ��6���	0�����rn����A�ba-9:Z��E��Ue�V����1�<̋��U+��VAebx-M�Jy���Y��OC
엇cU�9�Q�ks�H�og�Z�JeѸ�[�5�1�TLP�ha�y�:��~�+��5��\�#�����9g���Y[�K�/��֖lnnjX��!P�&�tk3��d<�ȃ���Ǐ�g���7._��?��9�9����Hl��e��	,��X2����zF����74k��������r�O�'����<�t�6�V ��[Z���lj�'�)W�X��rc�G �g9>ܗ)���[�_�$+����39)b]x�	����i��j�Z����B�;eRt�#ۯܓ;��_*�z���B�{w�g>IV�֓8�'�jk+�ɷ�g{�މt�C��"�o��u�K��H'c=� � 5%��ZВ<I�ֿ�1��C&\9���Þl�Cn|�{�]�*���<=9T@�鴥����ܲR���ʰ!�Es��I��O��,�5!/��j��~��?{(�g�5�Ku�{s�g7�f�}-�X�K��c�����_��ի2`�9 ��d����i)h!�`�+�)բfaES�7�c�q�ek�K��
�(�j�
�"7/���{��I�8�� ��K=�g#�e�I��K���8cVr��eE���"W.�5�w�kN�[+�y,����th,}e*s��m��(����r�d	 k��m���8=|.ɓ'�O^ec��Z�Z�j�ZKߔ�d�p+�`�zW/�����m�EO˺�EK�)�d�@�;�~�`�jN츎�&Y���&�Ə�Zޣu��%Y���}.��3�kG�m������к/J|�+��٘��]-����rȁ�g�hu̖��y%#�=S���6���4���!�t+F~���ֲ���훒L��ų29x mZf!?HhiHZmj����K����diř�ח!�n��&���s�Ma�G���~ː+z���:�n�0�<2��%��6%F��<jߦ@n��-9����b�j��9����ӂ�)��!��^�v���Zc��MK*s0����'4��D�e�ӥ!�yGs�dv&��s� gm洰�t��E˸��N�i���L��^���I<���&!��J�S��YZ[����i/}KV�b)��oPZ��8F��@H�i a%"�/�h>��Sz�K#�G�]E����z���|<���lY-�`a.���O�h�'(�!c.K7z�D��C��@8ZK�^��ܵ��)��T���.*ȓ��R�z>�5/Ǧ�R�	��Ը���c	�s�ȭp�e�9�zB�e3���C�S���b;�&��̠?�� [��z���j_��������'.%��𜭥%񡏹��EJ�h"�۹���4\wҜ�h��3��9{�)���S�m5�4{Q�=+KS���;�Lh!ϻpn	�rm�@V���)��4�R����ڿ$mA
�"����|��	��O����ta�hR]�$Y1ɜY�:춖�4�Fk#W�2�q��Sf5)�6n7�����1���Z���;����A�e`�6�Ǆ�zO�>�� X/��_��֥�%b�;M�S*y=]�I��
	Z�l����T)��7��_|���e�܅���-�P��e���S����M�H,��Ȑ	-*>Z������X���Ob���������o��%��6�׵���<����X�͹����yN�H%�j�$���y���k�kҿjJC=p�����DK
h�ε��!jv�Xǚ0�ˡM���ieb��%yq|"={*�%�=�@�t���t5.�H��y_L��Ss
3+T��S v 8���PD=�ޕ��9ܓ��T��	�LJ(9��R�9�����Ji����[�l\�+���C�^��I��t���� BK��z؍�W��>�<�u�ID�T�.=	�7�R���[�2�q]�_��!�u�2�j��<������Q`��-4|�9�^�� 1��<�e�1���~8
Ȱ����X&OE����À����I�Hg��ϻ��![�ݕ��'rr�/�4H0F'��0}Ҝ��l@k���X73�޺�/^�+o�%�=�<�b�Z���0��$������{v�_���ZL��z ��y&F�X�-'�J& �9 ��
���E	6���)I�ja�C�j9�&ȓ pm����Ҝ��J���z�l�vOÆ�WT������I�xH��Ǐa�9��T�'�3��7����$X4؀����;�e��{4h��af<�"��;���SC� hVo���7nݕ�D�5`��Ԣ[��v�2��m���m�=�m5�u��%Y��x�SV�YE�W��_�Ó�Ǳ��\ۄ�( ���08S"�ag3�I��Ҳ��+��#��"�9
�=�I�\�!�s?��;"/OH��:���c�j@���4�\�o��My��0�����Ҝ��ꥤ��h U��@��8�x��A��$��p(q���z��*0��K`rk[H���I�(��k�)�U9S/����ly�7��d��@Nd�N�U���j (��(��t���wwUvvwU>�����d`��i�>�,aku��΃��Ds���鉌N�tM,��%;��dz�n�2��P�J
��X/�<���tk�V������؍��a��$ѵ\T��4��)��y|?7'ԛX�RϞaYR��I�!+�ɳ�kF=�B��4@4yduF���߮9 �2^k��<d�p^����$��s<�������Hz��
--���.�A2@�(�|�7�Ƚ[�z���Ԣ�EX��d��'C���)��F�p�>�g-��(M�>C���@(��!����9�н�� )`� h�ɨ�)�q�=��xk}B%O���]�'��jR�hX�ֳ�o��4��n׍�Ҥ3
ݬ)�	j ��Im\��	�3H�x�)P�<���M��J��	/PPa�Zk)�$4SG_U(��&A��WW��uq���!x������Y�\�ؔ���pe>�σʘ(a��Qu�{/s�h�"3WK�{זd{���B���_�J��Ne�o���Y�u]��>y�H� O�d8�U:��Pm�(5<�a�d����ܖ��[r �.ć�# W�r�z�}+0�zXfe*��`��@j%�^��jU#|�5�7 R=y"�cYØlCyn��?bNžL�"a��G�$I����=�麶��-=`G��b!D���YM��Ǐ��$0��e%Z������&��\6���M�Z�F�D��������5������%Y�uSb��ω8ӤO�~�5�B-�MȦ�THR���fz�0���r�Ϋ2��OFS-k����w`�~��1��d0^�9K�a5^.֬�����$�3����e��5�y��<==���HB���$O��1|A/��5�C�R�fp� �l\�5�&2���le�V�G�@�^�ʵMi����=ܤ[+�u��n (w�9�LRdm�~WڻX�7����w%9;F�u�RQ�L4m j�j<'�ɳ�'sL\�+X${�
{�n��\*�Jks;je$)hFW�s_Ջ�b����s��i(\&Q@�k� _"^���>���95��^�Z�����u�[j��:LHn���`�"�"�ҳLX�:<%���r�*`�)��]2�ȗ.�����Ib�����ȱ�� ��Kzf�ӧ��75�����"#��}��k�m��҆��eb1H����jؘ+3�SkB6�/��{~�~�f�V����D�4I_���&9�a+	-���r����� �#����{}�9����ɐ1�L�����?X�����	��n�z ]�d�'=��S-��@D�/ۺ!_����f͒�ו�>Sf���T�* @�fKlMV�D�-w�#lG8����Ok�C[)�"�"H@@��P
Uw�r�����N��v�$1�J2Qu�ޛy�;߷ǵׂ+�9a>`�$��}��;�e��]�?�$v 5����P�nŹ��� 5��0p�*t��L�ld�!�r6�j�|��ᆞ��d&��T��DO��?�;�X���އ�t.]���A�H�w��6��%5X`}))�S`�FZ�l�O�KAS��ȕ��t[5�O��~��u�ڄ��8x��'���������&���Uz���D~���^��?�y睷4@ɇ?�����=�����kZ��b�sx'u�'RϷ���sJPIFq���8�ht�K�	�RSK
8������| ��:�!|�oЬ��^(�P���7@0!�����;4<$?:s���N��S�֝Ő�y����u����WwvdS�z�����ڹ:�>fK�j�ox(T��@i��u5
�Rҍ[2� Uj���U{J�&M ��e���/�n b #N1(��і�했b�N��qNʵ'�1���w�*���`��.~��WI����(�S�x�=S��1�sc�!������nh�a��x���[�o��}�Rf�9�Գ�F߳ױ�r�� ���+�S�l��Sǔ�6����ד��7nޔ���u��t�����jV$�es����H�j	H�k�#��ٔ�QO��������N]�[7).6�ۗ��}M�.8���#>�Wbʯ	�����ƛ�����rW��RT6��B58u�(�;��ϒ���7g�A�Ъ�������*�ƪ.����n��DZ7���~��7���Oe:8!D�xwT:Am� =A%*]��%h��hЊ`go4�d�t5��ܾD;\]S9`%!N�+)+�Օ�q�C�Փ �TP�z!C|rR��{��4�����,�I�Ӏ;����!Tr�ΰ'rR�2)�v�$hv� x��w�P��0�`������Ap�pU���d� DLb�`��7/�R���&GW������'���1aȡ�0PM�u��ׅg!���F��tP��6�r:�r��=���l6�X�x\oQ�!'�U��^mػ���7pf����B��9��vK�',�e#$��G��9B�7$o]�l⏁G&s���7��[$�3hRK��1��<	4���Q@��.#��*^D:��o�%g�>�����8d��K��"�9H�c
:s�ʜA!�^���&�9��'E%Ǖq�u���Q��#�!��rk��M�Qx��t�@5	��Yi��y���ٸzS��&!z�+n�@���dW��9�DT�!Τ�ڽ~C�L_O��^?�rx6�&8����(\�R�v��q栆x�0"_�٧�vE
��Ɔ�4Y�"~XPn�&giY�Ja5�Mt�t�6�vį�5��oȪD�c���k��a���_������?���`�5MY�%#���ҼvU�VKV�����N�w�2(��������-�,�d0̌��r/ ־z��&ؠd0���C��r;]��kr㵛�o�=��M/:1�u�38��f�.��F�� 3���ؕ�������v����?�c��7������d8>�������?���gH9�෫��R�"����R{��?���뚨��dߖj��w*�|������9��;x'�:�,0uu�w�2�G^f�/�q l*Gg�]���m�7}���t!dqޗ�&`�(��>JCm5Wjuҗ.�K9~q(rt*�
D7'�k��!y��Hq�=h"�mU���Q�����@Ѫ��S:M�3�[@b�x?7jm�I�����?�	��i`�sMc4[<Gx~E�%�ۈnf�4����ɋY
�;;��)��ʮ�A�����V4�fl@���>+E\�4u��F��2�WI����^��Ws��������M��l���vb3E�dg�$���G��,`Ѡ���kk�V�0�$pRJ�f���-r����m<51!���ip�WC�?�I�ޚ ���L���������{��+i/5�ū�������ܼzEz㡜�li�jK�ِ�:�&5,�(�@$@���J�b�<�հ�:-�T�v����%�G�nJM�6�z�p�)�Me���QyJ�ݒ*�ȃ4p�kAe1ԛP�����2M9��y�D�Y�2�h��q���0��P/f��1��.Rg����c��c�a=���b ���'��"�9_��������)���C���ʥ�-�Ns9�7��׭I���9�ԴM������p�73��2�[����A��+�=ʪ�]r�s>A��=���}1��v+���*� �|#(l��#�В�e��5ټzUfO�J��=�H����$�,rԢ ���f�!����In�*!)�VXj]+�݅��e�U8��u@%�y  f"�K��R9�1?ԁ�N3k�t;ҾrY�~a� 8�%�T�g]"��� !'�
��x��z� <� )�0���MH��DjFP�Ï����{�����(c�c��\�?Kd�AJK����k�8i"!$AWM�!��@zR���K��F���� nIkkKB��l�@U������5���l$�h?��HVXV�ˡc��h��F��|e)S���ڮ����Υ�r����6.C�I#h3�D܃>��-�I*�̰O�����B��:��ȇ���\�����ej�8&x�K��	2�=����bY��kU՞j�����s�E�A�ԝ	ߝ�g���J�^��1

Пb�I?� .6���r+Ȕ�����X��^�3��0p3hP�ՆFݖd����xoTXCP�����c�S����1���R����1tN��$ej�����O�x�Pf�Q"���ᗅ���ƴUuz��u�R­lO�>�n���4��͇Te���L����ѿ�������NW�]ߑ���o���|p/�Š'��H}�J���<��C�s�\ڨ���t՞&����'���q��5��_�q�PF�XBfpQl��������� 'd��o�����7�p�$��i����S�[Bܼ��~WK��8��P��AML���2$���j7��R�����h�?�K2PXT�|A���A��b$�HlV�恌�����!W5��a�YO��J�G�q=�+2��yY�DQ�C���c=�_r7/��H�p�>�S�P��Yt�:Z����~�o6�(p����Qu�DG>{ș*�p��hDqR$),B ���C5[�XI�_/r��~�ȇ^%���.��z�y{�Ս�<�Q��ʀA&<�9�e34̺�M4�q#堌a�SW)CU���C�\���}�-�dQ�߬ +�N��!�&�Ζ�74x�yM&���8|P,���֪����#HXCZ3��-�0#��rI_g>�R4m��JΗ�B3��ؖ�
[�TVU��`حpJ�N)��!�<�4��F��`]��Xc5�UOX�kaԃ_�1�+�;0�^BfY$mu�5�3� ���E����!��Q�t4g��	Ϸ:#�1�7
���U�L�.Z�H`ro�&Z�����LC���;S7�.�s����He$O��F�4��;��$f��D�޸.~KE/�o磅Q��D��C)R���c�2F���Ҳ�mf?ê�W�g��8l<XAtIȈO�h��n�Fz�k@�~թH�ސ��?�|��[b��`���c�9� 
L�J�Ӗ�i*�x@��0�Um�&E���).�]_����k\��A�	nz��d�Y���-����� �2:+��^�2I�0b��X��ʊg-lrO�'��2D�N�2�2�]���,�{�飲qO�5(K��L��U�=2��>��G���	�+g孬���H��^1� ���^����l�+d�wQ��.�*�E!��
'|��<+�1e�g�ٕV{�Xf�Z�1N8���5�X���V\� �$uX�7�Z��?5\:���ø��x^�O/�]/?r�	,�g��	Űڐ��?�ĭ�ĺ�T��^ꐉ��0�y���@�Ѝ��4�a0��rԢ����5��z%�s���G��	�j�%�hP$�9G�l� )����ˆG�:"��93헥g��T�v�`��#�{�̓�-��W�Z=���mV���`��
�ZF����>-�2�邜sg�c��,e}���-�]+�53�G�/����ɷ�շ9�;4�i:��t(G��r���\Q[�q��\>z�����2����m}�9��r1�Di&s��Z�M%_< ��Oõj��B@n-R�y�K}Ibr��#�֍�e���9����/%ch�@�~/ɉ��	j����͐h�^G�@�T.��hp�O�R4gԲ���$ �@'��Є-�J�6����nv�ݷߕ�&�K����>�`��$��E	/eW�LS��m����ٌ��1P��k�e�uh�x�A$!�w��������G�FX.�,��듗��u��4�� i�����J��y�MB(艗/�Ae���x��:<�u�����:0q�H�YoN:Ee�`� ����IX �Y�������=T�ߜV�0�>�|����
;�x�̌��dA�T#S�%�]4po]�*zŇ�3�kIƌ�����U�3c�.�qz���SfAl��l]�&��j�A�8�d4O�9���Y�YK��k�)cص�� �J��B���'x�j4:?�䠦I�: ��b��l'x2�)�pO���T�v?�AXN0\5�W���J�1�+�k�o�բ0�Uf��s��%�:��/�`0�QhP����F�פ�4�*T��[E'z���u�u��с�㏜���@�b�^�P�z�͵Jݥ��,l{cC���u�>��/�w5e�!pe������'n��MO���ΪX'�:`H��g��cPulw[�zo1�I�l7G�;��gW�a>��&Fu��W�~��� �s�j�_��#��$"�'�;�~V�9γ��d �a$��~Z��X�� ��3`jalX8�L�#�ֺL�Q$���x?K�|��畐B�}!/u2��B�,Q�Hԯ�UNZ^0q���Y�v�(7H��99���g��;_�A+0�d��V�K�=��@ܹ�ʬ�0h�><
9��q�J�LX��Fx�=	��|���]�uLL��� �RG�`�3iT8N�?����{���e���Y�O��^J�
V��\�T�S}b�w��J0)�<
;�cs�]m�'�PCS{"�P�(�殫�
1{��;���/U:=��"R��ļ����cAu�.]�jC�q��-�+�N���%o-��"`n�x��oIH���`��e~~��rM'���'2���88�7��p0i�.�%��IGTB����	�gG��h�QP�`u�Ld��ѮVu�f�������v��mwd48��ɹ����_�ދ}�{��~?�^�'?��O���k������o}K>�wO>��C9�2��H#hfQ�� �)�Bm81�����@
C�#�����3u�?K�ք?��Y��MI�8G���u� 7B�7�������֜g�bj��FS���r"��B��)�;�>��7�+�1���,�\# ���Tn�r~r,��B�ƊC��٣��;���:�tI�a�P��oK��!G�+Z�x�#y�+���Ʒ��J�Rg��"9`aR
�u$���V4umS|��6����_C&85/��
�\�[��w*<]����x��:<�C��+� ��,Ո� 2W#�<���sGU�F�AVDM8�P~����ۀ�r�����F���DXm1'v�n�0�����k�(VS��`TQ�dj�z��=���K���{]$��ъ����VAf��7��荒�
9;>�����ޑ��;2x�L��1X��q�jK���/�n�\RPI��`2�y~,A�
Ŭ�)Dm��O\��7��2;���`��p��.�n\#�B�-1gX�k��4I�ƁF�ba����=2W���"�B�iƬ�l�Ӧ�aRiv�4�9w�8��5��u;�H����m��^M����+5�����W�"	�
Y=x�<��X��9�A�Y���0tI���d��XN�[��jW�Y|%
�Y-�Ti���K�'���Ku��)m���A)�׊A�U]3r����`�ʈub\~Œ �5�y��-ʅu���]����ܰ>��8��$�o��,��Z�uBd6�Sx����BEX`�]E?Ӏ���W�j��UVF���u�\R�^�u�և(^_L��7�(��=+ 'NƲ���!bT��;��RE �$'�Jb`�s�Z��)��I����_@��k�@t��v̌͠�;����L@VBaP,�	q]&�~ 2�a�rM|jɈ	�w1����r�=�nB9_@υ��-2�� N�L���q5�?�{>�{QV��e��I�����}k)�W�X&(�?B��Ri+�5#XQw��'%hJЦ�[���*�^�';���ӻA��d���'�(�E�$�Tst�5��t$n6E4AΘ8��@bJ���0Y�F�D�����5��D��|厽*��F�_ �	�h�Cv!(l���� �c9>>���#99>W��`�Ot��������ч���#v��K����	'�ג�����^$Ӟ�d��g��8��`�p����w�}������6��	"��a�Bע��A\U_#A
8G�_���S�7zg+)BȄ��"7��4W�Wi�Hzw.���);c]��A`�?�F�GB�~��t>���#2��T�m���	�E�E|v�@���ӱ��e�� b�l�0%�����F�����w���FM�IC�a����
I�,䤾e!B)_������_�G�p<G�p�O��f��Bj�u�����ltkP���3�CBn���8�j�af\���
�����M�|2A$Ū�^�
P���=
M
@=x~vJ;T�b|kq� ؄e�z�G=�X���37�`�ALT,H9Y+ ��\|%��`o�@^�vC�|�l���4�����3��ʐYzC�]&8h!%�+�V����J4�Fڷ�0�r�ό��]�29ZC���u��ܷ �Xe�$�^HĐ���cG7a�@(򝯶k47|c�C��b� }P!O��!���x=Jp�Eg�x�"l�����=K:�JD�RP�Vu�1)�`&�;�c�0�yMIa�V��]�c��	��
Тt&��L�dF'1�?�x�E��u�y	�����wT#1��J��	:�`�X,�
J�T���+���������C6�@��o��1��Mʠ�dnyi��:�u��]�K��c���Ϙ1He�;��.Ӝ�8'��U�YA� XS��d���ԅs��@U�j�� D�%�֙�`�9ȭV�ED�
A&�~`8l��X6!����&���\yBt�	-*�iB�t���:$3�js�����q����r��Ž�����R@���F��zO58µ!�I(�$뎘��X��^����a�4M&�����I^n�����.��+?���2e���ac�A�#�l�	:U��uk3���{�hͯ��Z�͝/F���R���Un��8�&�f����_"MZ���q0�8��^�7�ǩ=*��3�r:Ѓ?(�%K���1dW�����$N+�3z\�I��gsVj�@X����`��$nJ���@�O:�`���g-\s��e��T�{�Ud?'ŭ��FW p#|��н$�oUa
}�EB[�"�4HX�ә��3G�j�!���
`��Oݺ}G�z�j��_��|��������5hd2]J�i	>|��1��?����W�os�Gv̊����^OZ�XUMևC�ٜs<D�]$�U(eGL�p&�˱�c��Kq�L�E��d���
���ZE���R�$��wdN��<{���!�G�2�d4�L�(v�ҟG�s���;}
�$+q��i��ա��#φ�ڽ��ɑ��>$H�'���0�Űs�b-��le[��f�vI+z߬�5l��uY /������_���R$��B�>�X1DK���͊�dV��Vk5�l���1p�Q_.�9D�jz��d�m;�gDE�`���*1����@KIq
�xtN�-İ3����Β��RlÚF}�C�#UX;�<��?:V��a�X�� *+��峏?�;�[Uinm�9u�끠Jh�h�0NH	��-R�Ćso6��s��LG�ah�a+���/�&�96(�qd���4����D�;!R4�+�0
RX�"+�3��G�@XR:4�W�.V �J���`�?Ϣ&H���R!�9bz�|��b�R�W8��}c���6M�td��Y��X��x�TҀ�ag�4}��3c $�J�ϣL^��y�1�P`	�x�� �X%��4�g���baʧ��;�X�ա.BHLy�� �s�W���Kk��rK�l)�L���c.���Ԧ�u/�/��9���UR��(`-td���9FW��Df2Մ�C�,@PP"�r���0Ey�fn���5rx'�O�"s?�t�.��ĳ���Y ��X20��5���&hD-,�p9̫�W�H�%�e�����h�2���e]�'�(s_��oٜ:?��^dƠ���&`Q�@�=��Aa���nIl�I�tҗP��@ϚG��{
��N��`���Kȼ�����V��s*�
ׄ[J�u��u�gf�� ZN�V�6D�g	�Q�Q����y�N�ī�a�A_�*x
��Rfͮ�ŞPaU��/�c�oq6\B� �c8�����T�tW�FC��,�
�T;ۏ@���\��H�?�מ���� �(��_4S�k6M8�Q�0K�b��HP&c�+ݳ&!`X%	��9�3�����ȷ�g���V�z>�)X� �����=�Q��an�'��d:ep��M��~�~[NO��{������p0������Vt?���`���M��&!H~q�8���|Wy�8�>�?=�A�8 �K�W����)�mFB�y/�d�~�d��D���X��G�SgK��|]l��$H��.�!	ab����E���J�{{/d��ܸq]�͘g*P�
��C؛���uD���FWj����i5�d�+�>d�Z�/X��e���j��'S�/�WYwX9[����by����� �KY'���IB���CTh�?/R?O���JM�J
~�`�-��h8�� K`�:��C�m}����D
&T�[�i�c��p 3��`Π;���U��dsH������(���G@0 \�
�jȥ�-R�e����{��)��4�����
q�-@iȪ].)p8��S���? N4���F�H�=?�O��)���~ɻX��&������B\�=1�
�ť`��Ӊ46;�2�P��ɕ4xUTs�Q���M(��3��h��ʨfXJ5R�"ae� pC���Zp%��r��cȮkR��Tǲc��|P��6��*�ahC	��*��EY��с p�l�>�dN%P��zq�@Y�
�ȝ�f[6tU.T;ӥD���ՑK��v���[C�֯�<���gf��{|�Ih�5TM���A0�s�:<G;��;ps�7X_�����H���4�,!�FT���,�I�"I����ߕ��A50F�+�,�#X}W13Rǣ0�+�5񬹳"%��=�~�G�u�#|��j�0��m�ʽ�Y�s����D��6��X���v��%\oTɒ�@F �fr�,�-��ݠ�����;-�zhp5����W��YS��W�������k��e'���뱙´V	h(3ق5\�qO��u*}��D���Zt�U�=��O�Z��;?��V��Ԁ	�K�A@��h[	I���D����{�.ށ�A�����zXpv�A��_!�.w]�4+A��<oݭ������d(#��-t��j���ւK-7r���<s�����+�(%k ��\9�Kܨq�(׵]j�Є��`O��Dbv���c�s�#n�?�	�8b0��j��⁎
MI��i�������#P���ċò�6L�:�;��{��u�(�K[�3p�3X�r�k�=��I��~���o����	a��nov�_�.mɵ���|z��<�M�t�r��-����D!��w_ӯߐ�_{S����/*�e�����_�Mn>V��1��n�p���u]���uj	LT����mC����C�3���$lT����3���� 5�$_�o8��F]�À�VHn�#�{�U��Xa2�R�;�Ɛ��f���v?|�g�q�ƻo�ҙ��s`��R�%��3H]�ޒn�����2�uXhC�=���	f�v��pT��c�Ra�e̋Ĉ�f�TZD�ʳ�D�<���~C�Z�F���  @߿aE߹�C��W��*)�5x��<Mf�����'�4j��N�	8<��3�lD��S�P��@/Db&���-���9�]@F$�4��B��B�R� �P��0���M�P�d;�U�t�~���;)��V��Q�m>�.�:�K���Y`K�3�+���*AE^�I���h 	a����X�d8��3�9:u���/�]���D�xtF�r'^�Wڅ"�&u��Q��Q�oj��lm��4�X�I�؍FL�9A�5����u�0�0٬ZA[ALP�D>Ҡ��o��Ti�ʏD1�ݠ��'td���6����FBE��D�Tu�0�8Մ+�C��>����|
�)%Fu��G@�I�n��Z5�1���T:�&�̥�tq�J	����.��ܐ/�}���xND�_螤+]��@����+�#��~�9E���Pd�H��	-um�`�Q��h5]�:<|BA�j�nה�)�/�2�uSt@�c]1�&��T"(���9�ﯤdo*�)�hd)lF��$�*9���@6�IH[,&]H�.�>�]Y�akhq�Q�����WaCy�%��A�JwY���%�d�ύ�p��~3~�=K6�`��u�gz���#�j�o��«b4����"���iZ��2��`{*+����`� Q���7�����' 
�׈��W2�ù��*Q:�e&KM~&���J��!YeC��&�/V5�r��0��tY�/eި��Հ<� �I
XV�����d�C��&���يx�0V����$��C8פ`2�ٚS��P��fil��e��٪��\�8�x��W��t��v��mx4�9@��yvt ���������x6KRPX@U�B;�� ������|�ZX��֏�%��R�/�nʭ;_��n�.��.�O�e|��H���A�ԯ�W�B����mA8��`��\�<�}�^�����eR`bt Y�ַ�%���?��o\�k764)����j��R�3��w����\�|��~̢�~C��O��;���w���@||O���+�����9ÄAq4P���r4�|:�E�_a.B@�Y��5~����,���%�K�<	��0�T��Dc=��,:W���i�;�p4H�o�6��®[dz3(x���J��iC�������@^�qYZ��1&�gU1��ة��`�ԝv��9t���%������t�`�.��WV끴7�2@���<��D��d�~�kR���D�z�cn��-S�T����ȣ
�L1E����W�����O�x��<&˰q8<���ޮ�P�C4��9y��FOs<e���FE��	!oՐ� �%d�.6�
�N�#E�M�d��޹$�,;����z��xrv�|��9M� �X]*��j:"N1ht��ȵC����\y*w��Q���OK?�^�"e8�J�@�ٮ:�C�y�����6�*�Bґ�=EȠ���,4�X���M�r%!<0�s���ʄ��q���C�02�EXHT�p�`!`П~3�v4[N�N�io6�tx&��t]���􎎍J�o�cP���RV{����z���Nf����%a���B6�]FH�^J|n����(2Kqmr`C�-�۴�&��05ѕtջvZ���Τ��>K��D4��S���U�l1�Q� ��9���iԟ����$(hn�t��KMt���T��>�����W��h���(=�Pn�y��: ��ҥMy��T�L��P���������|�$�NDQ��%�����]������ý/�s��:���Ԉ+f<�R)�V��W�l�G��h�a�&=��Q���q��*��ݗ5T����N������H�sP�Yg
P���KFU/7�H�B�G�����`5�:�gSG���
Y��hB��	B����8�@���n��+�j}��	u���M=��b"��C�! ��oѬd2��	ِ�:s;��n��D���r{p.-]ߩ���8<�L�����
�Y�� ��1;��S�d���/$��K�������x+&���}9�����AW����CE�8r���w�E#���	WFϾ���oH��D�2���B�$�L�Eͺ���{��[��c�.|�4��q i Ԧ1#��]?��pW���CY���%̝�=]���.�P���|��9u�(��ޣ�p,'���t����c(%]}��h@��J�j�`�������థUmA;�Dd�����Q����Z���#9��G����:�1ˁB�^i���BB�ѯ�+ǹ]߅t��%¹��L��Ʃ?�	xTYHM����-���ߑ��y�ɑ<��H���4a9��f]���K=cSҍ"��Ӑ�(����بI�&�s�`ԛU���	�&���ho�U��x��]��j�{�wp(�|���k =8?�_��T���ؘ��D�^�*[���H��H�@.��=Xu�m��&��ٚ�F~��⼠�&��\=e`��́@W�}`8n���<t��?���X�cB�R��8��-�^Sū>��8�l�hhdU�E�"��+�_*�`�[�Ljp"#h��f��\~GZ�K���k��\�D����D�;�`Tj�V�C��(� q��b&�p�o�m]W���R`���B�B�?:�Z`��HC=�H�(v&6?A@-X��dn��j6d�����%�������a�LM�Z�P�ګ�����q�����_�x���#�g���f_�f�	8Iɍ����b�Q^rت�����x��<l� ��@�o�\� ��KzX!Q�jQ��d�ʖ?��m������aO�Cu�1ۈdsq4�W��Z�Z�����Ph]hJa��뙫Ü��l�ΠT�����kRC5T���+Aj?�ϟ�� ����jl�%�V� Y�2:���D�&ӂ�L�����X+�C�fqm����M�2XA�ݑ��%9��	��N���k"ɲ/�&j�������K����b8HtW<&]�p�IF�;Ԅ��dO6�zW�t��iCJ��h� *�ֽ�(.��XV��0"S��$�'��
��ո��C���騯�1�UC����g ��*z�H�b�P<mp&f��r��B��a��BQ�z�%#}�y�`�WL-�21|��$�=��B�h㾢2��zt;�h��zs�����r��Mb{��Z@<�s�V�)]o�f�����g^��Pi����\~��@�� DD���G�5��יnP�p-��G�Y�01汕�����k�P�Ho��Lg��ª�d������	߇�L"v����N%��Q����\�w�g��h��åֵ�}sT��l/#� \�4eH��������`,��%��ͥ<����/v�F��sp�tv8S�gI������[�վ"'㕬 u��
{��h9/S����0Hrk��$���N�V�н�z��Xf{�kR��h�G�'�ŠR�����۽\Ya���R-��yS��Z�C�䕞�@�l]zYi�
'v$�!��i��d-�~�����6[���F��CM`/^H�Bp�#�C�XW�]1�R,b7Uut�ug�g2�dh�����u ���eKYL�^T��wḩx�������٠�	�Ǜ �dp��R���g�$T��6�Է	\gʱ��������nD��I��4p�?E��۞&�`��KK�R�R��O�q��woߒ��m�iB��_������NEŚn�HW��6���e9S��Q3 ���W2#�(�"m�]�L?ߣGO�����e������\#އ��Q��cW�]�Z�ε}��}t����{ W._f��9���1��**Ѩ8ʆΚ~n�1-W`�i29µb>���V���Š�0��I�|�١��1-D��G&1��	���w�v�s3��խkRow) H~�#=��(�!) �Y�ْ��?����
ن�ᑢ{"�iv�J�������t��s�M=L����0c�Ъ&$UKF�zQ��`s��v�8DCp�
X30��9t\9ˠ	�L��L���`D7����� ��L�4��	u�]����iBR7��	�� �엿�{̬��=��?��UR�/�q�Ň�����������;G�Cc+�\T|��
.�������a�mTqf��?tmFk�����s�o�� j�W���X4<M56]$���֪�ǉ)��Ւ�ﾾkO��ֹ\�l�9_��P3��p�������;�GW��y2�H���(��˙��\�zE*���Nb
�$d��$���R���P�=��&��@�?﫱�'r>>����:W
׀j�t��r��6l���l	V�p�tE�],��&[�ڵ�-�ب˗����i %�6gr�@L��F������{F�W8l�9o�A��t œ�r�oJ+�w�T7��k���p��H�	�ْ9l$c`�T�r��y���%�ݜ���3�����}�=ߓ���j�kz1 �؃��K�?���#?��. 0ZG�
&�y��'rwkK���"���b(XSF���L��0d��$�,"nO�F剟��k�������l��u}����L��RLG�2�٣+�xbD3�����.�c����'r{�?Hu�&�S�w1��'kHՋ8 �����r�ta%�U�ёJ�8��.�5��x����P�}���>�LF����n4za肚r�C.�r	- <L��b��������)Q�!3�s��׽�����fod�c��T�����y���z�2��f��{x"G/��?%d���4/)����0|p� ����%�zP�����Gɕ��.�7:��qи��Pu����"q��e1�JX���>�|An�ߊ3A`3[i����X>�T�G��Tb���t�����K�������&���z�~��zB�	�J��$�^��G���Gb�b���vB9��D]����V�Є�ڕ����/���A���Z�XB�$.#�P@��3$��;��&))EA���y��''z.�~S�w7��2��v��+�*d��b��T��6�{D7���$H�ʆØ�
t�c]�eO�x�<}.��u_^B!�� :��[�s�*��R?�����kMrS���'��9�p�Dr���}�L�& ��^�)�����^ni [���B:KO6�]�)l��~XaQa�����SB�MZ�2R;�ҳrkC5s/F�s������e0�3=c�*�V������Q�3�X1�ve�>!�I%�s��59����fP��:��Z��` ],��D��`��1����5���X��y5]��D渃)ߑ�Vm0m�H2X���{�ql��|��Z��[�3(|i"����@��yO���P��M�ښT\�,�u ���=��(b]3ǝk�58����=\H\5�D��Tש	�s�6!ӘB}A��&��BC�����p�"L��_6e��a6��C��Z]�17�B���כdЬ	�-���D�R���H|���x�f��~�.��1�a��"�yyJ
���򰒽J
^=�����������ه}��j+8��J�p*A�XHjɖ���7���2_1asY��F$�LH|z6oN@�LC���:�/��\�ЂǢ���m�<5�5
���4�b6f�d>�������ސF����vuf�'�)�R^��d�?E�|�����M��F�i���n��mD�8j������u���QqP�Q��@���Ff�B��B�4Љ�po�]�u����H���,�3��ꀩ�\s�qr|���PY�?��N��t�X�%����}tr(Ϟ�����KW�4y$6v\��KZ�x�`��Iw_��p_n�xGz�T�+�=�����k��&�ʍpXW�;�{�A��꜎��|YhB3�DAo2�g�ߓ�����\�,ဦ��b���|���v��m.e>:��{ҽuK��}2|�pG�}��ό�Ճa�X��W͕*�	�9f��)�zj�50ѽS��1�y/�`���?>9�u9�|�	pЎA�22f�߯ �]R;.�X&�<BF��r�ⱼs�5V��|���-s������ݨ0w�"Ι$4Q.0 �3�O�q]+��^_v5!8z������j8����}`r��tך\����R<�/���r����(B�((��K�Y��f�yU�ÉGX��T��eʮ���B�2���ny����3���}��I;Y��d��2�3�s[fc��a��1�ɸ?���?�߼q��%*�jG�<�@�����J�j��H�������1��' �{.GC���&0����g����'����д��2�0q.H𝾅%64��q���ၜ�=��I��uw!(B$^�Z6�CW*����-y�rh*Ѱ�~ '~
:͜��	���L���
;���$ׯ��a���pH�c(�L��\E7{K�o��T?�O�o^��mn��зz��uH�~��F{�Ά�Z�7ew9�+,��P�mh��ɸ��N���&����������B��J9$/m�q�y(se�L��1ɭ�Z54��Cxp�"u*�z����Ie�Iz�O�Q�UZ��/��<>ٗ�޿w7���;T�NW3V�1��y5�&�ϡ+���-�a,��GgUt�-�&�9T�08?Ѐ}�kGŻ��q�T�6�ψ��<��G�%� $��MZqW��.!=<:���S��z6�2���fL�p�i�H�y5���N��T�#�S})� ��9 ��fcSZ�t��Z�9b~M}����1�H_��Ϯ�l<��X}�&'���蔣5T������w������b=��Vk�\�����IA�t�(l� tzz,g�{�5:;�y���ο����s~����9�?P����-i�ܐ�&�/4A��.[��M�[�s��߰q��D
B9�2W�
��=��p��c�k�#A������D&��Ɓ�.X�d��ў�J
^=���������o~������Û�)�p�PmB������� �=6�����у����[��wA�	�wdj)��d��]@�0������ّ�֒���1+����'�K0H1RC�i��);h�O{T|d�n�K�:?���zK���Q:�j�S�f!�gC�zl����05�F��n�"��Q�	��,���S,��_�H����ul��!y��2Հtrr�����7���q��w��5M<Z�좵;�M4`�J�h�QȪ����C5nx�`MP���[��ޗ���\��2Հ���'2�`��H�?�6,CL�X��\8� �=؎��$gǲw��|��Mi��� �>�+�u��$�io��:+X��b_�s%��v���A�j�Î���=�:�r�hW>���L�<�dp&M�uR���aWJ�&�C%\*N���L�撎{��W���=�y���NW&��ƚ,ĺ��H�Ź��	$Z�ӣ@r�$u���TI�5!� `R���h��k�;@e��,�O�S�g��6�U]�!K���\�� �Jԅ��I�<�D���7��y7I�k(5�s`j5q흟A)U������T+��$V-DkAo24�;U0~�����r��s��Z���c仠��PqN��EҘC���כ'K��>����N*�������=����=*{`A򟑡j!�,gu/��(�Q8�U��YZ&ih���3s�����>z ��)6��i
S�-��(tVdLo�DkA@F3�&`��4P��{r�����W���:�[W�eN���s|Ĭ�(�ZGF)0��{�׊�S��{�k`����g���"�}=㾾�J̚Y�B�>g� �VW��	�r�:D��hO}���5P߼�{p犄��<q�6TNaR|��<��o��&��ȁ��S�%�=�T���_|$���x�Px�dP΀�wY^6�}�i����E_�L {��>�3߽~Yn����F+�{���m�����<�3<&���+z�j�P &��um5ѭ�R9����������ٚ���ĄC�8�c�z�c�Mɹ�ÊΙ~�vE��lfk�H���`*Ώ5!�.��	��3�&9:<�E>���rG�l��gA�?פ ���������l4u�L��T��j��{x::�z����4����p��Q�قX�T;n19��3K�+龑���X�*>ķ�����r���W=2b��$��m�ޝ�P��^C�/f%�t4�E�OQ>���x�|2%��6��~&�6��-�z��4���I�&ȳ��*T�1�����_��J���+Mi�o�h�WS�]�������L0S.����H���� ��R߉ٚ�7����Y��U��v6uD�������'r���\��%�����Z��H��R�D�vȓ�w\ڹ*�M� 1�r]�wߕ�_%[PPc�M0�GS�����I	Â�,��Z���@�6��A���U='y��0߄yD��^E���5O�ǫ��_���Ň׾�������������oLƠ���83~}�*���( ÝS���8�V8+�M�@�L���]�dEe+�‏QED�<������ ���O'"#&�pU4�,��(�p�����M���5��ds�9gE�L,���Y�C�jS����&�L=u�#5�MZ�{�A��OE���'�S5��#F��?� �Sp� xͭ��)%�����f�bpz�l!�����!�ֆ�c��g��ABG6c%)!��Q�hu�ql�Ī����w�B*�\Zj�z�G2����o�QY�z�;�p(�ј�n0�������7�L���O�˕�o�Λok��h�r�N��;oHW���,_f�*�;٠2��D�V�>�t��l-uz��-jN`@�P��U��7�^��E+j����~N� �V�2����Qz�$�z��/�ʗ��]�-���堧��h����U��Xo&�9�ԭ%o�������SKMR���2�@}���D�H|O����éT ڗ�e�52����08�¶�SЊ���>�!\��e��S�������od���r��d9>�"j��@�V$l�SDu����c����$���&��5c_b=/�?���+��� ��&��f�X1`ZRo:�9����ր�{��_�ٓ����O�76��һߐ�!�Jf^�s���Q�2�4�1��#*�
+��dJV�(H��1�B�潏����=��=�V��"�5t�
��2�\��+<��Z�BDL�߱&��.��Խ��M���P�w�B,���=	к�L/1�j�2��.e��vd����?��?���}�w�c�����GN<0��&P��T*�� `E�I����aERoҗ��'���hhh�?�p��v^B�D�S�uC��7E���R�����?�g?��,�> ���^ؠ=�e`<Yf���p.�˨��R
�e � �kbt�٧����/5�v�����h�Ǆ�-�L�^URؠ� *�0�~̹
(�"����Aw���Z��g�$���ɹ&$^�	��#`i5�M�1�Ո�슄��C�_|RVVt�l֪z/�ۆ��.��ĮPV����84��|Z�)~ܔ���ڧj#�~M5)�tlաa��;�#����yA%��T�5%ݨ�ÿ��v��9��M���f��Էvt��z�l>^R��q�8���x�j����9���)T�ëUγ�3���3���c�| _~�����(�_��hˍ�d#�ʥv(u�oa���~NG��l!���ϋ�, ��rv�>���h�����5*f$q����b���>����I����z5��0̀uM'&�$P֢,v�o���Kf S��Х�����ݔ��@�{�eqJ��g#9\<���b��ڒ�4�g MMje<�s8�-�o޽+�[7%=;
��ぉ��j�1s�i,�Y��܍�a�7�t��y�:���x�kxa��=��(I_=�����m���?������ק�|�����A�ر�y�91W�\����-+�! ��V����M�!`��0A�V�$� ���� {�D�^����xg�#�p)M�Ki�?Ӏ5%c�7Uc�}�N��р:��O����nʭkWIg�X����ds���r.@���M	�u�s:��H'X�74`����s��v�v>�H_���4�25�\}Q2��gUp�GT]�L܀jba�L��r����5��n��/�����t;�46`
YA�TeЄ`Š ux�14����4<�f�nc�}��|�@f��-��Y���GᆗJ�����-rB/�T#�u<z�=�K�/_e0����&8m�h�֨�Ƚ��b�&�2���l�\��Ne��{�{��ܸ�)�;�e��׶���.�NAn�����%?U':T�=[A�X8���.�#t��Oe�����_��?�N������$ih��T큁��i�B
q���}M1��z
!��DVT�悔��"o�@�0��=-@��;�]5��rfjγ�d�����Z��D���'�Wn�8�de��cX�#Hp>bk=#:-��rr��a@�zoj����?��?���������0�M�礦���6����N6�g���R�eC����X�41��n�;��llnj� ƥ�C�3��\�;��fXs(�r�07��p:�מi����^ߋ?����e�bO*�%?��+��LJ{a����!��;����6�5�*�=�$����aK:;w(&��p������� Q��nH{��Q�K���j��2���Dοx ���}�Y��Y�u�2�	�ȝ�p~�0ر�0�k�#P���譭����L{�%����c�X��Y��jz� 􊺟�(I20��EF�b:9���|��ߕ�{�t��t �`Q��H��gH|��X��S=+PE'ֻ�t�i��O�9��=�`��;�?������!ny��S�ȁ�#Q�1�v��B��zq���z�>�o壿�9{��6
�Ҍ�Q�:��L�m��S"T�a 9f��wz!~J������.}$U)�a���l �W�+�e3<�&��o-�i �G��4�T�TfgľK@X<���c�rƧ���M�l��L��g�4v���(�{c���|��-��z�9���c)��G���3'Ƶ���lPT�gimvh{�c_�2M<Fgr��ڒ1�3�'H�|^�|C�X�M�S(��(>�);\�� {ܓ���^�O{j�沬��z$`�����|8OF�O����{F����okb����>l��j0苿�I�[�ۻ]��tM:m����B�zt(M��s���v҄.A�:�$�!Չ&��k�V�����Pj�T675A�䫭����#]�	��g�Q_V�N���֗CM�*�.QU݋��7"7Џ�^9*5qT���J���W8Nk�f����zK�U�� �G�Y�����~������pF+d���ū���������������g�����H�T?D���S��(��<�%�sv�5�I? ���,wt������pF��J�f�.�N��`�+'�����F9Q�U�J��U��e�[HѪ���Y���J\k��F]����z��;<=��&=��D.o_��֦ԋ
���怳�T�Z�:^T��}�{�ϑɼד�F\�uۢѯL�{_N�}"slۓ�XL`�C�z�V<�Z��("粏��0��j��K�r�?���5��{G�vG����hĮ޸-W�ޖV��6�ʪ|�Fu���T?g��P���Gj��b�o,Ͼ<���3��Jv:��Dnt���N��ߩ0l�u@�6�OU�Z�ٌ�[Qc�ɏH�����?�o޽+�DF��S��=@u,	rPP;"@����:�~"Ͽx&���/^�uS�w�r��ߐ̓�əhUu`��Hḅ� �kZi�0@L��I\������C����9��Sy���FK^�����!gSM�N�e��,h�k2�IgS��j�|��d�Φ2�ʸw�v{
J�V(�������nlQ!ֽA1g��	+�˚ͦ�ia��*����,�tm�é<��O�����&�uu���C�/�4���:b0��Y�		:�~�{��7C��&H��>�/~�#9����/���!�G��WSG
[�ЖJ�F��10*�U�9Ձ'z6������i�]ȝ����viS�nE��u�k7����\�MA8�A�b�y)�M=}��H�����?��<���$=8��:�V�li3;�;�ז����$��)hRT���2O��u >2�+??�ϒ�s����ޑ�ѩ�^'3�u�o���ChT�/tA\��`�ѽ���~�W�Hu�~�t����f�ABފRD�bpx����KN�(�b�!W`G4������M�V.tT���VdB�����ID�4�X�O��{���ߗ�珤8�Ku>�]F�	1���FN���mA�[�{o� �g+zq�V��W{�����?�{$?��$����׿.���s���'zϗH�<`��
W3)=7d\��>�>�'�L~��%�_�I׫HUc�*91�.�`��2@�v6(� �����P��˞�h4q�gg��HL+s�[E��zE�:W7$F�h��ؖ��ս��t��<��OJ�	�t�dW�H�Z�5 zyrr"��cڅ��%��sM�5�~r6��������."�(�9���i,�G��{�]Ty���ѢG;��������Xw��� ̨�ٟ�]]J���B�<��ǻ��)m!��uOp�����	J4���ݗl_�H����tdc6��X�UP��s�h,��K}�c�j��1��̾��E��V�bW��=9NΥ�/���h7�7e`1����]#u�n(~�MA2 60tv����K�.K���	]��E��#���z���ė�g{�O�j�r��<��^6��Y_��^}���{z����Z��[��ݰ��+NYd>��E��H�<clD��pM�}_�4i��D]��9V��X��A��/���?^%����?�����?����-(B�Z��e��b�,	�u@��A�2��tjx�a{���ȁoA�_B(�M��(fp�qc�"��$��V���\�����K�zW�|56�S�w�-5F�t,��-	�߽�K��s��8
�0���X��4`�@!�s�m5��p̶p�zb�5�x68����\k����mi��\=x(g���ٓSu�U5��K���D#V%�P���_ v
���?8+�@~~_�'Ky�w?��W�������[7w��n"�=z.5�3��;��\���ggj�G2j�erM�ׯ�P���+�~��|��?�����'�F	+�a=`�t��]�[Rl�j��		-Z�)*����n֨<e�k�My��K���o������mi_��{�'9�+K�|K�ke�U(v�@��HIMj�Z�y�=������k���q�1�gZݭ�(q���^U�5+�*��[}�}/���c��
��(� 
�_~�{��{�����P�������E{=5x��AL��1`Kdd�1*I��6p,￳���w�4�����L�d�*H�Ʀ���9�R��t��r���FT������?�=;�E��ssh\Y�b��D;�<v[ۘ��U�����H�I9��ۦ<���˅���$F@I@:��L����rGi
�E1�8[�WWy��_Qb��I��#y��'�����跎p룏P�|Y�x�J��Y�MIJ�LI�:|nY��d3�����<������'�� �"L�>�d4��Dj�Q:�cvF���9�u�ج	51�ϑ�����;�}"���q���w���(��cv� ����J�BG��I�`5�!��\�䆕������<�w��@��B����V�Xv*=S��Y ��p���﫬%gx��c&U�o�m#�ߒP���@K �?�~G��,��"TG힬ҟrZ�cץ&{����$���96���{��G������(�+z�GtpUs�H%\�(���𘺖+��@k4�ҵS�+�&EM���o~�-yX]f.�Ҭ����O�V*�x@�x
�9ń��l�ɣ������Ꞁ�
� 3�h�P�FL(QWނ�J���W��`�$���;awG��%	�
�"�'�p	��DN7U���[�����~�}��e4�W��R�Ұ/ ;c$����B���>G���h={���y���eI,��U&m��OD��Bu�u�,�F�^>�%��&b��~SE-��9�|r�%w�����=ni%�]��<�dD�X%6�C�\HT���z���1>��\V�C�*Kd���a�X���������hE�-^��k%�N00L��Q��������V�*�M
Q�&	j��	�L���7�D�+%6�a���s��c�+I��(ǲ`��v}s���"݂9k�.[	zr^%Vn�/�PV� ��Q�j@��H����|7d�Pu�@�'&4L�/�^����a*�et�,�>:FCb$!:rJr��Ap�8��"�ԡ����Iλ(>{��₺��4*��̳�����t���Jꑚéy^�1���T�hR3��(�ʺ#m@�#��iNg(
�E�d���$�@N��!:*���Y�#���p>���嚎�CS�PO����~�ը3���>�{��~8�# _H�	zr��v�|��&�ذ�W	�a[��Ď���+�{u1�~��}�^T
ƃ+a�؞�����S��
���r�&`ˋ#tJ����3l�y�dY�R:�5Y��(�v��i���gj�e�m��F�F����%���� �i6U�-3"/I�+��G0���`vm	���HJuuN��5<�aqu�
�8/vj���Dۓ�A[+K\V(F8���>��{�(�gȦ�[��:Ɂ5B���AYҡ��a�1CZLr��G��RV��!�����?�{l�ax����ѐ�t�������O$��u|(yK[^7F1�`Q�3e���<}�_}vۏ���#	S{ _�j�(I��c��k;81��qjt䧉���i�PAx�U��1~ Y��7D��A��-l=}�+�˗��D~��I-[�Α��'�%����B�[���9zP��;���x����G��ᱺ%�PHRhb�i�V�V��Q�jN�]�)����5�F�a � �q�`���~#}k�1�߼�K�])����7}=4ĳ^��ر�?�}|�^ùF�z	�m;�(7��bA�r�Z�X��UmRx<�2�Z�C_�&�����g� W���3�9������v7��̛o��[�1{�2�^�nAX���z�	Q(I�����Q��q��!v<@��&��BA@eQ 1A�(0�Q���P�_�7� 9��tl!K'��˛h��{x(k��l��lb���X��&
g���c�XC��5)�?DI����6v�ax����&v7�# �g�2��S�VEH�	��9��H�#���B*N���a�]v,5p;&�b�g�ȱ<׽�>Ek{_���0�����VP��ffn	^�dP	�>������]�1>:Bɧ�JV���ÀH'h�����:���,�(=���c;2��a�T�<�|T�l�� ���v�P��$ы�H
�|�O��JRPę��[����j�����=PM|J�����']��਼��(yF�U��ѯ��%�S�8F���/��}O@YH?	���P�
�g��?��k��wp������ί�̵k���m��Jr���X���7��g����C��A��X��`����x�vu��C�%X3T1�� �K'1��<�h�G�� :�D'{��e%Ve���T�r�eb�PF(����JI����`�)����X�D1�$�#8�I�N�5����r@���H�
%?�&����C9��v�Әx��t6ϥb�C����WQ�ɳVE��
,�h���4�?,�70jNY��ǣ}�%� �i�N�K�T����Z���O���jX&�Y��p<R3z(=��mI�\]���y:��[�}����K�Ϯc͓Ώy�p`�"[I���P��ԥ��}T=d�e�g���H�����G�p7�ԄY�T���`<�,  ΩK9�5iw�;vk�dMwJ�*�,�(�yH��Z�(��Մ�t�X��D����.�{U���y�$m͍�������2eI���ϙ*G @�98wE�X02ϙr�u�'y��Ɯ�S	)Z�[ϸ�#~�����!�䴖Zs�|��"p�|���)|�����mR��5#�l-�{#7a��1�����J�S2u�&�w�Ĥڑ�S��Q �R;u����)�&���v�����+@�UrU�������J���}	r�����PNwi<QzIQ(G��&G�`W��՜��5��H�NyO�=j�U:�$4���~,�y]����%�U��u�R ��/�4�p��>8�&H�lY�w���흗J5�l�'���E(�f#�{@��[-{[8:����_n�)�ś�PYXE,�K�:+y(AQ���#�+�g8�p���g]}����G=�r@fǉ�O4j!���{o�T����7�!V@݂�ȚC9q|�"�)�Nz}I��h��i��R�7�`uI��u��O�����`h%�:(��q��*��������۔D���;�[M�t�����zz:s�ך����X�yj1n�7�`�JT�b�:S�)�E���ɣ�*�y��+%�*��J��UT^�~��=9��#��}���d�|�$A��&��/�� 4�X����F�El:��g��9ccC`ey����>���˲:*�k� �&�/��{�K��ʡ2�~׮ܖ�hu�,�XY���=~�7��$�/�cV�v=t�L5�KLEx
���N��!������1��&��h[;����P�
Ƞ/ɸ|3������/!' ο����GXY;�zބ�Q���ͯ�$�n���CNoy�&s��N�����Qp���,R�����3xm���t$S��1��1R��Z��sjK:�^����>����W�Ώ>B��� ~���ES-n��W�bG�3�x,`�h����HעOޜi�(@��R���u��vZ�LDV��� U�϶P��V��t���@�{�Id�'���j!t��4U���tQ2�X��Է�n�y�|�d����X+��Y�ՙI0����I%"}�D�`h����.̳V��i�f�(X��ɿ��X5�!��9�v)i�}���ǻ��?�Ӓ�$��|��(ԍ��SdZ{(ɵWʇ�Qe3ʽU^9K�x�	8*���/Ey���҅Q�I5��5��H�fǛ ~l�ؙ��F��ӂF��Ũ�AE���ҬQӑӸ���&W/�P����.bIhJ���&#<;�K���@~6(��r��Pn4N�𜑢���AS�m(0����D�����!�~O�_9K����:O�Eh!b�N$��*�痑䋘��u����b�(gQVM9�������Z��4F
/��ε����ή��l�I�$���mf�E��X]]V���S�r~��M��]�}��qIo�e��uU��'��fU�6"�*�$w�b�����/�8;�5���_
�})S�=�58�*���O^���r%��cYG�IO�x_�����,o�wY+�l�q��Ց }s����(��6G�&�AbO�'<KEc��zs]����""��c��žv�xMg�N�T]���E�Ld��7R���;��O5�H�[�D?[)�-I�{F��٫���灰���?_�&@_�� ��۬��lOfP(RZ+/���V�٩aj;�a�]���&45��0�ލ��3XN������ ���~{j���zU�M�a�=I�Q^����͓��'r@8�g�`�Q�%u�ɋ7חMO�� x9d[�&"v$ȫ���
&\e�ufjxC@���*FRݽ�9�� .��.���~��l�m�s�t��X��z$)8��]��'_b�9D9	��D�ނ�Eyߡ�duc���8l]��P�Q��6�z�����zOW\^�b]��7#���?|�Gw>C�l"<9Ѷh�	?���\F�^$	�)�Z�\ᔂ1��i�q����+�%�r�%��@l��)F/w�@�����Cm�,JtӬ��Ib@��@�!��A���ŭ?�	�2��bl���<������4B� :M�X�$�2T	�ĈU$��I+[6hg�p�O%ի@�/�ߋ�ƳDe~��X���{��� ��xtהC�/� ߋ�{T!h�8߮����f�vPP`{�ӑ�0z�E͚2��G�������n�캩���؀F�+�e����X0���C�L���}ln��������qkfE�^#������1Z���;��+��B�����.��X-e�[i�Ý������SU0�J}J��/5zSU�D]P�Q�)K��BH4F�C�?F@)Y���:�zÌ��o
@|������%1���G��+�3ΰ^�,"����z�ʟ0����e��3��ϕl�g����bSbT�X����D�w/����+�9I �zeO��JW���1��ȏ��1P5�c���$Fe˘��.9��:d�>��M����]4(��Y�,�^�*`�����
��	��X���Ũ���ۮ ����t�\�@��O2�b����U�����`�NpdU@�c�|y����u���J���H�(����l3���X��G����\8:��;=��6C�����
x��{,	X�s��j�K%6��l�}��h���I7T��P�1�N�M<Q";_�I�5�;U��,�wF�"�r�5~$݂"c�BX���R�r�`�P����K��!W_�r�C_�X�����$R�2�_?���y��1Z�[�Cp��Z+!'�޵�ٌ��RM�AG�;��3	e7�R��>y�n)���5����)0!�mtx�������%ϑJ�9���#3�Q���vJss8{���x�	 y��v���Y�g����jr���R�X���8��t"��q��z�!r��r�9&,�Lyv*{&C��-�x(5Jrf���Y�����������0R�"+���X�x���#���B��׹	�}$q����n�@�F�.g��l�I�$'�o9p�
=}��2Y�& ��OWk��UJ�g���J���D��[����X�?�Xi�����֙^}V֐;w	�lA;el��<�%��Y5�,����9}�*,1	��EY��s�&�J��v^��_AR�E��ey���8E�&ey��EV����J�I���G_�&@_�Xν�A��&H���͘�j�0r͠�jק� �!�Sp�8�NAj+�08V��&��\*��`M����-o>6���X��_Y�$?��P
�FC�dH�r��&���нГ�u����I��\�Ű&��q:��1�::�\����<��'8�r/�������.�y�W.u���a�!T}`�\\R���k�P�w���g��-����{����u(v��z��*��B��ܗa����c9|����/�0;�ꨎrM��-~v��)ܑ|��q��Q	�B�����_�#p^� A{�y�y��f�I��[*N�=[��35�f��T/��%��`����.��k��@�8<:��aK���ܭ"�]���Հ].�s2�ki'�J���h�S�i$ ��JMr�M�8y9�sT3���j���w;1��H����@�`@�9Q=�2�D Ao�I#[��M���t�&�w4�	��j��؊v��xK���K����,+��b� �*�7�`I�1��D]~ר9�V�+�$�8k�?}��ÊlN��Q!��K2�Zt������	f�Z�ee�	꒠������a�������S�44hyZ��j�cz��Z^7Z�I21��ɴ*ŧ���l�
`�ǚ��nQ�u����?�C�P�����!
�6֋3�Ge��f����O5+��ù,x�X��$�Z݅�i��k{ V�K�Y�,7=�J&�\o�g��.ݥ�d���cX�D$8h=�}Oյ���,��	�����P����N�V�բr~]�Oz�.F�
�XU1F%�.kr��fM�8�M)MVc3�<�G�9W�����|,Z�MY�ݜ�7Ƭ$�|��NS hK�24����Y�����H;Xhy=��$c����Bj$+�M��0��T��a����Ĥ =V��K��9��z2�>#O���$$��Vpy��H�G�Z���x?�y���$\��K����~�QK����.����j4US�h�?�(i
~"��Q�]�6��V�'�&<hKD��Nz��dsP٘+��>Q>Y�N�F�Q5��N�J�H�*{I�A>�Jg�
�Fbѐqv�v�����	isXt/��Rp#Ӧ����W]�s�������-��\��t��t�Z�(qNLq�s�Yh {9S�w[Y��?|���d:�l�g쬫o4{}#r��v���/�T��Y,�等�g�]���K�TP�4o�ԭYcL[ή�����wՇ�ӄ�CHwfr��y4K��vys�e�bS��0ge�v�T��(��L˽"�և�*���U�1�2�Qh"��Y[Q�׻&�Iut�Ó_~����{T������7�>-79���J�S�z��o�Q�s��oeb����4�����*Wj#�W�c�ct�����1υ�5�+�M`�����gHL�����]Ϸ_�_�G�Hc'Ł���hX�1\���ʮӈ*�T�u@4�z�O�k����6����$�n�!�Z	uN\��W	@kꡦ딘L�d��&#IG�C|� %�5�D3(W��^?T}�+Ai��N��l���myYeӒnu�dy(���~��}�|.���ū7p��w��&��F|����%�c�T�Q��P\>w�pn��SX� >:�ਥ.��L�iLFtЌ51� ��c�+�B�
�؟H ��a(+*f���Cv��#�#�ɳS�������w�}[�OK�ޒAw�Du���S����]����Fu�vv��)`$�F����V��$�bl�7����).�wa��}���v�CT�>f汲r�z33U\�$k��;���o�}� ��M��P�C^�.�?�>� ��Z�s�3f�� ��}IR�����S���q� :�
P�P�{�Q
�HCU� ^�E�TTI?,�֡��W��Pൽ��QW�T��܆�\�P�k�RE����������%R8�2��2���T]}c�h�V�ZWj�*�彺�	����P+G�ΩC�O0,�=~�_��~N?w4袞IP:`a(�q�JsFǢjLx��8DW�nl�OS���ib�{llx}M�P�t�8��,R�c:�b�ND��T[]{�\s����
6�*���dq"	�u��k8�eu������i�-w�njDƥV����v|[���v������1T75�'�ձ�Q�K�s��r+g����>z��AcJ�Fh�4�[�pS�9���e��m�9��g	P˺�u��X+�|/�k;�I��� ?�Wm�,���X�duB��J~��t+���#�UQ�_����wn�v���y�V�l�IꢼA�(�B^�\Y�.L�x��ߣ-����ut�F5_
�z����$^y�a��"��P����c��w(k��������#
�ݖ�M��B�EQ�_�k�`0N�����(3V�8|vO�gnO�ss(�F�ޙ5,,�!����*X�x��1tp��ڇ��ױt�
*+�d�ȶ[��ԡ��e�=/xfQb�	?8�0����K@u�[O�l�Z�� �G3	�2��9О�eM�z�=�l��V4t��T���Y��qj�{b۩�|P�{�=�) L�7:�[�<��ku��?XE�s��sj4q�T&1k�2��A"��1g����X�gz�l-���|m�9*��ƹ��5�Hd?G΂Y��4����@�~m+f��C����p��3����䷿�ѓG*�Y�\�h gyθoxB���lp�2�7��O�ʅ3���[��d:"ߑ�pl2Fe���)?�3��v`Jԉ�R.,
�5`ޱə$ߣ6r��d瓢 !Ms��إ%��*k�ؐ'��ʫ�$�/��6۪�yM�\��T�o�� �ݲ�B^G&i�ڜS��k��L�������,�o;�~��底�TlD��Iy	� �DL�|p=�C�*6�$�W99�<$��ӳ.���)%Il��R�,o�suH��1�PW��T��H�"'��3�3��Ζ*�mT��kq��<^�왁 �ݐY	J��@u���a:�����5����*�$Z��#h5Q��7��0;���oא_�(�����'���B��cI:�H:�p�jx�������oCN^��/��b�{,�]
]zP21���@k�z�8HǖeVrsG�p$PFGGH@K��>tF@N,;etG	:�L�\��u���?�?��_?�?(�o�K�4j<��HR�\�MyߧE��~Ǫ��k5�Qp��se��F�-+u�@��4x9����o�=���=h�尀�Ҥ�	8L�# ��x������;�����ޡ$p�ey=�O��fTC\��J@��g_H̀��G���C�C�	��	Ĩ�A
�dd}�J��"I��3p�[X9�Z[�>��s�=�����^�˗;x��3[-,��<�a��9ZfS_ݷ�,��j%I��Cp3�4�Ja@��e��}$6�������dtky���T�7�'axbfF���QϺ� /����KY�>�rw�Y��<��+�>'k��	.3(�ex]�gcK�I��U��&_�3;��L����A �L{�s*2�
�*�Qޔ|�7L��K*4�*��ǲ�Huj��f��0t���2�-�4	�A^�ʧ޼�}��)MhJwSB]��u(O--�b1C�4������`0����$�c�G��s�|�����w�9��z�X�pv�/�D��;�,�kE�-�
D;_��p癬�����d}�k��H�ҡ�Tc+�"���7��#����_��������6~# K��f��:־{o��_"{�J��+��ILJC�[	@�x V4e}�~u_�>@��ͷo����?��_l	��Ir⢶�����9�n�'1������ߡr�������}\��#��3�."�r(���+_�}�b�ّ�d�E����>�������G#/ r&�����ÿt�#��[�/.�҇?��?�)v�^���:�H�p���g��q[UZ�_����H�����J�NtϏ�H#�=�e����8s��I�(=���*��XĹ��H�xO�a���ჯ$i��$���T��%��d1�yI�y�Yz&�ͽ\��Sг��9T����a��X:��J'��,��=��P;fIw�����O���́v*�U�9UC6�	�����_<�؛��-7(�ݞ��pƣZ232t�ck}2�n$!�U���-��������`P�N�C�����R�<?6T\���G/1~�f�ꍊ`�}V�)!�	�6q��S̳*��Ⱥ)�J�o���p���%�1캶<k�D,���n�&2���U3�d��g��q�c�OG��}��7D��#K�ip9""5��&�=�o#~�������(��P)
���IMf��Ir|�-����G`���ң4]�ϩ�Md��?ET���r2��(�O�����k�����ۤ��ˍ<7W(���0�|��8;f.`J�O�!�<-�1���4�*Ęz��#R�&�HD95�3�|<�P\�($ր����lѩ�����:d�Y�'�B�w�8f ����WI�(���+)�$����mP��+䲾-��疤����LT��.��D䊃|�%�!������8{����T��]����!ʍ\:wE��ƌj�g�5=<TGE�q���*�N��$a����!E&G�c�ef( �Օ�=1�&=�)%�$﷤�Cٙe,]������P����p�����z�5��H���VR]�e7/ҧح1B��k;�,z����{yv:|}]v8$9��5n����ą�-��uą�vAxX�$q����v�1��{�$�'ou	��58sS�14��Ja�]�&� 	M{�D�0��g{��d�J���_J�ʽ��$����Џ�E�5]��x��?A��M,*��/7P_Z��]W�b��e���	%�6��W����œG�(����ρI^�P	xGcV��C�Y�fF���u������y�)��m�T�L"�l��uI���sk���^���1�G3r�fѧ�.=9���J�8c�ñR�Kr`վ`�5��?7y5f<�^�J����Д�KU(�@a�Wb���CHs�'�|��-���4 ���o��e�v��g��N/1����MTyJg�\����u�M��B��M�v-ǎ�3���Vfs:�p���_�+dϮ �/m<D��Q5��1��7�c�?��P�[��������,������h}�9��0{*�v���=�ud\�9�Y�=a�y�\G( �z�,�o��3&��%[��r����Ր=#�d�� ġfD``$xUu�N��Ұ����Ѹ���3��K��8#��WϠ��DH�d�,goIB���q�������d�����x�/�^R^~,`��[��H'�eI��J��4�hTW�cd�d�+X?|���}��m�',8(���X\Cin>�p3��Σ�����9�%�����k
���1&�T�^��pC�MF�8S9�3�h�k��%1��Jχ �5畀z��(Tt���)���M6�zӽG� ��:�{?�WJ��gX q�*3�"&ϔ����ȿ��\'y�,��쳜YY��f��ty.�s��S� %f��KB�E���94$�#5�/�z(q��7�3�����˵��~���	&6�K��N5A2p
����Fb(��hbr�]Mm�M��n9_��B�@?+�Ym���e�$a���j�GC�`)!/볨�9�$�b�+�+7�AO��A�;@�R4@� T)r5��P����<uНU%��8�y���#����1
���!g��!k~v���s|p���p$I�V�*�v����_M�c#�+����fK��­�*R�ĝC���3�Yy���0�R�ez.��(���\l΁��1�h���ݜ-t���}z�LL�L�`��Q'G-���[��G����k}���o��?�/	d�?��噊pf���T�j6��rf\�\���
c��:�q�u�=��.�F���ZՅ`���V�`��q(L�0nLUG��0�X5� ���R%W��rH2Q?W�D6#g�$@A�+�^��#��u_Lc9�倡if@#O�B򾙥�Ym}�ؼ��%����T�_�r�;OQ�k�Pa�	Bv�;��;��4'גժ��S�>�ߗ���V1�����X�6O��I�NA��A�`��_.�.u���G_cד��V�P�o�6��[oc��Mp0��4��J��N���uhj1�ڤ�bY/	%�$S^�ׄ�Q�I��Qޏ�'g$%A,KrLz��q0ؓ�hF�WA�D�~�/�Kd3�:��x��[�X>{ol�s�$Cxr��H0�ݏ��k�V��V�{H��E�L�]�UY�HP`ă>�r}�����;䄸��a`�\Yg�\���(�t#F��͝�eMt�sJ�/
�������
��1��#��*�vac� K�t(ҳ�Z�߮��cJ��=��ʟ�9M�b~���O�k�;�R!/k`l�fy]R�H���]z�|�g���� vQ`ё�s�� ��:�}D��Wo��[o�>Wǣ��B�� Iw��)Vjz5��9=���T�=z\���w�,U��=�A%V��v<|(=pD%�.�c^��
:�LgܭWX#�[�K�����'ظs�H⍀�j�,�c����A�I�c��T���b)����Aj�x����8����J�pt/4�H�xᬬ��"{�����#�h6��j���r�����僑�QA�x��	�o����=9�1�Sl�3�pM�0�	�\3��P�O�Qy/�З���'����4��q��e7#���ێ�����q��1���&�ϙ�n�յ�}�++�ka�rFY���L~Y��(�,'`l������>���71�t��(�gP����	�����x��':؎�@�W��\x��޼�@>ӓ��}�]Z���w�FU���ݻx��]�5S%?E����,�"�����h�������:�/ѓ*�T$#l��KJ1)40��� ���r%�"P<����QI@�*�o�(y�����v�Q�y����\�i9������SnVn	F� wm�l�Ō�vbZB��]N�:�kf����L�i�H Ni��c2��9쫦���Z���LR$���֍���/)w�$�ӹ=��v�����Q�։�s�S��K:�D����o>�)��]��]�d�K�J�����$F9�Y��FO�Y���hy���e$��gKY�y�J�JP�L�$�A&� 0�9��v��?�e6��な�E�O�0spJdb��@�f�|SX�1a}J�G�� ���9=h�ro�,*�+�ฅ�9�2
"3w�	�E��;�9R}���k��U3�8jZ���OA��$&MK�����t�*�?�Z#NO�]�iP��0Q5#*����s�lp��`Q��B�f����u4���,��D��;���ڶgv:�;=�ю�́�|����?�V�T
z�A�E]��go^����@[�j8+��@��J��1��`<�P�2���cɟ�ԅ��Q0�l��|2�5�)��o���2�4UI��OtX�t 3EX�a���
��t�t[r��(�Jʝ�QN��9�j����`�R��[��I}���ڞ��l�A��1��H�Pu#���I�NG����T9w�m\�r�rǟ���#	lݱ:%��1�I�2c�v�$���a02sU�Z��Wfe��VDǡ�L.���}����
r+K(-̣\�aqnM���߾�\�ZCP,��/`v}U�t0L>wU��\!�q�N�!�@1��jZ�i�gz�9Ӂ̩䬓Lף&� ���^��ju�ό�s�'��hu��5�ue�fT���iUy��c��_�/���|���+/�>��{�������e-Q�Z��&�j���	��7Q�Ɍ@O$�y��;��<�Ggۜ*����Ew21�\�f"�ܓ�%���Ȱ��������^����e�u+NZ-�a�̜`A�
zt0Tf�8��a�(W�,R*`����0A���Ԥ�Ij����z-�KU����>� z(�Q�5p�'���r_��n`��Clo>0-�@ɡ+�B��|�"����q������y��_��6���g����qO-W���������ɧ���H�h��à��{�p�	@]���+�Q]9�5IV��`�i�����qq�&.��&������-I�bTK9���n�gg�xM��&�Mru�5��vݞ*��M�.D
�T9�U|&�R~M�e^^o=���ڼ$|k－��\�3ON�㮀�p���~�T���V.\���'oDY�e�N��1���I�Z����\��,�\ؙ�ȞmP]ɾ��Q�PP׮�y�w�Y�v:�KP����?�����ST{�pF#�P�"�w$�Z:�I
X�u��"k��� �y�*O�u��U�j5���茕�1I�w��P����6�i\���j��_����px��#k���W0q|u�K�o���~3Kh��]~�^6ѕ�5)UU����4���琩6�y�r��5���~�*�g����zP�_@�H�S�"R1�����@΂#���2��,{|N��g��HԷD׈RP"3Й1sn,x0��O��PU�HAw��Q�r��J^��x��m:����?����9ץ�阓:��'�"�3(�R��5��W�=�_����`:�v���Z[��x�rvs��Y�#|�����r����4��s*���V��B����-�{���FV{�%c�LC�RV��X���z�8z���gU�N_���$�I��k*p�NC~�	Qd��ǁ���׎3�_F�3��NF,��ba�7(�F����Ț$��a2�I%��8�Nv���'z2�.�k�=U�X���x��9�.|*[���#m���݇��k��0(MB�G_�&�˂�)H���a�SEjC*s�H�p8���dw��u�$/�sN��|;Y�Iܠ��eS�I��d�Q�9�$AFw&qҌ��&�6h(��̦i$?�����N��]��q$�hʥ�po7$�]��s�K�b����n�5��Zu�R"w�;<�`ؕs|�1[�#Љ��t�g���P��0�E81�6�<�JGj��9�@�&�a�˘?1cgp�IP_8���U8�6N�^b����!�J�����P��4+w4�[�1�*>i4S%E���@���s���Ŏ\��**i��{�v��k��g)X_	V��!��rQ)?K�.���z���h� a��\2֠Z�]5(���ltR+<5+�{e٥`�m�F�,zrOά�ֿ�oq��M���|Q�?�Z�P,(�
�J倍�饆~A�Cy�d���e�(��Ey�*E�SI�XAZjP�	b�A�x�|�r�l���>F����BO��1�bg��ڇ?��� g����q���8B����f��>J�.��V��5�uY���{�Mf.J�g?5������dUȱ���J�jۘ�1��(6C�܍#�	x�UI�ϛ����ï���u�y���	꽱,��x����� �X.[��U��!eS=9,�;���Ecmt�$)���>��'���ʎ���˥�dШ�kB}Jb�e%C�������:�����C�M9��P5.�@��y�.O%h��k5Y7�����ޙ��&��,�GU�J^��%�=�S�bǤ��T(�`c��Z�E�P�$Y�4fy�ob���YYvh06`L�z�ŋ�zi�o��-�������'���Ԉ�~6���/�k�&�I\�����k��(}N�(�*���y�T,#-������}����aR�jTXYV�rӔ����D�����k�Ǌ:X)絓�
�(��<��4Hs��(*[@���e&%��࿥+,�Ā�g�G  ?+�1��|�|��՛o�q�6�=��� �a������y���1����Q��	�(c֕,,�n��1?k 7Z�r�N}�1<('��=y�@��O$q�������k�%��*K�Yo�gu$������y˫7�b�~�Dn��I����q��ɟ�%��̞����Ғ�d/e��J5��3�A�6��|�W�I) yٳj�IU��<��%A.��!ېdxaչeYfIPfQ��
��M�h��K"�f]k���+��홣(Y�D���>����w^+���QQ�;�"�z�J����)M��+<R�Rj��\�/8�W����K�>qz:ԣE4��i�븶���}�
���ީ<�)�0I �vl<Gj:�9K�Li����9M�}K�S�PL�^߇�nG��L�t�l,q�$��w�1)��ڕ�N�%R�9�W����@���n��Ʃ��M���7�F��9��x&	Jm��v]8����q;��`GC�lym�b��.M�,����0o�ٓ߹?����B���Qcj��&-�%�����g?%%�3:Ԝ�_đE���aӇ�t�;:�����0��S�''�O��o��5�<�I�Ɨ<ݼ;��ӫUMXz��j'tCI�%��H֖��5��gv��IO�zVz6᎗o��l��U�E(��1n�IgD�^'����Pw�]����$�ȟe�d�'�������qS���b�8�8D�جJI�~y��i'Ao���{9�{�JJ>��a@�B
�:~&�q��'cut�fsF��Z�Ԧ.�$�Ο©/y��a�a�~O�}	��B>6n��x��qG��JAb�)�4x��V�W�]JGR���@�� #B��)�簴\S~'yx���G=m������_�	���9��Ku���!������W~�� �<@�Ś�6�%��aj�Ì+����{e��X.���'�M}k9��\���7�=jw6о{�G���s�vL>�|U\�b����B�6�w��j�RP����+�9ئ�<�VWm7"��mE4� ��>��^��f,���"1�Rřga��z�]�7p��L�4dl(SZ	�"�
��(��ZҼE�;Ź%��~7%��Q0��o�6�V�¯�!�(Ug(�U��Z���~<�Ę�^��&���e�O	�ӋA�"��dR�j�
�����*gڗ�ی8g0V���{8|q(믤s��Inڸ�9��l{I�i�5�?#�C���IQ�!�]���Mm�)="ܐ�$���d�<M��@P��s6�0�Z��(��b�c\�9ˑ�XI���fے��&8<����s(}ﻲ^�b�-oI�rk�F�.�ɳ�!���<�8��D�Д`}DNU{,5 ���2NgM��f~6դ�&�LRU���r�͟Y��uI�� o/hc���mY�]I�|���u
�o`n�:��<��ޖR�t�FQA�O�����d@�W74��q&Ϫ]���,|r�#��Q�<�K�_�l�@ -?����1�mɽL%��Ҕ��U}g�;@N��&\9��:��WP�J(Rs?1JHN�ܯ�h��NiU��� Y��h�K�F���������z�n�����˥-j���H|�p�$FMf��އ(�,�&�=��K�H~�>o��J-B�ƁV��C�v �_r�
g����#<��ā\S�}��kl^bi-o\�����X��ʹ˸�����"��c-Lt�~��T�R���^��}>��ڢV�IX��QYXV�K��J��򵋨�_P>��7TE������s�J2���-d8s@�;QU3�[��p�v�^��\�1c"��:�w*�̺�E�=T�o��J3�d��O]Ki����֤�X��LgY�����1��
l�_�l
;�e�����ɨɨ�׮M�mB0-�0�8�����Åd��Pj�y�T�~��PI��/�x�]�j��
��<�"�����3-[J��P7?Z��Sϥ��'{��pe�s����!jj���5��EUv3CZz_��H�\j��z���5�ӐF�|�JEr����
�ڍ8[Nt�h�5J--hB��\��,}��ߏZ��!�i������9�T,��B��Pb�
N�B�Q���!~���_'i�"��͖2ɰ�Q���9���(��F��I�I�L-�f�]!�&��--!"I�Hv1��/� �ԓ�"�RpF ������౗l��Z�8*S��<�wjvSS�f�Y�R�ЃN�?Úu8��UgSw�&���~�������^�u��ƣ�H0�NLf���
]����*�8�h��?g�ɍ^�Ӓ��sz:|�`;�.�8@����F��A�����Rᇚ�l���k��6)���͆�oMp�e���vX���~�1/�A�U
G�
C���45Z���B��\�k�!��FK65��1�i��w]��m<A�ݕ?�QY����+��$����$pCJ��`�+���A)�8����Ea�"�1��&�K�AF@v�x��G/q���7�(�U���5{�<Zv+�x��>��c|������y�%0[�D>Ð�^��OUT"}�3
r����� j�y8�ã�?F���N�Q°&IO��?�{E5���@iu�|3�=||�?��I��g��FT]jC���`��c��� �<���l<�(��In1�������sx��a��M,\���"����0̝�W��$y7��.J�r�K�9/���[@/0
n�=�_{��kh:q͡��I����ņoNu+��y٣����? I�I��ܸb4B�=Fn4R÷�|��^��{]�Y�CL�*%�u=� :�Fnx�̨'ｄ�$Y��l����ܑc���/*s�}�h�j�� k��gTH��֡]�zl�Ib��PiO=$8����al�
B�I�ܘ�$U���y��51xx��!�+Z�% X�+�N��������s�|�F[��"R��2���k�Yj���h��٢�;�<���N��/�'�׉ 5��Q����Q�rQ�9������էؔ��k� '밶���ko�v��Jb����  ��IDAT��Q\ ({::ؓ���A%4&Z���&��^���+��sJt2�1�:�I��.@�/�w�IM2L�F�T���j�#�����C��F�F٢<��HRfl�	���8�Xa�G��OU���Z�*��q�>�"��%	��񉪋�I�*FC:�a2����&����l?y�%k�*2E8��j	��y�� @�����obR��]>'_U,5	IF�w����P)_>w����Ėk|���K���mm�![������#Ҫx8p6c<��t�^!������#��e9%@JR��P����[5�jp�L���2�ΘBM����[��jz��yx�ncI &rou.��lj�H�ʪ��x�>g~�����k�{3���������cy}�\�����T�Y���-}Q^R��W`�M_��u4�1��8:�� 5�J�a��c��Oմ`��4=��k�ǂIw*J�vu����@2t/�'Ngj�ߝZ�Ȼ���Y����p���1�Ll�Hǆ�
��885�3�Ν�M����������[�׷7���v�2�-���!��)��8��]�8�qر��t����°X�؂#>-fge�k�O"���i4$���|���&������C'5���5�L�9qlrf�Ol���R�����1.M%ju.�pC���GcґC��,'����~i�q'�����r��\��(	��FX�+��'�����D�Z�2�>��q�R%��Q��$UcȘ>o�q���3�鯘>��6���y�ͯ$�&��������������PIC�
:�)�'�_fZ>5r�֑��1�rfb�L���;Fm��"|�0v�N�b���z�AU��L��_�ԙy*�\VT��"��&��k�B�d��y�2��$kZ_�#5'�6e\f���SY>�彩6��!�2��߿��~F� u�ro��)����x�%爃�g�����$
9�#�J��-��G���c��>B��P,�q�O�����0���:��|�UWՂ�@Uk9$�H+!�L^���.�g�p��"2�e�$7���[o#C���.B��z����~�(T�j�=*;���`uѧ�BFh���'�ӝ`���h�$����'i�$�f}��&k�<OEGsK���t��� 6��DX�7P~7A5�2���e۞SN�g��W��W��	�ӵ��y��4%z{�T�K�+g�����?�P��*ړk�n���Q��cvf���~���!�M��0"uA ���i�J=����.���-2+5���	2TΠ
�g�9��D�
T�JiFE3y�a[ ^sK@�e�_^�_�7��8	�+�S��V���<�������{������5��{CW��������T���WΙV�=�٥��V�u�u���P[UVr�y�\O��&hZ��;9���.�;�%,������cg��R�� �ź�{c�W'������
0j���$Q�8�G��C�ac\c�c[�Δ�0�+�R�mm�G�F�$1���j}Q�wmN��R�4
l��䗿���/p��K�;�t�A�!�����|7�"�;���.a��8�ٔ�=т��Hib8��k1:I^���y�;�.}�,;F0�3W dJ��a_��b�����d{Y�3W��+q2�}=`i��s���M�L�)r��Nɬ�j�C�9�ٍ�H�h��5��0��G8�d�����@�.�'-}��C<��TbI��߻- �������,�h��$	���,���-,ɳ7�g�̠�|���m��z�A�#�H�5v$�1ToD?�/Kg.`��v�kH���O1'	�o_�;���7.b��*�9A���� ��̠BZ#g�8�OsG9>�R�n��sV��Qs&&RA��)V �e�4�X-_VeW�]4���Mbg����"��ӂ��;��µ�����I�%�K�#�ғ��7#q(?��'�8+���E׊��)�T�_���4N�.�78�hN��q�q�6���wFj|Cb�+65D��&��	��T����W�ü����=;|k�#��=3'�aB��r�nj�~���9cU�ҩܘ�W�`]�����бX�VDIi<֯6���L� ����M{��<���Y�V�)�c�9���@�)~��ij2�����h�c���L�$o|.�o�,�y��a3��vڳCC��(��ܤ61�W&罺����T��)AP�+���qT/�Y
y%Q%��d
�hqa躯�����ۤ�������G��?�?��K�g$WeSd&�ߜ�/�����Z��__��O?��_��X��ܫ��~�2nt�?]T�%���+�&m6�?��'=qN�D6!�B�9mcq���%fPiJ��|N�^ӟw�i���B*Opz}��H?U�|��99�T0	Q�/����CU	��'�nYy�(�H��P	t���m�1�r�4���Y�xH���j��T���
�s�(��̗�P5~QzRF��U��F:te��c[���8�<;�5�������R%(�P �
��N��" ��`{�w�s�T��  T
�)����ԧ�I3g�U���P��	�a�2�y7O��ﾋƟ�	p�"Ғ��j�W�����X�]��0�� �-��F�E�p0�?����:PB�����GF�I�*E� �<+y)T)z/���Ȓ�. 6��>w徏�z�ەU��byi�$�pá���U^�bmg�V��!�+��]$��Nb �kڜ�J�$v�cb�Q�5ZD�S9h؝�e�f%�s0��	8YX�2i"f<>Ƴ/>��_���	r��>�����
յr����w���o?Ǡ3B%[DA�־VP�
�醩!:у;T�W�i��U2�[ң$'�}譑
(w��8L�'�+y�%���e��;�~�9��˳���7�?��-��փ�z����'x��A������(˽��x��o ��cR��9l6�$�*υ��LʸW�R��4�hY��%2���u�"����!]�������~[�A�����Ȭ��[�Ȯ�E�QU>7JԺ�¨{" �T��V�=��KKhW$��ءUn&�0��;� ���:��ӵ�����M��x�ʡ��
"g7H��\���C~�$���\�P=�=0�58:Wӑ}��!��V���#�-. '��$ }�V�bk�����!�i�;��:���]_��+"+k6��1�>:FC@m~m��F���]�՛6�tw��}����}�p��5��Ϩ��qS����V�
P�8���"�G%W�� �N��I;�{=���;��/q�>1$�b��kLs&��z���_� I��[�Q�zksk
����}���;���`���K+(]��ٳ�J��G8l�	��H�����O6��� 	���R���1:{�xq�>��	�fX^W\2H�5���;�⳿�X)Wųk��u,ߺ���*
s�,�|�09j!�y��������9dfg�zU�RVԓ�����H��Eq�.	� Y��v�3���[�]���w������-�~u�' '���U,~�{@�"��F_S��s(��<E��ϧ3KZ�0�;��~�M>=L�K�1ê�h�f;M_a��F�7K<��DA�c�k�a�*dKIM�x}]��'{��$Y�]���\���)*EeV��.�ըF� 0�ik.f6����YqA��l������ �4��]Z�V�����k��xϽ��i�h4#Y��7�����߹��{�K"�c/�I��NU1p������)����9�n��9L�� �'��n�꬗��>%���|��\���q��6S��^k��ަ�4��Ñ;
��߆ug�UŧlW����u�f(�}�|Vv�R���1�rF�j��Ǆ�� �n�4A��o<�I��t���S�=u�"�1f�H
ҙ�4�	��&cn�{�������T���|i��;e\��?�ȅǽg���迚L�����t쒀0)(@�7*��	�>�	;�3��������˝shҿ�|��s͡5S5J�i�%L�����o|�x��ПE��-oNI�j�;+�y�f?.9�b:�.���8硰P�Q��A��G7G�ڡ���U�4^p0���d@��èI�ʐ�1P��5���I�+��3S(7��"Ip��2+����kV��-x��	��Y���ߨ��4Vzy�1�+Y�J�R�>�D��p&~�$��ϟ��S��5�캚�w����'�B�R9�-t�P������L%"�I�C�@k7"UnA��T�R���j���V%�D�����FxfUr��{��,�TmH�:iš%�Ǚ�D�lc����{�}�����?���˸s�>���a����C	�(����j�t��z�-��� ��&^Z?���ST��nO(oY+���SIp���:p�t��VB�NƕH��L��$���Z�d�����:���s���}$�r�� �76������=�쪫4_sU��|SnT���rDNT0Sn9g%*�a�!�פ���؋4p��=���Ԝ�g�?�7��'�ZM�w���o�]�E�5HE�j�'�I���I��·_�郧�z	���k������a( ��R�~��-1�����C��<��K��_�-�g*`�)�0��xOⱍ�S�7��[���͇�+M��#��`����bS^#5'��6��~�_~���<Z��\�� �2>��g0����hc� ��U�=��%n?�f��U�D�-p1ͩ�h�k;J'L�,�s�x�3.��)G�Zo����d�*[(R�&M����$��/^%wQ�����2VH��C��|!
E,��Jm~��p�܌[억$�̗Z���HKM$�0&�CM�����o�q�u_%C�J��l𷿒{ ��"^{�����߸{_~�1v�=�y�guYu��1�����;5�"G���H��������U���Z����S���$	ӝއw�L~W�������`�ϹI�mn��P���_����so��'����h�5gZݗ�b����$�]9��N���׉��p4����������]���%���YuS���,�Fb����z���n��$n���n��s�Un�a��5�~փ�-�|�)߹��^��K/�b�u�.Q!��˹|�������j��`�,iL#����Pb�$[�e}��8s��Gٳ�*�;c�����ܔ뵏FC��|+��*�l>|���G�Hl�q�&�I�|�I�fF���b����L�7+ ������2�����S�<w��2i�3�@�8�c�aR���S
Z(��­�c�LI���Y<�1��S�UPK�@�#yn���e
��vF�h�*�ɴ�i*WR�V�c2�l���Ƈo�_W���{��m?[�8����g,��i����u�|l��W�Q��Gh����@nUyLGrN�#��!�юRWXvC���ʋ�Ѭ�䘥m��$��uh����ή'���@Zt�<;-܄fި�����L
�ý�q<���,�Y��L �j�C��x7\7U�9޹]s˜f�a���X:�]K(���#�U�^�Z[��ڢ�a.&�� ��/l�+��-4�p. �/��˦mB�@��A�
����f��7����j���Z�gmI��k��30A�vD�|�����[T�r�f���P\b�	�>G��꥓N�t��낇'(���˶ٹQ�%�&��*�CL&�RaXF�t&;��Д����0o���6�I�Bں;����pm�0-*�T��34���;���h��8
���Q`<�b��7 O��3/}O���ݞ��|��X�{�AϨ��K�0���6��	p�Tp��>6��Lt�Z���}�Cy� ;s�\��R%�Cqnq~kN%Z�J<:d��~��h�hS�"���}KuRV^~⩣��WCU��$�<�7�֒��M�{�ǘ{m�s�p�ÿ����sէ��7�9sg_{�}���t���\�u���E��c�[�>F�b���d�<O+s��n���_r��}�af� mr��گTՔ��Tqae���s���p� ���'19��[��_C��
V���t	���0��Z�G�f*W7ܓ�GW�@�d�{j ��/�� 6��8���kO��t�Ӂ̅�����P�],{=�ǘ�W�[��^��'���%9��_��^Y���{]��`{�?�T���^�[����=|v�Gܓ�����G�B���	�0l�}P`�k�$��]�xz/*4�@�5$�������x� ��I�[ qpDs8y���H�+���e�䐫�MHe�.�=���_����.�ųhm>@P��d��$��\�۲n2l�Cj���LU�2���k�Ƹ��B6�-0��S�sWEUJ�*g���^Ӎ��� �'�!jϭ���5t�P�잀J��8��Y�t�/���s���T�sv$kA���7��E 5Sʧ��50�fF�(;�q�
u��nZr�9�.���+�ӭ#u:Ŋ����˱�/�n<�����G��������΢d�=�{������2����d�5����Vr��Pe7H��O��%'���e�.�>dϕ�`���<�4ב�"�\)G��Cl�}����F����(/��r���=��E�:�r�ڼ�]�Ȟ��>#��P����
�Z���/b��e<����=��L��=&�	������`�B�5/�\Aiy��x��$���7wQ��TP�T��3��H5�uXA��.���\�����d�<L�%�G����^��2��Ť_��������j
uA��q�Ȩ<�HǒDV�v�"9�|I��W�TVU����I����\���XQ���)�`��Ԟt�t=�NA�c
'[��a$L�d�Eg�s�1�M�����+6�;̋�������`�8�᫼�Z]鄛/��Jɴ0��؝�?�b�!7�n���]c��4�{j��dj�����m��ɚ���̺˙<��JEz�Y�ߛ��~�nsꡳYOu3��((�ivB�:���j*;��!�W�όQ�]�F�:<��J�R%O�������P+P�=Z��W*��Cs��y6��(���_I��:1Q�P&��m��]� �\"�!=�Hߑ�oM
�8�����~ �RT�[�K������Ь{�O�s��Eu����P�]|K������6.���ߊJ����ÉS��u���#�-j7�d�Ɩ���<��؆
lkb��������!�(f�������u(E+�'-@L���#q�<M�,Sdꙻ�D�g N���S�-ͫ�����2�T�5I�y�7`��4�)ir�V��ǀ��e��gD	
c	���L���S���J�j���$�s��0CSNxb��M���9�����c�[\:��V��ְ����h(W���;�ϰ�����Y���;�S�o��-E�9��\B�s8��$�o���xC�C�x��䰈�~�����w����`$��a_���<Z��̵�h�7�}��>����C�~�k�?����')����(Tb�J�J}��$/�N
�RV���}�$n8���k������ۯ�����ݿ������_µ�G��yD�Wm�qkӧ�P��S�$!��z�F.�50��j�KB5�e���Ux<����Qq��ӷ�\���Pe�"IHo9@���x-�^z�����{;=�r��##k'��z�"���aswޠ��\3ޙV��p��fbkT�Z#�6З�~4�eJ��to:6�{�� Z�� t�,�,�A�\��W�M@_w�m��ͧ8�I&rw���F4~ZY�+�����yW������~��;ۺ�Kr�+� �%/Y�v1�%5R:^�緧>��p���qrNI������8��;4z#�$�fK�\��2���p����� ���f�>y��޶r���.^Ks�ؐ��5WRţ�0TU�9IҲ����QW�ըȡ�J���❣St�,���� r�"Q�7r�>�&����x��Gw�xfE�M��\Ď��=l|ѕk��KWp���S,��Vv�:�g[����l�����D��`�kw�z�Ζ:�r����N���*�U�(,I���v�t�*(Ӗ�ɘ$-C*�I�0�X�HC�ؠ�����p�?Bww�V�(��X�_�$�:���e��{���&�}y��Ĭ��[��
��Xi�؞�B/��Rk�:F�=��>Tu/On���
����p��1���W�s	�_ZE����������%1,���j�c����+h�$z�:vv7��k�G}�%��I��~�����1�~P��Ғ$�g�.�[��?����k��L��q$If��:.J�b�F2Y���g��z�����K����ڭꬭ�!	�U�R�O��a�%���>��!^\��>I��}|;�s�;疁�ED�A�y��$^~�5�/�ӮW����K"t�G�T1?XQ���m�!o�-Nd����(p�U��h��]f����V�,����P<��4��X
�%I���؅���L��7�M��JCl`��L0B7`b�MU�%.Y`�;��S�u#flߛ%�s������W_G��	����t~�F����{��	WJJ�+����T�V353+@h4��/�����3	�I���w��N%p�K<#�>5���S�&r�Uem=�#����N��w�樜�,��&�(�F�քH�\d���^�o;Jsdg��b���[Ȃ��I8���w��[���(�
P<7�L�ib�3��v�Y�6�j!�w�.f�����N�x���9�k�}{@��]�ZL�B���0���t)�O�u I5�˧���M��׃{6pbU�����A�c�����6�	]����ݴ:E�d����� �� "$�f������{���ι�²��a>K
|O�ۋÈv�Q5��&Aw�,8d�D�7����9_��L��O�#��0��5�ԗP �T�����#��/�c�L4���!��8��%��l�-yT�UD�^��Q��D 	8+�ڒ�dG�l��&���}|��GX�rK�\C��e|O@�����^�-���<<V����;�p�� ����G;�%�n>��F5@'���	vn�`O��3	z/>���5,4�e=���?���<�����M����t `m�C�m�|���D��p/&EJ@#�O�)\� :j{�3��O�Ǡ���;�����q��
�� X<����� �wߑG���sɭOpx�dr��9�J�J���s޸k���SA#�}�d��ê��LbN��tTf�� L������^.`�u�h�v�
rb��nI"�n��ŋX��*�^"�]>��<}���#T�{�#TT�U/����#��X#�+�BZ-�Z�
�˄33�X��&MG�kH�&;�e:ې��wi��*zq[�cln�O�̳g���5�	�X>����Ϊ��⚀�:�$��	���\��æ��S���x0b��j=T�)��Cuȟ<���*;���a*��n�j���P�LuG�QyG"G{~	��_D���v6���a��8#�'�I�,I�/k�%פ�vQJ"4D�SA�V�܊���6�$�ғ�m���	P��U�	<�u�C܌aI!��%�]�� R%(�(<�sO~�ku(.=�u͹�sg��}H��g%��� �w%N�>��/���	J4�u�*��_�`|0j��rq&���s�⬀���X�sv#���ǑĄy���u�5��r&�t�=��ET���o_��
��-k���9)J��ΟAW���4Y���B�b(E�s8]�2ͩ$	ruY��$o�#��ҕKr�z~�I|iT}���u��(n/.���5	,v�p���o7aplJ��^6iQ��3x[�256�D��
�p�^X���޻��n|�ljU����$˛��z8��Ž�S\x��/��̯��Z��Uy�cJ<K�Q�5v���ߒv��Q�[Z\P�^n�c5]Q �
B���Z�9@�ʵ�y�����SY��r-�|����X�bY�ec�$�d�(/u��5�2����UV�YǃJ��,��&���J�q
/x
�,�Lr�ƫ���Me6 Z�v�g�g�K����������Bf��k��R��ĞT)�n 8�=#�|�wsc3����Lt������s�>�	���`�X�Y����+��U�N�&υ����� ��d�Wsn�ܳ������8�������}�5�T�r݉�>v��N]��5,Z����Our|w��/fEA�u
��#	��L5�g���T4��Y�#�P���5��hAU(��l�p��P��׏,��Ꟍ�	��S��)�̤4ws	���<a�ٗ%�^ο�u-�E�������<~kRP����A��x<}g2^��Z��e$�Rb�P\ofCd�]2��n��?V�C����������sOlt`V��Oq��m�eD޺�����f�*��C�Q�<���D��3n�>�D������z�J������T�
(��U��%^��A�����3��o�bz�O��T�Q�XB����QUŉ)8�H������O��S/|y�<,��� Ⱥuԓ�xt>I&�b:��yӒ y#M�t�H����BL�����PUmHoH����X�T)�����X��m
�PQ��{k�!�di���F|k��IX�p�<z����7#��*a���Z��l��7���_��d���R�x�,ݪJ�wx��_}��O?�ѽ4�S��D��M�8�I�C�X�R��|�����������P[_�����[x��8�s�����&�����<�JT��3g7O	M���m5+�/�w[V����%����3̟����2^���������Ď��`���p��/Q�"@{�AW�W��2Z��4�v����FOsC�T�Qi��¥3sn�6����:@l�f�T�م����H���g�����_ZE��\�[Bs��>��&�/HҰؑ��)v>��[_��q��\��V���n��4�R�;��C}_e��h��F���t$��G�z����A�T��א�v���{4cL)��ʝu�uʽ��W0/ oM���ڢy^��h���{�3t�> ���$%z���޷)��.�/|!�_���jR��a�?�h&	I��m䒔�C}�;��8����G*]"���6P� Rv)w�0�cT��*��L��L��,�j.	AZ�h�C�����4�U%nKR�l��9KA��6`̽�z(���2�:c`C�N�)in38e*�U8k��{Y�8���&�G�6�na^�IӔ�حc��@b̭O>�����w%韦
�Bٷ#�˲[�;��e'R��b��ag'��
�,W#e�5�c�X7^���嫺�H�3w�
k���������r���]V� �g(��Ǐ��\}<�l+ހ$|����m��c���w�b���U�K��u�:�,�&���2�7�x������]¥�}����S���A�I�<���cIB%�Qq�a����_�l�Α�s��r���|{�rڡ�u%��;>@�y��۸���S���+����5��
��Ԍ��s6�#d{�����Ƀ���]<+I�Y��XkVN:M����A�6�a�7�@ ��t�������mH,ar������>��>�s�xwi��9��-J2�W��%r�x>E��O�1�w�$.��pڕ�<fN�x�N�S��@9�~�)f\h�ˠ݂S�&��u&��Ӄ�@�ǜT�r�C��Q�h�|{��ت��3�b���5X���Խ̉wd�i0�	#T�HhaQYs'
��&�B�]�V��#b���m�3��%�	n5����Օ�ZHI!n�}�8����`��P�9��N����'~���O��̍JT�
�f?l��������o��,P��_��H[����Tg�I�i�ș�B's�S���*��:���;R�7t6l�E����Y����y!S"�����L�w�%�%�2Db�|!r���B�2�lX�;���I��u�����:���CL~>�N�eY�\�ʵ0��Y#�8�\�jKV��5F�a*�h*�V�u���<���  ��c��pZBJ��&�����]�{eaf|V��.��0������$o� p��I$�Ȇ��Bl���(�U����z�ɹ��(��1��F��`��(�j�ߴ,�$r[�u?<v����(��LмN���꩟��wy.y婜�>���a�ʆJ2�3��$+���\�=�&��˗�VR��r�x����)k���8���&�h����0�^zi�Vt��M2�7o�'�~���?�UP��J@F�2�:s��U=��D�C�>%A�NT�� f, ~H��t��N�`J�����ϧ�گw׷�o���:�#�X���*�2��R���fc)Ц����ٟ�y����^D�.��P�˶P��==����-l���ۏ��M���4^� 2��㴊^�D�k8��kX��e��
�\hB2$<�u�>�T ��67��d��iUPP+2�먱;���U+
^��u8|�j,%4����
��!���׷��w�E�?���L�@	��6�˦�st�}9��ܸ�'�V'}�F�Xd1.� 4�g�܌����!� G�Y�Pu�lHL�,|�L����=�sd���Cy���y�C���_�{���+�Å��D��E,�y�<���/�p��������� 姏���C���cU;U�(�33��ɭ�@���*t��RhHI;�Ϥ3T%R	U&/�i��&-��u$�����+8w�y�/�c���X�Ԍ~GD���$黇��-��d}=����>��OТ�olJ`���i��h%���uypu�ǔ��֖�ݤ,"�+ �]��\�n3.t��U���9�5�����>��_\�<%�ٵ�Q>�&�ޮ�Մ+��&�S)���D� �a���z�]#�[SO+�T�Yi�I�#	I��p�lZZ�X5P�XV1˴�ʽ���4�D��m �����]�k;Wɵ��}9��n�� .	|S.�z���Ҳ��.>���A���pYH&���z���*�FY��\+vg<x�Q�,w�v�x���h�i���T�((���0j49�h� B�<ӑU�c��J����i?�8��<�H?Ar��V��l�{G/��*L'�)��z(w��`c��a\��� ���}Tnޖ�+�갇:�rC���oIF���<Fcm�V�zM�pdMu�0Q/�II��c��tHI�ִ�|,ɷ'������Ý=��H���{#<���ǛX�ϘW�WZz��w�Q�%���¹����}�qP����٘R�=���}�[:d���;�&��"&4�dz.�h(V�#��LU�gw�`��]���[�
ƿ�5�ݾ������d�<Hwn�ђ�a�qr�G{����Qﴵ�2��_�i$r �P�py8<����tW�?p0���Dv�o��*�a�.2U���fn$���+��>���)+J�.D�*�Y��8�W��c��q��j�4;#=�rՃ�g4��]�0���/�����+w�����3�gZ<���?�$�*�b=�R��\�uFObmW��܇��v��l���<��{�����Wg���p-�T��"�>]>��R�y� w
I'׾�ЙN�)X&����ŀ)ϗf�ʊ�� ���Q�g�@����G<�@N<��>��b�B�s�Z��I�1�й�p���T�U�9��2~ �G���Ě�с$e#��s�M=�����J��A���ʶ��o����"���dY>t���њD@: �d�£����j��~*�N0���L�qD�.@>�#K�|-�rG����wYK�B�:d��Q�|rh�,L�@@z��U��CS��� ��e�8Z�V��{S��X�lɟ4�j[���L6azv<��<�F^�v>{�����u�������=|x��g�7ޒ=V8��Ï9���@�h���iz�,.*���*R0�nĞ"ku��Z�3�����L���A�<�TW��
�1�s�d4���d�rG�^�*��8Q��iP%FJ�ҿ�`p�&��V�Q�c�J�ټ�ƣ@��T"�-]D/A<>��k�@�*���啳�_����~��w�$�R⸻��O�HʣY$A��*.�-"�����M�T�!������Wcй����Y����,�b�>�\�g�o���Q�k�94K�}L��T��	�hз���TA��e9�S��|��v��p�,����r���j�ΰ�{2-uO��r�M*K�I�RM�\;mT�ɔ�=���M�qw��^���aU�K��>�Y�"�R�r�#IdH3�{�������>V��4t���7��8�MM�X�2U��^lM����[����~W\;dѧ���8a�5%���u���ξ~�����W$�\6� �������s<��e���X�Ãg��^79�8�N ��^ �wa4V� � i�
E��1lr(�9e�ҳB~�"�mG�y��(ଋ�nOiZ尢��t��P����OqA>�s�^�j��[�����k\ީ���E��㱂�1yF#����P�"�(Uw�Z������ؕD�4�)߷�2y�U^��d*�����f��n+�eILذ��YE@�3u<���tk_���
�t{}<��X�ao���K"y�:�O�S��۲O��а�1q��E��Od����(UT�Q�s�g�;4p���Է	,�f��=��+�n ?�W�e8���œ�3�:����Ħs�����dl�UR)8�%�3�=s$�q�Y,� V��(u��a�{Nc]�x�	!��s��W�'�~v����#�ܕ�֒���c�ߪ��
��`���桀`
 $ۋ:�F_�qo`�`�wh��kE�O����������^�pA�J�G����� �/����}���$t�G�N���hH,���O&
����{�n�
����C��z�H��*ݰ����1£M��%���P��@֘$��3*��;�x��I�7���
z��j�q����$u���M`b`�x��5�oҗ�Fg�:/?a+X-#����ڸ�Ku9�j�ϣ�z^���4�`�^bm��l��1H�7'�Fbp���,��$K�d����Ns�t��}�Y���	�����%9�E��)�q_�W吾��:���y �N,�|_�ЎĩAb᝘a �3Se�Tr���ƃ�vw*�2Kg�p���!7G�Δ6ybgZt	��뤻��P�܌��vb��Z���{��, ��<�rS(��S�2��c=U������w�N13uJB:O�FdI�}��X0�)�<��}Rq��T���T�xgݯ��to��SIz�gѺ�R�~�����x,,\��+������:���IZ��������Q�����3I�3I
Bō�'R-�ӊw k�xh��Q9��"�}�$}"w-��3���� �B7TQa�m�=6���`�����#js�!0?/��CkM��*
�C'���y��{��5�,e��7�z�v���ko����C��Aw�x�����0�J��t��װ���!��7�sk�ʁ�*��Wq�ZG�����������E�_���*	�Ь���FeP��0p���3����0*G��_�����b�{������rK�];7iŏ�Bkr�,�[�����P ��������c�&]�|ue�z�9.茏�ZRPt	T���.2.����:��
Mj��y6�`<B_>�.�s�p��pNn{uΤ2��)���(�8sf�W_AU�[���֓l��Uʞ3�Ku&���O�u�p��+Ӓ�W��g;n�L��S{���P�ߋU{Z��JKB)@�m>*�h+�\�Kr_�вV8��� 7>�6��[7�ƓOo ��4JИ��`�L��`����H�Z�1!�\9�
�bV��\�\J�5M��:�ݪ�P�5T�q+j,@u@M{��յ^x��y�%5+���>��m�=x��RUEb�}���Ԯ]Bu����_��^�Vѐ�1�)Ѹ�c�RAT��f�'��˽O���D��86LG�\�G�q{6�X���	#��1"�`�SQ�α���	9����$�u�!IF�5�^� Ĺ��sW�,����1t8xtG��X��f��������(OM��R�5�~lFc�M�K7�\�cW������c�W ���<+������z�s�
z��6�+5,U�hV�2� V�өĤ�d��L@/jE��n߱�ِ�K��9�Qs����*����4�-�rL䞏�)F����}Lǩo5HO�����D��P����L(Q������WW��Gj�%8#���A��ã4P��ڱ��$�>V#0*��V���︿h��Fp��a�*ɲ$�&\]�ma��s�CT8%�χY��K�:���K�>�� 
@��C�hX=����<)G%6c��CI���ֱr�;�eJ����$��6�U�˜�)��ZF'��Կ�g��������ܽ"���T6������B_�Qcv\+UTΟ��;o��rhΣ̈́��¹#I3�A���;|v���43ŭZ��K
f�b��91�z"vR��p �LG(kWM��>�ݸ��_���;F��*�"�*���Lh�k(�>!���ik:�Ĺ/�B��ܔw��f� �1�7U���^P'$Q���hf����d�Y��������V5/�s�r������2ڪ>_UL-p��E�3
N���'��ce��ٟ�%p]T��1/�Rdk/s���C�܇�#	�������*U��'%u��w*!������G�{|'��V�G?z5�qs�:�p@EB�,�5jq!� Ĥ �S�aE]ˎ�i� ��f����TM)Pp�0UIm?y��,�r^�ࡦ�T�#b��!�<Q�Z����C>QT����P�`�z��B�>guz �[n.!\�i�:ZǇ�}��([�%MV���W&�xE�E9\'H�ʫ�Q_ZDgiU�WS>L�H�$#�,m�@�� �ѾҜ�X��]r�H� �6�d*hh�D��a>�����������w�}
xm�P��>�_��?���w���W��O�������Gg}��8:�ţ��8�'6�A��u��V܀X��2�|��n��T�ә�`lK��)YɢZ�*��VA��} ̿r��s�����`%�+������*�̷W�Y�`ܞ��/`!�E�����XP�fTD�+&Qھ.p�8�����QR��U�SS�Z �����Ly���p`u�7���0	@>�v�R| ��E��Z Ԗ�9-�����{���j�V�&X��[�qj�O�&�9�A��c<?��D:92�,��V�d]s�a,`�J�Y@6G��i���\�zU��{�⭟�>ei��g�~x_ݼ���CUU:�{#	���P���7_�O���؞�/���	O���T66�kר�b��9턄�su�}O��Cwf��l�z<*@TP:Ks�@�����&��l��5b+���l�8]���&��
8�D��^F$AgI�k~y��t�!�L�����ے����F�cr�u�,='K���yQ%�c�tg:L�iB�Iv��Ӿ�� �X�{Y����6����ZH�����L&�و�+�Ӗ��jcN�ʒ�٦"}Ys4��l�m �\w@��=��)y�,������qO5$�t$�h��z,�\A6��T���Sr����İ�de}������Vmi52�k]�SS���s���f�"�v 1nb��L쇔�䲜�8$I� ��\&�*G�Yq�B�IvRe]�e����8�2��9Ȇ��ύ�Qɝ&( �#�	�,�)�����eKKT�-�w�1�F�a���^�T�ԍ�7�����b��&��&�,����!�^Q�'�Ql���H��V(�Z��̼��}��ֹ&�O5@�QV�����w�TJ���@I,��=4*#W��<��9�Z8S�)�T��P�ؠ��9>\H��$���x.ަ�2q�T ��-�J��U�쪰˽Ap�s$&�	Ψ�`(I=,h�F�o55�;;e�/�>a� N.���jY�W���dl���>,�˷��f�Bإ�n��&y��lN�a�����\%�5��V�����/���p�7�ŲK/{]�ה��<�N�ٶ�%��L�j�HY԰��Y��gr��g3�b75&%s�B)�LOc�Z�Q�rUQ��k���)��fH��d?Ԥ*��e�*_��G���n=�o%�{|��C/�?���e#�����-�&'j�3�ϲj�Wi/���3��L%dP	��Q�K�5a�S���
��#�'�5�1/��<���cd�)��#9�"�I��J蕫��4�ϑ'-��˕rI+܇GG���0�B��5��Eو���F.Rjb��N�an,s�C�i�X2yz.m�s�Ձ�^�C�.�UVmvJ�N�'*��r�ɛ�<-%*}D+�t����ϔn�F�����0�P'����|	��O��������q��[�������g�xC��{?��^|ޕ+HV�0�[���J���V� ;�?��IyᲝZ�4Uy<�=<'h�����Ifz�ڦ� V��k��ګ���_�ڏ~�rg�AϾ�_~�kܡ����ŕ��|�e����G{���k�>gεG����#�tw�wwɴP3��A��U�O�oEg'3�(В��A�j"NT��{��p~���F=���_b��J�Ϩ+u��E��K�p�*V����s��?£���w�����<}*�} 	HIݾ�u�N�,ieJ��9 �C$8�rF'������)������[AU>K����漬��pQqe^�sg�{N���}|�W��׿�{�tQ����"�u	O��w�YG�ڋ����|�u<��+YG����&׭�ݫ��/����.��<�9��<T��*[�%���Mt��]���I�Y%�<�Y4y��븺��k���e��QU�J�v�Q]�G"IP�H�YC����hy���A2@����:z��v*r_[�6���YQMtE��Ɍ5��( uJ��vdx	�%K���H�!���0¼�c��bIvJ��c<J�.@b�ڔ�V�Fc]�G|d���	 9�9�`�\�ʏ�#�H���>Q�xW@O�]R"���=I`Ē��j!� E�d&O���e������$F#?~�H��f�|V���Ֆ �� TBRK�J���(5;u
��U#�Y�"gj���sj����_O2�x�6�IHҕ�7N���b�d@�@�\�E�"7ߪ�#�bC~����^�����CaL�+���9Un5�2��L��%S�����<y��:�:Ga3�{�:�c�\iV��6-"Gmu�*�aI�;�L��AT���Pb;%%��d�ݧt<�A[=\Bαx*6"T�[�E$_USF�*ڱ�5����ԩt��%�A�H����[��3���
pКs}I
ď䚔T�-S%@��a��cTI0<�����g{r]��j�B+���d����H�ԄT,��^�����ƺX]���$S���y���3�MUᧈ�T7�赶��u�,�J-�-�/�D�l�����B��9 '��Q�m�~'�^Xe�܏��$Ɯ&Q���14	5��5�p�P�;%��.�t�fg,q�w�G6O�ͫ���F��(��u�|����-g��6Z��N-5��!U�d��g�-���%�H�ֆaXO��"�Q�I��J���f �-�A�o2�p>�8s�s<�&�:�Z8)���b�ܶ��/�i���u1GcN�*��U�N����md�@���8O����-�/���������
Z��9rC��#�k��}	zt1�\��$ A�$�F���U��kYP� ��`t��Sy)��!��u{�T��e�1�!��s�K: ����xϡ�fٍT��E��M�+H�+r��Ȉ�x�����É�x]P�l<ؐC(p%0�+c_�eI���ɡ�Vۈ�}=P����ru�^�O���.����3��_8����R���I�JD��#���ZX��"���/����{��$�~���T��7����G�؛t��O�����[s��7���]l~�!�<���OC}o:,�u�۠��Ԅ�|�g�����i���&Q5i%R�Qr�L�����=�w�a��G�(��bzi��Gm���y/��Xϱ�~������x��$:�����,6'Y�l��L���O(�'���t���F���ڨ�@\]�mH�jͰ��f=9HWiuԽ[���/�9�0zr��hJB���ÅW����#��/ᯮ�/���\B] 9�f�H	3hp(���)�!�$�d#������FC��p�hǐ��+%J��a<�q_����9�º��l5V���[���o�sy�V�b��%ʻ{�^1es�����?Up+G��Bibg1��dWU�#/6Y��s���t�����k�	������d�$*�� 𪀨����	)C첕ՙ�T�ʵ�Ȳ��^��JR�+�$!����Z;����N�� At�j_��2��_��8��o���RǦ.(�N��8�E���Ҵ3/�Nw�B؀5ct '�m|k����ٜgX8�z������3�:���2sВ*�N'8�pԕ�;��U�*�ZJ�̑���ę����RM��Jf�� �sC5<������t�]9bF}��j� �*��r����ޓ�>=$;�2M���8�(������]�Y�Ͳ�5ά��dJ�c@�f�I��q�cuƢrI�;U:A�v&jX���E���^�b.J:4Sұ{��l��"���aF�7gh�#؟FV���J����
k�:'��]>�$7���3e��&+�Z�����)��f���Z>G�!À�-�|�~�8����Э����O��,sr���g2�(�U�q36�/�uTG����S���#7�1�,Qnٽ�^�^�Yh2�*eDhQ�n����q���|�[��H��PfɎ�b�J��V����`�)��<��*QN�ܺm�����t9�E�u&��;G��]R���!A�P�(G���s,.�;��`uf���7�mrW1���}�*<p<@�x���|FO�*@`HP�����h	����x��@���ߥ���|��h�C��ĸ徭-�ܒ�k1�2'���f�9�&�l��kMZK\�5�*�R!@^��ț�H��f����|O9ʝ5xKgQ鬠[�bL�����1�n;�f�փ�ZGz��c?E4#���F�k/�Ui��~���}�֤;c4_Gk�)�+�3Q�G}^@��wʊ��ߕ��J�R��㣊>*?�7�▸�9o�E�cRD"w��P%c$�2�P �˿H�u8�>��E�t�.���x����]���H��=����ȍ�,.h`��3IR���bU�{7[�����ǜ`�F�'�ir��4e# �9����{�Vy�݌����T5}��C�L����d��E�4���}�g�`�ʖ�Fh;��Q��rk	�~��G7���V�x���U��e�Xn���6T S'����RI�Xf��b��^�������I�̌����	ꭝ<�;B����*��]������cٷ_~�{��^����t�7&=�	=�w�Ǳi��0#5�W���햂ǽnC�Mr�KeK�
gV�sr � ��^���������m��}�eF�j�k6Y'5ph+_͘���s �>�dv��I�JrG�$��o'��OЪ3|�k3���fG�������XI%%D6�^Y���8c./"���x�=��&��)�f�3K*�j�ǵ�:�w�Tf0<���>�u���қ��/��,�%[QU˩<ՠ4ih������&��F�e ��Υ���`�׶����xVf����B0�\��Y���d���i1@��4�Ks�0���5=ш�y3
:pP�
u{�c��1�i�f�T:S^CbgijG�5,J�ؖ���z�������s�l+E���O�}d*�0FĜ#�'�r�<�NC�`�I�����Lbϯ�L♤�k˷��ί�ɜ�1g�{��%
#}O�|��ۭAO�L�:~K;.m��Ԩ�qW��K'�k�@+Ҟ�ڗ�LP�p�8t��
�=���J��	����4��XS��פ�S�R��:5�@~q^�xNM�b7����(��m�"u��F�;�+K�j���S��C��H\�Ucúv��Q�DTJ�;��3�p�EE␤&T���ob����X �hMڍй�t��E�=|�4���ѷd�sq��=�b-'�>�U���!k��T�H�����s��Lq/v"	
�~�)�����G�^�����T�+��ꕱ5�M�	��87sz�yީA�ӛ��f����nHz@1`(p*2��X��a�Y+�S9d��l�;:�H�5��`��'���l]��P�s$у���!��HI-ZYE��Ġ��ڒobVu&�w��� ��N��IO�!~w�d x�L^@�OZ����xY��<����Π'�~�L��R;X�!�
�<�6p�?<�r���!� �r%�s�&�$pd�e�E�9h�U�2�.���$2���k��ĬJ�)��׶(�k�'����*'�,ԕ&���)e#{r�����ᢀ�N���?g�Z	hT��@2�����k�=�8�A-R^Y9ge.Ԫ`�dZٱ�24x��]���!D��Cy>��씪��(�|�iO��2���TC������c�� ��DeU���
�.?����rNq<Q��&��U^�T+�V���gO	�V�����*Z000$H�u��XI@eCi�<X+V�C�S�)'�� �����˸�ʫ��y�_m�������_�;�����-��q�x��zX���I�
�V���ِ2;��A 8�^5Ir=V�e����Q��iңswaYU�ldQ5�0e��ȅO���~��3�n�/��ho[v�;�h���8�v?y���/�$ {�Fsλ����'�s����%z*�G�v&���7z߼��r�]�[;y<�E�2�Qd��33tM�u�;h�zjp�v$�N��#,η��&�"��lxTJ��ߑϷ���v����P��{:J�$t&�V�^1/���;�$������$�h�͝Q+��4VO}����jq��'Ԋ�L2���[��?xO��L��h�|�JV����F�Z�@5���4���U^9�1ʦ��U�[�Ui
�ޫ�{����\��.k�J`ĊuzR��4O5:��8ױցhz{�Ԅ�%�b����9nQbS�?��u�T�c��b��ӊ��5�9qx�A�
6zf`UW�@��I"�l4ĘE�R�ј��%�](WT�ϣ��$�N�<���􌻩I�%w��)6�3`͋aZ�P��s��E�.t>4���0��ױ��!�zg�v
�s�X�����n6�(S�n�ۙ�E���c��4Ϣ��e�͊0fG=�qN������P(&��*���EB��Y����x|����U���zVD&)�Y�\��^���#BɈ.i��]zb~�S{��[�0���,��}[U�ה�߳��mFC�/5�xmi��i����T��wI�?���׮��ӏ>�����O��B��P��H��:��%��?�9��3�D\<L�&�-t��u�5-��r�QQ�~meg��PC�[r6a0�#�4�%�c���Ȓ�h7��O�x�¥*e0	0�'��8 xܗ�g���Ỹ����<��n/�X�8j��H0�9K@�r:"�c|��ob��)�n�W�4���Y���Y������hj������I{�s&qV̵����ڐkK91�Q��'��(�9\�irp��.�T�-�(?x�C���l(�:�66)EMdS��7�rg�UZx<��?�^�$A�{*���7ϒ�=�?����3gP�k��Pؒ@Kc#5�����fkj���\��?�?��O���3�{��z���pd{��Y1ц3��u$?<%GT�1�5TI%���\$V��]�hvs���3I�oJzyD 2`%zU�B���d&��(?�@myA�Q�Q���=����B:���] ���M���$/�|���u�X��
:�ўF���%����*AU,�ݏx}�2�Qp��F�ƫo���?��ʫ�@{���ε�?�R����TLX	Z�[���)E�7+�w�ѣ-���z%�d���i4Y`3W�hrHʕU�M
8����o��t5e5�I�\��D������˟���o�����=������k5h�{���9�.�[�c �gm��3�U�fz��d�	��2Lo�,�R��2vMuo�fs��w�$PN>g7�I�I?Ge�je�s�2~rf���q���f��kא|zXP��A�ʱĦ/|�fn��1��)�<���O�jT$�k`.���F]��s5�dt%��:�ݞt�[r�u�  ��m(-��=�:��"�1)�w@WMC���=���(���Z��nC��fF�Hέ�������£F�o.�|^V���[��/W[���]���_fM�ܽ��ieֹUgN�f��\|SVv$����C���g�Jw�Yg@�G�����U�{�JI9��8��Z�W��ټ�����T�qeI���Cġj�'��}�oy��U�M5�y�9"�t4�*�:��*��wO��;3���5�g�Ƙ������!W�m��x�ↁK
`B!��֋9q��O�h^=W��jzd�6An��Sp#3��03�&K|�k��s^�>� =��s�P�s��D�t���)�5I�\o�|����dF��9�S	�g���Á�Jպn#T�[�A�=���	F���aFmJU��ւu�}7��.&�����v��%R�r3��5Ў@�D@�Q�l���`f����wI�?����'���������_��d{��O���+U�V���T����o$��$��t
4p&�7�}���6��?+�Q=�����6z�%�DCM�t �a,�A_=�Ld��{�����)v8o�0�2����Je_��rh⺀���U�Dj�Eiӊ�cy�UP��3v�1p����l��/��>���U�Vj#l�`?j������s��JZ�I'�~�o�R�B"N�˸���1i5&Ak��J�Js���x������}�$A G�U*q�^EkaU���?|& ��s�
���T�z��>O���t�������&�w�ړ �A
���=��y	��*.^��3g�×ߛ�!;z��\���+~�	�pG�kENV�<@��,XYY�gk�4! 3v$�q��FvZQ2�i�+ژo��@R����7v�8w �KP�r��U}v&�Ԥ��y���}M�j<��>��dh�j{K�{T��!/�W�5���zq�N5�Z��υS�����5&e��:sǽ�V�"��>�Ϫ�]�P:����MT��u�4q��o�\_W����5�o=Ao_���"�ּ:k'��5t������c9p��6��Uai2�ÿ�(�����%	ѱ�^e#[�e���D�2iey�s�=z�c������0?�č;ϴMNjC(�A��y�V."�vSIM��0�`�9��G79|�jw�t�rTѵ���r�hx3f�^w�u	LLƪ̞ � h��vGhƖ�]٫�ro"�)����wZ�fs ��2����RS�I�$#���fJ�b�����C��fI��W�4L��&^=YC�4�#��X��h<)�����VfZP1�̳�j�����0�ra�u�Xe�{"v��Y�A��)⤎Rt�<����Fyj�0��3z����EW�|�G�cR����q:���o�G���A6�l��Ȍ]�(�82�ٕP.��Pb� 3�詗��;���̟N5��[Uar"k�:����6i2娫AV���z	TA����Q�`���!��9���V�y~*���uf.����貦��:���<X��kRp3.}A��3؛�IM���|�@Wt8�b�0��.�&ή[̎ωH�r��m������Z8�͙u�9��4�R`I�[��̬̽'~9���o���"TCH8��B�O_�ӝ�������}�K<��~��r�E�ɜ��jG9:��O]�YBb?j�`���$dy�K[L']�B>�p=>���.&��JΟ +��<�����������?���W����?����}�φ�~%pÓ~d����{���J�IF~�M7�!��
�V���:�$�خT�Ԇ�$���������0Q���
�?�c5ue?x[ )�9���f��J��"Q@Hyi+W��o�8M�!r�;Tj�C&%3)HF:9�������y����z�*V)�i��U!�=L�@�2�uPt8�g'Z��V;�Ε�x��1~���o�T�+_�`��j�TTrX���0�H��/ֵ����`�9��vWY-�%Km9�6��ߤS��t�e�����a&����ٹ���u1yxw>A|�k����	hЖ��}a��&gU@�踇�����i�ܭ�l�s$�=�a�;U
PX"��o�nC��<p��Ж�����/ ~�}D��i��Uȡ|���de剨v�+	K���	��6�#Y���%S��V����UU��!���;�SSMq��X��tAN�rr���B���P
9�*ˮ��7\��ZӔaa��^���ե����!p|�����x(��k/\�sW_�k �ex����Z%$V��L6���K.��CI3�� %���+�֦��^��G�W�֕g�%��+�5��7I�M��P����k�qa����w��_?�h8���._~Ͻ�������$;%I��%��Tb�a>h�@��ȇǪj��@�?��
����`;�@s��q�4Y唞ee����n�>�|K��'�lj%9�ɞ^X(_L吭M�IK����g]������ +!>��k�	�(Mx��y���Z��Uo�JZR����21�?�{����3?�Y���7g���Uew�]�j�鸛4���@��kn�@�@BH��\!I� (�D %iu�n���.�5�Su�o��<����{޵���ܦ��g[ǧ�9��{�w��3�������D�z�,�&���aT��V�Yߘy��gZ#Lt�:Y���S�,A���5�S�1ҥg܏�À��#���U�=�tT��τ�q�@p��z�
D&��,r#�$X���A���e�i%�T�x��Mʅ\�C"��/���-࿂u�7V!+��N -]�5G`��8ZL
zz�e�#-��6K�Ì7������*}+���^��8
`Dh�-�	U�"��߁�@E`c��潗F�m�v��y=6e��4%����^��uk�]MP����b���a�˺AǇ��&'�n`v��*�\�OH�=̀%+lՎ�`2�&�D0`<`�`�AE�W�bK���Z��v�� ��u�b��r>�@�������5�dc렂�L�(�P�)��ɵ$�j�X�]���<R��������t�lbK�"!pmF�04���">�<�?w?,��[J�$���^$/^����o��_�����NO�ޞ��/��C�
�*r,z��t����;�C#���𚍩��ٮ�z�\���Ya*p�m���M��p>�����w�ץ��2\C5E�ݛ�����[�Z'nُ͕ü�N���d��k���&I�"�����HF�ZN�V}��Ɨ4\R�q�ջr��MY��\����II���v�Py����p!QHЈ�HM>��]Rcg���@�*?t���X&۝��]��K�L6af5�I�bN�t`7���@�u9Y0��ƒP֮�1��.䫜2i�#&��� �k,g�����"��!Y��`]%q�%7� z�h�S{=��³��l"��s}�K~�;^d��G'U��b�L?wA�1�Q��M=�Cn3>�>ȵ�,�����e��]נ�Um�>�����	T�֤����\��ӼEn�_<{T�%��H2<&C+i��)%mä#�nO���:�%���#~|�ʸo������wv�İ,u3�9��`tn�-!'���t��Ӷ&)���~.̪���rr|)[���I��x�-��DΏOd��XƧ'��l����-�gO4����~*�p(���º%U����8���ߍ�|�I��Y�F�o<�����Q�3L4>��j�ri��K�έy��o�������֤�R�?xO����v{��Wޔo��O��~�t��� -�N���ԗ�~}~�vϜr�}a�a�h8�
���n�O�*�֘�*u��ZMYXQ�)� �^ߏ����{�'	v��|�ߔ����5����~[���T����ߐ�����ߒH�D�=G�L:��@Tg��JW��Z�!q�㚂���L��لUnt�(oZa:LH|��n���rS����j9�Sqk���m.-X�SuU� ��\��R��q>�ݼ���\�	[�W�=�+Q0Q$l�p"��=�6��[��(���=��D�Q%�����wO�9�GhXT���VK9�Dv�Id�Q,��A��> �P��䷿Ø�OR�4����}�/8�'�2c^`��o5{'��En�0�oMY�ۊd�,+��`���m�?�pQ`k�\1��f��~D��Ժ;����gs����>��'�{��q���nl�s����C�3���r9�q��������*�������D�8@_�4ʃ��^w)�W�W#?ܼ�\'0�w7ǜ[&�b����~�$`_'Ǘ�uk�ܫm�6�
vM<k�f���;]d�,t%`BG�[�b���P6^+�X��G��m�\c� �
>? ��I��������_�����?~vݘ�~XS�YMu�ڃkqpE�A ��L�a���!�X`�� ��{6���Z��R�F�ј� �bh!p�R�m��5�Ü�-�%��D7�d[�g����wg�fj��X�v�Յ��7=����ߕs�{`��!yi��Odr~��1+N^��w��A�ϓ�G~��Q����׀��o�!����D�����\���<r��(�P�����:
|��'��]}X�O��FeD��\�4�\�3X�$ɡ�h L;�{�Y}(2ֺ"�U�x�*d��W}�̃ ��.Ar���̑���z��R7�^J��jP��߽�&�D?x����Lv����sik��a)|�q�	I�
,{D���sVNQ��i��� �Ct{CN5(��.�^Ts�>��f l��|I�n�ꆹYV��{��I�����d	�WU0PҖd���\���p���S$:G��D�:�}��⚴z�1e(v�
G�.�K�8*�T�m��3p��Ȉ���V�P���R������$މ�A��P|������6v)3:�<�u�}��ڒ���y���I�U����Mrr��,7(`��'P�)e��y`z��i��{�EG��&&��I]�{_�
�m>X��ď�S��MT[=��-e�?�o�%������?�T.Y�ە��-���M����kT�1�L�'2�8��rLl>B�m������f��#Y��\�ÔA�*_�d�op�I��A�ʷ>?�,�h��4�F��$���G��{�G���X����Sy�&��^=����5��&7��U��P����<��X*VgpX���&���q�4  ���Whŀ����\.u��3KcHh�{2$1�q4�7��Q�I2����g3�$�Dr�H�T��3kI�h,�A��w���&p��u�lD%�<�GFs��)����b��:�4u#`�WN�������]p�J['st$�6+K�j�_�5O%+����"�p�P���=\��ln]�r��ŊI/,A��Q$j�y��㟱���H^	S7��MZ�Y:p�߈I_H�T����)�ȴ�v�]�1�tQ(�}�hue�ʡUcȴ�����YȬo梾¹VRpPM��i}R[Gܿ���s���dI�b���d�}� �Ty�E�>�9:r.���:�����445�@�Ðx�! B�������˥^q�F�^#��b#k���׋���@�Z`��{��`D�A�j3�$�pUy�ӈ��q�1�A?�wVc���I�/X��mЧ �������ӵI��3�\7�Ah��R���y��JNW�?��Xs��U0[,������H
~^�~4�ys6�e0V�2\�o"�"r�	hZ�&�:V����.�dWi������dTuK=T=]$����&}'%�b�.DTf#T��LCy��)��?��m=�S9]fҿy[^��;��NGry�@f�3����᝻�������D̡�Ɓ�&��?�/�{w���/w�����}�y�m)4�l롒�ٿs �_�%lg|�@�~�}9��}Y�"�@�A3�3�;h�kP�C�B�~��'�L�#0����JϬ�``a�c�fӖ�2+G;�UTK�&7����?W�b���I�֒��+��Cj	Oȵ��dz�Bb=pq��fA\ga�B��d	J�g��A��v���Y*I_��z�x)�l!�"yү=W�e�1���\YD�������Q��Hq�)���`�i��*�������҂�z��P��9c�k R�`!���΍ �4Ã�w2|�U�8�M��V٭����h�עr=yB�G.ĺ�5q��&���HFO.e��My�ͯʛ�|Cn�tW^y�"��T�A���A�^��ͩ���8�Fʌ�mH6�:�D�U�y���{��ˎS�<� ŋ��3�B�@c[��L�L���� �/��QKj��������gz�{����)�m� �>��M"�>vn�`0�b�7���0�.����$�ǐd��WbN�����l#��� .\���7v�
� ��L�\���rF�y7ӄ_ԝD��$���1v4M&S�x�s��g%��'�����f3�#�lv�ioH���,dVp�]D��g��\�玁3ǊED�K��ǿ$Qх��3�$0�<s�~&��^:}�5̥�  ���z���8c��H�5�F�Y���֎�lAL��Tث�����%���ee��7�dr�yn��r�����	��Բ��J��2vCB��!�Q�}Z��Dϧg㌼�P�V���[w��I�����F0�m�n�5Ew׏`����{+yr|"������1�wHZR7�$h���$�� ��yXҊ)�'$�d��~���?�ml��4��=	q8>�����jK����!WC\���o^��;q�D�8Yi�Oz��נ/F�7Fe�[�|�� �f*� I	�5׌�^���vp�d�kK��C\�����Wҵ���G�[u�>�T��^��4g�Z�T��Q�G 7��uX��q��?E�T���X�#��T��󿰡ER�n
�90���u(������5ap�Q����P*/�z0���17�Psp�k�!M��:)���ǯ��ER�k������[��/��\7��I�Q��2X�z1���g@�Ɉ1о
.�J?4�(��C���
�T��R����^��N+����HP5��̞��G��;��"H��r.�W_"�����Gy��ߓ'} ��zEv��ߖ0��;�T7���Uc�(�׆b��S9��ʍ�E_�M�Ύ���[r����(��nO�.���r��O�1�o?�/�`"!
����V� �_L��!�����/˭c/G'�H��>����t��X/�s�@�0��x�˨�6�jۼ���<ئ�Jڻa�vys�!�)��ZH, �j_i�B��Ar�I�t�	�@�٘j1Im���b������Ff��äR�s �٬�T#���~"�1�ae<�i�6�Ru�L�ٙ��m�w�8�@�pp���&�23����pH��=���f�|]$-HzvTP-��^�ڠ��*3z݀#�0�@V��!��2	���]5����1RA�b9Z�zK�޴��'��E]�}�6�S��ngS�;{ҽq(�����o�����C��L��,},ł��9���.{պe��V�+\%��j˂�����U��\�[�cDqJj���'��]f�<�;��p�&�R�rq�T��K�nDzݛ�"<~(?��?�'��W��M��w���`;����	>+֤ jo����\�'5<:4i�K�gRY����8�vW�[�ΥT�co@C������򕳥�740z�T��O4�� n0�|^�|�s�U����;���I����S����֖&-�MXҨ����.�دt�����D�{��;oH'	OD�;6)�5ϸ$򢚭��-w���r�{�>"r�Bs.�(�[Z�ѨUV�`���i��t���k�\�<�S�M��U���k����V�	�������㕎��q�;�|壅&^�̧�u��&AO��x��`�ʝ�%kȁx�d��y0^�gg�X��%2�NGҤ��B�k:��RӕDz����۟Q�.�X�9`������g���:,�r��HL���DO���2���Ϻ�+�-s����<�$�YY��FhE2n"³
�F(� ���T�VH&cIt�0���_9)V�% ���;c��oԡ\��I�E�"���)&QT�0��%W�� 6@ɿl/��4����6�G|��kB���T��+�?B\0[�)�؉ӄk�,�>����Ҡ�x�>���8.)\�ݒ�k��\�]��G�j����!�����ƌ����P�8�����l]���a�wb$렰��o�j�<$RO|����?taiݺ�s��ř\:���*g�w$���ER�������U'i��;z�ubA�j�4Gú
�MmZwM��{Wz�W�cU��މ]D�V�9_.({	�6r݂G��s����ʏ�����\�Z6�yЛփ'F+{�{����Hr6�d����٢4����L����� e�Alw�A�x ��3ڰ�����CZ܃���s*���>��w�����X6lŶ*c~���~$'?yO�?��b*-�s�R�`�V�>�	?�.�9|bs��K�&g?��t<���Od��A��U�H*��,���\E���^��aq�ԆD�*x�o?Ko�m�l�:R*Ot�,<B�P=��ϤM��x���ѱ(%œ�R�E#����*3pI@ĵDN�9�j*�+��X@^�K������6ojA������0���$K�o�ժ��1R�R��*����*K�Ad%`Hq�T����6�C;쐼��5xA�H��Y�VWzI�U�(��TV҅�|���+��ʺ2Ԃa�[��e6dw@�R�A �����n`�_~���4��>���}��ݕ�ԇ�6�>�������R�<�<]��-�N���'m]Z"R2�wxp(�Vk�Ϡ��	����ߎ��F�#�����(�,����dK�oܒ��&H.t���G?�g���ަ&����nr��+�^�^��9�&��X��be����ڤKϪ�8|y�.�j^�3���p��� �	��#;[���c:�d���z�F��N�B� T���'zy��[w�Ɲ���Ӡ.)0��R:z�ݮ��6�'��~q��
���&���f��O�r:�e��1�	�a�/4��$MT�U)�^Wv{ۺ���@��k��O����WzoI�����$l$ϨWDu�pKj?��-�D���̋9jx�@�K�z�G��t��Ob�-���@65a5��H��t\�7�,�2�*�kr��+�n��.u͎$�'�t�Ĳ��˓-}8�g������0%Ԥa&�<�˃I-�@��3��;�d�/ u����ّݍDφ�R��y�T��>z6��HǃR�:GW�B�)��CB���lK�ږYd,���_B�S�A��g�N����>8���Wץ���]��c?h�b2�x�ϵ�IE ?H�l[/֠���զ��y��#�:����\� ������|���[Zg�� ���0�|.�u�� �|��gD����W�����9���6�?�.$�¢����1�j>�t{�u�����Z���=�HSsb8m�yrA2&�>;>�Iy\��(j�첅�V� r�g�{:{ƹ�5!�C҄g��
� �X�0��vb�?|.��i�����$��5JQ(�h*��Z��W��")�5x�SGQX��]����t:��ji��$��< �������L�u�ϐ��l6xe�B��D�l�oW�J�@0�~4`�A{�Ys˯Y����*ƞU���L���-�����˿������~�}�-���2k�e�{�c��T����$_��u��j$~��ry.#�O����@�^B�rooG��w������H��K)�/�˄ ��	��� z�ڸ�U��V�ݘ=`R=HgC9���F��<8��r����u9�K�ɷ���
���Z�ր�ҵ�Bh~g�nJ�nh�"ʺ���[�q�Mb��TT���V<}*�?�c��ڕ����5ϥ]�# ��:,��	�	�TFl�Hnfvd� �ԥi�K�^�U9�u��N����#���BzOPe�T� ӷ �����!��B��(�j�\ީΫڈ�� ^�IK���l|v�&Mj��D6@�֍|�si�I�<�xp4I�����f��bp����τ(��5�a6&���i~p��;E;:�`��.D=����B��L�_�/�}���Ñt�>�`(Ԡ7��FiK�諚
h�W�E^����P�"$˧�1����uZlM{��b�����3Ҁ~��m���p5&og��X��4�~E��w���zS��Ǻ��z�p��5y��-��#9��X�h9H;fU.I��tb}^]��YI������n0��~�;J=��D�#C�4�؜\�㹬.&��V�۽]���~?0㡌.�r�ӏ���ώ4h��}�[/��!L��hP��K�\�o���������ا$�R��l�Աߖ�&�GG�i�:�&��`��-ʦ#y���&�+9�lh`��U�	&i-}.���^��y�c3�j �)Ѯ& ���X%I�����L�����^�έ]���IƩ�xI��x1ǽ4%$���!i;��F��O����� �v7�����@�ӇG����>�%�3Ȅ�\p�-�Ʈ~�����j����B��2X��$��1�t>o�nk�ޓ��*��2չ��������m�7uN����x�\��ř$:V��]��ё��o!'��&V���z�|!eW�Ȟ')����7��G�y���2<~.~�%U�'=������榮�N��S����hQ�`V��x-�a/�jr���<�k��-�7��b����ɽ@�p���,$���-�0Kq�ʂht�P�`p�3��iE=����n/�Ni�	r�8VW�C\랃��E�8�*@m����z݇�~Z�BG#Q�k_��R�"��k��T�aP���=��GW�b�]�*;K�Ҍ�j'�b|ۯ�, L��	�3�ۻ�l�I���w�r�@�k+��A���,�6�6��񘜴�r&�ٌc���5	�"��gI������	}u������<��_��������W��")�5y��P�!)����\��5�����f�f��;�����yf�N�N�[k�#���`�Ъ��Sׁt�j�8	�=�g�)��L%z�ml��pW�����{�')M6ZF(� ������^�{��h0���6�Ls !�b�|#�O���|�d&�ӌ�UU�f6ڲ��q��!�X��Ba��p��kâ�;r����� �U%*�Ԥ'��gO� ���HR@7�&	єB�D26�:0�	uɍ�`\��y���N ��R��2���|r
�e�i�A�nW�xZہ��R2��G?���L6��.[�R�1��s��\f�Jnm$:6���)m�k�aQZR�-36�3�c3���1Y��7�V�Q����6�6w�	�mb�S��K6~c�o�Bsn�0��X��;E��d�\�Lnt�4 �k�W��Q�jp���C�k��_<�r��2p�vV����1��4Ǻ!�� �+� �b��������`G���й��I8Y�{z���ߖ�/,�ώ��|&�(�N���J-4�gKr(R��CY�a�ipb1���� ����k�I	|�X 0hZ}��n��PZ῅Mg��L#�鳈����o�J������0��k�&+����r���m��ؒߐ���w��.�~����Ӛ�� �a��_�y=��^Xx(l̝�.͜����J�a���XjP	��D�!�1��}U��[2\jߊ�Iw7I"}�㙎�@���v4U�In�pgK.���C��J��&>�/~Y�K����{:�4�@�spO��ۧ
ԧ?��?xO������]����0=?����5:�w��_���{����e��%�ٓJ�V?msJɃ�����]���������7(%�<|$���w��>���y�p_�nj2ӓ��}з�-@%8sg���J���ܺuS?ק�����r�˟HO�?�$�X����Kr��ߒ���+�ɖ��M~8dF�M���"���F��+�\��E&����� NݾcD�9A�V���S>G����k�|l������3Y<�[��iY��i��Wߑ��ߤz�� ����L>Ryy)�xDΚ�u�lul׆z�ߏ~�}"��C���5���#�7����Вo�@!�X �?�A��LhW�M��N���0y_�P'�n"ݰ���w�8~X��b�#�j�K߼�9���pv��9�	sen8�8�3��+�#���#���-�Zu�_�X]SEq��P�N�u�*-I*<�;M�⺫q�>�~X��ߕ���%L��6V�۲_�E��|}q~*�?�H���a���']=�"��WP��`��.b��8�i��En0?H�bO��y���Bs��'��-W3���B����9�Huer�t��\��p?s�[#-Jds�_-��I���K7�`<�2��ڹ�\��Zh�{�8�Ѹ��'�	m�L8E&���JB%�z'-�R�C+���ϭ�6Ԭ�	�vHzhV����[o�7��&�/Iz��a������o�����k���ܼ��+���!Tjf��фP����H`��X��woi�?{~!�v,��T����p�ܶt#�Э�nF9�̦�*�F�96*���B���h%���"@������\$؛P�m�brn�.�)�76,U�a�z�=/�hꌛ<��4��Ԇv�d�`��,�I�KyC0�k��1V�,.�R���3\.s(��j���KQQM�tn�B�$��Vi�j�ee�2�� ���)PU���n���x�	��}&���O��)'$��p܅$4ɡp����M6�sUOJ.VK#��R� <Թ^�YP0a�N=B+�4V��D�Y�cw{S���E�Oq>&6������E+��(�3�i���c`D��rv�S~H�b(��g����Z�>�NLI���W���V�닡��d��&(>M��[I�v'H	M_bA��@2��`P���X�Yc���P�&1��_1���hM8`�I���S�M^�@ɯ��Y��R��α��s9��!�
��������y���^����L�l�z������j+�9ւI`-�G�]�ɸ�7� \�d'�dj��O-M�t�D ȋ��{U҃[���d['G�e����<;�/�<�K�S^��[�n��5x�ч���n�'m��h� Y��5M��NV��66�wdZ��ey�7����Y 2�M�b�{�R&,�S9ru.}~[�n��w�y�KL�a��"���įݢ�J��-tנ������K��oޓo�焯E�����I%����i�����ݓ�􅗜o��'}�z�t_8Zj�y&C����I3&��:��q[�����p;��|�1j!�\#
%���FE�ڔ%��V}�m�9"0gpԣ���֕F�ߧ�\��;�1��e�N�<�H�ֽ|W?�@�c[���}S�Y�$xyK���u�M��]6U}�X���d�և4?�uh ��{N��o��������#K*
YA�b�R_^H>��s��A0���S@�8�/K6h�		�!WW�<�g�a��y.x�:h������'Q��=��4�f9���R����h��V�73��As�����wX9�Jj���kr���V�^�k��x�WR����^]j���g-n�������������I��[[r��W4hO���m4f2�(.��}�#�S�٠>e9��ŗ2�0��uu.D!c�1`x�s"�Wt�"'���E������(��N�ݹ>_��_�׋�����ur~z�~��X�	�tf~?����7g[V�+\!^�t��_MxTS��r�ZZ��
�&y��$ �0ݬJj�k"�G�Р�7KЅ��[���~��z�S]�����O��G�R��潛��;�)�ޫr��KBi�L��g2}r$�dJ� lި����8���&_������Ma+���8�8V&P�t�^!v���)�ײ�,k���f�)��l�IGg�*r'	�JM��t��,�dw�J��Sx8���
���t\��U��oP�(���#��s�:=�1l�1���L�v���J�ÜDb�����2���M����R��Cq���o��5�jm�Qj�庡c#-H«�X��fnнGK�k��C������ڵ'v�h2�4���,�Y1c�1��Ō�QG)=�k��^#���g P0��� ɗpc'6���E# ���@�����qW��	���ev~$�O�'1 9�nK�w[ڻ�4�J����/Jq�!��r!ճS�<x(����F�����CqHu.4�7���U��]ۼ�7�Si�B���r�׆��i�?��`���y��O%���-������c�����������y��/����<������}~>��O�S��t��)�H$y�b����=H��H�U 3p[�z��P��D�����ܠ>��u���=����+�ےr��r���ۓK�ߖ:�g�����3y�I�Ï?�w����m�H}��͛|��Ls�9ۛߑqR�����'v�.50=�q�����d�dR��:S�ac^�=P2�t?�'pS�-�d7�����a��>�6�<�_xE�*SKY��@��5e3K<�%�Gd�a[6�OL�=�3bt�.j8븕
dN�/�L�H�S����p�.qs���q*u�s*�m�Ee��f�MJI��ճ�b>:�s��	��j&5)=�N����R:踭����,Cm1�i�:��ݲ%�WN��v�)���Q�<,���U�o��!c�2k��?�V��"�������H��!����Y�C��j]�tv
�}�� ����n0�L�tg�$��ڼZ.h��䨧󺷱E^����_��=8&�[ph.ɾWX_��~���0����ڹ�ƾ��MW������N��דY�$`��`P�*y�;�Gs�f��ɛ�4��epII��?T��/�EV�h�M����Pnߔ3��d6�Y����h��"Z"pN��v�
!.��\h2���Lƚ�ݽ{Wvv���9�T���t�[�R�������� t�}���n�-K�1x����ݏ8^	$Ť#�J�I���k5�w~��Ov�?jrZ�4ȃ!���6�Ll�Eš#>��6�)�l�x {�8uQAQȩ�@a%�	KD�8s9YT�#S�X� ��s�x�g]yz�]���Ld�X4ʗ��O��O~*��?���\V�0lk����L�zP��*�2�����~ )*,En*����KFa����g��j�����HQG����Q;�6��[�ZE��=׉�INH���Ws,� 
�b�`�q8B��@�2�>�wp�ÈƬ.T�a�W��LfI�'j�;���	x5�<Z�Ŷ�-�|k�X��C��RVxrP��X��Uw�� *��
	E ��̈���+L+H��0�x׸�����(1Ջ
w�����h�x��D\4�ˢb'�Gp��V�E��e���m0,_?cO�^�A5�1b���51X�"��x��i-]:QG$�ef$�Nܑ����!H�zLҠY�鵢R��mΤE�H�X �Ku\SУ!i~y*���DF�B�[w���+������]���ſ�)�AW�;"#8��$��<���e��J�C�^:�9�h�+�H>u}�8LG3m�����h�+|0�2R<�>�
;���7N��������B�׹��_�����<y�C��*�ǟ�
OI��}����O����s�::_���;zP���҈O�I!]���O�����$�x2��Pj \���׃}�:���%g���%~���cQ�im �����:�Mxc�9�_�+v��� �7���ސ��-i�{EdS�}g6<׀c*>�W���w�7��ݾ�����~��ip��H��'5BMJ� ��x-ݏ�?��gz��~�X�I�5�a�s��>&�]پ��&)��$�(fGr�\I��h(��G2i���`z \�Ӯ��>�`��1����칌�<�`�� H�:��&ݙL4����BǨ�[�b���fm)����%��~W����2�m�!�cɏ/e��3M�u��2��O��	x"zm;���`h�u��|��?����=vonw嵗6宎���Ϥ��ΖLu]�j�=��������t��i���kR�d�����e��&F~ܲ�x�i x!���� ��������<B�f�R�>���G�eG�px�&F�N��lnnI���y+I�ao�W�̩��zӳv쥅�yM&/e6�l<���߇7n����9�
�����v���9+`Z�jpH��þ��6���H<��&i��<��dڔcn����C?�Xa�XYG*��pU����^;��X�p2����sP����u�@w��R�'G�3��ߕ����l>�}�:'%	��Ω]�AfA
�@�n<�b>�ӳ#9?9�{���-}��~��`8�s��T���;z�iSj"�BL�8.:了'�Pg��.&��VBLqn� 3��<x�S�����:==����|����s��ET���F8D��׽���*י���1W�������A � �Y�#�-3��HƨN���	��MJ7��z����}�K��QK��e_|�HF�~����s..���\^yt,��7�փcy~!�~�~��~v-j��1~U��v�)v&�o��N��s�'�*bD.ʤ�%�1
�IGXE���X�]�㙺E���o�,�0�d�4���t8+V�h���D��kqi�!Brr����IAIÕ��l�tZ�_@�@��	b8*�����,��"$�;N+�1����@)�����GGj��iY��ptp-�J� �M� �V9�)xG����L0���G��J��ے���g,]l��t!s=d�|Ɋt˩��2���	T�ݛiM���iQ�hPY�}� ���3��ה[�	� ���/������3��z���ڠt*BlT���(y�0D%A*� �e -�2:?���Oe��J�I�ƫw������$�t��D�w�@����L�ˇ�?�H 5(���6� C&�z��:K��+b��JSP���G5��+N�<��'��;�>�k�����H�x���ɱL�=��饴$�|�<y ?�'�������-�t�`hZ�"�����p�"Qm����f:�NMJ~H*�NM�����I�x�s�ꐈSU)l�S�S��|,�?}O��H��%�w��A�=��|����p4�W^]�5PԈK^�}W�o|I�_�X�3�"ՄesS�-V�!;����O���q,��D?"3ǜ^ V��sgO?N�#ֹ��Ix:���|�X���E��Єe6��;���	�-����/� <���'�!as��w�������[�7t���W.39����������{:s3�"�:դ�+��J�gH-���Á,ON%;�`Z�])u=V1�d��S�i*=��r�A�@3��OI<4A��A�I�4�kB�/�|�y#�d��MS�GS�ʏ�����=�=f��-t�gz��ߓ[�������J<~*?��{r�ɐ{��ӑ��3���[��ӏ>�M̆��=�^�3=+�[�lw��������O���w����^�F�i,�>g$��AQ�cP�7���0ݎm0�p��D�ׯ{��IK����{:"�j?�	�l�I}��SHǴ��4+��J��Uf4�
9�UMxcv�SM���C��>��>�T�.�/Gi|��|� �e�>0~ �O��Dl�!*!��ݞ\�'��*����X���"�ɶ���7�L��pN���9B�E�#r4}D�,	[��� �j'�]S��2(�L��M f�I�����LI���Ij*tՔk���:������oI1�L������戩���Ku�k%GG'2��l<|���J��Y�� �̠���y�*���cR�b@9�t$$[��$�ן�����+����?�����v��"u�QÄ���#͊���5�8���;Ņ��=;a̜)����z���:�R��6�� �b��J�݁� cP	��r"�<����Y2�KK�-�Mu#8���'�'K�=� ����.���U�7<����Q����n��`�8r�a4�E��5��u ���{�k�r���qV���s��`t������\ɭ��%dW��&��qn��$~�BV�q����Ԡg2�iT�{Y �2z�2�-wO�i�B]��:`C��@=
�vjU8Ob�U�-���p�V#4��Y���_m
XHAXF H:��-�ۥf3렄�u_��$�).� ���P]n9�ϙ�`cF������b��G��Rf���K���8#�4��)�*W�D��ꨁi�X3)#T��J+��=�V�˃���H�W��葔ۮM⮚,d|�LΟ=���>���=�<�!�/�*�o��@#��&D#�+c�jy4�2�\��j���F
�\��`�$� !\��L��.[�^#Gl���_ڌL��k�N3���\>~.O���'p�D��f%@����AL��;>�1�&l+Υ��bV��ZG�$>`�Q��V?	r� ����	c*� s�-�%ge���/ޗo���+��l�n˷���.��H���)����[�h���_�m����Ko�D���I�G(AfK�hp��-�����ߗ��#�&�t�	<#�c��?���hǲ���^�#� �_4�>3U&�.�'�.����5��u�	��Tf�����s�:ng����������;���m��>�!ϩ�Mφ��翐����r��}����vd�&k�e+�ȡ�7���E��,t�������M�/e:�H�>�q-��X�'2����@Âf��i��j.��C��;��7u�rKl�͟���j�_J�-�^$u���Da<��ݞl����ޕ\�g��H'C�;�s�+�s�ˡ���CMG@��'�k��*��`|<���焨�Py ��3���"�s�(��������Jhh�@�f�s���ׯ49@ ����+_�����ے꽟N2��tu�����ѵ���j��= 	�;'Y�p�Ea��7oI�ߡD����>��GGܳ�=��Gv��PS܉��UFSB�(����K�M�Y�{k�"�A[p_����9��%/^#Z�n��1௸��Ú�Y%7���<sx��+�m4����%F��PkW�å@���ǈ�sK���b�n-������3Mf�T�m���	{�`e1�Y������;���G�?�15 
��~8�g�!��c��eI��\�ґ�����p���~��^$/^>���o�_�;�o��|��ͭ�m:�¨
���״�U��U�&5u{oCN6)�z�IƢ`�=��b�*ci�@+)�́4\�L�� ���3��F%�L-��S9]�a�$�R��,өDS*M����JW�i���iD��}%o�*���䣭gU��*�!x�+��k��f�Z��9>��N�;j�����Y!��{���
v�&T7c�߆Z����4�o$^��qlN��]�Z(X8��܆��P6�QP��݌�ܿD���n�q�P����V��XH��\ 
�e�aL+BЖ��:�P�>�@:X�a
�N�}�3+�a��g,wŀ�[1Az���Ul�Q7� ��ԠgR-���kE�@L��M���:�]��)_ ^���#1�yO� TC���[;<o<�tqs�w��kU.����Xx���׆�6�}�Ȋ�A�J�W����c��'R�>���S�����ޮl���?�r|�N�9jZ���z���ɋ������V�#+�k��~����"P}GW�05�JD���94	Ȅ�ѭ����KaP�&;�+'h�����$P�128
�Ҝ�ێw��H�uߕ�!�cj|�OE�s3�=&4i�9�2�3�R�L�AXz���g���?�0�H��;��a5��A���=�zx)���P��Հ���Ho�8pT�)9[8�0ǝ�MӉá���eS�wC`D����nח��-;���b&���$�{��#��%�	Q%)��E��[J�S��K�3�����J�	�N�-۽-i�F����	5�<�NOdS;z�� ���#΍()��׼��e������@��Q$�/���jb�j�4e�_ÀISE)j��[�t�P��۲��/�m] ���\�C�0�H�F2����0v�YhR��	"T�6��/J1c���;
MR㹮k��RM�3�/��vW
�I�1>���Ҝ���RJ�;J��y���NAV�si�N+�>�����pvD��.��4t:�X�����u��~4\H�ޔVԦ��d2��_qPt1R�Sis{<M�t�Yh����߁��Z@���C��m�D�sY7}��tOg�T���? ���9B�_�Ce��w�Ʈxe-;;��{�],Um	����:�`�-t]�����V:�+�qӡ��F��5t�mN��E�k �2>0�svL^,~"�9Y�<BP<�5n@"`c���ZeP*�_6�N�#{��zN�rrq��
�ٌ7�F��A< �j s��Dু}��x�8y֠It@LNb��Ann�W���ER��������?���?{�Ï����(;�rB2!���L�2�u#7����[�Ml�{k��53�U�����bT��-�1���<�Y�Y�fγ�̡�e���ݓ�v�� i���dt��ĸ\RSв�r�Ю#T#0�G����BN��U��u��\&E��o���H��_1ΔsI���E��gm�k�f�i�S��:W?smsw���$ٌ�X28B��+����~i�3�nj+��k��<k��g��͗v��)+�# �:?��,��ݞ��9����PL�ΐ�+T i�s�6�����}u5�J�����34�q��6��_�0��DބU�@�ͩnFHҪ�����;t�ё��{��T��B��>���k`��2���gp'@b�q��?& x���(�A]"����J��&���JG$_��UZѼe��B�	V�;gk/!$�<�y c����#���?`=���=�3����3y��X���л����/�J�Olq�E�����r*U	z��$b��H����7~�X&;�@�c' 0gZ��d��Rh���J�dDܚA������=����fW�9��mT����
S��ۯ���5
�BX����V�S:�F�G���ޓ�d@y;^C����p*�ም��2���G2:9���/;�l@2={P��09/��(@h^�z���/x�H/_���lh�Zɹ��|^T�����a�ѽL�9L�����@S���`5�C�:��`�3*�T�$�d��-��N|xk,d����]JW�����JjBE�68f�Zp��u|�w�(�F�:F��?��p�/��h�����[@h*�[Ҏ�=$5[���3؛o�
!|	6��>�ָ�4$�"��H3�	?�nW6�hп��&Tw�v�eֆ�OES7MtD���ڽ#[x_]��\�OH[��` o���b�k�F� ��Z��v�sxU�l$���}�_i�%�C�>�%�pkG�`2�Jt�If���t%�{���3�/��:��~k��+q���wa�=�}ao¾YLT������=�g�k���3_����I�&�3}?
sH���bB��&����yq<7r��3�X ��a��U�M��6��Fi�@�s75n�#�1p*t\���VY��=��7J�����yׅ%V��\gAL�1�ifF����>�DK` b5��X�(8���1L�K���39~~D�u$W���%�E�\�}+��Ο��p΢+o�w�]�EF[���������=�*R %S���/}&�WT/��������_����Wu}l�۱�@뽄������m �t��J��v�_�v�_I�z�X;����`��͖ܶ�	�~��A�Y��xH/n��͏� �$(�z��H\#*���+�C���GP�UjN�Pd�4�Euƚ�N��I�Ԭ*�~m�μ����7��ϧ�0\�&��1_\+��;����N��r՜�˲171r��x=�T:z(���#p�ul>�nW�Vʀ}^Z��H�:������c��M:������ܧ㕩��n�C3�*��P0�AU�wD��	� 1`@��ц����O��d�t�S�"����
�H�c�X��rA���Kr��sUar��рb��ԛo� u�]�y�Z6�F��q����2�kp��y���5D|t0�g� ���N͉Fd^�*�.�v$�Z�<쉆$䃣Q�_�&&s���Q�浟~�롾�U�S&��)H��~�{!��H��Ӿ�G���X씂�
TG<sT�\{
2�ZY�TAFv�L�C��d�AVFE��p5|+�Қ-���9�������U��:!��N�r�vJ�K���.j$�lYsm���Tr����58�ub���ah�� ��숭�d���J/��ⶤQjkܫNO��妤�j6q�t/׵��g����*�v�+�=���&M�V��#��$��_�f�-�+�ww<V�àcT3ˈP:�z��
�Y�s
8d�2���c���ٗ^�#Ǆ}�$B������z���2�j��[B�4jK/ٔi
WH�jr�k0�4� kW�DM�WU(S]�+�ذ�#�� a7��\�~y��j&��&
��>;L+MnE#�GX�\2v�r��N*sM�ۋR�{��W�q�����˷���q�{a"C}����]�$�ض}�#�͂L��j!��sه�yW��^O��[�<�%;յ�NcA��z+�>ň�tI����8��0A �����I�BYhpqI����k�T��ggue�����2�K7%��\����>�9�e�w����@�����A<] �"[^cX��S�����%��l�`V��|)��^�� Ҕ�إ�M�v�8��w5�~�I��Zm�}��c�:d�a<�hb��L�
���x̂�
�]g�����%�%�K@�t<�a� =zrr����ܐ��r[����1)� �96\Gpæ�	�40_
ke�,T� ݍ߫!�Ε \1���b�I�_��?���m�o����f��F�P pv� J?l{q�L k���J:u��sm��a����m�X��������W���iz�h�<IG:���;���8W��a�k烫�"+���a�LO�P�����>ŦhB��O��bTW�Ⱦ�u%S��߹`�I�!���7\��~֐�U^�ѹл"Uɵ�]e� #���=��J
��Ó��c��aUZ*b�����.�4%!�Rȋ�Jѹ��b]!}�z03-���
q�hN�=���
r֦��A�j����$9�A�8�g��T��y΂�܄�H��@R\~V�w� ���q��B�z�51��F<���Y���>�*�q��UF@n4�L�U�qƗC�z}��t"ٚ�K-m����`D��Az�:u.ޞ���;�Up�P�͟����k
�tƄ�h�r�����YM�Ř$�I�bj��G�H,�LP�����M��7]�DrV���)�44-����̣��$�0/���g�q�J��K2<jo�.�;\���)����3
���͍~�7 X�f��F���#< �6t���lm������*��_%daqA����*3,��(UPAlscG�iP�����<���;R��CI�������ljp�a2��v��k(Y,�?��p�>�R��.+����
>7ȵ9?�$�Kt�
T�A�L��4�oCBu.�Z���fP��J���Fy��:?u�+��Lu�q�e�Nȋ��?S�
�����-&�t@����Z׭�nGg+���`^j2��D�%����������'����KwsK��</��H�jz�6m���,)��1��"˩E2P�Q�Lc�j����k��Bյ��0�K�,N�4i>�K5vߖ�w���2���n�]��9��'�U�b��s:�t�X�aG?7���̇����3y�oV�**��5��Ȗ��o��)�U��N���x]x�K}����.T�YC�M5��L�:���^^�#�t�u�Y'����u̷4HŎ��g4[�L��F�hY��\�=�RX��JA�Ir�-�KnQ�U����(� ��נ��-�/�LG���Ը߱��!uv�y���
.,*y/�I��[�9�W� @𿊭W;|r�b�}���ލ���C����L�5��zXj��p��RE�쒅!Bmu�A�	��;[�L�W��u�Q`�x�v��l�b�5P�bnŽ?��+?ɬ��}�d�2�^�g�2�q#^�
�^$_�i����8 �1ی&q�`moT��YB��������C�8�=Ylݹ��4p)*�p��&	a
���Z�p�57��A�2HPa6�Uga_�Ae7ѝ]��>����n��!�A�����-��c���RO��A���'O�<{.�.�`����A$e7]�7A���A�Մ���޵j��y�߯�"�d����͸��Ѯ���J��1����Q#�v�0Tt�n6bln$�4�����8��Y1��Q��|�K��IR��Ƥ�%���� !�y�N E$L�c�@6�]�-����-r�-��E�Wx .�"A˪K�^u�C��2���&x��Xz�S�$q��&� c^i��\з ���~F��j�׎�y:��� ��C1%�����Je���("I���d��: ��A&0�hC�	��hKf^4�2�k�j mv}Ɖ>�$��"L��A�_;���[���X((�y ��O\������c��c��kГ�Z�{	��V�,p����04�2BgO���y��ZP#i���S9��*QKB؜s6����Cr����|T��"�T��	�Z4Q����d�`VP)k��5�(&5;�ػ��T;(����`��;���+�zvz��g���3���x"+�f�L6nޖ@��:�qD�OYꆠ�A��T$Cw����5;EH�j}F	�.<�	�&�K�~p��޶lkB�xy�<!wb�Oo6��D�갌5����6c.ie�B���S���~,����ir>+�ڗ:/�$h��j,Ê#�0{QK65)�w��o5�P]?I�+E&cy��f�IB�c�;t ��IT��~��H�
l�j�������>&+ݧQ��ڞb?�;���M�5��up`�6�ڔqSbM�6v6e#
��#��Fñ��Ne����ݗ��0m�]��]�\+��s}��ٻ}�{X�*��2==�r2��y{�¯�H���0K��&TVC�#�BL���R̍j���2�$����Q�`2ҹq.ޮI�sz��<�c�����tCn���C}AȨ���s�U�&lS��S9��EѬo�Q&+]�:���k�~��ŦG13�7���EW&����38�B�5pN�LBrB'	�����lw�5/�Y��1t���3qv�ˊ�)́(�m����6����k'�A#O�G�<ok+0�z��zt O󤡟��\��٦�Î4�������Q�з�.�a��"�/!��{Q��.�NG���u�H
^����6�v{6����9q�PT	"���3�BU��'0�,�~�;b1^l�!��B���L|9�ȵ��ܑ�jӴ��`X��Q��� Gz no���9�Df��$N�rm8Ժ���|��rKz�����y`�=]�p.fP�#؅�O�����A�ɷ���~���C�ip�נ2������;<���*M�:C��kTV$q^e$kz3�,���~��gi��b���!9�^�X�+����h��kD���|>�R/,	�B���ȱP�����Z�a@t�/fDƳO7���f��vsU�@��$#nI$eA��]�(�$ز�OXR�C��2��C��X���g���h3z&��Ș�R��1�A�s�n�-�M�

����D	ɥ�\�����D��
wբ�Γ�R2��4�Xd�Y�3��/��`��
�G7�|<P�A�A2��i�̈́c:[X�^O�%+�G�JSv	pY����4�q8�@x��D5����{��s+Mh=����Z���P��>�jYL���?��:��'!,$g�<xԣu).�1�7\�/�0��j>�N�c�]Dhs��Ԅoݤl��}�:�<_p(���P�H��V�1��.Z+@���ސ�Ҙ��� �� $+̅��GTl��� 恄`?���z)���O5���;�������7�%m]K}#�Ν�}���<?z��분�R��Cfl$�C��L��wxgߩ�>����?��^�ʾ{C���>�к'�{�k�ZP�$� $�v�5Cq!]�n�C�S�A�|������ޛmI�ׁv'�>{�9EΕUY�� H� 6�Rw��������?�_���EKK%��HPԘY9O���~��m{۹�Q (J��Vkq����p�ù���f�m��+������z&tdV�V��H	���@�G�ZR�:��|y6�2�{{r�;�޽�����j!|�� ����>hi�
�Xs d��PW/ʖΧ]����Qף�[N_=��_Zԝ��'@�S��N��^���X�?|D_u(3}��[7���(��]Z"�+���D*=�Y������ܯ��`�%=}�`2�����|x��/�#y��g���똎�T����ݑ�?�+�F���8:���%W#U.,]#�bݓ����p�B~�Ƒ:o�NO9�s)���	�|�F�#��"0��o��<�EU53����8��i@?� ��pN�����Q=$��Y�g�����K�+Qg$mK4Mt2�ltؤ�e������^1c�5���y��^泖�T(�;��,�ԅ�.�D���Zs1zƢ,+Gs�cx.KA�QX�1�"�x4�dq?jN<���(�ކ�Xm�}�AI����}�h[�U�,���
S�C�dK�\��~R�/�^�x#n�M�%R�	�-<$D~���StD�Bo5�������a�n3�7���B��m�7JW��~��)��ʂ2V#���j��K+�q��#�ܴ��5�BM�pq(�Źb
|Ki=����"T�Sn��X�P��G�P%T3�ݖ}��:��e��WpB�n��A������|�����]�xl�fЀ& ��s,�$ѕ���u�<������'�:��bj��r ��=��(�.�=��7�*��3co��uq0�a��^���6����$�p^��VjO����W9FdUt��
I�cY� ��$F��{��A�(�ҹ�M��P�q��d<�[�	6z�v��]+z$�#}Fz��R�e��S0�qX1J��h�U��n����KK�ր��QT��D���S�EtM��@|S�h=%.KG�,���^|!M�(g��0:�"���@�}��c�� j��Y����Lt��qxA�(ЀL�q��u�V�C�+�E�D�i��t�l3*��'�M0��/��#p�etҔD&��.$�+�|�>���p<k>�SI��g�Қ�xYx܄m����u�bQq�����(j��z�)����7����mPD�:�]�ԑg����8i=���~K�#�H7[�,f�
u �!aK��?��w�ZD~��)��i��	<۰�).*��� �?��s
 5G��*��r�����]J�"�Y9.+}�`G���=	;z�z�-4�Bqw�=`��N%<>P`7�;?�}imms��^ȫ�Ϥ��!bt�7��ŧ 7U����s9{s�z��67�m=Ƶ���sqK.{��`�>=�PV��T�g��>�c���oR��zo���9�rg#������Wr|r(S%$0Ӹt�Qs�'�v#���X�AB~�ܐ��/����S�z�C�`��S� g? (���YO�3��)��J�$4"lt�yV��zz�Z~���Z�^?��d����U,����F����sEs�ʛJoS.�������g�y�;:��
�����m�|���n}��@u0,���#ۘ? ��|�'D�I��I%���ȁ�	[�i����[��凳�u���k-��疑b�Յ��ѾIM�q�QERK�$)]&��U��Y:g1y+�K2��2��v.]͟�r�;�(l� D��b�-V�=go{.� ��(l�Mǹkt�G#5J����h��-j�J�t-rG��-��n����e�*����`��U�Q���Z�G7E�Ap2;״_:�Q�cj��X����qO%]A�9>����X`��jgAɃ]�'��߬���!�z
`d��j�y����HR+�&M�rd!
ƵZfWJ��ϗ� B+��]�Ӛ���6l�\����w�S(����\S�'��ϼ�5���L�z��)��j��o�U�M�˃��*�d�"�y��tE~q���n�Z�m8T�('�h��5�G���a�BU��	���Z�F
 S4$R`�FCt<�WǠJ2z�\v�}.�ᦜ6cYv:ҽxY6._a�Y�b��R,i��]� Q[�fK��+,��S*WS��@�7	D���yg��n�̍��'�WF�*��v�f,\�����~�v
����R���:ܥY�DW��'�7���*�f3P&Z�0�$������#��T��X�8�L7��k��QDk��i�!տ����y-�RG~K��A�V�ɔ��X�~�M�Q�t1L�yn2�yn��<'��3�S�K��׬�Hs(]1@'2�en��(d%�ǘ@V�h������L���T7�-d< <H%
nG
�Х�
Ȱ��P�7��j�塂�h&瀃�"�8bA�DK��I�nVל�KJ,�+s��q�BF�P�9� +�Zl�� �uÚϬ@�{�ܠl*�2յ6��Lm#jՊL��+��\u-�>�T_o�k\��hĔ��>���똕h�ԕE��7�e�@T��`@:���+��~$��Ee�b����{P�smF�s�?�Ҫ�z}易�����VG�	�o n Eqe)u�����������E7�A��9錼��c ���١T���F_vw6D�ԭ�ܺ$oߺh�A�V�����K� ��H�k�b<%��������P��(��"�&�K����W��'��c�{%�}=ϟ��\����p#��Ӊ0�
j\e}��|.�8����
�]::;l��ʛ�L����o$��)H�q�]��z�_L��`֬TT*i_Ѡ�w�l޾-r�<u���)b��53��5�pNAn�q"u1�p�f�jH�W��%�'m9U��й������E��>����*��3dXu|�}^�}z��M��T��g������U��zSq�sֵA�뱁���[�od���s�p��T�̧�
�p��eh���[��┦�_��
�wxΉP[��R�8�NW���oF�A�*�̠��l5�A-a)F�3`�M�w����ߋ��˂U�~dR�$����t���C�_?n�!�B��λY�M�+���G���-P�=�u��<��a�?b �4b�,��3a
$B�-�jE���d#@唃@3��5^��F����(�?C�n� {Q�S^P�M�o�(�=z����(>�����f� z5eP_+Iĳ�M��C=9��:!vw�$�V���A�f!�
:����g���>��z�Lo�4��AZ����L��^�u_�!���V�u澁�F��Q�ܨ'H�W.&D(+�9���
��0f+Y0�ѬV���Rlt,��}S`0
�G�:�ꌐ��>(<~�X�
��2���1w �·.�A'�W����ѱ����Pr��|�]y�G?���R.G��/����q����?cT/��{��}�5�ҨB��\ N�[��`�^,J����gj
c�
��D�*�@�8p�z߬:K��կ�0�Lù�-�r��;�'�Nk8Cmi1�neEYF�ᨘ���2��J����T۴ϊ)�%AB��jN ߷��*zV0��z�aږ��Zƽ�3��@�8��tu�`��ȉ:�Dtq��|���f��/���8��Q����G��qD�YJ���ʳ�m!�d�����e�T�:&��m��6��C������:�93=�43'	�Yi�Tqb��B�<Ҁ͏p�5O�@*ݥ�Q ��xZ�@�i`y4Du�M(�@��| ��ru ��N��@��Z3s�m	��2Q�U�X@�ϯ�H�:	�%:�6_�h���z�UY��y͗2��c�C��+��%��ޑ�֖�ͦ�������~�WB���L�s:�%��oՇ��׿��ӏ����Y�Ʋ��c�ltQrJ�Ћ��%=�B�t�b圗�m���,�X��W�.+G���j͈�I1�(]�b@7��t�ģ�O޼�o��	\�peT/ʶB�SЏ4&�]=�eokO^�6$J��%�ҕ!�7੣��c�R�N�kC�c]!+�s�H,�(�({�n*�B�UFE,^�	��-v�����_J���+�IMcs�e&��D�K��"���t"hh��b�V�|P�\襳7<=���@Uф�9�.�*��sL?�3���~�R��yNs��o�Zu���Y.f���u�� �0�u�`�c?J沭v'��:�h87�&}CDy�/�
o�����C[G��P6$��,��TE �i@%�#R�|Fv�߱70'�{�X�2�����>('�~��F�z����@�6�Ue��1\ì����r%��="��!��I��/��HSf��=��哲�j
�T��\�������1ĳN;i���f�ϱn����f-����f�F<�Lu���x6w��țp���Ìi`����>w��т6�;C۲��=_��X��'p����7U�7�L:�bΝ6J���K�e봐��
�����af(}�m +S��pA�v��T� G]DlL
\��d��ڗ�a��/(�a>A`�̷I��L��}0d����q���q��a�:�Wh����WU}����烝������b�N_��F,h���qر�xlD�Q�+E� �ŋ�i���^^:UK��:���Ĥ\�Ŏ��r	)���m0�(t>E�K�-2)�Ap\G�g�����t�?8�D�����x+��q�2�x��ӯ���~(�:T��f�E��C�I!����v�����޺3��U[7]�bE&���t�<n��s�q�)\�Y�mi=W �
�<W�]Xd�6{�hEn�xu���yuѓ��J�j�^zN�M
 +U�t��X��e�0?�� h�h~3<���w�|	3������� O7/5�@���A7��p��q��>�^�`璂��w6e��#��Ҋ�@Q`~r��e"��-���+c�o:���@��)�a�ѩ�NN��.�;�nn��7H�v;���>��뗲@��unwz=���}�ۿ&�~_���k������2\�em�3�o�+��ܥ��9�K*�,#��}%��I�#弔���r��-��
��Bwt�Z�=���H�z��/ɍ�(�n�&�g>K	���X|�����Sy�f��!;�����#�Wo�B�ĘNA�1N�%;;�����`)�����ɍ�|�Hw�z}�C��gr|�k�?��x"��m��$�ɟI��U�-
]c�����/���{<�B'bskS~�?��\�vSb�! �(��|!/��B���x�:���lܸ%����e��{갴���?;�����ʳ�~Ɉ>
����}��}u�P�����?7��h � �gR�#pxtd.�jYC���T����Jƿ��L�c�Q>us�.^���ߕ�ͻ2��O�J^>�O�}������L}����k�t�?�3��X.���\��xЗ��egK�G2���e2�lz�׬@��c�<bq{�r��E�A�BsGF��f$h��SgB��
��:��閙�o���0� ������&� n�����x��@�<}*��:<j{ΏN�V��֕Tb�d�P-G\��ц*�U�S��,헅��� �CI��%H�ff&�^��6�Fg������t+n�g�����2S�i�Q���7����ʝ3P�GW������?�4�I��� 
�Aς�RZG�uC����T��E�ݨg��:�_��i,�i��x>k�Z2�#�`�
�K��/g�8E������z	���A}�Р���ԐDA<����+X�euj�|�"5����!>���������e��im�I��/2�p�Q'��v�(�m�,���:�o���!����f��(��� �J�X�T�q��9(���� �@0��(XL���~�VX,M��fS������;�9��5�U;�u� �H��������e��g6��d��Ez��&��Vѳ@]P��j���/���l*Ij�g��	t��jp�ԑ��Ҥ��B-�.�m��L��:��,�D���ަ\��#�Ł�o��n��-Z��`�⯯��wN�?�WUհ�|�_/|׿�d?�LRf�_`x��J�c��j4�������?��2I�V����Rc�Q�a���)uAE���;��?��?����߂���bE�!<\s����6�ǂ�;uu�Q�xꕣ���XXsh��`�w
���de��wJD+z�y��K�":� 9���s"��,����̓&�lE��RZ;[r�{�'���Gҿr�`QF��d"���"�(Ž0ll]|!�!XZgH�e�A���7�]I���rd}/��?���pz���'!X��*�UG�Y{����V�^Y}�;e7:5��[}#LDҍ}E��Z����A�D7�$۞Q�$�es��|�G?�����m�����Xƿ���T�����'��ɻ������Fӎt�fg��˯�o�M� Zu���?����P�{
d�3�XQS]�l.��M�;D��>���D��+X����r�Lئ���ɵ;�������ܖL4��R�z�?���V���גǒ��y�����?�����;)F�ݩ�.ɧ��8b=覱�#;�@��S�_ m`�#z�My8�T7!���1xO��;��:'/�1~�L��)=�wO~�/���y�D׷ǹ�y�����Ci���$!;��9<�cO7����T�|��n���3ٿ�=Y8�����@?��s���ɋ7����t�oܹ!��)h�f	:�1[��tw��W_,�ç��ؗ��wձ�d�i�����lJ��d��Kjxc��._����d��]r���t�m?�Z�ԡ{��L�~�cQȆ�����@.����ٖ�_��OOe��3��=�t�N�)⺥��*k)�}�̙_D\!��s#S��%7mp]����:����&Ot�.A�C[��7[��u�]i�m�]ؗɛ�r���������εr���e��M�Z]�{2�lsF���� 
���w6:�w�?(�E�QC�RS�b�Ѐ,p�q�QO��n�s���Ҋév� s�L�J���ѨZ�T�:
�)�	���M���!�קz�#u��h���хZ��
m���dP�*�/#�,[S�@�]-�I�r�2ځ�>n=W���A�Z�CԦ�v��}.�W`��L�#��7�d)�k���&K�^)�@U,�*���w�v�J\k��سGFeϠ��!:��ɜ��^��������StY����M �ҫ�M~��9��
Z�>��p6��uMf��QNS*]1��Z��^K�V(bG?'GZ.�!�Xǀ�t��������J�zL�/5҆�}�#K��d}�CЋ��s=�X�}K���3���YS �a-ᅶ�B�� �9x���:$�����Xn��r�j�!R��� ��5 mk��s�We�!J"JSm�`����s�+�:��L����X�������T�����\~��A5�<5�N��	jN�	G���p��p���%ܣ�Yƀ�X�iĠ1A�u�Ptc͍5Fc?��4�^a��qXb~�3�sDC�9�H�\���d��M���f�lD�im��Ύ�`(���������^�x���ˡ��~J��A�9r��_��:�3��|{��p�vM�p�[�������-�u�T�D���Z���ҟS�ς0��/J��f�W�W�i�ʰ���+,�N������P�Q� 5x(�+O΋��6u=����曞��V�%��g<�tO��B)]ݬt��5+E$�%��
B/��Zfy�:=>�����G}�Ŧ���8�ɸA���Ld^+"��@�4�RM]\��xD���R
D�f"}'�Y�9c칈�J�6(
, �\A/���Q��R, ���gMQ��<2�\��l]�,;�/��ȝ��D��{_�����a˥��#��]�O�&d-tsiS� �96K�_���yX�]K��ڢ��b���֫��"�4ڜb����>[��`Ps<T����ǩ\��g��[�����%���9ϭ�n�g�2�QA�5�lDtJj�@ؓ�|������3e`����S9�����KI�)���ͷ�?�S�����o�G�D7�^G�ݯ>�S�GP���X;
o���w�͚O"=�mb�Y�y*�:��R��5�B�<�J^�^v�k�si)`lݸ*���O$ؿ�M�aXLJ����|���3(R_�;�}���ݷm��i��Ғ�n�LߋB�P7�\������vc�7Kc>���M9{�|�v��ۖ��<ܻ(ݠ0'B����J���ы�,�E��F���vGZ�-F	��x��_�5�<]�����[zo���P["�<�L�X�g����r\�\�2�q���Ffb�픒�|��K�s�{�L�z���������B�В��	�:�.����4s��S�nlJ���$_H?ֹ2��FW���v>5Q��IsS�=_r��1���E��ED±N+V�(�dT�|'Dtҽp"f�|��u)�u��Ki���p�*"����"%XJ�L���X��2�c� $;U����q��6�k��.�o���Ӆ��O��kI�A@�r9�(L
�^e�� .�� �_9u��T�rk��gF���d�d���x!�D���.oHow�=Ifmp{���A�����܁�jj��u}S9��Y�Ud|k�TPF@���L��L]�-�Vw�f5
QӅ~�cQ��siW��\�n���v��qk�MGƬt�u9ΐŕ�7�9�v]��m��@�cNi���;3��>f��o�PȚ-���1eL��{�\�-��u�۲<���%�ٌ������u��F#��z���"`�P�#����l��V,:7�������+Q	F�]��T��OP��* �Ԁ���gc C� BE�T�!���\����'$c���t=߾a�A�����[Ka���Ův!�s��KQ3� WW�3�h;��Tx��)���/.Y����f;d���9S�y��i(1��(6��q^ga*�Y�c���nWZ����DQ� ��5u��TńY���C�V]���bL!�,��H�*ԑ�Z�O��J���M�����ڐ���%�t7Rs��d^p�QO�7�A�h�3��m��{墄����q�pQJ��L���w�H��m��Ň���봒���\�K�@���V(Z���(��jC���m�X״-���j�,˪y��?����{��NAUvG�r7���_=�f����t��t�.M���&��r�^Y�{��Oa�B�)�����e��*��J�^Y�O��T8�9�K,2v�#�]���c���ܓ V�@V���;�Ր�5����w�ua���@\�:��Q����ޫ\�(�R�1Vl������K�1�|#����5j
��g������B�f���~om� �`�Q삉���(�i�&�H�>�.�F<���<�"ک�|:���#.$��І�rm�9�Ԉ5����#B��XT���d$�̲�YW��.�a���*[ �<4�PQ�^_ҳ5ǖ*�9��j�В��k���O~,�?�����i��T�`L���oK��\�>
gc�����i��*�=��a�׹���ZGTjwMd���_ߣ�'�R�gg�Bi�C�Je��?�����e�:�s>,���C���:J=B��V[�V7`\W�S�ru
2��@�}�ʐEx�����ʍ}ٽvEA�I�q��M���-��u�l�"p��~W���'$�0F,m�ڤ��z-)Z�,t>�P@��,Ԁ혛�OCm����[@Vt0J��On,�Dk2oc{Ӹ�
��:g�X��"
�ZV$[�u�m�[j���2Ƴ�c9����;^�\������hz�`iaqX�fl�bE��f �~�����ڍe
�#��V9"IySmz����T6�m9^�dK��Ld
V�(󅌫Df(�n@I#�Q:�a5����$x9���H�O����D��B�
�^�xx�_�=�V�:.����B7��~�xz&��Pz=ݤԁf��%_����~��Q�ɜUH�<��C=Q`��3u
2]�eJG
�<��3Jq4A@BU�9�B��`Qu��\T�I�����{a���Zs�kǺ�����9��"P�tC�t�l<]�,o�zۈth��se뢼�:2U��o��Fv9� ��N�	j��Bᤠ�~j������z(��f
�b�F'eK�"v�E_�'pD�����Pͦ�� g�)��$���d����P����������-	��Y	��6��
��8���]�;�z ��(�m�N*Zx_��R|>��L��KF�g���{��|��H�%�~K[�Q�]u�[���ƔY�A�ׁZ�n�W��f��hpe�t6�2K�SQ��BF>�T�,���[YMT�����Z��Tiv�/�8+��:.[H�O��6\]���^eR��@� ԉ�i}�3P��̆ods�{jV�h��=v$���R���g��m������ͷ(׉-}Y��'쪎h�l�P�#�U����+�;ȍ� ���u������{>y�D�jQ����_�9�)k�Ҧs���1^Zy����!O��y�ڊ��1�����u�e�5$�A��\(f��!~�a�Y�'JF�\�4]�e�]M>�ef�G�נ��ْML�߽�=fs{GF�D�L�B1��q��{�1|���9vl����zM(-����b=���	����s	7T88���ܾ&���n�]�����F'����ߍ;�[��s�G~z;P��̂f�}��_A	����=Ӌ�wA,W��E��4�{�����eQ=�Ng�����/���_����t
����0�������^�GeQ�ȫ|�(�.ݜ�	-�'�+:���M~=��+KVqZ���v `j�����Ჰ���r
�YZ�߱)��>�`�޶�4���s �[���%��C���8k��(�z"�R��e"�kwv+pr�o��n
O��O�'�W����4�N¯.r	����߳�Fn�6�5��\j4KMӘU�a�x����P{h6�����`���p~��+��Q�"��ؐ�lh�=�:�y<U�~�9l��K�W+ ���o�_��#��M��'��>�r��l)Z���IF�Dh��Gi�jsW���������sC��L��@�=�/�$��|(���w㮴�4Q���Cy����z	��2a�	΄:���wi��;�>��E`QH�Z�t�P�
�+\2�Bd�����L(B����Z^���bM��h)jD��k� ��쌜�'��h�:���=����XqS��&7_�0�z���mR�}�N�A�^<����ȥ���>\G��|"Gj�&�T���q�f����3��|��hÀh�9:;V�`v~�@!�n������&C��>B!-���i�zȴ4���F/�$�8j�gK��6S��˃W���o�}�d�F�s;f����_��O�jPK��/��B:��d��5�����c9ӹ1���!�0*�g#y��syt����L53u�?}(O^>�ᅌh*�)O���W��b��:����^��u�������}��}ٻ|E�;9;?#�z��ܻ��$
P��OGG���/���.�|K�f����O�W_~� �]��6��8xx_^\�)n��j��֥
c�0B����L^=y����\��M��ZN���}y}�R�؄�:б^>},_~�K������cQa��{q�D^��c��~�H_��{��T��%il�I�=�3�z.�_<�s�YׂH ��c�IJ�Sة�R���}rM�G�K�@E�(���̦T*�AV�P���s=/����)�S�l��>�9�c��G�?�Ay炔�}I�A�����V���D$� T+i��*t�Q$Bi�@��d�x`����N^K���k�,ZM�3;/e�����	�	�H��/)������d-` ��'�b��X�z��I������+�gK��`����@�n�|�D��c�0n7ؙ�2�$�o�-�{��Z�[F��ؓڡ�cBM� [YYQ3�o�fXi��U�I�ߕ��!6+�x�� {0�Q
���\8�+3�Pw�n�Ο�0�P���ƙ¾�GHȈ9�9�u�}�7(#:{�?d��5�	�u��[x.0պ�\$��p��`� ���s����<�g�����?�kN$U(w6���p!�é\�yS�����	�ROF3sf�!�S��{t��|������]��t4=���\�����A��]gp��޺�x���X�q2Hx��tS��΂X��������m.���`F��5S[�g�b�l6�q�"��4�hr���Av�Ԍ#����yI{�����GXb�h,t��PY̨D�Pn��+"fV4mD�
��_���ͭ�{R#�laVX=A}�p̨�WY�{�9`]q!���ҽ���g��*{�(�*�%3���[�G]6	t�/��N&`ƨrΟ.��q.�w�����{�$��G�� ���.�?''��_��w�����[�=it���?Mg��=K��zq�l�L�t�1�r��<�����|t���h��N�����q.*T�s��7�㕓}#�����gU~Nn3X��/)��U�{��P�i+iI��5Pcע
�*��H��q�Idә>��~�V.0Pp���E��k����o(3�s^�IȜ�1�vӥGz�D�O#�9���b�YoP���� �9�]<S5j-ˈ�.A۵k���[x�R!�Ϧ��ک��3����O%�q�\ROz��v�ꅼy�B�/��cF�#ټtYn�����%��D��
��./��5������~O��kҍ�R@���P�ϟ���@g#i��Dq�a��̝��ִ�%��}aCC�8`֒^��fWd<Q,X,"�}s�BF;�����,M��s�n�6T��������x^�)�`��4Q�ڣ�6��~��N�Y���̈9i0`a�T`ȃ�$�뿐��-�������x�J?{,G�c��j���@~��'�w���߼#�^[����T�;��IwB��|���p�n��aS��(�{��A����9:c�5X?ԅW&��PA��ٙ+����+���,K]#��v�:��3�y!��<�cd�"2-�=z�H��W�m]/[[[����gO���3t<��1�}��\�uK�W.KscK7��g���s�G2_L�� 
X�ޣo����K������ɩܿ_��f�'[�P�KN� �{;:�ߓ�ה)+=���9;9S��Vrtt(�{_��ѓt���^d��>���GGGꈍ��rz�F��+� ��)�5�u2���������d�D�y.���Jv�}&��+��b�B$$��#� �6�J���_�	Qd)j{��	���/��)m-ϟ>���#���r���lG�o�^�4�eP
�:�l�Ц�m���^h�W�#�UV�u	 ��F;����=Ej�T��),�g�-`zޙ$uuN7��ߔ�;���h(��׵|O½m�n��z<�4X]���-����������trr�s��S��98�:uV�@���gݡ�}��� ]s�(k�T�F������	 *#��d%E���4�d6�QbH�q�dP�a㿐c3�-d<�J�q�*С  ��IDATqLA�`�#��P�ʰ��f�綽�I.{Vq�ϡ�H�ݨXU��VFG�~�q˔�."j�C!k�H�T���i�)c}R��R-�,����gm$AMeP�5���np�a_ B�+H�Mu���\a+�LS��P�Pk���)ru)�i(���u%C]m��uiEј��pFb��P�R���_���|�Tv�.Q��l��������ҍ������:��MgC]
�{}n]��X���?f�	��zaP�e�(I_Pm��`�]f�r�S�XQ�9Y 	@����N�r]�Vc<6��s9���޵�yC��)�E\�n5yij�L̷�&#���[T��N���u"e�/s3�f��,:|F�VyN�V�����=��_�^��� �U���h���`���([Vkd�]�S���4�YY�}���v��K�T�ؓ��V�{����J�����!eP�[,��o|�=��[�v>?y1j�=�ߞ)�nUY���e�=�����P���E�iȐ2:���r�zp�4�k�SOXL������]M�������_�5��X�Ҙp�βE,FmY9(�U.Z��
�ד������x՞0y�v�"�$T/.DA�����"�0��>�����Ɨc��3Y��*�ٸg�)H1� �wX�h R�Hɀ���Gd�Q�h����"��I���^vF#� �	���3,x� q�+�HLW\���Āou�0l�������wpm��P�K��z�(�B��Q>�����,6Q�rx�R�����O~!��Ǻ��2>�7OO��C�~_�z���TA��l!ղ.���RDh�]D�x�k�3�[�qN��	9�d�1jZg��&L���*��zL�鴡����Bdh
�(|P���[�XNS�tQ��t�"}��A$!'�0�c߰�.�򯈰T�a� ��_�h�ags56�1����B�/>�DN���sMZ�)㶜�d�`�D]��#����t?��?��4{�:��6#�=Me6ui�:�'��G���g:�[��1��mj��m�����l�s;U��ql�G�8ۼ���L����gr���d4�Xq�kz�d��l�`����o���T j��� c8jX�ר`)����]���#�6 ?@�x�{�æ7#������=�#m(h�CaC��I~���Dڧ#^60$Mtiݒ�~=�kXL�+�Kԑ����\V�6nud_����:kz<l|S<�'O����6��3&4,T1���8oiNAz�F����� I��mH��a]8���M�fK����A���+r��URC�g��Ȣ�c���)�i��Q��¥+�֝w$}�@�W�	�ؽX�;"�U�`���o���ye�����L��SqJa� ���#�~>�����dVdqz 2>�z].��mI�[��\�yCd�)rv*�:I��7(QT�h��t����h�3�Թ�U���?�
3�V�=�bb�p����<W@��/h+��gk�gɠ"��5P� �@a�S�u��X{)�QY�UU�*
�^��t�9<��~f� �����#X�L
4�YUY`�<d�@"8`�l�l �����	R�fȎ�u�*e-K��HK:A�	9����쎝e3�f���̗�>�w�(p{	+����!u$5R(j��@sB���Lu@A1���x܏�_o�+;��tFfs��2?8�R�]��J{S��+~�ւ�I��R�	���u�ُt�<=�Wo�%��ɕ�w��v:C��X.�q�v�T���;>;�c]��{C[��F�Y0�-�^9�k���Ŵ7��Rr������/ʌ����z/��]�R�[�Ы�-�b;/p��_��i|� �]�:к���SWB0�᜿Ҋ��pD}}$�{�xXcE�.`;�%q�������Mp��%�����V6�ܵ��Vc�q��*��M9����IŞց���! G"� Z)�-�Y�8���pjQ�J�*�@.g=�V�\�Z��9�����L��Pc���,N>v39�k:��$��������@��0Z� ca��.�j5%e%}6�"��z���f���U���N�Ҕa��F�r���/F��"��UW���à|e�,��;j�y<W�s����u�+ W[��:�Kxv��^������bN��绂Q��:L�K�#�V�J���{�4��"���SS��	z-�+��"�ϯ�S��Q�:#ʾ�*R���r<��@~�f�eQG�Q?b�?nOL�x踹\����,��J�"m�k����b��W�u��K5��F��3g;Y�}��&��4`�<��g5��d)_N䛯K��'��d�����-��wQ������x�I�hQ��
�lz_�;���&D��{Mv�b��N
�8k�Rޕ�}��$�������1���qCac����P��΁*І�Yi�2��R�d]��@�_�^�N.�E�`�I�ʹ1 Z g=`�`N�L��s���+���4ՄYQ�h
�/)xC=C��f_�a.O޺#_��?*Й�t�H5��j����eo�6T/W pe_^_�"�vO��D�p.�X�4��q��F�w��0�:�9����5��=�
���+�퍛IQ;پ��m�}㶴�v���Gғ]}߭;o�ы�r���8SgcGZw��EuD�t���y�L����y�L�
$�����';:��aq���=\��|����V��B������k׮)��������{��_�ן|��&�sZ�����V��߹�#$0�mv�����o~.o���y:������r��{r��m�o��R6{}ٌr���=|ຨ�:���`�(���z��H?����u��bx.�J�!����K3��n���?�qH�FU)��˕kWeK�R@t��]^_���a�M�?�o�%Who��5hQ�2n\�w�}_N��D<{DQ҇H�a@*��\W�#+�_�3j.��4zD�䀅��G��
�|��G���)��	�N^����'ޅ�\S���5�-��?��{_ɳ�?�l���J���r�PW�fAִ	'���<b�8�g�rtf�(
ۃ t2[��j6����3,�,�*��P�Bv��i���A!����a-3J�wF����v�M�2��~NP�	�t�"�^�F+*������+��c=U�sv���&*��	��λJ�tٗ��%H	�3��᡼z�r@�*�I���J7U���@lEnL=��H���`��=�7#�U�=�����Rf��rv|b5�3�1t\.\�,o�}G�^�����#��R������=��+s����'6(��,�a�NqH�
)�0=���6e��[v������$KR\���L�Cj�up�#�����Am��1�Jz��U�f0 ����#�(�Ep��S N6�WTؚ����W��Љ[�w�p���#ṵ���;Y]ʫ�(���_��͘���6���6�յrN��_vЗ@�#�ܜ��mү}����(�U䚑ՙ�ڶ�u�Ö8["�ą�Q�X���Ч�ʓ|�vT@R�]{-�<%f��=�j)u!9�Z�V���\�eñw��jYg��8�#<�ܕ	4��� (@�w�6���z�;z�_�9�;^��)��̧�z��;�#97"35��y�Y!��軿�R�"��rl����Vr�ϩ��=O�9#T8>�M��O]dK���W��Q�^�L�״��Ln8�g��s�_b����j�dU�RoVe�<+-�n��:�Q���sA�_��� 4Y�kH����E��ÂU��g���\Dpf�%ĒM�r�Mp��S�S��?�J�D����J:�� W��ܒW�#�7Bi"��Lɏ�7|N.3'�@&&u��B�����"0�k����:�Ń�(۶V��;8��V ���J1�{K���?�a�+9��Df�hc��P����Ώ>�+��9y%�/�2Q�����"������/�����PzFQ0J��e��<RR�l��J��Ɋ�8P��[�����삎U�DK��(-�=�@ ���0�n�<q�8R�!�͆iqN��YU��L�#j�9�dh댴'誇Vg`��9��UT��#-2�����
����'Q�g�u��Hz����@�/�ѐ�/_�,ׯݐ��Mz+QtA.^��`~�j/p���j�ϱ��[fJ
����g�i]4c���X�6��� �mss��g����m��ؔݝ�(Чx��
���w�8-�[4���n�{�3�h{:�>�;T`WbM�9�����
֋*d�2�qk *� ��=䁫��$nw-��w����1#�SEX'����|;;��kESeKO=�o���޶��{�pbV3�a�P�f�( N����6�0����ӯv��H���ݖ,D-�1W������f�ڔv�g)R�L�3�
�:��65���V�g\u��=�}M"�	��4�MK�+M���q��z��ө���e
����NU��9{�&3p.h�2�FL����ˮ��@����u�\���ȓ�";z��M~2y�Z?����J��J���ᅮ`�p��g9<x-��g@�P [	:��*\�
�Q���vt

�/,:jEL)$�7D�������:ȆMv�N�B^Fz%���h�P��|US3L0`csSZݎ�F�ס��5�1�&�u�G�<kP� �5*�u�YFŲ_�y��B�v,
-��e�� ���z]+��
��^��I�tW`�J�D
M���S��G�3M�s]�cچ���26�d�2��led/��X���^8�h�&��g�^�c:כ:�7��80���v3J3Ku�Z.�j  ӄ���\D�j�"��-F�u#i�
�韩�2˩����%��S�N����c��AW�ӳ#y}p@��V�E���C��ŪM8��-#���p
J����a472�[�&\$���G�����ўĺ:̪r2�Ś*�������\�,��)�e�<���ۿ*'�QZ�=
��gٜ�e˸/��ጚ�S�f����/u��koou/���^��Z(�.�_).���U��-k����ܟ� �,��$d��.�Q;A��ȍ�M: 
���7�F��XXm����8��I��&�1X��1�Q��w��a/�m�l��"r��B� ���}���i�oD���Q	������=���u�Ş����E��h���::�h�g�-=�4���:��9�c�"(�8��ܸWT')�=t��r(�vʜ>�-�Ｇ[�-��"!�Q,-$�Hur!�2�gR���i\��o��ŝhp���e'Ѕ�-��l5qq�(��{��+h�N"����Ӵ�-pT���=���[A$/_5�n9'UF0���`6�aݺ}	�۰��A݃g1��������.�E4���0��ӡLO%�M ���QԼ��L�|,/��\�vd�������ey}��<��Y���ܸ.o�}�ݼ�0�ȃ72|�R�ŔJ'x̹�Y���U=�D7��"��q��Q��s���1bSgt�o!��q)��1I++z�1���mCQC���@��cڃ'�z`t9E��1?h�#.�!�a��c�5�ΎLj�45:�%�(0�
P�9�u��МQ���Dn�4�D���E�\�:ڭ�m� :h�M���C�9|T�Ƹ~-Ӆ��ه:u_:E�(bp��Q��7r�k�q�������t\��$ ���K@�$�%8��2@o�F�CGIA45-+g�r�b|v��g��X���5h�g�0:��Y���8!+Ԍ��k��R�
Η@a����31y�p�M�
p.�.�����,e�EQ� ��6�Ḉ\�bv�8{�86�Q���/]F�e ��2��<��ٲ���;�V���\���d���'�M��������ĨzGnXء��7g0zA��+k5k�|Ye�Y�����ZYz�. � Xչ�	T�()�0�u�kp6��/>�X�lgSFjK}4��<9}~(�?�JZGG���=�`��dx#�m^&rz2��/_J�H]��2������T3�&�E�����3�x�TX"+�	.�ޠkYI7TT"�^��@3Ԟ��lg&_s�m���:[Ț��� �0�̮���.l�y��9\�&Z7{W�<���<c�F�B�Z8��\��@<uG�7��`=�X���ux=5�v�F{��h{G���O�rtx��&S]ðp8(Ɓ�|e�Wk&����R0��0�#u�A��
}�0�^:\�f�ks�/�x�ZTVY�����o���d������T�"��f�3�<�����������Ć,��Ѵ���<}�� �,e��U���k��w�QGn[6�vt=4i�<׵{�f�8���wu���^�9�kz����~��k�s��S�b~�2g�tς������E.�oS��c�Z��f�W.��$`:6
Ɠ��u�sq^^7�V� Q���cM�1��:_�v�ӆ�eqFW�����qY>�y�x5��+HP���{�1��2(΁�y �@�H� ���a��*P���c^7�A` ��L"�~Ļιᵑ��f�:u�ֲʺ�TYOƿj��[���?��~�F�ƎN������f��P�:�Fr�*rko�U,���iCx� e����� ���C�� ��Kޭ�+�f�d��*?Ph�UY������\��巛�9�[TO�Z�ū��x�"�������(��:@'�ԩ��"�).�/KSg
s���)A����bE�+�4����譔�Ф����Js`�����
�V�0�F-�(�0j_���~�̡��i=(�p���0��sIu�L���j����oa3u8��n���j�x��i������m��\�֙&㳛�iRȝ>{�J�7H%���L't
����˙�I$�����?��v��y�����:�{����7�H�mJv�B��!�_�B�ϞJu6��b4S�4��8҅�`�3������@������֩_$���E=d�Ҭ`T�E�Kt���㭧~I�v��l��7�������	."�%Je]4V��=h����@��simm�:�RM�n�t0��v��S�5�*i�:��B*���s�P�:'��Q�����J�0��FL�yQU	�+�C�Q ��/PK)\/�c[��8C	{�g?(AD�]�QT_�*N؎��m��c���qn�0ݎ:�VG��N� �<�\#)��,%D������ei�)9��#��ڮ�
�*}?sxJ��� =�l�φZ¢Bp�Q �FH�fs	�ۦ�So�!�2��*�k)p�,�e��x5�x�ѐ*/-d&ܳ��I�
� K� U�5O�oϤ��`V��l��������FVǣT`h���wY�Z�˴�AW[V(h�P!`���;S]�A�bs%W�è�����A�-nr �h��\��s�2q�Bj��wncg�\:�%�]O�!V =}�X��CY��r4R�v:�P��|���ѩ�u!����-I���ȱ���mZ F��:9�9�a���$Y��.gf����5�@� A����!��&�ˌ&	�fS�5{��s�c
�x4bMCTY���|�h2%�����9����g�Av�edZB���k ��Pn��}6o| B��-uza�!������|���r'������0g�h5�~�A�������<K
N��g�t��[3Sb�R��%A:�tH�����2TLu
0�@����x�`̼�-��n�Kd�P���֥��[�{��9����N�{�f�_b�R�[�O�P�T}�E����0�ԡ))�ڛ�����(��-�B=��[�%|/R�ե=� �q��H��}�֔W�XSVVA}�#EM���`}���_!�ګ��[��1�"�\����Vɀ:�y���u@�Ⱬ i��t�K譃�5�Y�W��'hd�c�>F��ѕs"1�snP���4�o�aE-h_����8zS]d\����[��� ! �F������4�T�f/��X1��5��Njs���9g[�Kk/� ���Y��`v삁��j���!���$�\����x��Ey[��=ţW�t���l�E�tLZ:<h�����!3�B���ո�EP�VE�t75O��N.�䒰��K�V W#�{�nΩ��3�Y�h��8U|���B/��|
�T,x�*���<���X+���0�,Z�*�Z(2�fN���<����_���y�C_��.\�<�	\H$R�r?�7�E����+�2ȊL�C�7�D�K��	&/*Ƚ:H'�n�G�b�A���?08R��+ez�yy9L[Q,�,����O�Ju�t�(8�{������rf���ҊB��
1���х1�tcAZv��B��6���UQ����!�\�OV���Y8e3\y��39NN��sccb!vn�4l[������#y�����T�����+��+�����4��MW�����ȣ��7?}$��4�V��"�DG�T�B7dNu��x�,����L1"��m5jUC�S�H��E���V�8}����=ih �0�\�h�A7t �ɘEkT5*�X=ҋ`HB�c���ʍW0�o�8&��I{s�4�q��s3��S�Ut�dh^+ '6W wE	���*��Qd*�+��D�?�ć��4
��^��j2��:��\&�����XAE&��lnoI[�:\'ӄ��pR!@�MyM�pw���T1�$�L'�$w)h�Q�_$�^f�ܼ�mӯ{C � ꈀ�p����mcW��)!��r�i�Eޤ@�<)tmz����H^M�D���DC1���6,���1�g��(�Fqg���q�߲D�8 �-��4����-mSw�5�/.�r���sD��A2��
�Hba3�s΁��*D�[
���u��g�B.���( _�9�]����0P�*�s�Q�5%�Վy�%Av��N���4=�mBf�m�%` M�����l9@�������GC&p Q8������ߓ%hy8v�uU�c���?�l�kBV%�L���UdC��Q���R���Ne��6�X@�R��d�j��Ao�Pbu 0��V����_��z�vz>K��T������A�
5A�������$8�)�|�Q�\T��9fh���4F�)���><�VW��Ύ���N*��Ek��͡����~W���׏�=�.��G�5���j�_�����X�����u�Eo�>;Pǂ��ˊ�q�t���T_t
�Mt�ӵ:C&�\J�1�&s����*q��ROK�r��2A�ޒ�=�ܗ��y�Z��Ƀ�gpX�CN�;@�B�mM�6[r��[2�����)�g��_F�sK���޻�T'�I��r�)�*��q5��$̮Y���b}�Yr�>|ߵa��H�[����cQp���su#k0��=����*�i�U&aU�Z;"u��y�l�\Fb�%u�t}^f�j��_��~��F��e�I����s��cF/�5/�䬬�b���Ndd�f2\�z�ZӒ����Ω�?�lR������ܽs��5��k7*��gt�W~�Y`uY~d�r����� �##΃s�Z������NA����w:.�_z!�����v���r�7+/U�5K`f�F��za���+2V`_��Aމ�.������+R�ne�����_Z�'.e�E�.[UU����� �H��	`�(�.B�Հ�A�,𠼡��#m����׷�������eF:8v��Bϩ��~G�j�kt���?s?7���I�׷Q~;_�kk�c���,+��̶��$I��hT~��G4������'U9����ˍ�t�B���]�M��9�\ ]:���9���h\fё�ta���͈��Y�1�8�8)Nq�u��Ԣ�A�#̚�3i�}޾��4��n�Q���n��͓D��D<�X�/|ټ�����i�Z���e����w��ï�K���\��6?�g�R�t�D*:i�t
�n�)�ȩ#�3t=V]V�Wy�6��ڷ2+��/	!��6���}��,<,]� �M!������PFI%YB�S7 ]�6�k�������n���x����Y��J�[d�P�W����5�8��ҁ^J�_s'��9���K�c� g
 p6�T0"f�q�!I�����$���� �����@{A����P�s�inRP�%#�΍�=fӻg�E`��t�^R0ds���=f+~�����cFfyߞ��%�)�do�+�jH����G'	M��b��4�r�EZGĈ5%c��"�������X�K(�����[/4�s9~(�A��=��������`����
�5ҿ�-���2�B?��B4,CT8����41��ղ)m�!���N(hE�qM��$s���X�'jg�s]�!�B�,6`G�E|����-�t}T�i�Iu�!n����ꜯ�5"$@ZFi�~����X���S62�t)]�7P�
t��&�f�� r�ˮ�st*C�t������:����zA8�{l�ڴ�����@Ci���m?�r�c����^G�F������
�0��}ll_��W;j<6����Qm���q�s4
5�%�|Z�뵾|y �^����9�&�_�,�`�!-�o&C99<`�r��x��w�����<;��G�Tm5@2d�ߗ.]�N?�y����Up�k�v()�)@ �sG����w��}�9�qabdQ�F���t� {����1��ٙع�yޤ�2��f����hf9Zi��6Zj��V#@a������0J졩�.�U�ކ���kt����{�E��Ī�DF�3��������x*��#��o��l�ަ|2��:VЭd�;�"J���2�(P��f&s{ux)�������\�Jê��a�u}�"�1tu�Nu�W:Pd �ΜQ��f�'��0%��
fF���˔\>��%B+L�o��`���;2Y_5.Jo"����U��a�>�K��z�Ez���G�u5�{�s�0r6�����O�_�3�U�)�J���3��Q�1�z�b���V����qH��.���/�|\7�]���R� p	 ��"#]
9��ֻ5�#j
,⤋�Iy��b�f���������و�-Z��B�?��ο�?dZ0XOXL<btUy�X�K��N3���ZO	��p�I�z����i��G�zhnN.�N��S�Bb�ɳ^6�]�;��� �������Ï���y������O��|����l!�.E�`f�d<�4�/�8T���U�l!�:�`l�E�7��cT�M� [(~�2�uv���DEc.�� F�I�Mz�fR��V,h2�IA���ui�ܒ߼�-������߽�����TȒ�4��~���?���LF�����=�a_>��I"WzfzI)�>�c�:�tFl(�������49�Q[|Bf���"w=�(t	������O٪�`�������tB�]�{��t/.�oI�z�J�ӟR�n�E��(?����0�{�
lu^��1��\fAb�})Ɇ0c3��#;B6v�` ]��p)=h~SO�Ε���� �"��w	����rc6�:�,`H~"�xs�[�@ʃ�pٕ�*���Mʜ�S±��<�w��� ���\+5�<X*#Q)������rכ5�"�5B��N�M@�h���\������Ӏ����r"x@�t��N�rؔyc��6�	&q�������b1�B@�@7u��A�,��iD7S�!EPŲ
�E2�z<��������5�P�Tvz�s&�%ୡ2ti�ICGL���)A�C:B���.p��07�{��l�@���Dv|a�� é�־�:F��4^`�3O�cP�,@��Ќ1J�DI��F�,��ͪ��:n�ϥN��A�@T�U� �~���,�pn�k�3��g/���P�]zCM4 �������t8���#y����z^�X�5#�jcM���@�-��)������&��0�S����w������@g_������{]y���<|��$]��0޾w_�V�9��Aqt|���\]�}G���Tnm��P�`p�C��h�ݛ7�{����?�=)���S�����ń�A�<"��U��Ɗ|��ߕ_����7t�ӿgl���s��~A}�=x�l�ED�Y�z{uG�{{��ֆ��ZҬY(����خ�(�K�jH������8NAv�Xh��լ�JQjp;w�(��P���nxp�Őr�ʰ;���#)�Rihr����:ׇ2hkt6���HA�4M4��U����:ME)�>��p���㵉u3%5�T�s�z�ԓB�%��fb���9+����S�9X�a�=�~�����`�=p�R#�����A�	��}��\���w���L�۽�A�s�^�$�����궯t-�t<4ό<]����� ��]�q@ϭ# .KA�d��	B��ͷ�{�)�ؾ j� /�D�]�i��_2�	��R_�0���� �'��9�9X�!<&h�	\p@R&�c�*��qw�xXO��	E�X¿�!����UR����_��<~��G����.��
,ث52�};���Q����g�!��cn�.4��M�R�V��TG�,6w2/�&Z�T`<>}�P�)��z:�5p�$օҞ-=&�%O�"]]w��ߓ;���ljB ]l?���Wry~%��Uy��?���M��я�u�<�]�����r��LKcI�D�{�u3��;}���)7,2%�{=*��K���(r���fh�E��w�O!��4ߋ��X�'oV0X62�A�C�V_�: �1��M�9+�����G��y�!ȲJ���d�&G
�6�h}�T�r���i�5��S��pJ��>��1��Bހ?T<��mw�T���	u�C1�"T5C`Du�R�E��k	<9���n�*�}���A-pϨ��k�W�=�:p�G�
{�ݦȫQ�*[N��j/�S��U C�29ɀ)� p�V�#dS#G#�L���;/ò*��5٦݁�:�t�5�7r�g�9:��!�B' �k#8b�jΊRQ�;��"I��(G��}�sܼ%V�"���Y�e&��E$V�� ���9iK&	�7��H...48JXER"�O��{;M� �@�K7#�J���o� ft@O������噬on��1���<���I$-�^��tCI&��Gn\KP�*���'.�?��
a�.��:y�Y�3rhF��f_��.$�ي6 ��.b}1��r�L�G�L@lN,�2l�^M��+锌'�v�@6���/���<~��sᶮQ�;������(��;���ܑf��59�cvK�����v����U�4)�}�仄�8'F�FҀD��2m�$IO��������1�c�s�r��wey���r��]�F_�m;�_��ܒQt�:�XH(��2
k[�Ԭ�[r;#��<��Q�(2�ggg�e�NUݫ*P���2�3�ƚ�-���uKT�����ĺ���h}#G0�,(WpMJ���0��膛V2� s��#�ɹ�S�<��3�-�������&��턋�+�5j�'gr��Pڝ�C,E�SY��±�,2�w�6�ot����Ä�a%^�	A�s�9�O����k��V�����
I��+$p�1�%�V,)��	��_�_sx�-:��sC܅k��	��s�T;�4���I��ps������k�ހb���戮�uX�ʁy����m�B�]w�l�2ح��cV�5	�,�NQ������(t]m���J�����-Y�7���ރ�	�(��س�&���u0�)��irO�'<'���ī��ldف����#�M
�������i��E(JY�a+��n6eݠ#ʛ馟��f��;#�-0e!:��?nu6����`,1�����K���#�:��۰*(&�u���_i ����s!�.Ԑ�+�@y���Ft��ߓ����R����^��gJ��Ci�ȫo���#Eɝ��@*��J�{?�[l?{�XƇdi��I=��������!�:.In�`�\�"�8߉��G�t��D�������<��qs�+�dDE�zvH�#d?'8}����P����BD�*"y�s+�%H��zM�4w��j`��wA<D�D~T��kƬ�����I�A�ɣ̂ l&hM��k !Ұ�CS.��D|�˕�S��⏮��,�o�����Y�J�*��~��I_]���\*nJ�s%�gm)�k*բ86a6�|ѽAs�I�����z�RNNN��*`3NZ�U��O��f���+y���}�]Vف���,�#}~���L����u���U�s�StT4x�u��I���~��9��:@g�")����i"�A ��c�{�_����܅6:;$��b�Y5�V 7��1��ߙ�M��i�ҩo��=���m_]񚤺y�����(̹1Qe���.����rqv.��5��d
�Z��e�2H>>:�zL+ȝ����-�ީ�ep���M�߿/Rk�y�R�#g��EfƤ@�ג����%u���`>�
�ȵ�����gjG����yD�N �{3�44|���N�s�����A��AfP2q$Sȕz�ݻ�?� b8+( ����3�{���{_��S���h�ƐepfnF����a��	�T_�*3���P�H�'�3� Y�+�A��"�1�{h�[h ��l�	��98�GOr]�w��ܺu��DS��^��bU�y�;RP�G���u�Q�̵U&^�d��-0yF7�%Bm ]�NKp�D����ʤrh�H�:�z:�ׂ:�d�a��a�<������G�C:�&�46�HS�,���М�k���{��پ��f(eH&Ǩ��:�s�J�$L�{GZ��f�� n�*lJ�p�� '�lZ�?9�"gNwK��;�+YkE}�	ݮ������ o}sM�nm��w�ʆ��.ܐtN�l�k�7���R��$8݆�5�3Cy'���*��*���/<���/�DK����]\��ק�V�z��?�qH����%;��mNC��0����s��F��/�B<�\��W,t�ԕ�U�}�{�Yʉ ��C�����a\.�Mj��أ5yD�!�F�Do8�Z�u}���O%��5���AS|��n�k>⭒�M�So�lˊ&����u�]]ے��GҪ��XQX,�Jz�.O`��Ž��`S�������6)��x��@׽x0, �D��'II�Y�`���A�Gy��&%�B�9d����pi�a�oV)XNXks"�F ��f��^} �1�3���Z���I�j� &�%!1N�����r�ήV4��^��������sI�/�6Le�|_�N�d�����JM'`�|d�x�u��&��̋1���h.5��T�$A��UM �J��0~���=b��EE�$=�i� ?ɚ�99��	Ƃ<x�E�����q�&�vޅ,�9��*��캕3�"$�>�۩��Uf���f��&�K�`�M�e�R�aQ�- ��s�$E5H�#D���}$����3=�ϟ�������k&,�@PVA�dJȒ5�A.��F�<օ;#�/�n[ʎ��o�\PZba1Of�-�H�G4�5��gzQ�-���os��'��j�pt�/��P���=Ϲ�3`S�+I,�8;?��\E��9��͵�63d.5pz���%1A&��`�-^�3th�rp�'�z�n�{O
�h1ާ��!��T�5�1������\�&}����+�	�:tW�\�y����Z���\� �4�4��@P`2!�|������N��3�`a�"Ʃ�5��CT@�u~���Jn�Ϩ�ZT���J�x8��59�$���x�zM3'kl���f%� 9���H�F�N$w$9k��T�������<T����~1�a�cI.:%�� �Q����4�b�91�z2L����<�8t	�T-�(A����)��:	� �ؔ�z5<�1���)��
��1������P��]�sK��dٰ�)U�@D����O���
՚�K١AǧZ�Lp��k� �Qh�z!�ɀs�%ƒq"�!��0-u�5.���[�e8w#(���n,�|N�0�S�4���Hl��Sa1�*���9���iOׯ�^_��X
ь"T<K\AI�	# <�K�"�x��j���u�lHF /��� 
�
��pp%�u��
�#
����z��ir��U����z��jn�9yHS��%�¥z���ܽsK�ƺ|��e��?)J�*p|L���yU�B~��K�Y��R�W�	 ၶ{C�<r��ۇ���~[^�>辞0WD<5qQ�spť�z���>)��ֿ'[Q�ÍfŶ��ˮxr=y��� �ׅL�^�nGI��|�ž��}&O=Ԅ��.�8R_L����S�J��8��ѽ�%u�O�`����1# @忢��4�-5������5$*h&n����>~!��T%����Tju��F��1Pk��S�D@�kw�(����󀼮�����w[P�e&�T@�o�k����ǷI�?��� �=,fV�/�@)�BV��j�4Ɋх)�I�2qn�/%�LΏm��LBo$������j�ʐC�Z?
��G��k�P!i_��+@b��<�L7��I#,��I��9x)����X=��W_Hxv"i{&-���c]L�S9:o���H��� 3_���b�!�V�zRW��x*c@�Xŏ�$Pu&r�������W�������-`9ɛ�x��bV�P)W� 2��/ �P�/�J7K)�X@#7�3$e�oh�W� ��J�x�O�*69��Ɍ���&���[�06c�f|�9�'��$��W#Q���:��i��%5��vGΏ����}p����X���B� t� �A��N��d�"ֹ8���j�wڇr����ޓ��ޓ��W�ı��������FD5H�m9<ܗ������n�:V���"�@��ݨO��ל�qo�9�L�WϤ��=�b�{�AW�޼���$+X�� VT�܁�E$��r�Kue������P�!$������P�#�8;������q��}yyN�Q�N9�.5���ܼ��O���Ym�s
tΨ�qvr���R�!׈�� T��a����F�/R����H�:�I0��"���6:��_�|Ic8�����M�x�@�p�ք�r�XW?ݐ��7�B�~�:���0 �T�3�P9����0���o7 =l�jR���3�dw.�n�ĜU~b�	r�[)k���O��'|�0�H�J��I1�uSj5(�7y7�vN���^-I�1_@E�)Z�g �En{�n��@�
�fJ>�3M�9eBw, 95��$��͊4kU�P�s#e���O��!b�	��ƚ�JE� �{MI�"�Ip�okb�s�\�7n��܈���.@,\�� Ht�f��o:�\�ާZ�L�â��G%�v�u�By�cg���Y�@>�U��FC�2���qw��7��w��C&�`���Ŭ,.�ܡ�p���9q�i)�y��Ҡi��y��%(�tvt"�p	�ĺ^.�0/�,�'L?��E��
���͉���������<��È�VI�.�����b�:�UP��I�ߖ�`M?�F&�檡��ZE��i<�?���{_��6��.)����#��/������w�e�]m�j�dݔ�T��<r�2�����+��c����<�/��E��P'2_����y��<~�B.�(��rsN��c]�����u��3ľ��;�����+��e�����q�rv�H����Ҫ�Zz��J�ڕLr��ԋ%�}SZ����4�Yҹ�c�Reer�M��c���CY�Gd{j|,��Ѝ�����7sk�qA���?���k]Vc՗o��o��D����B�u�!FxK8�"P����А���ɔ;N���/4"Sn�N2k"f���o�^�������C*�9����T4��zC)Nt�`?�>3���sy>>�䣘(��+:IHdt�㜐P$�g��{���М�{��uQ��H�b#]�������L\ñ45�C��Gy]L��O�BI�̱XŜ����a��D`�Iu �EQ�4�C7�I�O6��������5��� �E-99g"@%� ��t�\=&�bn���@�/a7P��
,ep&�2[�b0�@�J�膈�v�W�Q7(�sg$�tS��)T@�� S�	`EX�L:U��i�3MҞ|�%��di]� �G�\\��h�zyѥ����&"]Bkb��4a<t( <�?�v�=�>}���.��ub���P!,��A:%OF��J�ڋgO�}��T_��{�	�\��D�S�_�z!���Rj���u���0��Ak2#��T����/e���/����=�`!(�5`5�T���<z�����+/4!H��Q������P�>~�n�k��_?'|�xA�L�i��5�ڗgO�e�K��Tr����+z�&U��^�0���S�&A�.��+ʝk&�\t��|��'Oe�AaA��)�~n��s���LӀ4!)x���#n��N_�Gv~z�ab<=�z�PQ8[���:s��I��)~)��!apc��Q�f4��72��9�@�G�7x�̹������K�GЯ��t$�̛�c$ѵ�g�FÎ+ F�AJR��� #�F�@(e��(؀�	 ��@�K�*���<O׬SM&� ^PA����5*�1�	E0��HV�Z|=b�,���K��J>z�c$��.R�;@�
)��t-5osQG�5��f��e�l��3����Ғ&����z����ȏuPV�Є��H,X���X����I�X���R��C�gkze�y�[���ܸF����'�]�(7�VHC�@zzͦ�9q�Kg�z}ϛ]]�4W%{�R�>�Br]�6�`�W�tpI�$yͨ*�j(�1�'M���}��)��m�*m#I��ץ� OYHr;�и)�`�	IK��)/�����n���;b�9d���[|f��ϲ��q��bʹ|9�r������Dߎ/�Q,����e�N�;ꍡ�]@��
��"��p�z�t#J����[L�X�~>v�'�t2�[�X3*�^!���	���EþU}�E:t�ȩ�*L�V]�e>)4��E0]ϰޡ���^�A�����@���ƪ�[���"[���{-�s���y |�Y`�e�Ǌ�ƕ�L�T2@�Z,��l�Ƒ�\� 
O)T8�4�6)��>��懍z�u0����x�(�ƛG��?/̚���hµ�<
!���O�0X4�<s-?Q<9 ��#�s s@2��3'v����U���.��5���@&8LPeO2��$gc�.m��A���*5��P0E�$c�Na3jB0��0���P���j�c�@���9o"p��V�@ ]@�wN0�BF���ZϬ���l!�F���jYH2]0 q�@dUga��d����谛3h7ܸs<�`,�k��_
�(���М%C�n$Q��L����P�%� ;aq�q�&��9�&z�z}��|qr������U?#��?Ă��`� �>d-Mk��-o^K�Q���0ƪ5[�&�F���� !�"��(J��2����M��)`�4��Ns�i���2T{#�U3MF�Иj��02�EYY[���@�+��O=���I
B�u`��5*�t�@r$���/�����ٸq��\�����bM��n��,ũ5�=�kW��JS?-�)�!���}CTω@�i"��t���Ri5�֨r�T����+���l��d�ǚ(@�pDxBS7��jz� �8��M�332䃫�9��R�}-�p��B��-��x�~o�nF8�����u���Ԅ�{��{:�����xa�X!�P��>����X^�x��eo�mw�s���t\��<�l����T��|#=��d$�	a�i?��F\ERW��b�%Ϲ#p����m#�����n���+&��m�HFLD���IGe>!"��.t�Zt��&�K���)zC5c�Z�mؑ.��	��Q_�A[������ON��W����xS�ϭ��AW	SD07��fTL �4"aQ��A��/^Ƀ�~��[�� I� z�<�y�G�?doR���V�ŲzW�h��Ԡ��ўtON���N�*�l	��jjk!aM1���_�z}|�Z��(\qs{�nЏ>�B���?�!�b���$��c}�̞j=$0�N���jIFz��:<��A� W�G��ˏdusKʺA
eT��5Aҏ _�@�L#r�Rt];~�	��&�Cc��1��[FI�ïʚ�����HJzWu^BYi���Z0?��������0�P��h�n��d��ǂ86�1����(h�I@�i"3/0��$�*?�P$�u ���֌ vjB�ɾ�[��=��W�e�^'������9;,���Ӓ�!:�o{Y�i<'nq� oA��Z������K3�[��s3�4�������A����U��Թ��x��o� Y�ȸJsǙ,���S,ExOP����4y���⺊C��-a">�q; w�Z�SFc�9 +�I���6�CP[�X����ԫe)����$��΅�a�&kk�TuC�q���df�����q�<,3�J�	
�Y�b#K����1-p-3��;�&�@�����N����/<���ѦdU���oʍbl�؈��#t]E��c�S����|�=�Q�䶹֮�l��94�A�u�[s(B X����S��8�qB�[��3���(���p�P�!���7'�,�cV�i@������J����s�P���d���0Kl��5�N�$}�84�#'zfJs\<C�ȸ6�@�eR�~�Ѕ�,��|d%bx2�>�!�)�Z�D�B���2d����g�GQ�G%�Lj k��܂�~O5�*�=jBB}*@�F ��`�B�Р�2q�y�!s)F)�U]�t�*֨>� ��-=�;/��D��N����p��r�ݺ4�7u�d��Gzo��C9�����r���+=ה�Xn�gc��3iMBp�Y]�+�ּ"�}2NemG���
���.��f��'rrp�:�����Զt����b�+�9����=i�����A^csSVvw�A���6�kxO�œWҞ\�1��i2P��*�]پy�Ȯ���/4ahO��2���ǵH�4������U�v�������H��H�t���1]�WVw4v�i#�R]�yw"m=����z�.�,�B]vwn��jPWM&���_��r��5AE}Mce�4�c���TK���|.Gz�¾'�t��]����8W�Ulȴ�#�;=�[����u�ԛi��iB����le���D�5Pż!��cnDR��	c���o����X{�ryx)մ��:e� ����c�����&N�qr�  ��
e-k�pe���}O���c���V��b� $�9��� rC7�`��Ī��3����tƐ�B�4E"Z4IH�E��<�J�u&���J�^=��|�K(�y��|�'�����z>�&������wޕ����I�?�Ӓ|>B��"���?I���������/e��#M�^��Ԓz}y��4^�ߺ-��u*�i�&�م��`'G�޼�����J���}���F�%����[R��C[ha�rI�&����d2���W#�_=������_
�P>��ړ�HS�2]�5����'-7����x.�7�%_��-P^1��I|H���S�d߽<�����3�	���p���0���I�h�q ����@Z���tA��s�����g(��=����NRiN���̥�Io]�r��utGk�A+��t*����u���J(�i8E�-���*�����ir����&L����d���������1o��j������}/���:3țs�dE9"Yʮ!�iP�
���ϊs��gٌ)���I��κ �(rݕ��yLP3f4w����e	�\��9��������B���~��;�3�Lq�˦҃-��B�_#
��yG޽�y��D�F{H�[��-(���� �- L4Y� ��>m���)�Dѫ<�(��F�kX$��B�խ;���Eh!�+��J����%�{<����}q�UI�3"��,�'�b����� �qW�~A��Cj�)3L��K�<��DSŚ�F�o;�����w�����_����~�����\lG�&3G��X���o0)�'r��ؑT�@�`Ui����+�v�*����ɣ�lң��D���!��w=�Y�o�gR0'p���ܰ�*�_)���`-�Eϓv3�[ �J�Ӆ 2��c}�T�LMs��㌄�p⒊BB�h`�Q������L�!H�9ө,}[��Bb�9��X�_�SM��2D��)5�x��V�;�`*lJ ��2r���Y�Xa5�<��ꦃ�; ����/n8C���[3�]�!;;7���$��Ύ���Ç�%<;#�t�K��ySv5)�P+�-y���_>�\��zCX*��
 �oucW�T�~b���SoU��^�$��'o���j����DM�/j��;:�;�//��Kק:�b}��;���;2�%2����=���O�~�뽷{]�Teu{Kn��.�X1��1�ɨߑ����쳻ITכ7��w�'��DtzNXE�b�K	�_ʼ?"	��Q���ܽ{�AȭU��|���}�qa�Ǭ�"��޽��B�\�t8��7�W�/��'��R.��Ӫ��͛�%�`��t:wֶ݀v��p���s�������;zÚ�2M�j�[+�씊ܕ��9�+py�\j�����ipt��P��k���%����S�*�����5���zL���M�\�ʚ^�R����I�xe��������hR�ݴ �w��Sa�$�,���,7;���<��H`�4�'���@�!g���#���Ȓn��S'��p�о�=N�^5p2MJN�>��-c^<!ݫsY��T[MV�_=�J^^��}�o~������a)d�;TF!�Jo�ܠP��(�$�)Uf��{ν�z�弮s}$��P�k���@�����T���O[�g�&~�Jӱ�@�՟.�]y��W��cncs]�Dl�겡�\k阋�����|����x8e�k:GX#���t���==��Kyx���Րs�Z��H��hO�����R����C�q(��K��Bť8Ҡ��\�U&k;��������������r�b�xyk)[����P@K� ��`Ơ����E^���v[z�E���{��؅��Ye(e��g��,s��xs+�a�Ge�����:>!aHEB �G�Wr�a��0�Wf�*
Z&��e����d�;��u	�E��^���g䁄�B͋�<w��e�9W����&.���s>��F>�]bA����`I��8�'��2H_���A����������q�V�V�?�!�M�_�&�k4��&.8�2�Lz��&t{����7��P+�����(:ށ���e�kcI���4��W��Q�[��ӗRU׍rĤr�= A�iB��~R�gz�#B��� u1�iZ�$>f�{rս-Ctf\+q�U���epͫ�&����_�o���/��������'�|�����-f�BZo�LK�9�$�!3j����L�:*'+&�M�����u\���*w�%Ķ���xY���j��x�?ѓ&��[>R��y��,[6$9�C��D`�?O�
�����M���k��T��ΉMb����v�,	J\�a8�đ;��R�\W=S������j�-���3�k�U#<�Q�DHbvj�'dKlH�CA5�D�II�zlC�v��*��T �L��T=�����9q�dA5f<Հ�V����A�֦T�WIA��������Χ�H��b������$2�`i��:#��i��կB�$kkk�n���8/Ȧ2m��7�t����}�g�dS?���*�R��|��n�P7t�r�o��hb�&�&0kĸ����H։!3d?�V�,A����`ky���ȍ۷䫇Od��
H���TuAߺ���^��#bJ>��_>�����Zxs�?�mm����P�ܻ�AtK� ��ӈ$|\���-M�6�C�Ҕ�wnK�٠�IBXZJhZY6�2U�J�f��ܑ�|$:I��]7@�Ij=ǜ�JЉ���Ep=���9 6��f}sC��+��M�W���deeUǈa���`W�{��i�_�>6��۷4���vwJ�<��h�o"��dk>Cg0��w��X��ǁuz��}g�=F0A�$T.]���
��|Ɣ�ID0��,'��Y��R�8¥�3�`/(���q�R��}0�K��C,�>���֙�u�]����g2-���5���ڱ3�`E�{}Kv�+���D���ϙl�����.������>�H���� b�?�l����'�F��.(Tv�yIz݁t4��/$�7D�	~H��PV���Q�`I�;[����r�kFC�e�T6�lG�C�8bo@52���'���)'z��wde�&k:>e�����|!g�30'�؃��?������u%Q�N#��Z����#�K{Z�J�L�4�r����N@�
0Η���M_D�*��"\g�˩���6F� �x$B��I[���%��꾈9
���M�t�$S]~�LV����=SB�L�
�qT��R�QH�G��b����J������l5tS�J2�&b�p���v����D�,�TÂ Z�i��K�����V�Aw�}����K��@l��w��t=X���[ܟk�A~_�ҞȏS"�?��$�E��ω�Γ0�PKjp�P@E��T~ ����'��P ���\��n��u��n�g�Ԓ]|e\�l���?��pk�:6<����I������	�q��u�����l����&LL߳��}A�J��q�LFW� �\�H��f�!:VGÞL���C�۳��j+0�zR��̯u��^d�&�������?���?w:W?���.~Gd�_���%vm�����3����a�ܹ���)?�ZЎ�<�F���I/��*�a[]" �Q92,�E���hXYL�. �V�D����t�!��5Mg.K��X�j�!�,�<G겻*Bn
Bٵ�EX̲�u􋡄��|��Uei.�v�0��F��8N͸*�LJ k�h0;�s3\Eэ	]��7� ����n�zo�N]����7\�¬�W�^��07[-JrF�G���BU�����P�@�B���U�ЭZ��@��PT�"��L����4�y��9�6wo��R��h����ϻ��4�hRfx��JK�Hj�\��yT�Y�4 6Й3BrRԅ	�F��}���}�=)�?�NLX
���'k8b�����s�����_���#��kUՀ�J(W�7ꖬʭ�w�!�{��T�&S+++��
���{\��7��t��tKFr� �֨KP*������z=�4�?�1��767�� 2�1�Z�Քw�O_�-��G���A{mm�p'tɞ������j���#�nh�d�C���6�jt��ql�Y]Zk�T�@�A"�t���66e^��+ P�衿��6:M�y�=@��Bm��p�&� ��! `�F������=v���e����B!X�5S8��Y�9z�"�s	����/o@`�`<�1��!Ԡ�Q�k7��2`6�\�s�� �c]8}�Jm����}	s�X�.�@_6Yߏ�G�A]�b"��s�_�|jwI:�cS���(�}@R�BE��frHf�ŠO�g�`LiZ��..e��S	vt�L�� Ay�ICY��4�9�9i0�� dw_mM�c�����������e~H�g1*�fc��kQ���Z�Y��|�II,�s_Z�s�E���$s-37�_����5�1���s	p�{l^;�����}�f92�G������vn`�	�&� �O0J¢�V�J�&| B��^���u�Q{1>S��#/
L�u&������VhJ2��ـB�'G2�6�0�s�zN�} "瓳���������B`���A�ȋ��w��=~��HT�����u���L ������X~.`��yKI�����J:�(0h⾵������s�y�4��0��\&���2���%�y�ZG#2W@�:�O�U�s
 .��b$�#��~����ul�4��c/Þ����ӧ��ye�9�5D@BР/��u�4��NG��ƚ��u�-ȵK�����D��~�����5O����>�M
�����w^��O~��`4��8*W����;?�-@�)�jw,x�����6�a�ߊ������l[q�耇}�n��pB[y���l�
�t(���YT�=4���^�o1�-4^����%0��'��' �B���I��Eľ�.����IƢ��Pp�+�kyf����p�H�bA��[�W����ೝQ���:�z�؊�0Xq�*�~U�>�IfN��d��R�A*���a�vp�,���_��Tj�nIA��V&�#�_`U���5�5�$�3��X������C�NY1+�@p�jh^I�7$Qd�Z�n7R����c�������i��5yhR��*X�W�VY�5n i)��h�s���\�X��$+ ֻ�l�� o��K�Sk`�=��]� �uE�R�0��V"���Qf�\�@�p�A ��cE?5M����ln�H���1��Q�ҐU}.6xK���p����>�/s�!@d�O���PzAAϻl�MF�/�m� �Z�X��m�>���kj��@2w^����A*����`�R���ߜ���lol뽩RN6��� �����\�����U�O� �"�����J]}n7uU��@yR���W�i��p4(�0� $Y/c�� 
X�PE&�1w��b�s:���+�.ɞi��N�,�I8��\��m���:����2�U� t �6hʃ��:&t�5������T�p^m��ҵ��Jq�T3��h�>�/<TB���C����|��L%�1WF�0.2؀�V�츆���`���@�P&|3����&T���#y�wO�wߡ(D����&Kp%�b�&�. ���kT�0F��Ki_���3M�_Jv����B����6g<g�HwFp�E�#M-���2���m��ƭmi�*2	�v�N^�6|�Z�{0qDW+7�<��4�̨.��^'�hhlN��:�b℅��&M��XU�\���w��l@2oL�l�����?�����V�"�>2)��јt�����{��eQ�L�đW�pYY��VH�*0�J�Lǝ�ʟ�����T|������5����}>d>s�eY�V��^,.�񁲟g���S��]W��<ξ����/�~�"��c���2b&T���X���(�a�Y@�x�M^���� ��g���	6ާ��u���o2������8^`b������	[���Vk���)��5YݺAN�W�}�I#�eSM&��|�
��d��6��9�ʥ*�ze�>��N�l���eI��.-.���0��>����G�������%i^O`BǺB��[-:G�]V�����`9��V��j�8k���f��0L���>ׅ?��%>�k�1��V}���3c���<�py\׆���N�7e+�2�V,�G������\`����9]r���5�c�(� �pA�򋦏���*�n����]�E���m�:�$�W]2��c��Jj�,5��*��5�K������	G,*T�e��Ճ��~�H?k��2��?�{)Ʊ.6W�T6�=.h�ZX�B��ZЋ/W���CJq�|:�da΍��A_¾3�Z�3'��IY]�PՏA��^R��Ͽ�ϋ���!k�$c~	&�cn�<�����U`8Q��uc�(����%j�t��A�h��qӄ+1H��s�f4�ڍ�`9 �"�B*Ő܇����9+�	���f!�̨�!�D�m��$[��qqT'����Q�<Je<3��@C��K��3���u}�ghI��T��G��u��1�&C���n<�����f:���k��b4�p�R�X,��>[��3�FUx*}h�Ca%0	c^kj'΍��c�����%�p��A�������ƽ�XB����>��H�������&���{��q����]�B�)A���+8X"7w7��"@@т*R0Ϣlx����".X`Ь֩���'�|.k�p����l�V	�I�ߠsfJ�x�ꋦrf�^f(�e��ϟ���:G�z}o8u�! �eM^58�8a �n$�S���E��1�8b)��ާ��K�h�y}���%I�V턗Tor���E���F��5Oa6�,9��ٹT!-�.| ��Y4��*H�stbRv0�st�5`�b�.:��D�fhk?�>tI�̗B�dAu⦧�i�M" � �USSM�C3PC�IU\L���ZW�T�<(���C>],�]HF���{�$a���`�H�nl���5�<��HnQ iT�4N֡�]ܘ�+�u'���1� L��JbәI�z�װϹG�9�cHMLE�,��)��E�
9��'���w��<�f��^���>Y�߻���_{����	x���6n����k����;�Pc܃����g����F��5k#�^��C�7(���������=����<Dt0��q%1���	�fl��P�]� �����[Yݔ��ޓ��cv�����ב8À�G�M�`p� R�_�J�Ά���:8�<���K�]zKk���ۤ��׫�;���x�ݘx8#�zY@�2�����t�#sj �3�2�.��, e!�:(�[>hw%�q�q�܈~�c������/��rq`"�XF��̜cD�+�����##���	�pĂh�׊Eǹ�@\�ɘy����(t\ 8FfԤ6��,u��k�3d�k՜pI�
���MꝠ�0����0WJ��g[2�e)7�X�Rg�}n��'dG�d�s�HW�י�����1���,�-Hx�!1��� �p�<F�é	��T���|�u_jY�`b��d�`}>O���05����w)�y���z�^Eʅ�\��Z� ��9�q���d
E3���;2���z7�5�)>�%�2%��+&"�%V{���s�x&Q6�썇��Y��:%�`{0u�����~~��e������_|o�N�T��E��N̫��MI��t�E@�@����4ωSM�9$�s�L�u�t�rqy���EK��`����l���¨�U8L;5D�}=$0��������H$��M!T^��P��s�&��	����~�[�L��l"C��Ma����\�Q�G�<��7��1�^�ne`�A��r��s+"@�,��m�X ��K(Nb;q쾸:��)�`=���*"����B���A�V=��e\�Pe�i���b�L����_z�����?�-���~*��5=��@)0��m�cLu/�z����V��Z��%V����r��̏N�y[�V�\��1(���l�1a��%8=v�D(I
��Xי�ί�����a2cg
N�	��\��}|�^n8�}��~��ptZ+�I��T^�-����!q[�6�c�ꘊ�J2�ˀ��8��]K�OO��X�M+����J�r�V�ʸn;���*��A�%����cL2T!"0��:; �h.Mn:.�i,E�u�W�ߞ�?�c/�id�*��,5�����K�S3���N�{l	A�dJ#���Ui����\���*��0�|olOp�����4�B�=N��S��w�� .���K�f��e�ND�CN#L$w=��;7�g�\����A�� �������L��V���סD�^T��%��z��3d�u?ث��x�= t;�E^�q2>T�<���#���N��>퓑��Ѭ��Z yB�1�ޜ���%\RA4Bqt�q
%E+|%z}g:�g�`�+�ۗ;#E�C�K#ΣB�c���߽б)ꩬ��^�$,�4����dHsD�D��@_7�d��be�U���8-q]
������:).��||�|C��������L&��}Z�r|=)`+�Z� ��νX�x�@�K�<du	�Pˠ���]��Q�k�x�Q��u*�=;�N��<rq/X|�W�V#~O�oT�F��$ �Q@<P���*KY��f�
l��U��d,s#Te��.���m9�`��t�9AV-�m��%",C�/�`���V� x�x�J�,�i$3���l�
����k�A�L�C�[�Ѝ�\?�L���~�jg1pվ���{CݜG�&:ʀ�8�3�"�B� }��7{�i_ʍ�ˋ2BKƮ=�c�(�&r������5�. ���ф��9�����YW�@���C�2�]'T=ڝ.�@�Ž3�8����*1�ب�@t�xρ�?6��Ɍ���
9��%R�	�	�/��#�4b����G�؏�==Ǳ&�<Fr|~&{����ud'u�I�l�@R̊;6(ȑ�u����;����e�0� ��n�w�5���'��B�~@'Z@�J�@�ڮ&�|JAy�׃�3��BЁ��-j�^���hRv$�W[��H8���<ѥ@�	�������y�捬n����TC0^ڗW.0Gz��zW��}Bрs�,j�s)���tgSv��@�ԤI����|F�?$I��Zl�t�?���v����JN1H�1p�~3�x�|f0Ab�	/(,����pj]���\�E��|�d�ư�!M������=�"���X�YO7�5������?��+I_痎G��83��h"�_�����w���oժ�����AA�g���R�������)���,����S��6�H�ɼ�3�1;�&�N�d����o}�;��g"�����*�\N49��ˏ�X+�O~�S�@M���#�MGl��R^�w���LNu��阂�7 ����H1�W��Z�J�*�J�h$e��܂9,A*?���T���akH�ܮ��x�H
���-,f�=5e�qOk��E}}C�ɖ^�mM�劮o%��^ņ霐"��� !tV�:�,ƺ��+�G��;��8E>�D�aC~.���q�Ċ"ajjpV ���r��a��ڞ�^1�r��$�.Ɓ�e���������h��R�X ��f����pd�;�א�*���l�[���������\�$\�����:��n?&|�r��doÏ<?�V�۞n]"��8F����MM��(zE�Ɉ��2t��84�:���H B�@Μk��."ɨ*�Y2�8	�$���n�� �(� �o5j������|��C�\�چޯZ�u��R6sD�[�n���Mi�Nu����d.�I�e���p�i����o|�|C��F����ǃ1�}��"`��-�������%m�b�[m�*���"[G��-*AZֿg�!�csɿv��������?Y�����ѶM\��Y�茲M7sFH)[�>)0	�@��x���ض�LT�� A~a�E�/h[�x|��$7��.&3��n��^����
���T`jy"L˪4���b�I��PG@�c��TX*HW7�b��u����仸�r�c`l�����sy��ܺw�A��[G��5�+�mA��𛗯(kZ�g���p"�}��iP��g8������䕾��[;z�4�������ryv�����kU#��{oh�A�.�}4�O�x��`�����X��dk{�U����D.NN9����p�c{�쩬�֥Z+�1�Xϟ>���}���/�K=�{#��{�6�0q�=Er���1�RɈ��a8��0���u�*�;�L4yzM>JL�uN9�.^�x&w�ސZ��k�d൞3�+�z�ORί����ӏ�
#8T ql�����ݍ�ϟ�w�7�C��hB��4�Hk���ߋg�����l���4�|��\t�R[mZ"���ە_��Wt[^_m��5�I$?�"g��k��Wz-v�h���A�ӗ/�ߕ1���ޡ���9�p9�sp����smcM������u��^�*��oe�3�����Y��Brm�z�_K�����ɳ�CB�(uq#u�L�U���/T[2@G&1Gx�JIǻ��^��jY~��ߔ����5
դ2����B�RE�B��㢉 �b�Zi?$���`Tad��$����grS?�q�"g��Q�қ�/��3CH�J�U]0�ĸ.$�꺌NYU�ɽ[�%\�����z�w2� ʇH�t`,Ԫ5s�u��I������!�ͪ�տ�y��s�<�d$ѹ��S����-�Q_����a^���*�Ϗu�hJM�0,A>V��t�}EJ/�LL����\1t\�L7��51�Z����H��&#�k3��Z��j]�u�{]��.�A(Ls������&�N8�L���N`N𜉳���9�0�r����-8F����DƗ�,7���@j$�j����j�a$� @��8"䛹j�竡28�?:Ņ���q�g��-�5�0i/���\�!=�ĺU�W�w��d��Ä�a�\n��n�w	f���e�{�p_����<�P(,��k����|����a�ٲ(L�ID��2��zM*�ޚ����G�(��J�I\�X�`R���#�$r��"�ɧT��$0�s$ϥغJHR�Ʌu�c& ���X�5��l��ӒR������\�����50G<9kR �"C]��0�����<"�1���T���'yb�����e|k^���=�d^�ISh�+ry.�
/ �J7��%�")���̂�b������EΣ�UjIo��nR�B�X���G�#���O���4��_(�p6=j�q����L%t.�)�@��랋��ڢŉ#��|�=�%u��Ȳ�o�:@F���OdX��xe@�oH��ҹPY�D�Ϲ�]�����z?�u/�^^�����H��H��.��DN4��k2� +�1������ѾD`�����/)�י�
� ��/��Nw@�~����׿�EΌ���H7����rzrN�Hd�%� �|DW�Սݨ����)��?�͹.+������>�@*�:%u=�	س�O�� �Z�`!dbtyy)�|����m�N���/�u��詵S/ϯ��'��hЕZ��F��o������Fnӝ� ���$�KE�4Iz��.��,�@����f ̠J�AN]���D�./�����݀ோ1�D�yA`����U�
8Ì��ٳgk0�s����{��իW��ن������_$��&��&v��5�J�
��'��R-q�����NG�; �����=��q���&.������R�1���~��n� x��g�����X|C�	Ӕ�1vR�	��꼩齛A���W�����5�hBFӨԙ'�{A�qOc-�,��7dK� C3SE38J�T=�!e�`I^��!+e��3�p�qE0V,�q9��P�<+n�ߕ�NK����i�{���u	f#���䦐Q�.]��&�u Bxh��7�6v��6�/]M��G���	����Kzu��V��|b~+A�2��8'�BB`
$r�UM��B�C^.g�h��D�G��'�Uq$��\����3���s��jib��Q��iB���� dh]$UK@�_�����g4�?F|/HC�Wstz�d9�Lh��8������,�b���	�*��Wu��8���RY6��PZӠv8c2��z�Z�=M�~�A��Ll��5CTJL�C���L_���HQ"75ND6�� �����X�H:�Q�uMK��↾?�q�Hs���FJⱍ���(�	}�B��)��x1gw�H״����6�Cp�����)�[��^\�V�<�t����ԥ<�ΣrYv�mn-%F���=^O,�
�p�y>����N�B x����r�,
y0EQ EI��P��h1��i^{&E��,���>/�����m��k�
�5���uJg�z�Ɨc篤���'��P�iM�����~ٽ���Ǐ�O%o^��b%`'��Gs&�຤��q�\?oH�!�F�h	9�6y�7��/�.���(����mR�x�Ϟ��Ϗ�d���T��0s�i�W�f�� �8��L�u].NN��%�JL����ÐO�A��(-� ���
��O�#M	�񆕗�bO�~���.H&�ȹ����H#�;@Є�kn��Ą�7��uc�bzA���xJo�"�|���;č���*̀u��|�łeAHj�\A��Qh�Y�ΤNz�Z��
���i�YU,�)y�a�z�=��(̨�R'ȐGo<b���B���~F㔂���rt�*$>ib����م|���s�����e>�d�Q��hjb�d��A�X)�:kg�p��@���gY2�h}Tҿ���I�p��� *ԇ"
Ȁ�c#V~,_|񕜞sS�q�Zv��*�f�$@�㳧/4Y8cR���\]��3�4�Cv�1^C���s���q�3&��+W��{x��4�F2H��}�;����!0@���� ����dHq>�j��@�b�"gz����ׯ����S9��h����۴���k��)�fNj�>���3�
2x��O�8����Jϡ�`�`H���� b;9�D�KM�K����C�������T�:�H�� �;Ԥ�Ղ��}2��K~ ��O��UK�ޠs����t�j2��G�!�w��� :9��˴o��e<���7r����ԑ�V����3�̉<y$�EP�.`j�8��(jJ�N(j��3�8Wz��5���X	ul��s��A>@���!��Q��R�>�H�zWr�A����r�Yg �`Ul$�H�㕺�|c�� ���G�2?<��Σ�ե�ι��\��H�q���	���l�V�������/��/�=���Ƀ���<�ڑ���CXL��T�ziUZ ��.��"�bQ]�蕾���K�4Q4i�5��w���+�4p�pZMS���W�E5d��+�֊��H_����/����0tu�Md4�A?ۑ(3�N��⺀q���W =�:�43+��o��w�c��ߛ�6)�5��A�V�T���`$��H�_���H2���{��Ay��7tB���t6��dfJV��0&�ҫ���[�? ���d�Snև?�yt����B�R�����dk!���
��8�]��G����ǿ��}*��9��T��Zo5�}�S���ɏ�g�q���H>L,6��8�����~�]R�&�u���~���I�[|�0\����������B�����gBX ��I�l��!���\>t����D�v�b��5����D(Q���#��3��m�pr��c����q]EU��	38h'�6<|�\>��|���Υ+3�S�!����蚑��OI�Tj:�c;���h�LVLf}�8>���p��ߛ|�|�F���}��y���J�]��H-[N���d�1��_���\�Zc����(��{o�$Y�]��7�<�9Ufe���U��"@2`�L+�p��6�h��� mD��i4�"�F ��Q� {����9#c��ߤ{����/�
-�$3�5�ˢ"#��������S��U��b����X�9yu�ƺ��ԃK��d�\yKV_ĵ��JLX%k<��M����l"�Y@j�����!���Lp7Փm�Θl�@.���U�����xܦ�r�c�E�U�,���K`�T{a;Q�|�N
��%����z� Y��yE��(��r�æ���Z�Kqr��&*�Ɖ.5`M4�C�P&���̩p�r�r�` �h#� �g@Py��'�n&d\�u0��ZLA,����f��_�z����C�Dp��A5N��Y�J�f�n|�I��r�
|o�Q��X �4�^gMv$��59ju5H(�6�7��c�4p�xu�0�3A7;���ͬ�rtz���%ٴ���5?wApK���� -�M F�#V�0�@@R�mu-�4� �C���0zu��Gw͚-������Q���f�4Y��G��� "�6�J�����#��稐�!�N��qt[ ۚ��d�X�;>� �s0(еz���D��ӓK*A#!�S���@���VC��ltY�/Q<���T��0[�^�S]ϠS���$����Ŝ��:�CG��o�J��LB�0�5Ns�����Ub�C��9ESFd�2�a�8O$VIcgWn�]n���K�x�D2����c��*ÿ����_Le��J�I���ߗ���m(�6F�����(F�fs�5������?�Sy�W?�H�D���^׶^Gܳ)��[Cy�� Qt]r��m�҄�'����ӏ5 ]0�[�Kg�4i-�����\��;o�]=V�ʾ����v�@��[d�"m����ӟ����?�#ib��T�z� �؈��]�L�������7�%�oݓ��&u�䞞�Z�sB��Y~�؃8N�,F�.��	��5�G4\�� ���4�Nmd뽁!s7�ND�N�Ά���HgS��<��Gr��C�k�~[�.�
����B�`G�3�x�Jc ��GE:Om΀�S�|�sӗG��}m��!@U��HmI�처���]72�i2���n�R�D����	#s��L�#�q�ʜ!Óg��?����K�ÄO]A�������O9`��{C��{�O��>w� nyVݵ5��RQ~��\�E�����iT���X����Gj�U�-���u�9A�������TmИH�T�>[�KI��hK�9"ȇ-�z H�x� �׷IYkP=�8��C��B���BX�H�t�M4A��_B7E���[r��}��������>��W'���.
�-f���� ;ݶt�X�8��v���p�PJK�|����z��p�QU'�(���_&�����g/���/Ƈ/��l��!���N#��B^��,��ЗF�& B<qi�7pu���F2�pF�D/�D�cR\G�b��&�h��r���:X���MրB<�qL�a��A����"�y��(�����gM��&��X�]Xq5�}JZ@�u�&Q��6H��P\��qH�ƌ��+�0�cd�V��(K7O�ʡ	�0�A���
�O�3
H8"�aEP�Z�Ʋ`E�8SX��`���a��S�z���"4*Pf�cP�Du� �g�*i�~Z���8B3 �JI�(��H�A�A;n��`��m�*^����=ka�3������+ÙC�7F�Yz��б:	
G��ST�Q�S��	�������K���Y;T�b������Wl�p�!�|Nx�A�"�+�z�� n�u���t��TQӕ��FDn�L\��$�D1O�"ZP%ɪWIWZ��U�\K4��UU�B5��fP@F-}�2n/]RN@.]z�&:t@%�6('TCS�Z��U��A/�1�N��vL�\�L-���kbg�%hS��*l�樔q=5%��0�2C	��a�#�\u?�P��g��Ӗ��H+<2��m�zX8�27zXH��+2ס+����yk�m�o�+÷ߕ���z��?�'r9:�8L[g�LNFr~q.��wnlK�I�R��|o&E+%d�!=�M���-&� ��%��<{��|�ʾ^��n�I&5�y[����W����'��[��"�������������kB`J���#��L�ܝ�p�f�I_�ZU{�
Uh\g$K��Q�+�0�gr��<��OeK�9$�Pxme�`K��R������}���3>rz�
��ӟHq���u"|J�3Smգ]/Kt�t�%\mz���j ���\�f<�����H:v��v� ��Rx���E��'�qC��%>:��:jZ���(P0��`�	a7T�SS��P������,�@#sl��T���r1���O51YQ���w5q�pv����$x�����]���M
6��-�Lr�+K����G��@?��c9��٥���#}�&��j'�Grq�L�O����y�I�kc$�c�	�3��n����[��s�e\�b���q}f�z�@H�A�|���}:�o�/AhB�����������DF�\�N����G0aR�'M�<>/�(l~�͆�����`���٬B��3*�h�� ������ղ"7h�j��C��g� ��s�P��:6ғE�:��uM��/%t`�F�G)w4��u�����Y�� �C�|��]��ý������ࣷ?y��<� �� ݵ��ĵ�|ez���1�W2܃�tV�����ژނ�Ƃǰ��c2d�Ku�D)�a�r]%(��&1
�@*ѲҊ������ss�#�Y��>�`���� X�D�b�(��E5������=��d���C^��Y�`ؓ���4�`c9|���`��_���)���TBa���}2aE�(�ॠ��aG��� ��V�g��/���v�`
�xA,�
+RBWZ�d,F>6�/
T:�T������$V3��\0�����٬a�o��͆+@�*���Bh�g6(���&X~$������'�si1<*~T���/ ��L5�luc�q�ة�r�<0�\��50�������� X@�2pxt13@� 3�u�\��Ht��e�;�&C �)T������j0@6�_�m�ƊI��f�e�9y�Kb
��I#]�����!�Qa�ꑉ�`6�/����u�L�0a�ǳ}�[�A�x�Z��	�}�Q0ڠJ۪Cl08ȍ��;Yepo
�d��âX\��n&�T�6���h$�;���pR�T�M���a�i&��A	<����J� E��?7oI�[�y���&}C���?����Ϊ���]Mձc�8S�AEQ��d!tL��,H�88��`�ඇ���+`�ɗµBP��+
�e�÷����q����鵆4�9�~�]y��#��jR��^����)��d1�-|$�1A#`+�K�m��D�Bq�+M"ƚ����cJ�
,�L̡S�L6��ї��=M�z��_m�۔�et�y�kz�B_ ��Wo���3��0 LL#��q[.��llc��z,tw�4c��$�H��[F�Jm�$�i���0�Ѩ��i0�ܖr{�D#�l=����aK����kvL1����)
M��a�"�N@F͕��z��S��\ƅ��"eᬳ�%{�} �w�&m}�B�8�~�7?���#��D���?��7e��v\Iq(z 6�0e^ت����]��1h���t�"�I��r5�d$��hr:?���K9<<�Kt7�&G� ����zת̕��hA�8����O�O�U��,;��O|Q�kj�����k�C������'�'���|��7�;a���)����0�U):����i�+����a���a��t��^e�g�sA���k�}Y���D�fn��F�9o�.\�V@3[�B*f�-+ u�V���*��pu>��W���u
*�+_&�����������}���� j�bB�?J:�%r�떻a�V��P�↭�C��P�l�Љ�6�û]qW��pS;��[�E��Νr�)���W�}@�1�fHB�Vغ�P�`�JeS���Ϻ�YL����g�_xmkI��7*f�����Fwo[��QG��p��@�~��>YP�xy�R��RFx+�p���������;sB�ru4�Z��J%A�?�C��%�2�y��x��� �� ��P'�`׈}����X�x�8b�0�
��a;\��m�܆�Q�f�[,@��;��0��]8�&p���؂2:>`����0
IT]�ή�}:!&Ox~�����B�J[S�=8(���Ħ�ïax��8ܐ4!��cb��{� �a*��0�ɨ�R+L@��p��&O���ֽ�ݠ���} ������Яy=v��(�!qT!Q%ì���P}/��=�1L$!UQ��q��K�:��)J��"xǽE�$�VF���w�*P����&D73c���߼pJߡ	�A�6�� �2ZH��D,���ޖ�3�gH��峊S1��F5C�*��m�������\ցMEiCf-��X�Z=�@��هdkS���d��S�����;�f��J4�ї���ǀ(�	,"Q�p1��A�`ف��濱�����r��A��H�f�c�c�$�%�1NŹa��P1oҾ3�3\��$�mwm��KN��(��V��`�/iG�M�mo�ޕ��K�\�KӰ<n�){�_����:L/5I(4xirP8р=¹a����Ы �+�AwC�����2���<�AVS��y�ǉK�1�ٲ�%��G��Wl��d�3*	�ޢ���4��v�.VW��۱^K��#1���Yj5�pΧ�<w�gۑ�X�H�9ǂr���񃡊�]$�K�,dN�����M7n�����@����R�Y_���V��_��ÿ���*-��}��S��{���>�:�p��b�B%shT^qx���`��e�5����������Jm�2�L�a'���	�e7�,ᚁ����Z��.��~��}W@������D�P��Y�իbh�}�7� $ձLu\�g><��p���L��ύ���Y8 mm\���p�k��,c��`��
	�+�W�Ά�n���BvW+�jEƤ���XO�-��Nuz۲��˖���x�95ve (��j��"��f�Ot1/���z8���Ǯ<ූXU�S���%	�$�nЗ��w?<}��������������L��6(H�96Y�i����4�C��P-h.Q=$}�\�pCTm���JB��6M�N��i��kF(m-���h�І^Q������?s�f�a�ך*���o`5������08QI�/\2��빛�_K�f"��������6���8Ѝ���-�n�͛7e��E|P� �;&
	Y	�X�i��rtr"��TF��!�#������뮪�b`����ʌ��� �+W��-^H��+��+c<*�EU���Vy1$��?����&���F;3c(.�S8����j~�*��4	ڎ��\`�'h�"0d7"e`HZY���~���a���h�3�A^��` F�����6�@����v���	��XX��:R�fE7u�G׎EkC�X�!i
d+[R�F���r��31��Z��~�{ �9U'���uop���}�[�4!��p��i!+��)\(�R�YPpN)��!qt4��S �dG,f����.XEx���ʮ�y�Ҝ,5L��i��I^Pm8I,��~Gs#6�d!�Ha�յ�9Y��p�6�K���(���J���X�ןz���8/��L�
�yn5г����TW����;k�Or����(����sA����c��Y\'>(!D�H�\���3I���GuQ�/�)�O𽷭���59��h6�����H.50)�6�)6���Kv!8���:�L�$r�64 x�oJO���\��S�q�E��/�^O4��}�(!E�"9�L(>��.���w����9x��d���gk���`�!��v��2 �%y�E$��:v�O4��y���׿-���w�է���_|O�>���)�����j4Cء0�$�!$OHb�w��ΰ'�^�G�ȸD	���p��D�\ꑘ��	�Q[r�B��L��J�1�����[,Τ1ܑ����H{�0���JA���/��)0����J�"�\z��{Y�N���!��t�-�.4�o��=w��`��̗�o��u	�!֬ڌ^C6����ےln�Kx���M������x!��O�-������W��C��W�QL�g�=w��LF�I`�jk��7r��H_9��������G�(P0���߈�������oA�TsN�\����$4���� ��-?\�bB]59�C�n?�E�X�#$� �*`r��7�8Cv||�D�=��yT�M����yt��i%����H�Z�4�+,�	� ����v7���{ݍ(�%�F�N�%�gS��m��ʼ!M���������&����&᠍e1
 �2�v�U[0���>(*.�%n_�YD'X7��2p�R`�c���/��_�ǟ��?������������}r2jv�]�m�j�ו�:���t�[R�s���8Z�Q|�@�e�KM�UԚP������� �� ����NC�������k Z�xS�qd���kV�73�y��@m� �]5}5���RZAK�vS ut-�W*+��i6�����%�Y{�W~��G��;�`S����T��q�Þm����۲��-�7��:#��t~A��c�����6�[�_�/d��0�U�^͘H�I���ތ�X��dP�����ҥ��`vEQ(�`�ۤ�3�5� �8l4����e՝��BoXT�u������p�!٦�?;�͈�
+\c@V%T���1��T�Ak�JPw��0v�"rj3���..f��kP��Eu0p�<�#�g*��Р,����v�:,fk¸Ǆk-(���b��4i����)7c'!HѠ\�&�q1�(Wn�+�V1�� 2t |n�{@�0@ib��\��%��D�	a��K*Ñ��]��P���X��A�!O�{.�[m�:j���ރA%]dR��5?��_`ծ��p�6Ǔ񹀗@u�t��%��U�K�B�?,�7؊*�))<QY�)��������O�)��0�����^�(G���I=h\C�X�XEuÜ_��a�9�]P��zb�[�w��T���	���ԣ�����!I�kD��F0��
 �b�#|�䅼��u����{�u��y?~��|�/�T���z�8&cvNV+0G���-7�_����o�������<�����R�N��49�;����;",�zO7@g*Cw��]�N��O��і���P��?��nK��-��<���}M�����L##����+�<��9[g��1�z�;ߑo���ˇ�}]v6��֛/����=��mi��Y�*�{޶*����aM����-���d��W��L���^�;�~S�	V$L)�i�z1*c�A��in����y������<�����ő�YS�(M���3��H�!���o��tol��b��ls���r�K��)�֐��h9!���O̎��r��"������f�����ڈ�^é�g�� �K3��}nH:Y
���n�ȣ��r>.��<�K�L��~�k}>��\��c��}�6���\��o�ϴ����6���B�2ˌ�L:�v���a_?CG&����YN��N$�i@9��`�s ���C��g��l�����)�}Y���=��OV䕯�8��t�`�,D8�S$�4��:�/���޸{W��?�}����'�=�/��$��_	�M��H)0\�X2�P�R�
Ax�Q���2��X��:�A�f�l���BJ]t��Ӕ��Y:�� }4�X��M��ꓗ��\^��^l�7�����_�{S���7��k�JS�^72+��<��P�arG�6��Aa2�;fZ�L
~-h�����������Ɨ�]8g`�@I���L��4
5���\�)��6��E�D�/-zCbG�h����Xe���,e��@�A�9������Gп!Ё������3z�>��VG����0!��U����&`XBЪ_KV�m8�<���aQ�Y!�$\+'FS�	�҄:=ʙ���^(;�7�?�=�d&[;�lL,�i`8��`5��tt.�l,�jrvg�kV6Z����I�Ր����, j�q�8jQ�6E��{G��u!��*J�_<a�a�&3�?o4�xNoY�R���>��Z�f�6�x� 9�4��g�xJFaI����'��F."v�Υ4)W���]3Ҹz8Ia��HL��l$�p!��14����?p�u�)��0��`�'�7��%��� V�2Kb��R�A;a�b>�1o641׃�z0E��1;)�����E�O��+���>�	������s{GD�@����j��1Ɣ2g7�{��u��� IX58ԉ�(+*�\��׭*]eް�euOi>l:�`2�\��D�n�����_K�Lj��~�K2o�]� ��T���L�A��z�Z~���a�҉IA��	�ĘFYIf.��XX����drVh���V��d&^'m�-5� #�v���/��;j��^��3�9;;� ��A6�%�'��t ���Ȓwt_��n#��nnj�#�ӱD�M��P��*�H���S�-�����l��l�g��ƘeZ�n���]�C�ysG66�y=���@fP�ı<�;����4�mno����дq�u�e9�=�Y�]!�K��pj�V�0{�>FE�i�LN�s�uL5��;2ؽ���@VH�2}~��eb.��6QTS�4yO��oQ�@��*zC�J��UC�L�ᜍgҞL%�`�Lb�xЕ����7nKokK�UC�U�<����P��i6'~
�ӹ������S)4��MjR�"A���T3�,S����Ӱ-#M����;>����ãs�̐X��-f4u��W�[kh.>3�ct�M��/&�dwt�O����X�}� 
��i��Z40�:�E���Һ8����ى'l��U�Y�A����.CS�W��\s�	�]7�jN����';�Qu��%�Ŕlz�߻�	���7>|_.'c�Fo_*�j��5����$Q\������5��:�a�햘�X�M0E�L4_h���Xѥ���(�S�D��b��E�&�K^��5(��}s_��6ak����e�&Kv�a\1a�f�-a+�A��/��_�ǿ���睿��G���G��c6��kP��jP�-j���������sqes�E���ԋ�T��W�n�bx4N&<
� �ΉX;�?W��)�'3���,�q�bJ�-J����xkRo��%�) 9���b�D�%r�H0V��(���篒��W5,%�+������U�
� f8�KW������ 2�M�$ll�%�5���;��}~�\��$�|K'��ۃfL1�Tb�tE���r������)��]��5�U_	�>�%���[�����������}a�� �@��q�@t�8�;6wL�!N9<)G*]r��U�.ַV��s����D�͙$Qf�j*\;��4�� `G\� 8*��bD��r@�jLZp�NGi�&S+'E�W1���B���쒆�ێ� 2��q���rRxI�m� ]���ے�UG���P�ؠ�c՞�5�Â�c�8�/h��8$M��  v-��f�Ib��m��N-(�6,3�?|����37~E0�09ځ���*�C=��ɋ1.5\ײ,�Z���9ֱ�j����I����֕J$L$*��\�� �a�K������Nk���&�G��s�n)�5 G��s�f�}����l(Ү5���`7��&������D�:FEj�-�$��qG�[g�qt0` ��ԋ��Z!1�xF�ego��Y��d��uc�	�>�Ya�� �qI����	�̍��Ve���ǩ&=�^�,D���.�si��t2��W������/[	�H���V�>CW([��j �J���ƀl�D���/GK��)��&գ�����B��lY�~kS_���d9�S�e��My�[��vO�E��k���y�������bf����GzmO�$|��(j��.�`ź� �W��Ct�������,����
�c��~�[��{��m>����Y��{V`S!�=�kD�󂝘O�u�]M���D�3h@��O���`�ՌX���B��Q�i��z���G���c��zAi�z��cqu�w>?Ũm֚W{5�"�A� L�Z�,�{;t��к�����ikr{_�~�-�ވAL��!��B8��g����t����NY��j��=��V��u��]�t��s�8���,c�2s���R�>��D����v��M�5H���V�.� ��eT�jn0 �`��ǗI���ctq�9����$� -"e���ԑ,gl�a��m+�����(XK�{C�1��|���`�[� �sTp��^�̌2����
��+n>#a��9[��/9�����^ҐN�&�W.�ҏ�WJ���� �Ћ��C
EF)�-*�.�`I��� htx�,���n������y&@���sY���=�g�s�U��J�ʲ$2��Sc �N�^��D�0⬾b�tYcɎ<*��Xp�3��I��J�1������}��ye���_/�{=�(e]��z��U��V�b7�L���JXa��<7�;�z:�":����~P�sO�ZXu����f���[�}��U<_����A��nQ��{�e3&��A,�֖^����@F��|��F�/��&�W
w�n��+
�u��j	CJH f-p�-�7aC��$B�z�UdCϸ����0T�!��mo9�pi-f>.f���D��R��d��)�E.�g=_P������:��u��G�_M�'���VR[C>P��J@Ř��AN�7*��o8x��uIA������x��<XU��}P���j���t	�?������7
mV����Q_���A�8������Zf���n�< E��.��i�,XB�׶k�B�ian��|e�X�o:�1��, �{����.@�g���mz7�\�N #C���_��]Үt�JP�E�	*4v�Q�,4�pO�s� ���M}��R���!�j��Ӌ���P��:}I�-jn���2�i�.�`�1�� �tvqp1�Y8�<	��Pє^�+�V_ڭ!?��:���酼z�BNN��uKd�'rgGd 7�c� ͅ��	^�0�U:ϥ�IA����[�����9?9�z��&M�A���Od|y�m%]�HL.G)1�����;���l���P^>�u3�=Mތvش@��,\'k(�Ac|�c��ӱ���P0�O5)��@?���|�&l/�^E��l4��9 6�s�	v�t�_8��.a0{{5!�]#b�����`���[�m��$y�7�����ώ7�uM����m��Dr�k���]����C���a��Q�W|��wLպ�����G���S�v!�Ιp���z�z���"��n�g�q�J�H
�P5
^�dWJ��a@3��O,�j�zQ�f���f=��L~��ˤ���*惢,�`��uLB��L:n#�������wx���pF(��Xu�S@J/��gۉì3�F�%�
6�/�c)��8S�/�Lg�P����c-!��fCY��q��N �{�q'!q��$�2y у+�$kCc?�n�U���1�@�۷	˸�',�Ng��L�x��29%��SV�H�dU��N-pΌ��ȸ���z:7��o�%-0<�(*��frK�Y��W�����U>�$I�Q�,��ښ􏺒�Ԓ�q�ZYa-]Y�`'i-&䶮����؀l���J9�*������
��i^i���l�;��턹��-q�۬@�R�2L4�����^���xN�UL�Q�qiB1-5�:���m`�[Xo�A���`������-�����d2^�����]�pؔ�wv�ƍ�ֽ�@����kB\�v���syu��bl�G�9.�"R�I&o�sK����?ؐ�������d\Z�D�O�YH�a����uk������v��k��q����BC�|0Q�"����"`C5y<�k:�`��kz.p��,��<���+�/J7STv���*�ơ���c���!��.��;{��t��Q��N�aS��eo�|�>-���-�V��i��`��|�]���X9��=+
,�"�p�I�S�#(2�����Z!!Ab�g��X"Ȁ�njp��$�k0B@���@[�� {���&��ۛ��,�8�=�o~�R[R���ؾ�q���hx&$��wY��/Ĺ0����}{�%�����0��i�։e�3f�3hVjۚ�Ag+�+�7����
a��nnd�@�fbC5��'���ޤ)�|,݆&6-���?@�d��SBj����L��@�t�?O�usK64	h]x= K�ֽ�dj�zo�i!i��p����g�������c����,�T:�&�6jk�U��a:Ib�u�
tH����c�E�
�!���t�<�Wta����ªw�E�X������rg��&�;~����|��a�u��l��s��tv�`gM�<���{�ڌ+���-�^�Y8����^�6�ݿ � ���?\{��������X�IՊg�n�Pי�*�ָFTu}�A	�6Q�W�9�t1�uoE.\��uys���`Ƕc@'����_��2)�5|QG�h��8�n8�J��=N��$ױ8lv�*��wd%�zP�a���q��w��6�IH-�8� a�,��Ѳ� ��K%^V�f(�U�cZ��T'���h[mX�� Nz��������ֆ,^�R��v(�,�ܤ��)�Rc�ܵ�����>ԞWUB��<�`dǓK9??���Cih 	�|5��ّL.��l!��j'�y# �яr�ĈK��BGV�0�p0i�>O�<>��A@( &@ٿcR��Ie��s�� �Ԫ%�.Au�d苬�z無�5��O0�1�M^��sY���	+5a��'Ђ^
�e��5���d��!�	�-[V3E����u;�c�.uiU����t%ϟj75�䢡N���r��d����4I+v�m���� ��)��J��?�ӓ#�}�|�[���~_�7'.�lI��76�X"[�vIK?צ|��<}���7o�%�������?`p�P'8��5�Xj�·��鋗�=����gpN	Oi���^��r*�;�|�ݻ��or���#
��A5A��� NW�W$.�[;Q�A/BQ=��5����^C{wD�c�6l��d���3�M润�R����f�Y�	�$"u�S�J|h�bߌ��.(���!I�-XQGP�$a���\}o �ǯ�z��@�'�� A�p�I(�S|��;A� e5�|<��8j5�^��!-aG�M�c��%��Z⃤U�7�e�����z~� x��̩KS>�7��i�Tm��٩��<^����rHQm���#�g'�I����s��x��1��ϩ��-�]�]��-��Ӌ��t}�4�-穴62�5���dL�L��q�:u�w���fN2�����/%@�/ӳ�8V_��4���H*�V�/cBJ8�K��&�]��c��1��5�)�׍)�0C$y�3Q��2�����c��������l��xАM�n���U>��g�szƺf	[�$����Kݳ3��q�tk�;�� �qrz�q���ݭ�<��	ӓf4�t��.Ql�<�|�X�����.�틵^@�( O$�\�g�a`�kT	�y�TT��j������ux˺(a��\!���|��(�%6G�'v�<J���[
|��l�ͻ��:�^{����_}���Ǌ���JHP)s�1s�	��Fi�.�	�*޲����S�sJ�'����޼\S*_��u��D�z�=�L
~�EZE�Qh|�X!�m<�XHZ��f5&��UY��'�1A��:[��=����N?��eX	� �-+@�!XQ�k�|���k-�cJ�1�H���}�r@�)�g4��'=2T��9���|�7�!���<;:�m�c5*Ӊ���\n����>�a�����6`i�H
�m��rÙ��U�XN�g���P�-�pe/�R����4�!G'ÊU���E�9hV����^�>�	Z�ѩ!���,�UT�#�
L���lR�׉��^����	��|jA�������Տ�O.ٱ+o�R��,��
`邁��-���d�(�Wb�Ѻ�S��uH����� �j�;z�#��O�������z�t*��t��?����T������5�(�r��kI퍽]��ؔ������6�w#i��x)/4蚧�W�y����]�b�?�egG�����j���r��x�ۗ�����P6����p��g�����=,@�Rbk39��!��n�ا>}�X��K1@Z�u��i�����=��^���������������r7kRu������!`������յjÀ��U�3�f�y� �
e��<�%� �9M�n˄	C�c�E�`�ѣO5C�f�1y�z?���܌��X��?��/�ɓ�/��5�kȭ[����k2��H��#y��TN�ǲ��f��';�mW��Q%�p�5 i �'hg�	è����yV�������%�B��r��RX��7_�db�3qnJ�/^��gO��I��ޞlnn��NK}I��<�|�vMf� cSK� ��&�]l2�*��'S�_�%ѿ!�oBUT��������WO�hrԑ��&6,Mt��V�Y�k��0���&��'���$���?jR9��NC�|AS������m�C�'1�z���>�2᫘(!�Yl�:0�zC�S�^��&���O���c�.��o��W�څ��6 �lJb�L�MWߏ�#K�Nc��c��'��Z�L�JBKm�56p�K�ѕ&3ehb�L��p'D�p�p�XPXjүy�|\��d�\Rͳ�2�0^>X|�=�9a���gX{������+������p�u�-�0*d��bU@��ڎ�EG�u�o),�y��8tc�ĉ��JE�@L�`]��N���DWE�
��XN@�V��U��;9�5��HS�ߕ��O؉�|I�:Z�Fd�y���שjڜB�c5�11��ʦE���rdUa����6!�2)��|Dq�h�P �Œ*6^�>�q����ȗ�QgcQ��\L��p��Q��}�����a\��nC����h�0,�k@MR�WW_3�8�5�)ɍ,�&&�"�'�A��YҒ����E��E�+n�&{�����dԎ2�KK7+�e�a����W�Eb�����k
�U��gurh뵛`0	���j��r��-�~KFq*����u�0�v��E�.Ϫ�Ll��a�q��A���"6	8�8.v�:`�8S]��^)�0��JX~>����AQ�fe�?�(���Ǽ��U3��AU���xЫ��C��0��}�@�~p_��%[W�"W��������5SԖ�0�/�D��d0l���m����g/�ɣc���t+c�`E:Dӈ����l�?q�A��h�~��q&�H��w>�}��l&���ࣟ�A����x@{O�P��f����3��G?���44�|t�����ޕ[76�=h�������Q�S��ς�gg�!o�qS���Ć/?��B�����j��uX�Z��:j�����}}��y^�x��K��OTI��w�E�ָ�j� C��s�N�*�r>������q-�+	�n�M�� .X�����ooS�D��?|���4XG`ՠО��u�svs%`}�s�>�b'�3R"��7%jv�S�J�jG�V��y����~�%o*�K#"@�pE�&>�*��Yd��"M�H-!�� �IU���j�����ϠrF�T�B��뽽��kk,�<�Dz�-�mlK�F_�6�F��::
��`��-.'�ߠ�����Bm7�B���\��"2�b�$��FQ�J���Un��ґ,���T�&��޺��3���>BG�=�%��C��'}��h&��cypx&�_��"�Q� ��&���>�9���/���s~͏�epkW���{w|0�Q$�@F���RƳ�d�h�dY���^I����ݞ~[[�pY��u�`��LP���l�Ͻ^O�Q[��6�m\������A���2͙\��$#�İ+���G^��/C�����B��3�]��A��59 �X��e�����$��Z�6�bluf�B���j��a�b0(!:K�d��=m��
���64��"�j���͟Y��'�P������m��dW��{b3|B_��O���d��0�'+���2�tL�ºF�CFպ���"tr|���݋/;�� ����OѠ;0d�����'l+�9E؈X%#Àe�6��*�n�zJ?	����Fܔe���UqK
`H��Kk�y���r�iS�i���Ԡ5ڱl4[�Gw4��j*�Y������ݑXj��3`ur�������9���_�%*77vD64��۔�U�0d���l�7gd#W�0>s���݂�bT���!��}n4�����������^���Ʈ���t(�ٔUT	�������n7*�5Ԡ�F�Fq*�����r��&��3��P��Sv�
���4��e�U�#��u��PI��pVe�B_!Z�u�TO2�wx��	ѹk큧�AK�hr8XX�.jp�A͝�-V`(<��Qo�ʅ��b*� 
���"��!�JGu����h��t>n��z��q�X��i*�?{!��/ϟ����f�0��q�O�����m�������B�<~�	����n��ǳ����X~����я1�eJq#ට�B>x��đ�G��/�ŋ�_�:/�rz2�=M:�����PG|��P�d���*s��v�+����6�fz^����2.�yǎ2��u�BVa=�� ���bZ#2����^=1����{�����žBp�`���PeC��-���j���E�Ve�-ɪ�[ T?naԱ�<o�,��)���@���������>�X�O���_���@D@�$�:�%�����<t����`S(\tC�C�66�j`߫R�Q�ע���z]�vW+jp��f3<�{��==�d���H=l�r������-M|��]=VcO^���bJf�V��k��:��Z��sۿ\�z؆&��5"y����DU4�j��f��34�^����;���2��[���� ��k�=��e9�`��{2u�y�� ����R}��T�G��,%���-�
�3RrSt�Y�䧡��)Yk(����sټ[��M��/��l,Gg#��.(Hh����s��0��A���P޸sK6��"1C��H(@�� ��9��t���@A��A� GH ����\L�.�OIC�zUn�Lt1S'վB����f	�OPBm�If��uU�vk��l��Ya�ead
��x��	gd)kX��=2]$[.xgG n�~nF�༂;��D����/.q���8�?�Z�⋈���Bqf�c ��Y��{	 DKK/�h��BG��]YQ
g�hB��!�f�9���%�vp��A�&g�=@";��*/�i[.�L�����.,�X���{0��������4 ���� � �Ebd%do��b\��_&�gg��7n�����%�'�p�����ߔ:�� x��J+E0\p�y�mAYE�N�[��2d�VP4&��n�,&VxF�9�X��` �Swon��#��:��3��i�^kp��+o�o���ʽ�|�72SC��`Cö�~�����F�L�mwK
�B���NNdvrjU=��K�@�
{9jT����-�%�
|�.)`�4�+UE1"��Y�H�x�a��j�/��y�Ә�s��r��T���kQ����~^���u�A0>3D�@A�@"U�	����IA)���}��i)p�9�:��:��+5�s�"H���� |<�p���rW	ZW��s�SX�π>����2���|�I�4JM�6p�x��N��iN0�r�q�rQK��B>{tāuޣ���w����	�l2�gO��g�=��Wc5���''��v��1�	������!�OgE�x�]��=��1����u��cC:�R3]�ӥt5�}�.a$0�3M&OϦ<�9m8�O�518g�I��?��A��8�"Y��n��� �@� ��X�ޛ�/�L]۾��g�0����񮾍I�֛3�ӗ^��\OY�w,8�G�ڣhaU>T�	��Pf��a�R���h�,�bHNܞ�]�������OW[��fn�U�]KCM �f�g�T.Rf��޼��x,#�f^��n�O����h@����#T@1�F�E�ⱁ��`�T�A<*��������N9���S�!��G(?�^AG�z׌�X�;@U�M��⦞O�	�Y@�h����5�;
H�	.�BR���h}�^ߙ3�Ƞ�-��vwc�#3qER����󍍁���2P_��V\W_9��f�\r�{]�$(2w4�@22� �=��B�����h�� |�_j��t��!�F=}M�F�O�x���w�T>|(q�%��Si�z���h4���BN+\��ނ�&67�^��^��×<��W�d_��3y���3=�mM�����#y��c9?;ֽ0ׄ<1���&˚�WT�,���ZH �L#���@�tt�5(�֍�j+�)n����� �v�6@sK&�|a�k���t0%�f=��D�²Ͳ5t�b��Q�Z�V�/ĩ?gL����Bah���\<����^�H"`��0Ͻ����&K��ОY}<��>�����lׅ>'˫s�g�����P��7�
F\�D�3ŚHž:��N�@�WZ"���u5��4�A�V�8�Ʌ�';(����~�),*��p�U��~�s��2)���Q��y�W��8N��'��E\cC�k�n7W]����b��A{2;��5������͛w� j�g�a����+Gmp>��4Pc��1���47���N� F:��+p��D���)����D��򀡴v�C�$'`���+��[��~{g ���%<?��W� �w7�P�Qo8��} ��J�k�K�b�JG�F�ۓt:S�;"��uw(w�7��16��v[7ҥ=�L�j,T�CO3f�IЁ5eT����gX�jC�ѵ�b�6;�|���v�ի��˲�~����X./@�֣XQ���6�[K�UL8lx%e����Xu�U$i)m�:�X�\�	4��E�QN��s;W`5D,�62���~�Z�]>���n-�;b�n�m�������f��{$���h�~� A�<G����?�ዏe�� �!(�\�e$ga�)`p8H�`��6(�Â�*�!*�D|���lr����"�8;�@�h�X�I��6��`���) W"#}.&�\�!/����k~r8�$��"(k�;�pT�W��~�;N[[�t/^�h�q�{4d����/�C�D�n�/g�8�py#�#B�)t����5i����O��#���M��up����-�]W�ǭ'�+�C%x-1�:��{jSC�j ��1�*uF�pK�����&�m°ln��
68s���S��П�^ٹ��r�t-�$��FfpqN~cs ]�q��w�]^'e1�����*Ϻ��<r�eU����fh�T��U� �0y�t���4���5MtR�NJ�Zv	{���ϟ����hx��� ��i�1�����Tж$蒀�Xʊ��]����ᆼ�5�Z���֎t	�Il�� ���_��z�5��J��#=M���:��vI�Fi�9P��0��i)1+A��K�w�Z�"i�@n�:r�ۖ��9�L�&� 1�:81*�h�{����k��݋g/������{XYC�n�#M�$�b�&��нx��y��rr~�����z��I�G��Tڝ��A�q�u�xB��$���g��Ï�����.eЏdw��:�nz��G\cl��Kt=�ʖΎ[k��$�jE;���+������v��x�p-��|����bvV�YXw����e5�V��:����L��+C+Fn�w�����}��~>A��.��'4���(SU�*��t��,t��e��m���"�/�x��ø�Ҽ�)�M��ρ��-��R�4�'�h�a��S�i��c���Bd^[vSpn+�c�+��F5�?�Y���$�"Z����URP���]���ڗԾ��,��#������Ͻ_��S��<J�|Я������Q'|�Q�^�@qE�zy�=���*���
�U.����+2�Q��u��
�����ѳ_��	q�eП�t}��"L����2I�g��A�AʑE_�y�j�S=f�x0^-��%���t?˖o�������]⊣f���+E�
�����d$��Xة�_��}	�+Zˬ&wG���~mL�c0
��ơ_�i����p' J����㭆����u�0��L�˱�Ki,��"�i 0D[Y~��Kx��h�n���4��������L��ܸyK^�wW�-�UC� zhzA��b��uL8EG��,5
V_�3e�DUdb�N4���x�ba+�L���q=V�w��%	r�˓O>5� 7�t5a��̬c�x����z�����ZxF�Ґ�Ea3�`A+�04�`�-�dQ����s�+��8�u�T��8�u���C�H9�����ܰ�d��Ԃ��j����[℣����i$����`���Y,G�a���s𕘨��·|�t���� �c��L^_�xݎ�TVWS�qГ�߾+�^�I����9=z��0u|�u��^�y��5��`��2[���MIr�sc�XcT6O����L?��{�ۧC�?��A���}ٿ���s$�Ǘ��g�tN�iCW5����z�{��j~����Y.,���q�H�T�����&�R�&�iN�(j�L<npK-)�9!qU���X^���Z\Y?� ܯ��Z:Y�0�&/@km}�|�������չ&ZF�k����u��R����z�_Eu~�jN<p�i�"�2 M�>��m���\jtąP����ben���}wN����m��I�|�(�)g�2qG�ZJV{�٣ʎ�rU���>'�c���OY�T�9�6nX4tX�Ҹu ��'�����%�-K�@��1�Y�����6`.��fo`�X���@v�544��}��58�H��3�L�<db {��3W�6�tR���J@aI?���x"b�H4�l����^6���m������E�	��r$;\D+r�!���ݒ��\�tFZӶKz9���s�NL2�Y���n�]W��~��8���P�U?{|2������@z�9���&J�n��"�˼k�@X?����;��C	�6��g�	�#g�*��3;\;+������J9>��Ǐ�Ɲ�W���4@�P�-#n��b�5��.�״�=������z�9e�Z��Mt٭�d���I\��H �Kn}�35��W죚��d�� 0���Ca�@d��!����an� �]��\H�6
ٳ2�uX� ��'\�U��PU�A�����@?���+���y�����C��1�	��)�gh��Q��b^1CEHR�e����+*�a���NAyz:�G[���Y勝 +7�����KS�(	"��J��j�¼d�Հ�l���]����i�/�&��{�8��it��A��-=�����/��%F֬�AuAj<G�ޏ���V��H��Q��<P�O>���-=\�*?oh�e��&4ۃ8lh��уu�@��"��#��G���YG3c���:_y�xE%��롯�s� "���V��f�B��k�fE@K!+-=��)S=݁V�%��P�d�zo\�+Y�ƒ�ǲRGwrԓ��pi��9�$`!�1��@���*����n��&Mke�t�.��Xىl����u���ޢɳ��|�JW7Ws4�&���6�X�\~$�O5D ���@Z}���x50HfeK��C~�w������5�hҁ`�
��C�VZ���H�L�!uC���Ӡ9)r��ka=)(��������K�&|��P������T.�����{���~��!��k2E�xi�(�^T�-٢$CK�*WeJ�:p�G%�N~��s0� (D�MS� ri]���t��*X���pqB*WY��y(=�������(���;�|�6�ׯ�Ra:�xE-*�%����_y����{ty��tl�x��U��d L*��߁y�~�U�p����D�Р�Ͼ��臿��xnU�f!�nn��{{������zz��7��]]���5t��*��ѓ��i`�z&9U��b-��ǲ�5�[�5�m���W�L�����MQMF�0��FC��-�ubv؎NN�Os�2Ɯ��L�����&�7�D^<?���,!>f;[�vƮ�������>��s
1�-�
��Nq����5���?��������:�HJ��Q=�n��������[B����_^�N�_G��U�<lg��%��
}uؽ����=��(M�Ø�J�i!���c����7��h���lO4��K�$@���%~��")hC���j2M�)�=��]D�&'�֨�X���ރN�2��XR<��g����
�Lxb��&�_��/|�1��);7�~�ZL
6i�/����=�:Ȃ6sa 6,�H�v�E��ax��!�uo%�e�&�h���܏AQ����6!YI[ �C-Mʻ��$�֏ўh�t~ę�"!�8;>�;���������1���%�mH<��S�͐h�Tv�k�p���K�����:N�N����;�Hf;`��=�� S<V�.�Z]�����&�mKLi=�j��ـ��ܸ�������O��u���e� �ʩ^ω&.�_ɏ~��$��:(���+�;.�y�"���6SNn:�>T�q܂xw\c��L׺X���ڀ�_@&�i�T$n�\��\5�~v�j�e�L���_kA\T[8-<S����0u���
}W��&��t�>��hLn.#w��v�Q�?f�f͜��rb{ܚԖ(�P�!�>Q�~�Pj�O .���W˜�8�X���Wߕ{����fW��ة�5sɎ�m�c�uRP����wش��Y_���I .g/�����g�~o����-��z�{�a�^st�0��Q��M_�`�cp-Q��Z\}��W�0�qoP�!����5'�۟k`�'�A~R�6A_��N���G�2�s)�၃���Y�`� ��ew�f�E�����3'�Wm'_%7���?s��?�BX8V��9XtKNZ�҃�;9�}{(1�>E}(%�3)@�ؼ��o���{��o�{FA�h�!��,��]� v2�̘�{�\�R%����UW��b?��Q��3-L)��+͉ j�!)�k4��Ԥ$Tc��'b�ϛ�(]�=��8'�O��ဲ\&jG�jj �&r�b,�n�.��ߐV�&S��S67i� ��n��픂�~����rX�zRP}6�����i��~9��35���yEZ��vC�F�!�8骑�d[U:ȧn�&-� O�H�FT��@�B�[C�Q[�P��B 2+�I��0�>`2\����S�u�(���>]w�$�����q͆\I*��>t�]e�bq ľXcX�[�%��#���Ή'Fe46�7CPV��bqh*�6k`���G|���:jQC���B�x5��A[^�{K��!۰��;�i������n���P�ם��˟�ɟʟ��K��s��$���)5�~ o<���xv|!�>}%�^�d��N���#:K��[r SȡU������~��}F+x��[rp�m�l�����d>
�Xa�*S�<h˃�o1�|��t���ڔ� �����^��X�[W�-ُ\w)`%����io}G�JR(ru�$��A���j��@!�H�;[����\m�<���&��5Xеغ��T�#)��b�����\9g��Օ-�i7 &G��cR�*��*D����Qi�d`HA�o:��v��k�󦊷uKpL�߹������,>�P�  l���Y݆|�<�/��s�kc3%g|�f[7�s	�.HC��	a��(4	d��*�I����wڜ��+�d�%@d/6���ᢩ�2���(���.؟%+��UW�Y��&��Eo���3�K�Pd��V�ZÈ �y�����a3��& ȋ�}iA�<e�����@�$��0� jht1�:F+�z^3M���%`��$U��H���\O��&k�G��n�5�����C[�}��u\�f{Kvt�jk�jF:պE��k�K�=&፣���?V����ް�:_�[�����27 ͝n�O�(|�������@?����9�ؒ�~�\���p���J�� ������\ 4�u�`����\���^_!w�&������zXlf��������Xx�*���s��������p$}�n]:H��@��7f��QG����zPpQM#$Ȗ�<��&C�ځ��޻�ֻoɻ_}G�����{����иh��e�0Z�㓵-�9¸�?�)(��Zg/?�����+���ju�Z-�`@(\��&��.īǸ�3��6���ߚTǸ���6�2fPkܲU*}��>h�p�PI5�o���ɕ��W?��E�6�\�7[����#X�J�Ln��ksX��vda�4��f���{CVw���..�幸8���l6q�vi�JJ
6_��/�Q�� UK0G,2���o��*����*M%K��,�jm��	:	�9��֒�� ���ٯs���BG�&������U���z.��V��ʎ�l����Vb(�\�	��;{[���9�������ޛ5Yv^�a�Lw�7��ʚ�*L�d�=����
+B?��~r���bK�"���l�a���%�"��y A�@(Ԑ��|�{&����{� �;�dӸD2�2�p�����kmˣ�=��5���h!s��°$�I��d6T0�Y�6:�̞gSd��%t�ri��(=̦�(��g8tȵ��X
'{	����*tf�Q������3S��F�VO���R�<h�k9�.�ϙN >4(�&kVy��Ji�	+%"��ܱ�, ͇�}��qy�V���{H����)�f27�*���^� ������ʳ��1p�ę�mtt=�2�`x�������An���$�>
�]S��I�"��@���~`�j���[�WoHG8���?�}M���1��7�zvl|��ۏdww_��L��&�20���s��z(�����H�N���u��擄�a]�閮�����O/��t�g�j�j0Mu$w��&/�xK6ֺt�~�+�z.�[��	7=�&pe���krG���ڕ��s�A�"��6+z�Gv�:t�.w?���-���m?����0+ ��g�(��+��W�����Y�B���j;acOAחZ!�F���1+�2�
�I����`���J�U����%s4�If�O<�V����2`o��\��
��oM�#q]t���M�6�L�iCIWn�H
�o��2�1��H�7'��g������N��WX4uX|�cj�`)'�z�搬���%�F���VIh_��|��9����Y �+����3���q^���\���_+귁+w�
�d缕�2Υ�i���/A��!�4�}�&_��Di_�$pŅ&��^ݔVw�v�P[z�{Bm�u���"�A�&㚉�G��5�����U�����M�C
q�HY��aFc��VK��n)K�s���1twfR�k�i$;ߌ�p��T�/��Nk���"�%5�OQ�T�S�`_����AǤ?���'��#�K�w�@"� sQZTk��ێ^�&D�±\�ڔ[�_�/��Uy���I��l�Wb�	�sl�buB�"�����w~)G��j��8���]��~��pz%SW���|�@,���zeu�|>�Gl�A,��81q.ͱ�2Ft�������	u�������o�kp��q�It��
�j ��^26E�2�� �P���;��?��>x,YԖ/���������F�(�ۓ?�g����X��a���8��xt�_���W�#�8�84vڂ��kK�F�d'[V�-�}7�{���û�g����^	��)�;����J�o1�*r�{�>� /=D8�Ȝ6���;Lׇ��q
Z���\�����s��l2��¤��{�)dE)qG/F8�aBaT�O����0Mi�� Y)��æ�{ap�۩3p ��jV�c}*C`��i��c)3V���~�bfA]�i�l�{)�,6g*���+QY.l.K�2E��*	.X��9
y^�	+~h�����{��\�d��Tv�t�3 ��Z7�������/��g^�j����?�7����J:�S�����W^�ϼ�yB<\�����1y�������VZ%�Edڱ*	iH߄�]�ٗfPA*��H�5�}�N2nz�<�f%,�A��/���l�a����J��HV�nhU����nXIly� $�;�Qn�2X��
+����>Z�TЌ��ǡCT·���|��ٙ���Í�4���3��}|�x�Z���Kd0���	I�8 g�����\�~���@`\�&�ȣ1[�d�*伣S��C��Q����p '�X�O�e4LE}�ԛ�������������ͷ�͟�'KQ�k	D�:oݟ�$	 @`D	��T����7���:�M����=;��O(^���kp�:�hR�\�N3b�6��u|t����f��y�u����k	���޾�Ȍ�P/ǵ)�i�ze�k'�w���u� gBH�_L�\�;��[��+�R���8�^�<|_�-���_0n����ԆA}��
���H�����n�>E�_+�:)� !v��JV�9�FCq�n�%K�i��y�qL#!;P(�dj���
=��+k����4�k���v���a!%�N�:��v��w�J�Aެ�� -/�jA��I��Σ������X�	�0�d��� L��DN�H��!y��sx�
Z�$\,����	�}t��8�ܫ��(tA��vU��3��\@O'd����
[j�S�S��B����D��1�/ὠpXa���V$"�X#-'��E%��: J�
!�������� פ{eY�B�P�����'�XHM�s��U��_�Ͽ����9�9���Cd�J�,k2>�>C�
d �N�O���r�_괖�GF��^w�Wz��H����<�w0��B[�R+x݋{�u[��0�[��#�꼽w���HgZ���U �jv���T�/�ȴ�l0&�\�(��~tB���q0��o���6�u�;w>C҄��\Ʌ�㇬�L49y��w�_}�[���=��Dk�U���APV�.�bE:&T����}����t3Q��U�*��y2�
�Bt?���u=ת����̨�qM�`�w�
��r�m��&և��1cF	�D$����� Q*]���0��h���LuMl���1A"՞����̼ϓy<\`]��7y|bR�oV?��:��Dq�Ć,m@��� 7r<㹫Б7�4\1�0��j�#�!Y�Z�,��rƉ���I��<�}�nN`�Z���{�%�ݐPh(�"\����0,`�ɬ��0#$�
��m��(�r�:~�S��`8(Pƀc8j���KQw�(vf�!��Gu�*��i���<#�}
Tr`���7�0;�%��,`0�>��Ҋڥ[�xo��2�[������,h��:�k��Z�D�'��lP�C���xt9�� N�N��@"�hԙ�rS��@F���t�5���+]Y�\�Mp&��2��Fh2a�(�{��swY���ŗ?/����\ݒ������Gl=�+_���x]�pK6��d����O�J���t�rf.�Y-t�)$������-�l6T�؎��s���0aJ��_��j+Z�Yr3h�L ��*R�v�Hg�r��W[��G���l���$(S7���x?��qLF|5FU�?�$�VJ�u�Ni�UD��|�p�V��4��&�����*p�&�6��c]�-X���L ��j"TD1DeR��@�����#���"�����nS�fU-/�d��}��W����hVLs99��"��I�����T��ɻ�?�G'MD4��VH-�غ?%��ʪ`f�'�H�_|����Z'}ޮ��mK���������j��G�1��k+�����sH���G=���݊��S���W��W^�.�KT������/�zW�g�Qf|�8��y�'7nnr�Lƅ���c���k&� ��blU�).c�-��4��}�2/Ą^��3]� �@J?l�	]!cZ�9ٔ(��Y(�A�������d2���}_~��ۤ�m�}m�s�Ԯ���[�k�~��V��z|G��~7�E�	F�� Ȧ�!0��$�1�)��$욞��Hs�Qb����VO�D�WǟY�9��f��>���pi6�U$�}!�V̽YG�*��1r�A��#5u��ӱ��P�B�V]7:��F}�+�858��*�j\��Ԓ��0�Y���g��ܪ��Z�P#@3@p`��As��m(�2a�m����S�V�>@]�2MXg	���&O=�\��)�C�l5���  ��IDAT%?�@P�j��f%0C�b#O���3�,ݪ��]'�+�T�0��X����Oq�>�%�d|�@W�E�^ȝ�V@�n>l����ݒN$Wo]�/~�y�k�/�0�� "|v8��Ϙ��ζ&O9����c�����-
��ov��d�و���D�թt4]Y��dZ5�^�2�Q-��7ޠ-?9��\�D��H6�V9��������,�δ֨���*�a�l�@~��m�|
���
(5&^�# ������wv��C�/���50�5Y�?�Oe��>鑷�������&�����:�ҠQ�}g���=���ߖ����LhC��v��	�������F]l��4�q��P0[7!#� @�ï����6L�I0���ۡk��Կ7h����4�o���	Ʃ���.PXAB���jW�v)�q��:�'�
_��~tt!n�ӝ}B�0(���y�tO�0�-�[	DQ�u3�zWm�^�2&�U����B�
c "R�Mv�B������̀�=~C�`7"[)�CWEr,����CPcUS�pYl^:���
7ri�����ma�����MI�c�z�
~��s����]��ბH����9>�7�Z+��%�WE`������%̂�Yv7\�F��kPg;��*� ���'���t���6|��#�#���9��:�Ta�<"k��A��Z�Aq���ӥ��X�p��K�խp�l<͒�� A� �T����}*l�ŊkE��v���e��wC�{q �99;���Y�D���)-��x4�<?�ʹ���7���/�!_o��}�,���$jx���ߐW_�~�����'?����㇏%�9�Ϛ�4�ٞ�W��sX���GH���WKǾ�I��r8���UИ��T��;_$g5u�h�#	��X�"�����6�`�3~!�.�=�C �V����1��Ԁ"(��a�pɨڹ�)���~�cq0�9>�����K"\���4ϫ���\,���M���ݔF�6$�����u\��D���8(p�N2
�
��y�̐��M
�E{pv"�j ���:C���t�,��r19�ӳs�u�9��2�4�n�/5��S�G��!t�I�齟ɵ���y�-wt9�Nupr��B<LpLK�MM|o�խ�=�����?��脶u�ʆ|�w��_��<�����?��?ء�]��jIǙ���խ����M{�xG=ܑ�f'��9MW���{>��,(Zsv�8�������pp�o����s��,�k���Y�åg��ý�����,�f�յ�U{׃N�:�&^CZτ��4��-,�9�A[aiJq3�P [Ȥ�jA�-`�{S�sX=@/PDb����n��J�N<���A�T����q�`��	���3V�7�vV��_�p�N��� ��	�s#x	���b�Dmg��e��Ȱȩ�ތl�7�HBB2��DJ��|�Z԰�y�6ր*� ��Γ���c]��80�Gx(� /ߣ�re]�F�E
DF��R��n<�y��4ɛG��n���>�>N��^/"�dk/֙��.\Ry*���#�.꾈r�Ud���FpѲ�Ӫ�C�Z�E�m�Y�Mt/]�}Md�#�FO�����-�7���myr��<��LZ5yymI�66����J��M
�ԟ�rv�O�4�0P�fN	+�����]Qr~�)��]�-���(f�j2�xӶ�<B��H?��s�u��ec��U����f�b[�	<�Z�$�F��/(x�X�Y?}O��@�LV� �{zO%�L�s?��8Y�د��ZB����Tvv��6ҵ�:jA��q��F�c�4����lmnܴ�XN�*y`pI�d�k��/�~�
`87t��rg�I�����s���5��`�Nl|�Ӗ��%��./u� P�$4���L~���E�Eac�"�CM���}y��_���]±�o��f��[��ns�BK)7nn�W��e�{�%=����	c�-xm�=�-.,o`L5���o�ɿ!)ؚ��÷�Q<I�|�T��#N����U�_5�0 ���yX�.0<�z����yɯxܧE�b]K�G��S�3��aм��Kw��6�7��0��0+�I� ��X�ִx<�1A��B)�*��5lN��̡=��q5�Ȍ6&�j2�I�l"�$����i��
@]j5f���M��&l q-j���j�z��_+�3 ;~��Q��CV�45S���6g�)����''O*A�<d���0$?%�q��iUm&nR�h�H�R���ɀn��:�V�ל4���/ޒq�)�C�z�3r���scM�|�U��^��7w"o�����}[~��)��0D=ޡ�֩P	p�D�g���߆[-8��}BV0�xG�F����hN��
��g���?o0:х����L��)�l���&����I�g\J�]hR��aDv��9tOBc�`����m��@�'~Z�nE��o/Å����~ y��(��Y_�H�^[��嚌G���`,�S�mj�D�:�Z��zk�[F9��Y�N�Y�g��z��}��w�{(��/����j]���)7�l�jx�ɓ���C��1��hX��]M$�Y�'�<JcM
������N-���]y�������&����"+ ��ڵuy��W��A�L���I�y�[��rE�ܹ#_������r�{,?��{�d>�����0�H!i�p�2Y�X�W?��\ٺF*^P���QL+��A2 ���X��U'`A���{�<�YQ��.���/����3\G��6@�Ȉ����NN�e��I_��6uUmSO�JO��f��A�u��CHq�Y��� +]��� ��.�tI�HEQ��Zh�I�A�����,ml�n1�9;<���?���TmE�A1��1����%,b�
��[��t��Q��sQ���h�gnJ?�\�k���Э�����ǧ�$[d��j��j&�R���a����b��#�x�K��Ƅf�chPE���$ ���Y�dN!0�Mv�C�)"�n��� $+����KG`��~��|0�
��*�V��ՠk��FFB1�Š��Ψ����y`��3P5�i0%㬇�GG�H�Z'�	��R��A���ڕX�z=�M�\��2HG���0r8|���r�%�m�z~K��������/�~������#�{��k���J�+�k-�.ץqL/h��s�$r���0"�E[�Ð{�Vs�($�c&�EU|�#z�|zx��?M"�.q�la~f�>$��iC�������-��u�;�D�]p��_iM<u�XgVl���3�\����Ys@6pQU���Τ��2IJMz$A��nt�)HT�5���hs�|>C�s�`Ⱦ�6��ϨǓ��V�n�s��l]f���lȤ�p������Ou/�Eר^P@��HV����e���Zh��R#�D~i��0�v�{�8qi��`�H�p�X3��F�����套^�[�n1֜����>������+{;�Y�7�?�L_z|bR�oP��?��^�2�����q�t�5�zP㼦7 �UB(�8l�88PĶ=Y�[�K�glhg�ڕ����J�g�I����	���ji����A`�Q8j���.���������DL�̪�g[�������P�"���sK|�#Ь5��a�	-�����"դ<E�~�Nc��ˍM)��i6�hY��i R���q�@�A�Xo���)�d6�u4�l2��n�d����L9����4�c�]6��O��p�@��%rƢ���'����I�fCb5��_5ƶcF"�Pj��������=
� ��`9�pglZ�35L�����pЗ�G��F1��|�Y��"��eݜ-�_��-�������'�?9ɥY�� "A�g�t>��+�Y� i� 28G�;C�P-�a-*�Ԇ�їA��u�"���Z�y���)c1�"�U��ήTĈ>%���a�r3#�ShY
 I8ϐ�Lj��sc67����u��
�3����^��TA�"V������{>��u��j{��;��jP��zE��O�@>��dp�G�@��2��OGF��d�&���$��q��3f�[')�q�^��ub�A�Ŵ/ׯi�}�,��cz�s,O���#�Qm2d� 4��3ѫ9��Em��Y�:��ܼ}CVV�Y��_�d������D��S�H�����{�0n���A���[�FsU�FG�7���Xb����}��~.o�y_��Φcu�� �7 ��y�����t9u� }��1%�d�36�ZӁ��C�P�*����g�c1����d!��C݌=ߓ�q���
�1n���zwYV�3Y�����^[?���څ����z!39U�r>E5�61�s�r|��4/.���%1;N!� �iRHS�5�P��M`�O�/�
dYn�$�9��1MJ�����߾_��i`]O�bMG��a�QuoF��`�YҀ���F�JM�4d6аx���X��-���ځ}+@�]g�TxB��lE���\�qe��X�P���F���jȒbm�fF�\&z��3�^��``����c�����8L�E;s��J�Y�eUg�gH!��l=أ��}��^ݏH4pOF3��O���>94�a�B���s�
��Q̒��r,�>����Ui�b�\�-�t�ݟ�fDۅ�/mDq:���T�9�|��atk1�@�&S�(��u���©���%�d�c7�+K��d<�:���l���~F�rn�f����[�S�º��A�	��9�F ��{�r��Eذ��1�<�b��:(��Cc�>'��<}�AQՒIP-B��	;��QJ��jv�ު�Mp6�U�@X!Ӡq���'(���p�|���?�څqɽ�����H����6?�� �&�}��@��NG��NUT����� pd$i��iu@K}G��	_��b4ĩ����N��!A[Z6�IjT��8���fO�ʗyؼ�����'S�-��8h��t�dgg���un�A_Wc����z�뚅.k�ۆ �~J��,�q#�hT��E̦ǌF;�?�a�CN�A���e�����1��>+K?���WBĕY�/�+�l6�����^�>�	���3�㘅Q@�*�B�P�`����qrV�k���xr�����
i`|s����h �AR�E�T�� ΍c���O
de��KY�7j�w��A� i��Q��//���F@A?	±��\�eNK `��N�Y�]��?�@�+���a�|,���\�#�ʰ�&��c��������]��?����P��AL��(�f�����1kGF��X�
5�#�,wT�l��NK��H��
3�9 ���㿘e�?��t��$%����:�@�&��Z�ʇ��M	��d��-�	���>����$�q2G�ERV�daP]��aM4�/�9��T~���\Y��
�	n�,b���܏�F�`T�f��^H��UO�o)��	�Pe��9+��g
o<~sR�l����+��r>x�5*��k_)h|�TTC�en	hC���x�rusM�5��L��N	C�`�I*̺��npz��PV�#Mbr8���X��	M�����_��.�^�%�k�rpp ��w(�6H훕��y&y��ż�Y:�(]���K�~�@f��/�'�V��^�&���_��֚:}߾Q;���Y�ոDv�O���]y��y���\�O9��(�zư�}���k)﾿-�;����1��RԼ�������bXW��tn�1ʫ������x�}`qU?3i�>t��ip`]тZu���%�Z��pq!=���`a�B���ha�����	j�N�����O�s�gFG��ⅼpblRV��8r�h��Z����u:��*��&�,O QA�?����*�k	1�q�(�B�{f\"L��n�X���Dx! 6���v@���q�6e}�ܹ�(L,&���i�X�N���;28J�hJ�뱦5B�0��F\#����W�*�ڠ�&���9�����4Hi�+G���4"���}��AN�t��:	E��%mݧ]\@�xz�W�`� ��c����3׍�.��-0A�ҕa�(b�|��V��0
=��O5}�!��9߳�j��ʪ|m��L�pJ6d�Y��`ux������}�!�r��#�$;��M��i[d���;'V'���(��X������+>�[� �$&����m�f�f	:X�+]�=X���ޖ����	z�$�\�*�d�$���+r��(��;�0�fD\��o]i�N�������66/���3��
��9�S�kz�`5�m�Jrj��G[���&�W��Z�10��X^mj�ޔ����!X'Ɵ�"�d�	:B7�����C1���v�#VO�����@�#t~��^�Q`%�]a�>����Hx�a:�fӞ��ၿ$�yn�"?rc|BGpFz�)��"�(�x���p^t)}��9.�-˿��S���k׮���}|�Ň����tZ��Q����0�"u�; �W�G�sQ`Nݢ�{ft�_����!���s��j�9*v��A M�0��<x��DH��-B܎'���3^��gCIl%{�J�%�WlQ$8�4U���]m�FA0��a4���m��VJ
&�oYԭLʟ��h~�N���/��������>��il�a7҄�f-����yd5u_i-oL���������tm����ш?�Za~Q����{���V���D��ĄV�>.���dDCF���L7�PFÉ%)+`�-e�@�E@�ckrU�(��ȼ�Gᆾ��YjbY�?�Gip+ҋ�v\m���0�5���JQ-��h�7n\��^U����|��2�ʓ�۬,�V7dmsS^�vUV��Gn���[j<���=��d��h##����GV�fe��fSo!�">�<���������"�JN,Q���ED_J��2[K��	��	���;+vR�n}f�P�u� ɝ�-��ԑ��x�a��2�С�Z������/R:�s����霽�6���xIvL���m'v��k1�,�go�U�q�u[H�gʭ���W�YIs�a$�` ��?������Sӳ�k�֣����6��#�b�C��WW�#�,g�Ԙ�`bp��<�ޗ��s9>>���w4�ن�5k�Ђ���|�+g'�z��!:�z����)M������t�	o(��2� &���R�����6�������w�A�d4���~V�"2��,�07k1ϓAv�J���x��*n�Ğ��9� ;�=�X�y�X1W�$<����U-�7V�����cF5�d2��9O39ՠ�� 3M8n4QesS��E�;@�t���œ[��Y\0fq��l7�3��i���Gb�<�@���S�� 
h��չ�NVU{b�|��DI]T�.��Lm�xЗ��z��`��\ꮀ�̴o���AG�经5y<<W���#��pM�7Z9f.83F^ t�V�( (7?:�VəR�w�M�.Yt�_辙h�]���Aa�P������,�.&��H��<��w�i�: �q��+�Q�9F��(��YhSX7�0����N��g��hUGq6x�����$�$G���JoI.;6��>	2<�3�G�#O���x�@�d���gL�v��ʽ��օA�4�SIm�����3�D ~�k�5(#)R�VS�A)���Ì�S�r�A���w�+�Υ�KW�����[������'+Q�ń���%��egI#%�6�|���?��]~g X�2$Q�/���?���>��f���Ch��ޗ�V��b�̸^�(�r
��蠔֑��Y_����[^z�s��[<}�4���i7�ޭ���:��x�z1�r�Ǩ����Q0f�)��Jsi.��!�Wi�^ǵ� <�`O������;�����w
tw�f@9ϗ�Ɓ�b&ela�?��-r�5	}2��u��ñ,����.f����_���<�Ɗ�@�"�������'�ꟽ����V{��
��V�5#�10��MՃ�@�1Ո��puH�G���7�,b(�/�jcr���W�g�9&4���N��5������Y���Z����C ��Z���7��Ο�W~���+/��~����@^�ngE��>'���W�%M��\�W�ޕ���ɷ�����O�Y\����f�m���;�fbܹ;@X�nx��0x����������ڇv=�h�%(�@���;8!4�͵�.���*�1�Tg%t���_�,�Aςm?�{�0���Y`�s��n��{\�(X8�g�>k\L
��������m��w���Ȫa:����r �w|'�sz��g�A2ku7nC<���-���;��ݿ���r�{"c��XzL ��P�.�Ǝs�@c���&�M+�/�������p����6���?�@���w�y� ��������zcI�~S����������F��u����AR���S2w�k� -m�P�"�[9W��ѷ\�r>�\�ޭc��,n�!�պ/�(x8�+��j�Ʀ��_�`r��uUR<;P�E뿦�1H�BoƩ�h��:h9-餲$*��M�D4����">�ҙX�n�����k�$�Q7�Hf�,(dd��@'�+���;�p08FɚL�K10;��!�6s�MT��g�I��

���ß�T�������A����k��t��g���!H @Wʮ�y�*Ѩ��x9}d���-P��d
�L_��]�R�3M���O�?�!�!dciMJM<��l�����4�o�M��*'��Pr
�1\t�ʔ�h,��#�Z�;���ɒ8[s��׳���)&�M�J�e�ʡ&k����wC����9��ܖ�z���B���Ξ�{r1���]y���<y*Om��α����L�Sַ6���M���,�k��T���I�����^'dֆw�
W����*�\�����N�v�	��E`�}ǎ�7\B|]W�`��>� �ߺuS���74H���?tE���TI֟ �1
!��C�6����枫}�H��H��,0QM�U��4���S�af�08a/{���)zm�nºB�Y�|���h�y�ާb=;Y]��׿�e����d����F��Nu�c���QtLɪ�6M�y�9�
V@�E!��u��Y5�wE)l�(��e`�Р f�f��d��Q������#�9�Y�E������=�纪�(�{�V�-Ԓz$P���ɛ��W������C���'�>���H�����Og?��O3�v1QOF��A�-��Dpj�eiA�R�f��h��F���=G��Pz���x�g.|�;tC��;N��	B.�e����rU��j���pa�������z�9��|]�{垜�˓�%�������we|p"Y{]�>�rx&��~SV^�+�~��)kr���rr< ��x{W/y,����1Z�@�Q�*���TꃅSn�����<=G������.݋�U_}�_���;'7,,0���.t#��\V`�T������W50���R ���� P��˰��u��UY<�}!)�Ą�w^�UCgv���Ow����T���P:�I8��ت>��ͳ���m��뗺�ji4�apF�h���c�ȭ��}yp�}VeF���<��k�	��"pA�7L4#gnQ��d��t g�}����C�pPnUP`N�s�;����8e<.����
����(�\4Y���㇓N5ul!�.�c�oj����Igl��)!�2זY�?�����BG(pC���5���r���c�d̓F�'�=�Z������'�a5LΑ�=׵s�f	�T�5H �p��*����䮫�C�l9;hT	��FUrt>e�2�'��[N��9*,�D8Rۚ��2&g64o�M�T��d�2\�x��Tp�(��.
�n:�-	�<�ߑ���o�����M\�!f'�x� w��D�@�ա2}��}o6�^�B��X�4P��MMX\W���/�c,@�Mgn���D�����BN4x�5;��c��6a	P.(�ꭋ�� @/�G�����=��}*Ћ�,�IS���i�>�� L`��hQ ��i���_?��>��h�ƀ�P]?cp~!C=?PÃڱ������c�Ԗ�՞��.������?�����_rVeoWm���4��j�Dj;��'���ߓB�yP�+GU�.��}�S�?;��=
�a�x��ujq�Q�Kc�8;�w�~G~������^�3R�v�~q ���͍�pvp2T�1X�̫[W�_���z=������.����
��37������F�H=|�X����C��&#Qf0G�sQc�^gɆ�مi���P��{�h�A+��o�)3�ND�$� [C���LB(��ޑ/|���ګ/��n�`�2Y��z����p^(j��BȣSE�`�rهU>)2�.�����( ̗ �[�$ uW�E��gn� �����y�`<֚6�|X�0I~S��R4sl�� ��*�^�"v��V�#]9uILC�y�74j@��<���H��C~��iR�;�h�:�(jMǣ� n�l�Si 0���LB���G�>VQk���){G�V�)wvX�)̩&�E��dAb�R`进p�ø���P&~2��Ѿ���5�y���&�6���L�y�M��_~Gv����?| ��SY�`�<Hq�$�O.��`_^��o��������	��m,K1R�61P�v ڙ�?TB҉)N&�����!�Ȃ���c��+�����L�d~�M	�p-�Ҩ���yA�����#t���M8C-���I!iY%��	�!ЃmB�]A�~��#5��uh��ZAhfp Mt:>�Ah�4TP!���Шx��R�"��&.���W��p�y�sp8ˍڃ�4L&�?����S3X %q���`|#c�izQ����!���H 1�kF���!�	�T&������,�d��?�۳WKK+La��#�"��P��3 D�{:�
�p�˧�F�UUj�l�Ӳ*�MV��0��h�!$��� �y�v�9�B�ݩߧ��n���d�t��_�&��҄�<�������	��@R��*�X[���y��lW{��X�p�
������ػ4�|;��oYҦA�8˩~�h�=�!��Ն��Sz�W4`]G�����;ʄ��V#�wA'`w�?\�qd�2��������@Kʤ�:�ޒ�ͬ:���{|>�'�wd�։Ԗ�ة���uT?s���Ԃ���ױVi���,t��@9��u���:���Y��X��F(��yG���䡛�V\����]�����L��S]7����U����UiT�'�>�ȥ���J0��++6���C���r��m��v���xh0S}��ɀ�]K��^�)��&����\F�EciS��ޒ�Gʅ�����<����ܤ�ؓ&	�3+H%ƾ�$����f�;N��kR�>TfAI܉�znz������5|�xOF�;�%��?�e);m�ḯ~�*�]����<�կ��j��cI�/��
�� vX�; ���=$�u�� �g t�P��ʪ&[7�dem��:��h2�e�I�������w��h�U�^Wdsm���JtA �E��C�6��Y'5#9���}��x8�w�KS��]UӋL�I����Ċv��H=z$�nO��� �
<?-�of3`����/�'��m��뾃�7�։�DuO�iY�
��n�ssz��fB=�^����T�q�1A"]�������Z� ��9;&/�{H*�����ޚ�W�q
�%O��)2{&��g3 Q\r�v���G�i��L#~
�������_���~�a�Y��%N��E�47*`\wtlP�bic�`g�Os�d�w�B~k>`�V>}��=¢��G0
�Z>�OI)Wk4,+���:�FI��(��I�qQ�U �H�앜����5Up�z'otg:�r��pI�Zc0�
��Vui����?|�����(��@�I�F9&orA���h[���o�D�������;�8���p��,Gm�XOGgL,Pm)�]�9<�ýc:ܘ�i��C��֊Cq��F��!�=��:�38y>ʲ2:�%��Hy�x�K��� ��g���*���^�\�^�U��c,-�
����j�ap�y	�,	�~�P���Yz��N�R2��[���|:�I�g�h1hG��p�Gqm�y.�Z�M�D�tX���8bĖ.b�ɩH5� �T�3G)��$g�t`�"��i����3�� �B���sz�Q���ᾀ�XQ0G�1�(6��G@m��`<e��]���p8#�,W�d&G�G���.��vF@[
�-�|Pb��{�N��a���_�pÍ9/vQu���Q̃۪�w��W��̫R�](������ԥ�x�0d�:�� �^u=�+��k���ۮL�i�P0.�ҟ�d6�#ꉂ�:n	�d��k����_�{�P�v���J��r�ė��U:s:��0p�tH&��yN����X��s��nݾI���1t�c�e��m����@��e)��w:3a�=
�si^$h�Lk�,9���S��z^��2:;e2�C����^�!�Ԗ��1a���z��w��g������(�]��פ��Jx�X����c�A�?dGb�`2ѧ&���@S9���	f���?�¦>epv!g{{r��j�����ݽ.7^}E@���P<�j�X۔[���O.��'=�)g0\�H������L��D���TB� ����ÁU�ql�ģl v�*V7�D�̶�or�˟�p9���^��j�x������r��T�{	�ʠ�]#��&mM2(7�j�>���Y���V����bN�&Yo����4
��u�����&D��@1��H�M �,X�t(��R�����,��܉HL�?	#/i�?'u���CiVQ��p�<�}5�?#mfª[[�I]��|���rUuR=B�Y�5�=hTt�^�'6�yG܁�����`-MR�VSMF �	}�BƟ��7��&�>u��s$��h�K0I)��x�21aY#�(�C$��,��q~0�`�]��'4�p>�zw*�� ���@�)}���z;�l�-�Z�����6�W�/��y���ǧI����Ԉ2N�8�j^�o28���6�RV&4���'�q�{��$8�8)/�	b<\����.)@�U@o�ɐ� �t�Ea�rd�,��6!�ÓC9A�0�a͈��&��L����=����}g#�KcRJG7��7M
b���'���{���P���8��t�-AK��
�z��ӡ@EP���sa/	}�m��9�N�@��� �s�j=��q.\/�k�3ӎ�/a�Q��݋"�Q��/��e�*rj��ߌK���1�����P�K�o�X��Y�'����~7�/ٹ���S��@ܵ��6yF*5���p la��e+���^#�NH�[o&���o-��!\S35u0�Z2���Ĭ�v�a�nh� ��E�xǨk�HI��!0 S����[�X� ��J�x2d��Uέ�RM�&�2g��=+gz�}����𜿖5ݿ�9��e��X��PA&˃_[�1�ʹ��!EL4����g��p�ؑ�i����?�>�y�F_Aלqx�3�I��W��Kg�h�L�W]6Wץ��1#$�F���N�39��y�� C�v�S�G%�{[���6���a�Ht�В�@p���zO0@���6��`|�	�� X<G�׷�5�z�e�����Dmߐl(��%�,/K�貓�!p��wrM�ԋ �Ix�s�%��féP:��0E�wG����h"ؑ��^&���\@U"KzK�Վ����{uX-�16E�c�6X��������/�C;���,ip3��%5)J'Q��q�� -�v_1{�Z4���`?�\i�͗��l�2@G�>dpz.]�PL���ҽ�*�&�%��Gغ��vj��{�4\ѵ>&,��-�Mv����be�m��-��H�j�s�n���ӤjRXg��ja�y5֛�M���k��$�&��uY��6$n5�&p�<�P�w��Q��I�g�H�#nY�V�<o^��{�_�_��Jo�:��DN5Q"k�2�Nt�^�:�F�z�޲H�uG��VW<�r�v��{	�%���|�7�+����l[R�ע�8O
�v�-�q��������?cG��M������|iD�HL�8s����H���w�D�^$M��q}���k?��l.'㡌}	 �q6E!'�ǮmQ�.�7a���U��̟8OM+L�В��W���^�2�b�sK��}�v.�(.S�{���9�'���a�]�A<9��������b�;�Z�5A|\T6|���1��䓱��O����Ǘ�����������p��2Z�0RɬNQ�$�9)����F����\�6����|��`K��0�I�X^ܰ��.0�j\�j.�y�J�pbN�ft��&�t�aO.pT:pt`�QCt��\�R��z@�k�Tn��FY���GC�DF�>h`6��2T�3�N�L���/V�{�۸������f&2�=�Taw���4xÛ;#�-Q�dxam��p�E`��̫6j�s�a5� �����:��0�@o��b!@[�<���>�Y�5�ď%���]����zG��ղB�)^� �g�;-Ǫ$����+�t}I�)]c�ʉ������MV�2�����.n<Љߺ�%k=Y^Z�5�ёl?ݓ��ت��me��cy��Y��޾�����][[!cGMR����P~��/50� �����F3V��PA���t{` �{ﶾ�sr��-�u�C,�����C��=frb/ M �BvL��*M�'�ɀ%�ZJ�r��/��E���=�<�{��.�O�Y���kv�UT݄��C�k����(�{''�:���H�0s�a|�%,(૮�l9�ˆ�+�3@�{=2҃ )e�=$���PhU'(
)�P^Q.T<Gc�{�����[���g�9��0M<��@�*ڤYF�c�Dfg�a��f�0��d1���EyT�ޭ۠4��a��FuʿCBt��r'.�Ķ��3�B�P��V���lP�&��։��ySmz[��f��iA�	爎X�"=֞�=��@7�� n 9�X?3A ��Wm��������dN5w�_��,��0 T��ޓU��<�6;����-U���1�ϑ����[�ȬDyc�j����I�'j�&��/p?�>�
*��t���9H���?�Q�|�&Vq��cʸFZK]2_͊S��#v��d���:E$Y���7(;g���d���K��Ĕ�0�������`�Y�&��}��VL<��8q���~�AS���X����,7nܐ>x���1�$þ5�k�gJ����
)t[`�z.*dP�����|��X���q�zO0_�SD,e"D����o8�0O=ma˜*�vH"��0��8��h�
7��'=C�!s?��;���̻���]��g\ge+K���H�yYHL�#��^�����μ�m�̳̿��iR�;���������������i���)k�C��8v,�F���Yͫ���X/d��5%�*�8�kj8�CS2����S��!� ��x��rL�W��P�N��`_�0'�EH��IQ
d�I��|lB�c���47�J�R���s7 ���. �����Sf��}A�ظ�]��jH� ���g�J`�ꊧ�Xo�:h���$�K�	q0���gr%�b|��"IQW��1x�2vt���O��K�o�}1�[����� �k�9rk���s\��w^p}��sr&j�0���PVxxV�0���`3��(n�yuU��}E^���r��5�����ߤ�������ܺ�%���������Ǉ�Mg#Vvǳ1�n�|A~�_��wn���cy��#���WduuUN�����r��+�w�D�{��~v��D��5%��#R��X�P���?���yS�� ?��8�p���n*�8�f��}�!h`�#�n7e�ԮgdB��<�&TD�<T)�B䝴�G�^F~�M�$��&��A��n�^�;{6��s���vۅ��b�ăp�0N�y��#�&Vy�ܴ℘h
�"��x�~vG���=P=�"!pU� ��-�^�a6�3���2C�cf����;������60u���Y>8Y�D �]��#7ס����r���5��BpY̼�4���p��d���!ef��èo�=汐�����bj������dS�#M��+7��p��9�]
wqn�t���1%�\7*�8,��S���S�7{��qc@FC���5v%tM�|5�]�2�dJm5�s� ��5z�*+��
X��	�����9�dߑ��}�`__�.P��L
T� ���n�� g�2�ݖD��z '@ؿ��`LT���jH�jN2+z����s��ڜe��,kR���t ��gM�32��e�I^Z��T���`8\����R�!t���{ǖBi�9�Y&$Թ�bW�
��e"t����h6=��no�#��¿Q� �*�n-�S��2jZ��$�0_�����T�9I(f�`8,8&#Nr �e�����1�@r��H6�c��^u���[S;�&�����\Nn�=�=W�,*!+�4��� ?�p�.�lq��0�c6'WΌV=��/�
uFZ�m��s�/��*�E��w[�?+s�j��Q@{Q8�_U�6��K�tSF��"�u���%�⻾������jާI����?���������?���U|��'�����R�Gq#�#�;e��Og���M:gb��ǩ[�0�����&��l0��0���b�uc�2���sV��f�K�Fp|c 3NX��D��.Aa���:S+�g#�&jLR���T8�"�#G�R�cC�(}��*��P�����Z���$M�sb�ZA�F���"���UI�(k�zV8�TX�N�Ts�����4�$e�ie.�d�'��Hⅎ��&zf8�rU�r���N�w\�t1��S.��{f%~�Ú�C"P]2��#�s�p!a�

�^l]�mI�-̄54���ʨVԛ5�ch�>%/4*�)H	��eu�)7o���ᶼ�����G��j��;����@�ܓ��M�2�S�4���bz!��@Ndo���&�����.�y����Aj�$����Z�FMd(�NS���/rM|�{���z${�R� ��}�ϱ:I�@Dmb"Ky�0�5+R8&	�n���ׯô���ﳯ^>{-�0��3���yv� �
[�ދ�)����V��A����aB�5D����ݓ��(@�/�e<�Xm@Cϱ��ˊ^��FG����U)�:����t ���\�k-��}h�Y��&v�:h=�nNH8p���weI�{u�K��!�^���Q��X��=�sZXU��i��bn� �}��A�ڨ�Y'�I�1$�z� ��nAH�~V�#���p3]w�%u�{{r��O;q���d�ʺL�/��Ǽ���B�}]���+v:,����t��)�����1��lP ���q��T9+����h�����MѨ"vmS��0�^o��
��(��\�Á���PU�5�w�H#aI���=���Gm�ݕZ�����T�?��`(1�,�=�X0Z��)�k�d�B�=}߳�����'���IG�u�r��5��������7d,u�LC��j�v|"O>���y��T�'��{�~jЯ�4f�j��V�F�b�4%�ݠ��Y�����ڍ�r��M9?y���X��6g� +a���?-	�1X�A�P=��Ϲ���l�8����-�9����a��Z�>н�lEj�����pHe�Fa�h�]e��hN�L;;�rz�v�n��6���zĚ�f!H�&N�+eA�a��-��*"	\`��~?�=��}'�ߣ��Y���zVv���^���,M�=��%T�u��� �;�%���=��#
`Fq���%�e��X����B���)�8%�>��������?����������׶���^-�w뜮� Y�������M����IBY:J-�kg9/qܷ�
�)���x�99�[Eý��������!F�g�&�砋@@גF`8��O�]����`DJJ

���.���ϙhڲ<�D��hL 4��, X�C�6u`Yzi��O
LC ��	�5(�فka�X� X���Ds,�)SV�_m'N����ط0sV�]�m����$O��wn��a!���=�&�g��"��ߟ���G:X�"n��.���ϲU���N�Y�n)A�k�!Y�	?��Ȣ�{dm}���
P�`E�k��H^�˯��r������=�s�y&%�otv�o^�_�)���O�o�\f�P��:��u]�Tq�ܹM��T��D!fur2��8��0���H���]ٸ���kPť�fS��0��i`Ƚnr��'?����4@����h�ǑX!��e��0�+�#,cq��쎥����V���Z8�GG/+�[�[���o{ߣ<l.���,B�H��|q���Ѽ�D&O��G�2Рnc}�Ǉ��!=��k���$�>����j�)�ڡ8
'ʪg,3]c�/&c9�@�X�S�CCT�-�`��q]�4ڲ�j�
Zp�*fGg��{�X>N%y�'���4�4����Ō���hO�5j����$����c�h�K��`���UU����$i�����PMxRT�1��?9ؗ����=D`":���/MM"��IU�{0��`{Oq����F�zG�ܺ��i�j�;j3MD���� ��p7����2�c�@��>r���q�?M�0����-t��k��&��fBx	����eiw�4P�Y�9�ݗ��L���h�;u	W�%����u�5�4�Ndr�I��%H@Hƺmi.-��S���J�Nկ�Rs������@��>�b ��g������$H�ʃ��&)� �vν�?'���M�J*_c =vB�H
Ώ�d��w��?��<:?��z!��^_];Iݩ���Ldsc��Z�m4c�-�a2���h��躽�%_��ވ���0oK��P���H����o�r�R��(�9g�\`\�jf��X�L�*�B��� ��i�+�'fX�	�*:1��(�����ҸW-��9`&���������٭��k�{t
��)����nn���A��w
��".616?������b������N�ŷ<�T�s"���nI���É�\IK�ϋd�/�����Jq�7^(5��B��T�~��$\'Ɗm���ץ��^ ?9x'���Ӥ�w�������_������Qo���7Io��
<�`l(7U�Z|`�Z����Jzh�)�n�����6�U���ȉ�C�=38[Y�>SR@�j��C�Я�O�q�3{TP)R~9+���a0<}r1��g��.�&i�6����U%��`!�u�Ԟ�a>GP,��"w,��Х���]�"�Z�Aa*�h����#)� (<���0#�Ư�u�Acnb������U�1�
��� Ӽ;�{!�g���A�!��='k�,e��p��x1�����E�3�&$a��IsŎz�����Cw��E�:����0��ў��q)k�]yᅗ����#7�o\Y�����ǧ�m��P\�mZ@!܀����������}� �W֍�>H^��� t�uٺ�����c8р$�j 5Ġ0�]cY�{��4nȵ�W���L���x�I��N}Vpũ����Ċ�=aP ��R��*��:8�U�����3��v�@{�+���U���|��C��A�TU87�΅;�b�gB��ޫ���>e��X����Y1��%��J��	SN�:+ .!(mю^��H�&����6 i	������r�+�F������4�D���\�Tw5�\¬�^?�i��g���.��nߑ��7�"�@d�R�/0�
�@�Xz�lid���#�uƽ�c��g��uY�Ρ+�l�ku�Ȏ	��y�#=}���-���:k�k2�&T�EWp�Dϩ���j=� +W�h��`!ઇj�dD�D�Z��A\td��KLf�5Mr4qʺ��䲪k}�8i���;��$n�백ғ��.	'0$
{�d#2_���KҀ8�K�mH��6�Z��.u	���Uh^'z~5}Β�����$?`��?���;а�ؿ�� ��_�߅>�X����z]��Ů��s�kp���-р}�`l�nG�~%=��z1k][ݥ��V��D��&1�o�+[�܋w��iSd�U�^�+�o]�V���#&"�3F�HA�+jLH%�҄��ݛ�3�'M9>^S{>�c�30��x���bq`���1���8��Ge`�;��
�D�A �����
V�
<�ű���Y��Z��n1���QNA�m3.� ��:����.&�����u^��Z��(��m@O� ���0S�AlWT@2-nVVU{��fEyU����pӀ�?_�;Nti� �a�Ů�����d^4C�A�Q�[� p� �Y`�?�-��r!�eN[}f�U�$��|�w}R����ы.Q�|�|��?���oVV7�����?�ⴿ/��6:\:�Bm�_�3�@QuX�B#3��'#�(1��j�Ƞ��t8�T�$��L����V	ɡ�Th�}.���IT��8�f����A7f+�3�f�'[�K�c�C�L�<l�I>�����e؀��Sbȳ|R�"�J�p(��1h�l���J-�;���R�VGB	��9�0���'�����O.Rˀ{n��5xu�PiT|�P���T5�i�Z�R��U�	�Y��ر���=F5[��\hz	l���R�0�L�r3�4p��@�0G�`$��,��KBp��$s�� <.�fP-�4c�*߆X�0�H���� �M�4y����9%Z7NU��5sC�H~�9�{�NO�4x	��d�?74Y]Z��`E�o=���mtk�y�����@��|�+_��ٱ|��>g>���a��|W�z�uuCn�ޔk[]�������s�?�,)�۫q���QS���>��)�8j`��k<;�K�9�M6�p%l����US��J�32�瀢%����-���4U��K�E��e����o����W�d�u&��I�7嫻�T{4� 9 ���h��!��]�zԻ�����>C!G1�#� C�0��Tu��]zw�����3��.� }��}o��s��{�e��}�Mt�8V`�g\a�e
����C0�| �ZI,���K���B QJ�1ʛU��.����+��E
1/}ֺ�6��k"˘$`��ѧ��@��X������c�_���h�4�P�y�P�2D��
��*u9��:�K�����?��o��l�H��廯��k�"���o\���5�=(�20�:���u\]���ߤ��w��0Id4��2$*Ը���Q2���G'��7ߖ�������lj R�Mft�eu0�ߏ,������O%��������B,�����dJ����H�@�%G�b�~���Y�>'v�:�������{�6G���3d��˩�u�=ac0�+���� ��8t�r�@WI�	�!t�k�\�ϼ���-�����b�x��z���~�Ӏ;�`��w48����~0"=��jC���lH���x�zgL/�{ؕ�IG�Ӯ�g��)�o\�^�w�O���3��ؖk7n�+��풞v�sp.��O�)L�h,�VIjC4+�t��ﵲ	�a>���l�E��G�.!<���J�0��m�H��6��vn:1Y��o�鼣����9��ds�Y�,>Q ���;=�Ss�08�V�*�.+�����TW6]
�h%��t�����S��65!��h�po�_G
�7M-X�u1	�/ ��#vt���*���Il��a:X�%O�X;�)E�'�����h�Av��A���U"�O�]S��>��(�J�vx�$Dq�)s=�gj��� ����������m�uP�;p|�[ߚ�����_^�qe7�[�юK}���f8D�������9}�2�!'�E��Ol�	��=Ѝ}�ﳄ�H���7��8c�p�]t���H��bep�"�����M_�
��4�N�9��Qː�S:��:^p:�����:�t돘g89���q��G�3U����,ן�.7n>/��Ak`�*������=�����"K�&�;��&���p$��9�h��J@����
B��E�&�˭n0f�"�56�R��/�z�4>�������ɃsP��g2�����3?�c1 ��b�A�|�.4��?�j�B�#�rsfN-�r��R�BL��j�P��Q�eh���?��s=+:�`��З���X�r�ꖼ��m���l�&l���}WNN�dy�}���t{��{z+��cҔ^�r]�;���E��RS�����/��R�ҌԤ��2�-��;l����G�D(tkM䢍��/f0�����mŝ���{��*�g�#���<�w0���M�ܴO��"��TlN�qb2��2��%i�X�Ul�ԉ�LC���rE`L	r'����H����9����D0��Fh��N�ZQ��RK4��:��7�U�'��T��~Wvչk����5��O���s/���[��r��-��(l����+n������ ~>Y���r�3~P��QCcqd6��,٪��ڨ��֚���ր�#<��k���Z�օ����alI�^*Z�t��g��)so�~�{1���f�tf(������|J��R��{�GVh��dӱ�q%%�0�~R�&���M���YI��/T�:g,�J�R��u	�.3Xb��
�4�[�l���ݿ��=�A"!�Ƭ�A]���fKO&�%�a?�a�`� �ӓ�������{�r�>��=���tu?�������)`�S�Q�騝�?<� �'�bȽ�p�#Pm�p�^k63)��3;J��m�(p��������s���&v}n��d��wcL3_avp����;`�YeC�L�;`:-�"A?�*�m�MӁ�2�Q�/��a]�#Y[���Q&<[�(w"��ALM�.�����i����:��!n�na|�*Y"���=6�C�gp`+��K��������*���S=���a�3?�Z?H��W�w��D#��2�|� 
�/��M��@ݥR�"�g_�#���K�ۗ6���eߦ���Y�`��Jc�2��#���$̠�[2w�(k�0�pr�잝u��i.�>�R��)��a��/n��A�/.�l�4��^�Y5RA� ؕH?7e��uS/J[-5iD`� O�ћ�Dާ[\�F�~
�Ԅ.1g�S���$��i�e���|]�޸I
���m������޽;��������:{�Q��0�����(��(!�@�Ah�[x���6��e�ED.:��6]d
J�3x�aTi|<��m���;z^����~�b�֢��E#����B�s��97�̺3fN&z9�tkΫ�{`%c8a�� 0��+F0U�Rl^�v��~�Ɗ����<z�X>��s����]�ږK�ۺ��:��J�����~[�֛R�W�Xjh�pE7�'�dw���W����<��MB�?~�������ǁ�;'�	��{"O�>�kW����\�(�N	Ш�\�X�M�9@-<+�L$΍]�,���"<L�^�.<��9��=�tFu���߀3-���ss�+&#��=�`HE�@&��<@����^,�+���,U���lFM�.����&��:r8�j��߆����u==*K���*-)�E��~����!�����}yzt"��,_�Yj��|�X�y��(8�I�,>C��C��BYx�����a(5�<�BŜ�؂@I�6�q��R؅��5�a "�c!����)�;�f�q�s�+V���Q "+�*�, \����������4t6b��e'ޟN=�Kh�J�΍y��@Zy�⎞j�l0������4OfI'�L)���҉��$�W4�'��cm����ڥ*��)hWV�X[���5����ƿQ+�aߡ�����4�]ĕ�Hf�h�e�
�9U�>���=��;?��W�_� �AW��ָ!T�Q���'	h �_"�/tkb�:O����?�XpD�@�b#]H�&�Sh?}��=fSsoF�Em�q(�s�TӮ􈪺��%Q�e��7����ä��g.��_6���e�/���x�7C�[�C��pw�  �3<��^��:5)�m-�U�2˒;�dfpR�&~9#��y�e����x��.)j�� ���c�)�F;��wq�ʪU^���l�PI]@��p��9V"�py�K����[G�� ��	l��I�SL��w>* C��n�=�RP�����C�V.MVW[ÓՖ��m�#�
��*f�8B9�̝Ó�3��]��P�!���{B<%^=B�!��BP��{����4���ӊ���M��(;ݺ�2Im?F���������ּ�A��,�T��U����f�����t����1#���.b=�Z�9�$(ꚭ�lnoʆ����-K�Q475-Jk�*�A�`F���Ȉ�`�+6mEE�b�E',�8v�E���Zc�	�I��;��̲�~lߴ�#�索���}�yt�a�?��柙?������H.6�~5����Η/�]�7��tZ�i�rco��I5�0I�+@�e8��Z�z�M����H�H��F�|�e�cn��)j���.�ƺ�A_n-I��$�rvڗ'�#霞�!����pp�N$�O��T�Ï�T����w5`�G&�v�'}�#|y��+�>/���H�Z+,�zm�KW�U��L>0�;�v̙�B��+�/<�s�tAo`�5tc{.�s���/b�� �
����
]���=��ͳl� ��c���SP�� P'n�h�c��4@�R��:� ����r�8y8�`Va� ��J����h��>T�k��Q;q����9~�&S�/�(4��*3r'���<�5��)"���p0멁�D�q}���A��H )�M-V�Wk�|ޅ>��9h�Cftb	q�� +W���&��Q��39}�@��=�@�@֖�R��JAw	8�ڬD��vO���~5s�sÌ��%��"��#�>�J��Yod�Gj�z:oG�Aېh�t�l����؆r9�ّ'}$��?j"�ZP@�R�'��+�f<0����S����*d�	Qs�>�*h]S{fC���u]t�+�s�M���oɛoG��*I��؃4�cpú�8����-�S>��!�DC��'r��H�QG�{_�v�JK���Ԛ-Yn4�71�J�H
Ĺ��E?' [M�zs�A��5�$������wP�;#�]�kP�g~�-.�A�-���M'+���R�4Ofױ�\d}T���/���Q[���W��4�xM�����ꎩ�xO�^e�2!.�)���� ���b����~!���nE�?,�cLO����Hr1?~Z���m�ގ��i�%�A�ߓc��w�bO�c�6L���A��Vc,4�W>���Ws���X���_9�A�v).0��|����3?��lFዊ_=�
~G�0���f-[]k��IIm�)%Շht�������o�l_>w*��gM6\L��� ����tldA���M�l��3�U�0s��S	{Q`ɰb.3�8��y�5kh�*��E]I{�ԕj��4G�Djѩ������(����Ȭ:�{*�$�͜ݳ��Y�:\kA>��d�ƨ\��T#����̓��13��nb���=�����Y?2��ƥ�nb6�RC�,�@#�R�T��B6L��>���s�L)���n�e[�s%��}?H����D��ם��>���'�����Z�_�ȭDm�Wk$��l4�`9�2!�6AŃ\�0�c_���}uL&:�M��c�s./����!?<<�?���RՅ�\�yE�V/��x ��:�cΛz�Ad4�c�c�;��^wD�M^g����%���ռo���������Ӧ�q�Qu�@#'nu;
�p :H�C��Y(0�'2�g���Il��7S�:��W�8qz&���U��܂��)�
%p�I����](�6թ<��ϵ���TgaC�HS�*P!�.ҡkM�=�;���C���<dYJ�E�U�I����"�%uP�����9Ȗ����q0���ىt�y���:�'��\Ǧ΅L����{��O��L$h�������W�39�<Bg��`q�qӧ�Tp�	D�)ej0PV@��T�ȱ:��р�P,�ُP	Q'��?�#���D�W��F������_�����pO�%Y��iI}e}��r�p�����4Ԡ@�^
R�@�:%-V��,*/�ln�uV[�<2}6�r��ʱگ���}N:F��M�Ο�@��֔��6�z{�������/4K�^�H��AO���d�ޢA����wd4K؆)a�, y��ަ{�vVEP�B��p4B��S1���d%��Zܗ��ib��o �H4 <�����/K�[lz���o�aO;m�<~�P>~�C9:8��~�ʵmY�u����Z�*�h*u�j�ˍ-��)j�Z�r��N�rrt���T��M@a���%U��B�����Ω��兌��b�-g� ڈA�e�cW�F@�w�z}ڧ��=�]�P��������[Ѐ�A��q�4�@�?�t{{[nݺ%�S�wj��@(cR་R��@��K{0%�Z.�ˌ�y�d!FӚA����ޡ7������>*��3M�*�U9Yc��o�j�K����S�F�D!�8Uv�E$Vs��Y��`e;�;����	���̅<��Lr��:w6�~Xj�����ߟ�����̿f���#��!�_@��H��Tu1�5^�z̡,��}v���M>��4h]�ށ,��,b�"��g���"�4�����J�)C652��i�D<�3�G\�&ڙ�2P��ɞ�q8�12@�-�rT������`��̱���eP�l�{-�|�1�1�Q�螞��������Lzm5�}�wNe�>�q�m2������&F!7[��l2�t�`5hᢢ���Jn�3E>K얹
��W|�� �Qp�ڏ�����
ѳ2�^y�ߕe�α���A�������9�'��J�ݼ���wKg��,���MB0�r�Җ�m4���Kܜ�z�m�Bn��|���dgy��$�J��+��B��ݻ����N��m<����!�'c��#�Z�4��s��;.��ɁԪ1�E�f]��������M6�!{������d:d�2���?�1��~�-�~�z���:���w����;*��,����xg����Zxǹ�_�	�,S�p��*����W����"�ϤE���B�|��*��d]��ϵ��)nGTN.=u�������ઇL�tBAJU6j*�R[X	sҽ���aV璘��ߕ}]����Y��!�@ǩ�l9��?~�P����QN?�\��3��k�(D��k�ہj0{��T��D��4t��$���#�6,׵���l��5H�6��n�Q'���*�j ��tJe��c0c����k��H��S	ώ�b�b)2�,P��K���֡ldx��^$k��e����~RN�ϣj�j����`XǇ�sׅg2����P����R@��
�2:.u4���Lw�D*�j��E�jm�q����1�Q�%������Xelmb��'�g24g�>TάOb��G��IK��V�����ȣ'�ٷV[N������|"��۟��w�K�jԮ���n[���3�-�^z�jaU�����C��WH��?PGv���\�Q�|�e2�11�l auM�
"t���?ّ���mP�s��#ׯ������/΃s/Z�>!����r:���\���<W�;��L���Ч�=����`��µ���������?g2���ٳX���:�5O�2�M����!��2(�///�|�=7��Z!�8$ ��}�d��ے��[s�g��}8��f��Ӓ(���{�ja���k���@Z�JҀ\FF��=��df��|�`���H��*�Uo�К�h�*F�11eA6c�k'��Af�<�vX�cB���������r�7�h�7_�#�.�R��)�=b+�a_.��@`���s��������i'��2�b0Q�Ԁ�DSi�Eˁe{.d�B���)<b�
cJL3L����VU7�D���;�� b���(Xfx�P=�"ʛ,Ň2ɌA�"���̀�H�śrה�;����MT:����]k��讴u5h���jP0P�\��Zk[���t��H�>]3�`/
�����`�́������.�N��2�z̚�}&�ѥz/p�^�ȟ��ۿN�b�'i18��FU�U4�E8��y~]Uaf؂l�G�U5\Ss`�1|l��s��WZu�$=.��{����5>�G�kp����U��	���w,|�ܾ}[6��J�R��w���w���D�B]�A%�GE?W�� �_��S)Wj��|v��T��@�U��������쮎^E�uݘuuM� �F,l�:���=d`]����@u U��:9:>��Χ�7f�4 �Y �il�w�l{vs_ܴX�g���A��4c9	���D�gce���+κo��3
d�)�(ī��6�O�����ɑ�ײ����$+:�}VttBc���uӱ��*���Sw���A��%u��u���fT�ٟЙJ�lJW~4%����~���0�j�:��;u6siT���d�:��RTG��N�F9�udDu}@@�8�{�� �e��!����hՕ,2�pb�+�S�]�X�R�N,E+}0�G�(�CW�-A�ٕ�ei�6T���s��*�zK�HדH6��4�VA@D2!u^��С>y�1��X�~]lh�@��^י^s�ϵelu*ϐ�l�+i�/�+ө3}t�K)t��9��Ϩ�sѹYpn�W1����A9�X��P� �'��Y�(��VEב�-��0��0Z3�#�}�%��U��*���#�G����(aˤ��5�?}�#g�n��GS,2��k�-�|<`b+;i��<m"T��l<1a)�E�l�dcsY��[������W���Xܽ/�A����f�#Ӗ�~�<�ۏ��k�uk`e%��~N$
g�)�\d+��P�H�"4GO��_>x(���W������o/T���]�N�*z�`����1�������N�����dH�*��߾�"�fE��tN��'(K���'�,bY��#����֜���ԋ:~`r"��5N�j�d��yh���� ��yz�j����	L03CO蟳�LP¾���u��ϐ*�L���ed�&�{B�$����@�Î2��e�u��(P��s˜��������ߑc0�V����ߗ��=�b+�%�\���L6������&P�����H�W�Il'aS.y2�s[;-+�j�G�&-uN������[�Fd�!7�^
���Xz��Q�.W��!o��+U�ow��_~�yWں���{O�Pa�v��"ު�p�o��\�s�`�S�^f��y2����3��8 \h�;cF��Z��n�e�䀹R����9�yX��e��,&���ӛv!�aĀ 6l�L�^�c�mp<�	�F���^t䳅,й�
w��K0�/�x�gU	.��j�:�1`��F��`)s���m���g�)@��\�����7�/�ݪ��8�OԏA�`]�?ܑ�k��=:=�ý}�������(3p�;�Ie����XY�&v/�{Grvڣjx��	S:>>d QQ�m0L����rC��4�|+�>��/>��+k0Y![R�Xv��&��q�=�T�K�@%r	��N�Ii�Ss"�}x1`[d}ʲ�oAA�d�L�c�8�{
��͌i�BI��<��:�E(Џ�t����^\ �^ׁ���C&��:�m��^���TS|U�AK�V5E�l:�p��\��<��!��FĎ�<�lh��m @�����^^��Z]
����S 26�������꺀�$�o �<w�5Qϔ�
dj,)d*
�L]�T-�l��0�M�p�5�@�2F�:���F�W.��	���!�tFN�)���πφ�_�4�E:U�U����<���Y}�=�kT.pydMs��Ux.�9f7��W<tp�t��h|z&���Ȋ��z	i�˄M��L0�����,p�����TX1�VU]+�"����`��G� �`���[o�]�T������y�ϥ7�fxv���孨��jp�91%��{�Q�c[�5�H��-aa�5��	Npf�'z�rA P�"X��R���^���G���"D3u}3{�����i}���ƞ)�΍hs@卽�9�<�)�Ƅρ��?����_ܕ�����ή�c	6LG��L�`�g�ً�������~!0���Yh�7�j��	H�/0�qL������$��@��,����AA6�=Y�%�����4��E�S����2�C�r��r�����49l���G�l�E2�N#�dԣ��9rA���$��L�
5�پ��F�A_��&i���bn��S���H'���X%�1Dzw���}S�3�����o�1�������C'K��O�c���G���> rcc�8�%������d��f��\p m���%��D���h�J8!�v��IL�m�~f*�",r0HdRF�F�Y,�L�߇n�̔�����W������u�|�ey�{ߖ�T��������ɣ�:���Y�0�d������u��]��w�)���UL��9;���I�q�����p����NPg����X��ω�N焌pL�ܜ�=�_
��ԉ;�g�)W+З�qJj`����֬�4�1Aa�<��,��ϡ8l[�����9��`b�����d����XfY�g�S.��b�h���!'s\����9g�ێT��>�n��eo����y#K��2kT�k���ޓ�<�����JN�R�65`�rN x�T
�p*�Gm���A�s�Tj�3�3�5���s�D2�X����NuOuP�㾉KR�A�B��j5&��P����U4h�C8��Ӊ�x��I�R�\3"	������+BXL�[CnBa�����g��_�X�A�k�3���"/2KY�M�`6��y�]C��8�!@LФt�yU JUY�5e�t&-uB���AV�U��YW�#]W��wu��"�j�TRg �M@�����t�j�N�H�3P��L#��)��ڈ+f'%$tP���љ,j�} ��H���u&�����4*���UB5����YǧF�@'Y_�TE��L�q�� Ղ{t������::9d�`W���6���Z�|iYB4����	��X�gR�����J�\7�G8�>)'cRA kfl&��[RR�re�,G]��ź������ȑ��!��K�3�����l���[�8�$M*��������B>�4�r	LK.3��Woa�4
*��*�$&�1�MҩUBk���@��@��~y�Z�V�.��	��x��s�
��Rr�r\a�����vdʨ$�<���3�Rm�)�U��|�5갓�8�M�2��X
�e���B#9�mqN�T�β�ƚ6,��*�����;T�ԩ�>�����<��O���-���We��-��@��]��e�� �!��\M� d	�9�s�]�W���)<��G �,�纏���=�݃
)��a9�Z]����('�vߏ�/#��$az��ace���ع��Ef{��t|^�8��,vC��xǟzB�Z�9���X����_�Q���*t= B?&�20���jj�#��b��>(�$TI�$� Q����}h�YOB���[�k����ߍ�x��n}��g�O��c2ɥ�*�7�J_���Xl<^�(/bȽP��{��̭��p�"l�S-�i�H�-C�Z#3���^(/�Є�f<F��֔�����/m	8㷮n�ֵ+r��\�iV���TVVr��m��ۑG��Bg�쌗�̝�����W0�i&�Uk>R������[�����iV+��a �h�O�Pm6������ްGCGY��f���Ɇs�
!�K�c�)��;�;#��<�C�p�$%�{�W���/�}^.((�W��:f=*���h��Y�ה�?�=�ț{�%b.6`��T�AfxA�}����D�J�4��1O���g�M?3#��ѐ0f*I6&��ԁp�}Mvjȡ�"�M�Vc�*Mbi��6����,iP�lg�sՄfcY���c��Ct��zԶ�� <sI<�%��%�kj�
��SH��8�Ũ��yL/T
+>�t(��=��3���o����cp��:��C���ެ֤��=N&|O�\�z��5�Gr��wW�l f�'�"6uܗum5��M��D�pj�;�18T'��  @߿^�-�$Cax�����cr����Z]����������L���^g�R�����k�hHY���h%!VV^]F�	����J�q��_�U �t�6�z�����:@AS�_��Tƚ��I��ʪ��������"{KV�K��.���Q� ^��Xf����!@Ɗ�� ��Wsu��I'OJQ�MC\�Yu<z�����e3TR�ե��cP�d�SGR�y�Ւ��-�:�p6��3l!�%#�ڔ�4e����y��i:�z��~������5 ��g�:T���Q��3Z�\#Nz`�'03�6�`�����L��PVS�Ϩ�=\u0� ��{$+YIm~�2�coWJe���]ձ(�� u�>d��bw�}K89��q�>����I�o.g��Y/��i[>��<|�@���S�{�Z&=��q0v�,Ā3e�I�L�Bc�j�U���S�g4��X�g"{�D3�3*�⼘k�Uޙ �)	��Y�X�\�2<.��R��"_ܽ/��ݗ���Ϡ'z+��ZҠ�V� ��&)PJO�P*����k���d���Ȁ5��F��zfɏd� �2��� �MO�	Z�����H���L���$��=��w �K�h�Gq`p�8��"&���5�
�lF9]g{�y���Q6��:��)�F_�����>�~������7�$�*A�ђr�)�h��9��BstS�9'4-5A�|�џü�0�g�����mbT�p��!x�����ϐg�����o�,�0�C4�!#TS��%Wn�(���w啗_��_z��p�(��u��G��we�'�z�C����9�dRA}�3�0�{E.3����4'�B��u	��ɘn�m�-����^����yЍ'�P:���.ůJ5� Kz�1�c�LD�<l+����~�4w����B3(0C���td��y@fc.�`t��EX�ܳd�ZC(��ޤ�ř�+�B�2�󰡋p�Y��BP�G3j��Ex��u�}g����,YΣς�S$U�v`l|��.AXfp5B�j�����@�bb�$cP�y[�W����F�<����p�!Z�r�Afs��I�UÞ2+[)�ظ6��!�5@�M�?<R�P�-u
�"5�qINO:hf,'�z�@%*�������M��	-K�l0��`Dh�5]����^�|!(xV��l��d6w-(0���=�6��$~�X`�"0�W�B'8�[���������+j�	2�%Iu�=��s<S����̂$�V��Z����ɚ:+u��X���T���ӡ�������N�DL���p"��rK�͋R��dv�6w��'O�$���nݔ���������! >R'7T�{(W+�yp@�B�T�+���Oah���S��R>ؓ��G���;��Y�ކ:����7�k`��s� 0����B���X.]�$/}���˯J������>?4,0���F�e2%E�j�8[�(�֒��M�����T9�j�1�����ϙ�/�b��o �`n�~�2����՗n�����(I��1)��t�1�S�ܚ�͙���r>������!'-������������� ]�=4�t�Ŧ �:K%��a��+��%�YS�Ӂ����&��>��� k��e��玬,H+�����h��2`�F��4�s�	�*�;	v�72;֞��6(G�y�ʪ�Ɗ;ֿ�f����P^����w������4,D,�c_�Q][&}��s�x�ڞ-���(��Y�q2c雲�5�W�cOS�F��ht��0	��up�/;G���ä�Ϳ��LP������9U��^zI677u�hKP�e���&u��b�dI0}cd��0r��e�2RS�?'�%���%�ÒD�,ܾ�5f����܌2��h�e�Kp�q'���3�LS&eruD��4�ܧЇ栲�����t�h����m�+�o�5��A�o�������_�o��O�~ 
DD�h\�ɰ?&1?ޡd?�E&�y��T��-��L�5�\	��'b��<��3�M��7iD3@��ʪN�n����nׯɕ_��kWuc~Yn�x����6D}9x���G��g�"������=uj+�>��jX�0
zn`&��PCV��E쪿gҫ9�D�,�ko�S�x��K��4��de�,�F���;��A�QMI)v�n(G�gp-nĉ�3���F�����bǦ�˿��n1�Jbeq���6��\v~�x�����j��[l�7�[3����! #ȅ�_&�q{�8�f���p8�p5�f3��ׯK�`N42ˀ�ʓǻ�
����ە�۲��D�8���FS�w����A
�����:`+B����H��H�����h6cPs�"����:5%����s��.��ꐽz�y���t.www像>%4	�Q��w��m�y�^{���G��_��cD�z���\�o|��z�I����_ȗ_��F�粺��׺��v������>��L�Y]��=iv^��;"s��"#T4��X�.��i��q��iso.hq�mt9Ut3n�If*�̦��\ϱ:p��:�e�ߑSuRz:nh{��"���Z��*h2,��ԁ� lB�J�Î��8MG� ���U�S��0Ό��F�	O��\Ȟ�u��/�D�Ú�ݔk���e�ۯ��>�����AQ���U�(�g�MC�|��	�V�)���3��7�]Y����O��G�I�T�:�j�`C����/���<���n���������5}�$��d��d+��PUO�bZ�R�1EvQ���^3��J��K�r[��+Nw[M�QT�����jP�F|�k�O�ޥ�Wd��7DZf{1�}V!!?� �$.���R�L��ς~'�^�s��e��uy��'q�!i'�PV�c�vՎ�Q5�\7g��/���)�lkE�����[�O%Рe���p  ��m�?���'r�O�h|W��Tڀq"��CnYަ�kc�.(��J��B7_������ƺ���H��K�^��K�RoT�/��轥i>�@ �����Oh����Cy��P�Q��u�oN4����|qnㆪ	`�H&`�
�
��앂���u��N��Ĺ���J��硉F*l�G%��n3089=�~O�[V�I�$�&��t��:��8���'dB���!��*��ҵ�cu��U}���h��&�s��F��Q��sĜ�:jP$��<�u?H��*�*�	�(s}ڮ���\�B�*	Y�)��y�~��k�UH���oi\A#�iN���1+T�~�	���^�v?5�m$29]"�WX	��Ld�ib(�`Q��Y��A�o���~T�?��_�������E�;X]YYcsb�Xg��FL@�sv��鳄�a�|`�ϋ�Ɯ끣Ģ�r��o�3c�Zҿ�T�4=DZ����A�%2Re$	Q�H�k,W4(���r�7��N7����D�>�X�����O�λ��;w>�6�S������E0qX����8���H|g-�!�R5p؄M�:؞[��@���lLh�C�YQ7��n�qT��@�I�ME(5�*U6��Ł�q�6	�`�";�3��	���M�)�0(�F���C!�ȓ�w��HV��5xW��2�������3�����.[��+ �0���{V�7M-B�f�+�*�K/�� 0�3!C�8������?����E����Q"��_�ÇO�����me풼���r��%9>=Q������юt�G�h��7^��o]a�o=��Tʱ��]�u���*�ĘN�+�� ���[̀=x�tq^�&�fU�z��lm�3��l�o�fS����'��U~���*)��l���.���[����{R)r�������3�8==���[o�F��Γ].ɛ��&7��&�/o����G�e�0����	��ּ�܏��E]]���Zr��M���uM�7��1��L�U%��7�j W-1[�s��تC���2�Dyu���U&�쏳Ut-.#P�������Rh�N9�E!N��=�� ��ڨ{�}9W�n�}�Ա]�@3�x�F
Xf�b$Z��P
5u�VW��������4�G��c&��`�'Ý�l"�&�k��_4!`�I�4*��T9^�rMVW6��8!�R��SYɞ5�<{�;;��`*�����"[۬2�8���gCpyJx'���G5#R{ѯ�`�^8�FqYi�Rl.K�޲�(�9���~��}{VH�k ����g�6`ć���;øꚞ�b]��&���n�`��i)�;>L
�کTY?�@m���L �uhP>
\j ����:sSKT��p;��+�L
��z]��~E6��nR{n��y�[�3ٺzM>|�r��P��PZ��\���ZZ�-e1���.뺭���#j+,��-( d$e���ΝW�>d�T:'���)s���:�SN�f�0��䴧�0���ۖ���YYYa�������8�q�=������b�a��+��kN+`D{8S-��AC�d`�K��m�\���}s�M���Dm�4�)������/P� �w	M�3�G������9]��T��ç���!�<B��SV������ac�ׂ�)�<�<G��&��yu�}o��To
������m��(�t8�%�`8����'Vea�ei��	ef@�	Ӫ�	قCY�����G�911��<0x���3��,��24����k����:(�->���o�?��_�O{��j%sx��$��z�ȻL"����3��Ձ��v8HH>���L�$D|��#��5�ԠQ�F���6�L�56��`‑=2�w��Y����s7��+/�Ig���tR���#y��'��{�û�X:G��da%V��v(}��%cn �������s���7
�q����-Ge�1�b�R?���^{-�#��	V��FP�m��׌7�=g�oC���y�aâ�����(I��!c�>�p!psB����,���A3���-�Σ��O���=>�uW~��jQ�`v�&7�hXs�)��:��y�2�H_|�9�jceK��6����]:����:���S(rp�+��ջ�h��q���(t�D����/��ٱ���HO�����n/7������兗����Tg�"��)�2������՗o˝Oޗ>��:!5���O����l���/y�������W�����es��~ ���ސ����7�#����o~󛲽�)��t��캳�8T6�%�$��I��Y߆s�������������⅔fAAv^a�ڳx��si1(d�0� ͜��񪵲:$U��!�xG7d(<Cȫ� �2��(�g�t=l�潦7���H�����_͑���r<�I[�j�M���Z�ձ �U5d�FKu�'�|m&��t$X��9�h ,V5�)KRBV2$�
� �J��	�䇽=�Z�4ig�N��	X�kF����Tx�!]��!M�ՠj�,�D��;���OX�b@EQe����������P��`|��C��7D^�ՠ�af|�E��22�������)և���,���9E�g�f�Ī�mu4���xp�x�YD�kX���y'%
z�>�,���YO���X������cRK�'-�X��ɬWՁ�zC��.%�H��HÞ�'1!�[��h�'��`��ܗ>�7�P��`T���\�vWvw��\)ʫ��*K��?��]��N+�c'�+���ڞ�ݐz�*��}9;����6�p��\(�ɬh�8��C���l7�� :8�\�߱��$����"@	��#T0����:�v�^��I)!�hk$䄕�~7����"U��t���{$)M��EҊE��	���}/�W���Yߏ�$��L;��ϦT{�tT�KS�+��C/F2�%�,��}"ɓ��a��~��P ,f��y�xF�g�Q���:*z��D5����6�u������a�gBF,	�&���3�{��<��s��?)��վ�$O9=�j��2�0�dI�ӊ�oj`��)��W� ?I�g�z
l}�;��#C'b6�sMy_Ç~7��������_�<=|�z�&J�L1KQh$V�(B盵�~�Ν��m�>SĮxE>�9^�\�`��L��2�1K�h D�K!6�ߑ^4]��1�XL0�W�E5B(g"��#9x�HV�����lH��v��M��h�ԁ��b���Ξ��.Φ�kJ�yX l�㉐)1�p�5#ΌifF�ԋB-��o"P�a��f��9Į�wGc��(�$z��;2Q'���Q��H�YGƃ�����K���G����i� ;)�*ݧo�eY3��/2���_��̥ԃ�J�v-�ü��N�w!Fs�*�����.f�{��9L%��5����y��j��R�u���/�����~Dÿ��&W._�����+�cF���x�n�+{�;򳟽�sĠ(� �Smj@qE�I,��?���q)�uy��o���%���Y~��"7�ݔ�η/�P���n��f�%/���N�|��<}�T��uC��o�"���'��gw>%u!�S����:�/I��֥�\�B��X~��ݻ_�
����X�����ç~���'7uM &Ef�|�q����ѹ1�A������;��=+����/ϳ��-0�@�"��Ԫ��ŨN�_`�V���FxFO�QڒH/�ps,�M�dK���ƚ��+6G�~A|�'����N�i�6)0���PLAe���^�!��Z���:?F�s�F��:�{g&��d�ky��������oL!���)� !�N�S�, �	|r�6�ǆq�y��F�e�-�4�jc@���@p8�e��P�tϤ�<!�c}�)CA��T[� �\u �{EdT3�<�����'��*��C�F����Y!�A�KL�ڜN�$R	:�@ncs�4���u�J}iY�X�Л��J��6"�u���!4Zg�r%�\�=AZ05)4if��43G�
�����%ttM�#��#�d #�S��R�F��Q����"y���d��`�x��ϱ�V��f��O;��D�|�����?�o�-f���NX�;APR�HM����%]Ӻ�鸎�2[�
�nT}�Bf�G �o%ݻNA�)F�j/`�q�	�5m����;�ב��W��$5z�|@�9�a�x��9��ȒĒ qhUP9��!q��N�$ Q����X�)R)���^0�s��Cf�/�,YO�8� h��y�5U2�.�:&��W�7fP�����G���O�<��*�/&:����p�ܻ�O�'M��%LV��y�anfv��G0��#�3+��mo�ύ��Ye��s��|@��D!���%O�w?�/�>`��7�7�t���}r �:o�QY��R��y���~�����n��X�9��x͈��˗�ۻ���5�}�.w>������[�����#; L� r�A�� ;�����]!>�5g3� ��4s���h����3���<�xll	x/8��预�o�5CFI[{8��/������V>���l=wC��^��R��>��~]�^�!;O��Ӄ=���])|xG�t�f����.�Cv���WԨ�d8 ��"����5�.8E���3���W��v�\�DQG����A��.K�I�P��rzv��E7����C*����EВ�ܬd��4���cNz5a��#ʲlJ�rNi	���_���U ������m��A~&�ɂӿ8]LH,�n1 ��h�X��*<�5̊�OG`�(P�8�kd98��D�џ����������/�؆W��ِ��Q�R-��t��[׿�"��n���蘛���^�+W�Pٸ����Q�7�彏~)�J,��r��SdZ��	�����>+���T�ӓ�5�� ������������!�D�VC�e�q����l��8*�<HOJl<v�� <�Ț��m���DĞ��m�L7��4�F7:c��T���`�ߘ������ss�\��lyN��)�k>9!��20��T�3þ:�}�a]	�Q0΀ޱ���j�$�� �hs�S�������:���H��G��R4[���#u��sM}�9۪/I�XSw*��d�́ŧS��hss[����˺�ӑN��D�UH�	Qѷ`H^2���G��:�L�� _�Ժ��:	�z �����όf�֐��~���������
�M��l�p<qN9��$����8���)vCh���=4!���� lY��A� f&�Y���֖,--�ρ�7��T��Bu�L}��l<��`�P�OM�H,�9�+hF`&B*f���qn��`J�	�?!0L�j� Y(���[݃Syx����.�Q���P�Ӊ��F<���I�lD:P��C]ӽAOz�6�u�|*�"E��:�����H�;Gz]9<���J�q�g~� �LH���Ωζ)5N�H�aN1�7Zf�1����D`;B6�7c�F�x8���J��O�5��Ɗ�g�ʋ�skP�F���p~�^p^�+�^�����\Y�VsE&y���3(���h��J�@��V��F���q>f�����h<q�ѩAz��Z��ҋ5�F�T�P�	�(6�6�'��#�O!���� ��#+��� �P.[�p��{W���ޏ�Y4�b	0�#B�&\[-�����V�!���U���@�Б����C�w����Mx�R�'��5�X��^3�%��Ϭ������Y]ݖ��i�Vt�Dc�f�pZO���/�1t=�̪	_W
~G�0�.�CW��􂬛	 ّ�`��Ѱ��$�$�)�6 6��n�0gà.�T�pޠ#�<�o޽m�(�Y�����Ȧ��J�����_���P��ŭ���C��ӟ�'w>�+�m�p6�d�Ҷln]�ۯ�"��]]ߖU��Wvw�������B�c)&� ����%�Q�02��kZr�P���=�^17�4�������G�"���R�H�a����D:���yw�Aܑ��T+Kj �Ѝ�-��99�S(�@�1�����0w�5O9
�nL��	R��Fұ �57������3�n�$��?�FfV��Z��$ҹ��9�3]���g�+E~��q��s/R���7:�{�����L�.�c���g�F��,Ӡ�^Xr�������duyI.m���6ݑ��_�o~�;R
�+Q������*�v��R}�Bv�~����nȥ�kr��P�:=y�[r_���ǻ�75�Ц@s�h ��%'0�FYsR���'�h�����FQ���֕e�;�o,�{|B�P���Q��F9� �+XqU7�b�L��e�(|E߭c:��K	U�C{:��y(�hh<�����e��ƙ�Db�@f��{H����,p,�����7]�*�O��D�Z����K݇���}"O{���15�A�:��<^U}K7�u�)�z�%d�t���,��?��^豎��X�
��B�41�t��ڋ�~���m�֋uY�u�� ˮW\V�8��4S��t�K+�_|@��a4�~>�:�}�ፍ.����x;�s�� ��l;�u֢�ĉ��S���Y�#�؏X�X%�ն��B�Y��XA]i4d�ڔ����])�Z�4N�k8��	���ZqI�G����b�N��Bk�B,76�hذ)ؿ�PfG'c�Ϋ��8�2����1�
ji|�Xb���;���M�:��Q����y���?;Yn8kA�KB�4.!���:{�B�kV�V����X���E�������Si�UE�)x�%�JǮ�A,��?C�8e�7`���[���:��c]+}ON4��ʨ���u2����|:�~O�yv(j	�:h��J:f���G�.�i�w|���Ʉ�8�c<3����w�d�i<�z(�&�8�שPnJ M��2�H�>��Iԯ�=il06���,:�\���^�AأI�9a�yܬ���5uX�$�g�B�ԁ�&�(���z�h��՗Y�뽣Q��){bLPw%���X�>�;��Nfڙq �9���4����1&��y@N7��I���Tű�4�Ab��$��S}������;qI�1������ �i�5���g����[��}*�R���'�Aq��yYz�B��:0�ҖA�C1�����c��p��ă�D~��uP�[zA��D����;��yl� s��.��N�j*�9�/��>0E=
��^���CYĉg���A��B��%��)y�N�,'�����HP�D68�z�\��ח����}*�}�m)7���\�$��M�nT���)�>�x*����;�女5�*� �t�v���3�:Y���\�-3Q6:^f�����ln4��r|z �;��6#cP�4���Mmww_���}��ߗ̩�Yr�.�᳗ sVf�wTK���T�捜���\���܋U���{�s��h쟋?�����
���,~���^&|���ǩ�	�w����Z�:�� ��ܬ?��r���p�/�j`vږR9�k�7���������Odw�H?~(�^�,o}�5��������P��QC�vK���r��>�Y��QA�����'.��Y�����eƴ�M
g��� *$r�ƶ��֛�����XchTEU��2�cuh��MRڣ��x����a��s�ltw���4/�8A��c��p� ��,䖸�]V
�ķ}^<<ReqܟUqc��*�82<�{�� �PwT��ޣ�x 5uЫA1Uwת:�k��WJi�7S�A�0}���p4$m�� ��SG�g=�>��d�
jV+eY�ʂ:����),�ë�@U�^��ꁼ�PAnYǠ����%��"a��ҙMF�	�O���40�В�X�( �ҩ:DH
��A>::���)�`�i�A�\tM�pspMu ;���>(���!�$����L�B6	��5.l�RA;7J��ԒD�J�5�q5��j�U�K�SP�0��t~��~�}G�S�>�|g#��ʻ�u�:�9�(S���u���D�����Ѐ�s}8M���Q��K�� ���a�)G�IE�JXE�m̊]�ݡ�Xk4�<�̲z��k�k]�E�K�Xь�����FG���~z������8�ӽ�9���_�qH2����\�%�suP5�K�G?����VmU���������D���C&*������d�AR�5HP�9��0RY�S���q<.���,PMN�]�U��������,2��)���,b����b��D�V�0g�Z�z�,�����m]ֿ5hJ����Z%D�	���y�����dcm�A`=n��E$+�J��ʝi$L~g��9�+�|F�଴;�OD��<D�:	�3����S�ɼ�d�iFtngCo+Gf��� $t�;�P.��@��ibp��5��,ˍ�/��KפVi0q���%�J;����y�{�	&���E#|��:(�-=ƣis:���-N�E126uE�ŋ,���$��Z�CcKjJ�`"���W�+�c�2�g��R�Y�l.#nt�2{a��:�̼�6�rEV��ȴr��r��-���O<%�/������ |qj���c]�d�/f3��x�V�u'�,d����Y�M�&^�љ�;��h>�/��Ss�o,��ظ���ćP"C�����xC�� ���8
R;T2��.B�B����Ͼ2~�p�E�x���p���Ï_��� ���0�s}	2*�p�de*� 0���J�`o��,P�)�0w+�ՠl��;��dR����QQV��+�Ʒ_%��ӧ��;�Ik5�?����o�!��Ǥ����;r�{$+�kr�ŗ��ݻ��[Y������������P}3��?<�{�RBI��A}w�f��������y��O�ߛj�X�"�m�8_	����#�����̤��]"C�nn �X#;� ��g�Q��	�s�ȹ1���Ul�g~.wyq�|e.8�v�y���Q�����Df����i*h�Sǚ��R�?/J�Z�KKm}dd2� �UF��D�˽���ۛ:q�e��2)����J��j�sSë#k���ד��Х#:�ԏ�c�I#�9�dd���ɏ��+ ��Q�=�,8�Z.(0ƚ	q�4	�����P�����הC@��v�ލ��(<�K-i��r��[%6����~�!�yF:o�tH]��U{l�g�C'B�0�����^T�(P����F�bA��k��t��-������_���)�LT��Q;� *�"��x倔�O����i8����s8Vh<���[O��P{|>�������e��������i�0� k����5��YG>�������զ���.��K���������ݟ�#�O4	���*�F��j��G29iK֬KO_T{ڇG�ퟛ�"z^��9�λw��Γ����Ȏu^���E���3PD@	gPǮ��i6���t�Gf3���_��<�?h�\ꡗ���֦�u�T�����&@����l����(�	���?�nE�\�*-���TC&t$S�,; �{���_���wh/�n���>>i�m�XMџ�oN&S#����y�ZTR�B��,<�n�Ν|	�#�����é�g�Ee\��E["�
��|1�2�� �q�"�q��?M���J*%�r,7�]�ۯ</�����ʫ�K��sk8`E�U�$�rQ~�(�#�͹i�X�������A�o�f['N٨��$�^�A�
�
0��gg��2�����	)��CČ������G 66�-�y׻%����
,��8J�̸9����$k{�k��z�D�S̕�7�������l�5ei�)%(�J�%�ƌ��.p��MPRLSL帧��Z�t�Q腅��+"��sYN���2�0xs��3�P�20�����i��Yu;	��~�ep*��np�v��*J�H�`e&TC|-��q�l�CmQ�����i��_�v`��grr�obѰ,����Ξ{׹�v����>K��=��4����8&�g?6x�����e���I��/�lo_Vǩ/�gglG�XmTt>�T���| +p�Mzx��x���LzC(���ۯ�7 ��ZuE�/�Rk����ۗdK�0{�nF��uS�'|��򲬬,�Y��|���\^y�yy���7�������!X4l�&� ��g'����@��`D<ǐ�,����×����>�
y�Jd��T\έB����ǎ�������] �������G`�Aq�	�k�7x����W8��!��D�*�F�^m�V�)˥�TA	��΁yG����d�� V�h�)D������R;�Z�Ȋ:�-u֊hl%�Д5#|�9	1.P��U'w�P�ug��ן�4�����ޛ5IvW�~��##����ZQ�$ � (R����i�zZ��R��<�˼�����	��ƺmZ[M��
� A ��+k��}��=�.���wo�L!Y[�X�ZA&2+3�{�ſ��Ǐ��z  %�`,�E�1ԅ��HC�����u��#���'�� ��U���9
���	lw�촽��5dnN��(1�}h�vx �;[��@�@:��I/ӦT ��uT�Og�#�LF= �� d7�Xh��ut-6u�����H��
l��ߎ>����zG� � �CI˩��7&�c!K 	�LH��O�{uP�=����B����_�u�bB����}Y[^�=� \���X_�/PfaQ��ˡ:1Uo��T�JEώz����D�|�9����\�n�dY��:i�}
K�d Fr��d��c�!M6���;�Y�P�����$�������5o"�{���<�_}�Kv�udq��~7�쓢�L��n-;3J�Y0"�m�֌g����dБ�{�v̓��/ʛo]�^}]�%��\�v~�s����������C�f"�j�=�1C-�l1���7:nE5����Y0k1o��s%�gv'���*��	�S�5	8�aI@c��!ό3�E����t��u��a��cnI�N�1 �<C�e��.АR�{�����������9���3�[6q��l.'R=��e'�[E��Q/�ڙe���%=ÖeA��P�s�	�5�u*�Ӛ?�Q?�.��D���ъ]�����g����#����_���,d� ��4��H�p�t��|*?X�܄4F�|��9�I��4Zo�A�d!�����e ȿ��y�	��E�9�Dp���3Z�G���� ��l�B>��x��o�o��,_:'��D��6e��M*!�X^���2��J�����n��x�H2H��`b*=�uP���3�&"q2�JO���q�iGCf	����H�_	��]=������0ST1g�Q�&Pc�Z�9���Z���R��f-A��'����Mi&cլ�=��{�g�B�b��`����Y��g�]l����E���3��fQ�b��<�C�lF�QoZr�ӯ��͹�\z�[�?y�T��>S0�S4�,)������b��aY�G�v�6���
��ͭ�^t������zH��MN?$��^���˽��1Cvhqi�8�p5Ϭ���������%y�ko0ʿ���kYACc^�5qpx,�/��;�x�hR���XX\���-=�1[�V��[P�cV��:=M+��*lv���"i��%�7����+g99'�C>J�Je�(�w�w�˨I���d1���9�i]I6�l^�;���P{������ pU���9�Ou����F���d7��x[@t*+���i�K��]�{U��s�\�@IH�vK����.g�*z��u�E0!�I�1P���G���ש��H�y_�}�L��Ǳ�X��Ǝ�WӪ"�-�a�&.Zɚ+2�21j{�Sp{��O@RN"m�qf� �w�g�뀺$A��HtMޖa�*]���x�͎N����4�(]} ޟ�����3���M�����&��BoK�V�Zբ�<`�J.��� �{j����כ�v/��a��?e��xj���gun�:�LX��E��%mR6C�S�� Ͱݥ��k/^��;�r�=0�U}=l3��U��e��(�*z�@�n�_j���������9f�ׯ���y%s�����Y�|)CV��h�t��.},��Qo{Sֽ���*/��r�)ù@��^w ������	k4@�k��V�������EI����W���>�q��%P�qV��o���ږߒ��kjˤ�S5��	���q�ժ3�!�S�~7A@�u�3�8�	ڞ�^�mq�}l��"��`��#zd��eg2g�y�.tŎ��#�,d��Nm`��s�Ԕrͤ�M�#Z�e���B� c <�3���ꌙCb`(tu|&����}��譴q�9@ɳ ���璟��A�!*�@��%uv�TLꫣ�׵�Z$�7B�D
CdT^\����N벚Iv�NRIS���?;�7��������˗u�TM��� tz�� l�"p�ɔ�!�t1��xb�Cw��`�P�+�͗w��M�TFғ�E� !�E�7}O�_�*��$�X����W_{C��[�%���x�����}��=��FA���d��_�9����x�>����������,j�$o
G�=����{-�����fE��+]��%��G}6G�������:�T��Ϣ:��=�����>w�"*�L�E����4L�7�#JE����U���/��E��}OF�s���cqz,��/>NֿL__츋�i8�%Y=�"׮�ױOx0�9{V.^='����n��ѡ~dE�^o���V����/���rO��NFo�W^}���	B�����uy�x��_?���P��X?�#�֮��T6��rpd\�?�\�񭦼��ר5��ٳ�r��#y����lC���r��yy���,/���o]d&���ǤZ������M���_�?��� �Ԭ�p�ݺ{W�
Ƞ�}��r��ʔ�/.�/$�����ۖ۷�e{���b�D�_��\����� =�V�����{���C��\��x��*3��~&�Y��w��n!L�L�)�f�dI(z�=ط2�uΎ���G��ڕn�oΰ%�l��T<�0�6l^��L����@���$$���kA�,.P����O����㈵&��@��t<kw莥��gaqN�j�����F�21z�K�
�'�t��ņH���y��}������,�7�:�'��4(j�6�>�v @����;��q��-��bv�MAC��j2��[.��b�"����jKJ��6�h* b�ד��#鵏d��9��'���W��k�� ת�V�����E���C+��e��m)�~��������`���XЍ�6�A��|����wz
��h7�H�)�^�{��Jx|`�.)�c�<Ն*V�[}���'�4�	�i��FN�������k�/����������,��(.b��LZ�����:�]���ų2�O�/PQ0�I���1$��'ԚB�1 	�D|G3U)���'͇��ľܾD�S<��z��L�ʙy�v튜_=��׃����D���_����c��ԚyI}�s:m�ꖦ�}ϨA�jD�z2�;�N��,s���i���V��;�?�� %�Vx�GNV�\uA��d "SXC�0���R�K�,�ȷ38t����&쀞BS�g���s��b�,�?��OL`D\�oG#���Y�.2��H�!�N���}�*����f������}�?��g�࿑G�������ƍZ��k���NG�~/�������J��H4�b�wv��}�ޕ�/�4���!�p���~��H�NF�BG�-8;S�ǎg����	<�	�.Joڬ�Z����	P�mRKKGN=�*b����J!�*���X���厦��.^`Qާ��X>�����;2��*%��.�c��C&ek��B��p�!2J�z�N���X i�o>p�)H����w������FM&�1y�����b4g�Zk�!?�,
�\��(�z���E����`,�jSj��3��_ �T"M![[BpS,��X W�V��?�M)Ap�ҠÉ���x��ɦh_|^vmy�ɽ��=1�o�����WuHB�T� b�p[~����D��u%��\{�%Y���:h5L����O��)�Cvٞ�o� hI g��`>�~F���@D�f�s╆�F�����~�'x�O�#y��o�������ߔg��,�b{{�N�깋�?B���H'�Ν��8A��F�:<|�@�[4Pm��"ma���`u�b�j���	G����c)���`mFj�SQ66�Y��H�Úd���
:�8P��e�=&��@rvP��/Č��,�G���,5� ��>��ѭd__��c�?�P�NBl҇ј��g 1�=�J(*.ˌ�Q�)M�)� %�)?�2�؄
���@��Ѩs/N�pwGn]�L��fv BD-��!H�ڣ�fdr̢׏&^���Q���Rd	z�t@r��9���f��w�3W�1��L�9^�_������g��Y���V��C�a��g�Hke�t�Y48S������ҝ"�`�Z
Z�������2J${� �z�
,(bJ�(i'��D��z:$ê����g?��,�pUfV.H�NlLIאY�,Q�:HPIy�6�;	�'��x(C(n��\�V�muiE��1H�{W��
(��(�U�D���-Ep�5 �
?����i�hn=�����a�B�6e!4B�q�Qϰ�g��@Z�o�A���:��E��/�k#�;G,��ڳJ��km��e���]����[`$t�{/�SD-ԍFÞ4�ڿ*�k���="&v �QS �q�B�M��9>��&F�A��&Uo�����&��ǀ��.����(����N'ݚ-Se���F�-��e��Sਲ�7͖�߂[��F��@E�� ?��8�eF����6e��S�Z�WJ��[#�R�<�d2p����Br'0���c¢m��A���]={��͹���g�?J;iR����?��/r
�=q���k��?(~��7�s�FH/F�]2|LC�i�H=����S�i���=�;��9@'³b�ׯ^��ޫ��iv�����~�N-�}��:���ӥR�=�Z�i�:���H����Hm|Z�&�L���ϋQ�b��U��:<�{?}N�G�����A*��-�x���'�(�Y���~�^P�>�(C�k��꘍����Zxi{�\�s���+���z�R�8�_���P����]��P�ܻ>:m� �[�*G,��P� �lU��S?�:���� S-Fs2����-��Cw�8�4g@�d$�xp���'?���~*�̍Dfu9b{���uo]f.�J���Ԑ?�ݓM}?�A���M�B/�'3��z �̚~e�!�^�5��D"{U�B���Y���0�S�ъ���ۈ !��3)N?����\jD�ٞ�fPG�n�t�ܙ�c����(�},��p⹧k��Fe`����Ws2��u��
�'�]���E:�{��|N��:䗿���tbu"Հ��?y$�����
jҨ��w���i�.�����|��M��zO��>~*s�B���r��]���FY
) �v�{kVvv��}x�*Y�Th��t,�[2��쀉C�H?M��AU����⃏�<���,^������qj��'?�����E��,��E�Ɯt���G7������ѐ��F�{W���8�kvΰƑ����]��>�<��7Q����o�y�aM1b�'�zp8E2/�[l�ɹe5w3����a^糖՞��!yȱ:;���=���>P	 P�IT�XC�:���-����4[�:�	e� B�T6��RQ��57�l(�[������w���ˑ����9fu�fF��Tl�HqJ��=�@AA�c��Z�Q�s�ф㝐�l� �j*5�-#����C�����tE�j�p�P0�� PQ�b���3T�<��Ps��P֬��Xl~�/@�`�͗_�ǟ|(I��!���*"�z�{�����L]JE�%�"u
�`��oW}򙼠c�B}Y�k:�a�t�&�t�V�C�3����~bs��#�3���lE�{�R:�JK����%Ԝ����Cu(��IO��<f]߷��O��Zj�ѿ�o�2BtX_��B(`b��d6�7I����y�fo�-�6�.�c�(N/��Bv5.�wjT(�0/�JN�0V�L�d�a5u�HM��]r�y��Ԙ�ΔX��g�I�g����¡��E�h��9'���z�É#��7����a]IHAv�$���y��t~+8�}����L�g�:+�-��u���YPx�&�H��H�%uj<ٿM5�s�ۧv'W�s�iB���5����DtoycL{^��u��j"��q�(v�k�F[�'ε�!,��v��N:�O�?�7����4K��d�b+�jn������6鴙$E�L�6�[�R�FwôRH�?��r
���vW�Q�ryk�[��Y�S�Lǭ(�k
LKx^
��#��$��S/Pdm\�4�)�e�� �GP6ص�h�� �F_�����b�YSO}�D1z�%���y������;��6R�I��$I�F����Z/Nݙv�g���j$q�%�$Q}�Z3���O���J��Ȗƃ	Z� ���p���!ʭ���}u�x pxn����P�)%�Qp�Zs�yl��#�ZT���)�y
Y�AY��ƖS�Lza�x~�N@=�`n��M�������㾌�m5�Ǥ*�yF�����͍�><:����ln�X��Ԥ�°���1�u*�̴>����y��Cjxʩo�ϲ�eD(PO�7�[�G*���H��X�:�:wu�HaRw{[��ۿ�;�!����!���zG)�A������T)O  �C�I���S� �����gY��b���"l�V�S�񠵍��tV�T��d� ��������#S;\�X���������k���g��4�?�NA�o:�Jz2P|��g@2{Ϣ����QJ�ț�fl�΃e[By�Ց��?|��a<*�_5�5_j�68��
/�����K��J"4�I�EoK,���ܑ'O���� �������QxX���0��L�މ��+��Q_7S��<%$���]7Ru&�D�BP���m���/�H�ن#�R�Դ�z�8������Mut����=� ���c|��ɾ�#�cS#FX�㘀���ف(�bR���x�a��wYtLĨ���_q�2J@��*�{N�l�xj�t�&�-ȥq�8n-�ۍ��r��j��F��7[�@T�Yb�+�E����eW�������RlAU�AY�f6�PihF硅�eK�Yd;+��h�lP�z�):O�L~Я�Y��hԨ�O�0�{��KE�����m�p�ei�/A���搷MB�+����W��!��2��	�(�����+��'����WI��'CFg���ݞxj��W�^�����B�r�*K��z~M��y���5�t풬]��@tE�� * �c�����Ӣ��4 �`'!��i=ܗ�FYo|"��Oi���=�BĮ��� ��i���X j,��-�K_}S.]}M�l��[
��]Xk�-C0�B-=�m�X�71I\(Tu�9	�ml���#�;��l�dk��UЕzB�)ѹ{�+r�)��&k�p���;
�/���Y�Ě6Y�AC�F��@��L^���G�䳧�7�g���!�A1�J��2�5;�!n��dv��Bp�k,:Nt-�7
�+�܊�掦��t֠T�[�`\��(�v�X��TyƮkp����`���5�m���R���GWh��'���G��{P�
��i�S��Ȣ����;�M@�E�l�W�Nؔ�|^c��)�˄��.5�)�)���d��F�}'�J����~�^��Q�b*$��\E����[�b�kI�V�٭�~��I�(�S ���Y@ g�����p��t�A��S໺/�`���	����e]��C&�%@�g�c���,��b�e�',U�?-G�%��)8:z4���;�A�/��H�x^?Tw��\�v���<���ţ�9v@ݾse����1�6X�똞z�0�u������	���T�٢��9!�G_��8�@�E��{*a����LG�w�b�,��i;O�,��;H�&͠ת^�/�МV�gm2�w���!����y�u�q�.�إ�q�Z�(,��;Jk�ʆ05��� ��<�}׍�5�&v|4�a`D]���"#����*�����MVThtu
�e+="�90e�)@뽏�1S�|]�=�T�0jj����o���zF����R�}&�����!M@\$�'��2ך��@��o~�Y�46=����v��@�+t+�F��3j�O:�[�D��_�������HW���r�D�1Xg��N26Ih9/Fֱ�	�S� a~t��C���<8\����L{ތԔ�S��z����bU|��;�/��y�u�V��(�(SL���UxdDT������K
��C
�)�
�0��IʆB,���m|G��u#���1���l`6��k�\�Е��5a�7���N3�� 9T��^W��G�8��RH������p��CF�j�R�P��9���B��q =t��x��]6�f3}F����Lt"��L��ys�G�J���qz�O?�����>��i>�' �Ԅ\�n ȹfCV�����Y8��t���@e�ߑ#���9<��)H�ǔJ]�+T���~�AUjpJ��Q#�DfL���橁��ss��=���ZҺ�
if���4a$[��7��/�]�?��?�@Aّ:�7��3:���!��h��ΘRL����t����%9�wWvn~.�2Y�5�.�z/qQ��Ԕ��deeEf/\PhVή�R�Y�P�<=�R�@N~O�h�%� RV�3T��bʻ���;��'谋�'�F]�_� /\�jM����XO�8]}�knNΞ;'g/�Io�����@�@�FvV��Zٳ�٥:%+�b��S��#y����五��$���a�����}�����(���#�N�%����Wߒ�~�_�ٗޖIXӹ��lv	��h0�'�����;r����~Kv�������uu���l%�V��PG$D�u�K�:�ő7��Ekna-{�c�y�@�SѫT�>F.��V����%�&��B@Bu�Ւ�vx�����b��8��~�O�}�eЩ�����i9�m��ϙ�.ڃD������k(��d�ٟw�L~�4�* 3ؙ80�-�9�8�<�)�~$��'#:��\�h���H��:IZ4?�#��y�0��sMA/�9d ��SH�������ޱ�=��q��s�)m*�d��ב|�Z]�p���>��[���������z��W�4�}ɛE���57�l�����F��%9x����p<�:�	�P������\���d�;?���XR� �F ��Y������;y�4M��"'"Y�v��u�z9A0R#S������ʹDkb~�E����O|7�iRg�U����d���~���h^�"5^*h�3I'���Xq
�]��_�-l��z��g!M��7DwF�X}�	@��R��(��֥��59�f��1�6����`�qI͓��bӂ �7l!�3�G�H祻{Ɗ]�������x�%��o�������?�����{�s�K�z�ey��_�z�"뻲�xCڻ�2������>yNi*�Q�86PZ��],��	��o�Aژ+D��qA2�wQ���b\s����F#��	�����"$D����D�>���9�_�3�R�^4q���l�O�t�r�Eq�\�q/�5 R��_���T�IC�=��a8����S�hթJ'O~OO~F���˺�ёN7�=N�?�}�ac�4� ld�}�'�r��b�A�w1��32\5�В��
v*�QPL�B�#��W�� o�N��z�֊_��FC�f���Z��aG�qH���cFz[�e��M��ie���<e�'ꔲRE�8��Os�|ܦ��b��4&'�#d��u4>���.��P�(:�,G�ɗM����$>�d�0AZ��^8A!h�{d��b�H�Ia�}�,�j ���l�ew��P�U�?q�z0,%��(U�2��c9�@��ʔ�RR�bw�0A���9�eZc��4��(Mz��m:*e��A�p��H�j4%Ev���x˘:l�K�8\ ���%FA��m�d��!�G�z��b�8 0����d�I�C�x��ʲo��V�q[mBE*���Q�YI>�pb٘2��sYI_υc9���X#���E٭�_^�5rS��D��ٖ�m�08U(@n��WUЊ7B�([���B�T�!!���D%
��3�Q��R�$��$�Y4o��@�H�39ģ�L�Ǵ�Ȏ�	ݾ\��H8��cޗ��`��Y���e�ko�,��)O�j��o[��"={����9��P1@:Ӓ�+g�Yk1ۅ"�P'}v�.�M�H8G�ּ:����:L��+W.Kk����J�Q��V����ο�:};C�d���`��S�Ш}i��z��n\�����R�Li�F��ű��{۷����N����	Y(SI��5c���<Ӝ�l�;��4g?{ϢRY��Ȝ�$w^̡�k=�Lu�,5|H�t��u/��!�eTh~^��8{�؞/�1"eA����a~��2Bs��S���M�A��QIN�؃�k��F�Ĕ�'N��Dޒ*���[ �(Ħ,�>��B�˳�9���A�|N�{|�S0��/�I�?��~S\'D]qS�d<9�	�6�(�L'���M�Xd�A� ~TxM�O����B. �ƝJ>�gD��A-LDqq��Jez]����Z�G �$v)+�<��0�L�`ÒK���є+f���`&���&J� H� jH�.2��3�i�M=���q�p8��,� ��CU �ʸd�IT��ⸯ6r`?�H���Nl��L���/M_q�2N}v�ٸ}1�8c/�c@�a(!����F�#RՏ��ho�:��.3��������c4��dU��W�}O.��u��ِ{�ݐ�����=�u�hI��pPDuK8|��}�9�)=m�N��\.4���3p2R�0 9��K��o<U
Ⱦp��IV�i�R6�0��ڌ��n{����Q�q�Ӫ�WR�RB��t��EĿ(Cj���B�b4�r�^Vd}�!xޣUƣH39����X��욃B�,p�=��$^�{���ˌ�K�s�؀�UF������jͬ�مY�A�C�
@��p�\�����nG������G��ن,�]�~�KW�ʥK�t��Ec�O>���0�͙�|�\�|I���`
���>��Cu��p����[B��ǓX��ސ����1��A�Ϋ��$�.���7�ȣG�n��P`�+�F� �h���)a��yzm.��CV���9=�'��wNI|b}O����^qE��C�ɒ�D�(0�.���D\"G��l��eGT*Cp�!��F,���Ќ~ȼ���g
�!g
�8�?JYvЁ����;��\@
al�,ZWW@8wfI[�w�d�2C���sء�A���ȸ��8�%\+���	��������+���q{�t�pGƷ'�z�i�c�R/�2���DPP2��n��i�8j[�8�I�+1���+���~f��F��*S�?���A�?>����($��Qp��y��6=u޸^��g�~ds/���,--K�\r�x��;t�!Y�X؈)�5���).C�.����
��Z2>�׳o�g�:ܳTC�5�����S�u|K:&����M=����_�Y#Ȝ��8a@�
sbS,�D� �746�η�ko�*_��W�\��Ɠg�������9�2OE<�?�WC]n�4�u��k�7?#��?m]o=A�#(>�b�l�W��j2�$�]<Gc1��G�(��#���|ɥ�s�SȲv콐X@�l�7�rN:gnO`�2ӌs�9A!gN�>�
+��^v�v)��E
i��Ͷ��|e��`��w����X�L`>Т�l8�8�3;������d��(�.S���0�(V��ԄX|���1P�%�tJ`�����t�Du#�G塈6���zd{��Nv��j"ͮ��4�0��^��wz�O=~�S�H��������U����Q��
ֲ�g�u6����')����i��/�9:��AbRb�y�yvj�@��O��2S�fP��ySyq��KV�5��(��xFur�{�M&5c&mz���6�k�,�=��!��ǈ�Ix�� t�̉1
�EY�ΦXd�wY����BШ�4��D��j�8�Ӌ�+뾗�9y���!����%�"��ay6���r�\F�Td7�+x�#�j�V�c!$�1@�0|�X�:|��}�u�3Y��,-��}x,ۃ��"��������5P�Y_�_~��ܻ~S�l�膂c�h'��������_�f7�d!��T��V�Ο\���)�X.����o�+u�7[��P( ��a�[$�t�A�������cd)@p8����� (Q\<V*z�?���4fm(0��Qb�H�}������u�L��A�eܸ���M�f��V%�F���W��(�v:�P\#�ߋY�ܱ, O^+�/+�qp�o������wO�9��p�DK<ِ���>���K/ʋ/]�u]7���C�(ةVb����t���GABS��;Һ��{��u�����jY[U���i��lԴ�tQ��sp$��nPq䕗^�W^}��5 �ٹ�ƻoKE�ҟ��l:v��e6H�;ڤ"���3�4wA�%��+��jU�|eM�\>/��<�Oߥ}`@#u��_��di�L��$�m�l�K��;�A�g�R(L�H�4t�kj��E|Y� ��@�-)���X �z��[ι��eTWA,��	���ޤ��ӑ-�}�Um�-.���'[U�BYA۲�e�p�u�ְ7��N�@�Ǵ�d��O��cv�*�l�:|s8`��P�ѐ����ܜ��/����Y�ߕճF� �Q�T"d�A�]�������I)����@����o<��Ύ��mF�kj@�Å�SN�D� `�������n������ ��mC"Y�z(�+���A	+��u#v�ű!`������
��q{Kn޽!��Gr�>��C�s�B\�w�v5h*�j�~Q�Ԝ���g֤���5�#u��)G!����t;m�2���,3	�=��D:VI�_��4/�zE:.�N��ok�8o=~(�a���������d�"&z���P�X�: �Q$�74���뇂�k�f��9ǝC9ho�P�,�i|��#o|�Mu��S:�KgV����j#�@
����c'�Ϩ-� ����#�u�`�_����U�\�b��y�	�igk)�]-YmJ�hGxo�t!���%@0�@]�A%)ǖ}�$c�0��[�t�B�j1�����{?�i3y��`z~��f�+���K\�v!�3g�R
y�ud�p�23f����Wf�lh�$w
����D$=�̾����!�Ԁ@t��~"}��>b�M�{��W<6*8δ���:n�AaW��H��i?s��eU
��tN�K�4,QZ�|�,�e
�c�c�	C&N@l &y��0�YT*� ��oOG�Pɞw�0�.�S�;��<k ���;S�p��M �X�@�5\H���W�L�N���yj��8u �1�υs��/dM
@���d��`Bk���+;����}Vlt#d2��&:��:#�75 ��q�R����Չ�@�sX`��֧jQ)���;�ό*���?�������$$	Sg0�
���<�nj��A��:�[7�^Y�*v��x�Ã=����@nݿ#k���lK��PV�|C�z���r���ѯ?�޾.w�ݓ��-�;}��pUX��s��*�>���n��q�:q�
i⺮f 6-H��!q�l��m��A� ڞS=��u:��n���h��/s�Vpl�s+
�v7%>lSU	�H(�`l)i�d)ߓ����-vr.f6�ەԣQXx0ǙT�k2�� �����}{�(f\��P��M�B���N��vTJ�Z��s��]�C�x�XA�PȲl>ە�q���ڵ�27ߐ������d���q��ğ/;;[���<y�.����ŋ八�䩮���;�޽s_���_���~[6� ��Nu,[Ow���m�z�X._Z�o�ֻ
 ���[�)���6]�������3�����b�ٹ���>1�@:T�u��'���*�f"���9O��K�f���)��rr^�4�������'����F��FO;�f+�/�ԝ�8��6�jB���Y��z��ї������t$=$�b�ZX�=X �A
eQ¢����}��t
L$p�8�S��J�F���;��=��W�YMhSb��J��V~/t�6�����ǿ���G�8��I���5&C�����N�n�Y�
9��,������=_mp|��3�p��:<pX�Z�"�M���P�:�Gp�l����`��Z}���:oJC�*L@�@1�Qh��X������>�:�P��}��|��o�#���q�.�=t�Ԅ@2���0d= �Hm��'O���������>�1�n+@��N�Tk�HU�L� ��g����eYXZ!�1ג�ʒ,5[��vifiV�5����$)�2Bxu	�ٔ�~�>jA��CZ�(@@Gv�d4��N������&a��}�����N�9f�|��1�����R]A����A���X�[���>P�t"��bXw��W�n���63�����91L�Y!�	C�֢�Y�1��bM�zz����
���U�z9X�N �O회z�@S���o<��Dp(��/�2g���ĝk	OL������,[]~�5 %%UKH	�.b���g�̩�i�.f=�{��[���^L�����������Yp.�(Ai
�a�������PcaNiKjݞ�Z��6E�=a{���{/�ˢ�J-)������������h2M���B�r�Ӓ���/�`F���;�	�i�R�`zCY�&.�̂�:t$/�,.��}h�U��V/v�x��r�C���r߳�R��g��&	,ߥ�?/�����&Ӽ &u�g��6�(sF�dnQ�\ˈ�:���U�Our}��\ �Pb�غ5�bʸڨ�P��v�^1� �*�-B�)*`��(C�_FA%t��q� �X��P3,U\���,%��9aQ^H+67B�g±e�c ͼ(;K��bE��nmJg2T#^���r��K�63���.{��<�ޖ�[�<�����RN,:
K'�䜹tl��m�����̈�0��^���D�qc׬u	o5[�����٩����7om5��}͸c\Y��<�}lrP�f|�ԏ�̸qJ\T?r�͘�*O�A�jftODa�{p����af�5%�(�3,F����� d���_��Y��it�N��M�Bd<gd[X`�d+���~�[���{7��~� �Hj����t�h?\_��7:rt�-��y�� M<v{=:�����4m5���Sc�읯�'uP �o<ݡ:t�`g��rfe���ڬ��ʧ��)��}ݷ}�uڤ]^�zQ��9YX������e��9��*��H)h���q��2ث���k��E�@q�J&�s����F���N�)JY~��� d�)۹s)�	^t:<ߓb����0̯Ϩ�hA�����]g�8
�G��:Q�r0T U	��>p�6/�x��PG�W6�b`���*!Z��17�sN��a\ 
����!g�cFHa� (��SE�"��:�����Y�������9^ w=P�����GlB�Кi0��N���>P��A���0��>�u�-�������7��������١�SW0Xb7ՔŬ-��u�����r��Y�.�O*�釟S3C� ��걐׃,$�	@=��j��ξ���R�y���x��q�{l�TpJ�)����%�R��uW���L*;{G�����������cQ�D��&搤�����������W��+�����QW"�)�����-M�����Z2P ?DW�t̠qZ��Tc��!m0��ȩD�F�CpM".��:��G�jg�~����s��(h�, dT�������|�
�!�!`�l��ESǰK>x��
Ќ㡂A�$9�!�7ۘѥ16PJZX�g�v�\��Nåc[�E��	΂��Q��$.��^c�1�i�Z�e3�p<m��e���mZ�PH?��2�ó3����c�H6�KG�pE���:\Y@	�.����1��+�A����&��.��yH����G�*�1t�@
�Ԭf#q� !��!@�΀�$K�@�)�D�U�Vd��WVde������#�z�M�h���S����`r�2ԏ	�4K�Ǘ���ۥA���L����}7��s�s�/��< AjML+�+Ƴ���R�ZJ�EB���|^�d�����A���#o<��M>Щ-TF�SS,=�azv��:$ ���nb�4l�ʕr�'/\�	��G�_@%_��0�}T,��M56]C��%���Y��H¿)�]�8��L���r��dG�a��y
�=p�u�]��~��R]Lb��8�֕��)�u�(�x�,�Do ��-����,F
�%i �X�^H�5ρmD�Ag�b�1�t�E��� ���;e���xe ��l��M˚�9A�qƍ2�:�(u2�.-��AAF�6�Q������T`!
�kqfFϯɥ�^�o~�=r7�-�۩��?3��N�w�dggO�ݸ%�ֿ�ܹ��a�>\O%5',��7�΀i:6*C�bI��+#���ЦS�3bN�1q\j*;D.��>�hQ��7�t��F�0�	���¨)��ef�a@��l�N��A��ΐ����u���fҩ����;�䤝(�,gQ��d*��~�5yK����S�|�s$��槩C���4��!���d�N�g� ���X��D�	�Y���W/������57���<��u���p��̯�`�?���K��<����A�A�h2NMd@|*ˀ�C�� �
':����X�Z5A3��)d� ���� D | (`/��(0�K�+褭R��H�X{F�Eғ�-s�ɶ�c���H�1O��������9Q�P̈f��/f������<�A
���1�@�
y�]���`_���DPW����FU'�H��P�IeY�iҗ�"��Af�xY��e�kr0'qE���Ð[d�2� z� �>xp��noJ4�H��ޚ�W�V�����h{O�ߐ�>�����q�������uPս���-G�m��Fg��eee�c�L߃�:���hO���,Z���cכ �̑��l̢v M+�LU�Aw�@��Fn=ۢ|����n�f�Xw\�ȩӘTc�5� �A��N�5�3���مy�#���eh��㮞�C;+��8��r͊2A����=u��n���-) R'@��&C���S��HD`�ő:f��O��� ����������%�d����^SE?���%���H_�Dv'�45;���H�
�w�ȅųRO�'��
��Il�z���w�S�|tW:;�?Ӓ��M�����G�~G�i��E:���:�(��kU��С���j���ҀO���5\�7�����d@`��t���È�c=��������غO��@F��jU�DN���\]�g{��#Ms�
qL��L�څ��?��E�p:�P��˧_F�-�r������?������eg��*e�3t�}H��l�}�9��Z]�gL�)Ȥ��	r���;c�!ȳ'��2���"��L�$�ذgtO-,-O�w�AȀu4A�u]����/�ϯ���xG�y�mYY]�����l\��~��˄y`���R�m����	z��K��[��+�����ް�4�g�/�T7<ug�4(��D�0�Y���|��iT�A�_G�
�9=�ߌ�{�1�G@Y����L��	f�$Z�|i�	�]xʣp)S��s���`L��=� *'�B/?��p��)����^���I����	�
�ni�R-Ŭ�N Ue�^�ޗ����A�����=dzJƨ &!�zӔ���Pg�6��g] |2�:��K��A�$���
$��4���`N?�2��2���r)�MF��{��{��0I�I
m��S4vB����j�P|���ݾ���=�@9%f���㲂]�aSPFc�Ztx��d�%���80��H;�3�Ȅ�a3z(B�G�`Y�`(q_?��#;�}��4�ܵ��?�������55F:*�2<�U�)"ʟk��қ��S���9:������� ���a���
u�U(W��G���1X��Q���$�A¹�8c\=���
P�x�E	�BK�X��e�@�s��x�l���EÙ0F���	KJ:�Q	}5us��U��h�ܙ9))�l�A~��5u)��]�>�Tw@CdJ�C]�n(�*�!���E?L/ۊ���d�*u�GP�ѱU �A*�LD�s�F�"<Y��Y쌬8'�X�P�4�iK S/z�V3Ƹ^����<���k�,��C���*c��jIM��gzh���[<�M��Q���Ն�+X�LJrx8ҽa�,s���6K�_!5��۷>בʱ����J�nJ�V�Kפ���"㝝�n]��P��D^�ڋ���nA���<y�%���΁�eZcυX��j�����^p�A}db,1.����k�~/�"Q��,�sv�����^��3w41V�3�
��e�,QL� �V�H�_�L����f��J�_�L���QO��$�  ��IDATJ�T����+l@�Z���;�� qE7����Y5������g�q�︖=�R�ɩ����29�ژ��ٙ�P��1�����ɭ_��ƺ,4��ey��\y�%i땤��>(8K���i_A�x�|���H^}�U�q�ܺyS��o�F�|@e���ߐo��wYk�����5��Ԓj�[/��A���Ȭ �ӄmv�{���!U;gR���)f�Z��ČsOm�X��˗_�+W��:�<y���{̢ϫ�Y�p��0?�����k�]�x���EY�X�.�X�yt�����3]�:�[r�V�'�'4>��n?�vU�fmYފ��� ���fdz�:_p j�i M�� 7ޯTya�L�yr�ke,u�����#��_�TJ�#���R��vE�}��)���l��d{x(;�/=}���#�=_>������y_�^{[�j�N �pv�w��Nܽ;w�֧�ʰӑ��� @�l�?��~擧����S�zc:d�U��M�����ё�OU���ʅ�-�;sV��9��y���-�Ϟ��c6=[�����$����BD��p�����2j	�7$b�ۥ���O�Z1Y��p���Ȳ��e�6�+!81�z�|u�0�Qt(�m��8�&3K6156�l�b�7pR���)��EY/��L(�B�*;�2;��!��P_��l[~����&#�:�Gt�k�W:�9�$��e������M,��8ʠ���l��[��υ�]�4O\�=������<����^���ɢ�J5�c�i�3�`\)Cd�cm�ߑ��{���Pffu("�i�Z�e1�1l�8V"\��pE�x�����?�y���B[��k�M�/7n���eO'�_����Bľ]Խ���; pz�H�����wB��%^M����G��|�_s��l���9�SO�(����s�n������ I�O��M��ۉ��ѿ������2�'��W~�o���?>P�N&͐�t�c�\a?����~������a�.�,� C5����.�BCW7��cѩ����X@�}B�����@������S���N�R����=��@��4�­D��+�s��_ ���c���@O8��@uW�o\en�����o��o�-���~���޻)������xC=�Ϝ��_{K^|���u_y�<yp_�:m��-u�Z���1�UM� �%P�"�P�a�)R�OȆ�T��,B�bD��d<��7���sa>F�������*�� �Ho��:���ECOZ�9�{M:tA<������\[;+��P���dX�J�zoC�u�T#�&m���) eC�9)F�3��]#�5���5=��gF�p��s���Ӕ��AѸ�.lή#�^�}�=Ms�5���\�̈P	uB^B�5zw "���)�*��Lj�ɧw�|�b�*"o���g��:\"e[�B�"E# �aO���w~��r��+���!9��+D����׮���Jk�F�t��K��%��H���Ui�S�����ޑ����eo�X��.H��K/_QP�ʃT����}u.��^;�y�M�]�g�]�"qc˄f�)a�9���s����*���sSp�N;f'�p�9Q�iCEg�tT��>�8�nܡ��߉:Y���wH�E}X���:}��-'����CLЩ\�=|�t�������^��NZ�AA�C(tJ+X����')(V�,r�C�����e�̂�a$5�Uq�-M5("Łu�=ؗ�:�  3�96<�VG�H^}�E��?�W����8&5݇�����9�F�`��C9�|���f����:ǌ��a�hcJ�'\�r��������������'��!A��#�w��Lo #PX�vWƤ�T�M]�_����?��}����ݻ�������_���.\�?��� �%�v�pm�+o]�"[�RPE�<�ʽ�-k��һ���������W2�uP;�]�S ^	cY�|E�K	#����Rg��D�9��<�5�2�F
H�YSFA�z��מ0��~��#;�U�T��猥�?�~(]=���"�zO�>��g��`;�N�+O�����S�~���ݳ��,�-���}�%cD�р�7��.��:��G�㷻��l�P�X�o\� �W���ҙ����ډ�j/$�K%P;�ݛ��O>�_U��;W���Y\>+�F�{�0� `���3��R����h�=��_[�b�H]��w���]}�=�2�v.[V�Zߊ��S���2�.C�S1�b��Ha��QU.���K�+�dNC1��<_�)@��u2��N�Sr�>?2�04�|�5�j�t�@�t���5��6rà�Z^�����NCb�\����Y��x�ryQu*�3�gч�/5Iņ����9�?���ͣ�V�����1�;�?��΀�����5s�S�ZX�Y�Z!E���/u�QN���0�����<�q��s>"�5z�S����������66��8��@D`1VJ�hht�#=d�Љ�1R[)SRX�����9�������'-Y�
���h�D�|�Wz���xP��o$ֵ2��n��rD��o��QS��ZSd�@>����;?�[9Z�� �+�:�z��#���y�dW���7������t�wͣ׃�T�IXmHYA��Ӵ�+�	��(�I��Iγ�2�k2W�ndO���� �:ơ+�F�FF�$�4�R� �
���>S�VeV�IY�ИVg��F#��a��-%��:Tu������)���6h|f�u^�/���WFHRS��!��&�˦u��`<F7�y��ژM��Ȝ&����Ȍ��$�N.ΰ�i�I��x�벱���c��2,����r�ʢ�?8l˃�e����U���=�t�F�B�W�jɷ�11
2u͇CI����D��]�zY�����{뺾���Crx�#7�����Oea�)�Ν�o��;�n�s0b�����Y�������������ܹ}O>����W�}��r~uM�޾/�Ρ�*@
��^�LQ_�6%-Q4�(*�����B����q�\�읎����s��o\��or
�2�U���'���3��NK�[��V�Jk�G��@���@��\-��rF�r�R�9�%t���Ң���}��!_+�T�"����L �LS�R�D��ǿ�L�m�H��`]����'�wb�C�,t{�@z�JΟaֆ��ј6� �Xu�g��O��uK^�zM��/~O^z���O~&�uZ�Hv� ����q�ۓ�oW��4��7��ʇ��ˏX�Pa�0P>P �@u|g/^�JZc��~^ZY����[��?��-��|�����sN��vܺs[VΜa�}UD��`�����8%-)��>w|ܗۿ�T����'��>Tj$s�&���ڼ��n�ݵC/p�ַ�7H��t�N�'����
�+�g�}�z���W򤛎�돤�P���_]/�qOv�w��+դ�@��{�]��M������J_z:爴F
�j	e.AGLv��6«���h��Bϱ�:��Qح�p�Q�@���T��r��+O�	A����%�{[�w�+��� :&kkk���$��9�p�\�|AƳ���^��6���*���e����7�f8
�j{�>������#�hBz�z��"U��w�v���\����?a����?I*f�T��Ìe�����L�	���_�r�)�z�o<�eߡ8�$�G��5DP�L
�©	�3��	+���ip�� �&�Fj3�H��c���9Ś
)f�|R꼌}V!]�{W��/��_�_��ʯb/��译 @Z�m��z�b5u���8:��[ԑ�If-����< S�L\CPkt�N����S�Ϗ���_m����~�_�:���fP�4,RZ�FD�0�ј`�K2YNk��v���	�񴶬�ڑ�k(gM}�J_
�?w�Gɴ�6^
pBOֳB����r����E=#k�ˢoA�"Q��l}]>������J�pW��-�`��!����消\+
������̜4�2�XZ��aBn������
i�� QT�mR�H�g:�]:-@� 2g �d�JS
Lf�F2e�F�s<F�X35��^�"
�`����R�G����~_��IQ�L�=�ˎ��Ƞ� �4�ը�@�W,,e��Sd��$��\��X�sp"�І��&�
�|s�fcx�t O�2�#�F"@�k� �q��w��v&.R" >C*!�t۽C�����:R���sZ���X� ����y(I�B	T�V��^��\��*�����M�x���T���Aw(�#5�=����ַ�o[�?V'��3USo��UYV��Ƨ����b��%��
ƃ��Z��f��(W.�(��ln<eD�����
%g%��03 �Dߺl3m;e��!�,�t,���s�Û�Cq���=�y�$�T�����w�1"|�w�����h_�5��"RK*s�$�:צ���
�C�S���NĢ:�M}NY�Od�@X��L`���5LSG�F� ߜ�(�����5/������l߼-���s���>�ܬ:]=��K,:�c<A�H�Y5�bp��mn��?�9�J�˯��,,-2r����/�F\�O
M��	Z�=�G��Y�Z����eK� �!�7BX�a����z�D����<s�ї ��N[������ϟ������S�i4�:��������kZ.]�,cu�j�:�q����	��p�B��g[�$����B$��9.P�Fb�֜D�����eI,��l1�"�K-yQ�dfv���X� ���8aa��:U���r� s��Ҧ:��3Bf%)3`2B�B��QGJL���X�]���{�RV�'��:�5oLIk��%:����Y4�k���aL<u0��K�����o՛ry�����k:և���1�6���=ڑ��g�pւW��ey������i�4Yo���=p  M�@��f��4��g��3'T� c��0��Q�46��2�B�M�2.� �I��u1 ��r��Ŋ��~x�8]c�e8�NC�n�eB3�O���ASW���|�������4�u�|ؐ�z�DL��
�9�Ĥ����NL�Y��;�":����3K�^Y�r&a��?�%v�'΢@H�,<�r����`܍n-�W���?��x��-S����e�;p=x�%�
�I
CˆX����:.�T�%?s~_����)�'��ߏ����c��魰�1�W��(�T B�2��tM�,�80X���^e��bU}���z@��g���B=W@���ӄ��|�]M�qĴ>06]
P����_7g��H�(�J��n�&R�T����Z��:�����ܺ��C�M=z]��>e含C�P=qP&ѐQ��A[b�p�-?a��)(J#�4�N
8j�Xv��ʆc�?����Kq<30(,�8�Y^���Eu~zr��)c=���m��q+�RF����,�S'�K��z(�d����F{sXYL�PV�fj+֝{���v.�I�Z6d*��N�찊u� ���$��n�v�����à(i�
`TN��3`��Q�u�t��T4A��d�BFmj�8�huԙ�JV���Iж���Ԛ��z���W����c�zC^}�%���+��\��?��lm��Ls���� ��%�n�s��J��A^����\�p��O>&o�cOPSt���/�)`j0������JȦ^�����|��g �	�[͆4����� ��h�<O;Tá�s����es���Su�H��W��#'��Og��7 ��9�djA{]p��\D���t�2��
�}Y���GC���%=lu���G԰nSӲg���~�N2�E�2N&��d �kv�OE��HJ�
u�����:�M]�(@F���"7?����m��%KE�����5f�ڝ#���/�ܗ��ɿ�����,-/KW��'Ϟ�u;�*����Jف�1�%�T��eV�
��Ԗ�dH%����&-.'-_�|l���6 ��?������O���ۿ�k����E7���N��iԫ��8��<u�Rs�d@�<?O��V����?k�����8�¬l�7J�������e��*����M�Јpk�����������{�.ɮ�J�<ޤ�,�P�#@��Z�zF�f�җ�������0����[3�Z3��-
�@� A��ʡ*++��o�{s�>�FD&����V�2ü���c�ٛ�YԠ��ߩ���O�9�i�������е�&.a����8'�@�q �9
�D�3�����u�����LY�101���Z��{Q��g��In$�0w�йȨA����ֽ\����IY\\&������tC1�q����o��0I�0�:<oaa�Bq � �4�_�#}�}U.^�"�����E#�|�}��ܦ��GE.=�h:���0�E���LC�~��}@�_��ǂ��#u�6s�?�+W/�~�y'@-y5QH��G$>A�3X�U9������C}&�� ��CZ��I���׭qʐ�@:�I�P �=�V*����A�]�)@qv;}�X��|no�q����Ȇ8B�������ŭ��a�W�5�6���C p���������~�)��LӦ(�⌔Kb�}Ї*<<��
��X������i��䘁�<��0����c���	�.�Ick�k{:A7T�@'�JR�"q(Ⱦѽ���\�xJ.\�(��;"{���9�yxjqY���P����C�Qg����ںĨ��(}�q-P�d4f}b��5���ؗ���6�
�qc+�\���R��j{O�$:F|��ʒ�����s����#y��/k;����"sJ!T���ʠ:�bh�?�����
%fC����&���%P@ѐ�^�x���5�gR�}L�Y���`����N8M/�l|B�}7 NW�����d��+����i�AC�_�r�1��
�VnU��XekE�Ԡ�5I����ĖN,��mks_�#��ʙ3g�{���DqB�c8љ��䂲�mh ��|��S2W+K�pW�}������2��>x��{U�{�%y�ͷ�����uZE9h���TQN�
�II4���{�`�p���zKvv��ݲ��q��u�� ��q�gss[��i�!$�s`����`A�s��Lݻ�0_�:%:f����7�/���L����� �v:�M_�,e]W`����������L.�%MՖ���1��@Ǝ�K��i)E�`u�\f2��QT��/2�#l"������F���y��v�ph����lmHl�.V��cH����5+�����|�`�F�B\ޭ/���w	�t�>8�ǸB_ �CW�H�1g��U�Y��XHS�)Ǒ��ںC���ݻ��c���C�裏eso�g�7��<��ζ|q���F��L-�r���u���(����G�"0=��@��bzP��	��3K	� #؏�})����е��uYӳq��M=�u��r�K�tQ���3�;����(��Ls�I��"
l:��02�N0`�T,�/p{� �?��������{��G��,�� �\���V���|n����z��a�QlÌI? SB��h�N�7I隙��}g̰-o��}���Jco��J��� ����y��o��ן����Zj�|/������i6��szx|^`�5ӟ�yW|��,::���
�˹N|N����i9qr��)t�ew�HFN���ɡ�%7��Ǌ��˞uo<�&~^ʒ+:�l�8����u�:-&~��@��G��'7n�����>g��,�&LF�M��C�d�|E�W�\#S��~�3��E6Y��Gv����tx��x��?��&)�#}�|�<��Cn(%�H�49���u��0���D��$D�1�Pt�e��(5���:pF6�8U���:�j���3�@,�5��5p����А ���u�k��~A~�Y�G��w�����aOFO�Y���U���?��ͦl}���6����dL*�	��!���lD������0�����Tv1���O��K�[<˃!O!�6�*�����hr��
�L>�Gsuٕ��C)��fu����%+i�T� �QyP���mmC&ęb�:�OÉ�J�j(p�)�ڐ.A1*��uq��Ҡ� 6xI�=z� G&d���c\R�GN' ����N���c�+�Ǔ���shUmT�˅n��`�K��Ҏ�0��Gd(I2�ʪ277'O_>#�e9��X�V$�֬T~(�;�t�2�E���\NʥK��ݷ7����3�+'���6�����M��/�I�m�ʩSr��S�cw⮼��k�C���l�7e]�͝��;d�Z>Z��{�瞗����^~��-�o��̂�=1�����dskG:Q�uX�_,���i��(��#�����+"����K\�q#�h�`
�G; a0�č�B:�=�����`م�~�#�>#��16t%ЭBp��B,U�����M�g�5
"8�C��C\UM����P�����d�H��\⠑`*
4�ǰs��Ao�v:}Eu�����@���+N���h@G����5HY\\d5��s���_{���*U9�{	���u���-��m��0��1���팺7��ļP	�rt� �Z"�􂣻l�C/g]�O?�TZ�Y�Μ?ǹ+O����e�I(����MP�v
�5H>��0���k\6�HE�x�1��9'@5} ��L�*:���;�z�8T�Թ?;�(��g/_޽�.:go����r}v�n�#cRCe>���>�c�fd(f�V�g+7��Px2��/�1��,qM�O#
u���5H���1�9:op�c̓E�����Сj�.��r�C��y�˘���W��op�d^̪��+W(��u>��H�k�WDZ�FF�A$7#�} Ω-�i]�^�"�j?0w4�{��{�ziaF��r��	��.X�W���bpP5�;%��ʸ�3m���3mߧ�$L�2M���
�~���犮{R�{�J���1+�x���!Rː�.�{j�"+���g.Vɜ���@N �~}|@�QG�X���f���wAC� ޟ�B������d�������g���C�ZQ1-�K6�Q=[2�MՈ0(�c��C$�I�P���l�P��!����$_�G�P\���¡�wC��@� ���A��E�Ñf�2�Z�8X�<�efx����ò��,=�x*1k���n�ʌ�7h�� G_,H�A۰�Y6����2A �pQ�I�ِ_ޑ��K��y��W��ڕ�o�~����z�����}Sʏ�͵U����y}�ؘRR�
��Bn��T���t<x́'V+zFE���TU��C��TŃ�(>���D��O#�k�����H~��GrbiN���	P� unPO�dM�0�5 ,�
t~�#��О�.,x!��CՋqL�`x@�nr��^ ��-	D��j'* �h_ɱ�"��A�`m0��X�p�( �:���Ȁ���qz�l�1� ����A0<u�4&�����xeiZ>��M:��F��L8	,y`�æ@�c�y`lQb�=ԛ���������H�6$v���鴇�؀�g7o���ue2�PJ����$9iw����Gy��#܌&��r�t5
iv;���}�K}�m�c�/��j&_|~OV�˰��{X�Dc[��s⸣�n�{���m���!��C��H��9�\�K8p>��8���ɜ��'a��������������x��.�!@���
9a������6���q�\�9(~�o���&�02�n҉��~���@Gb��F�0���>�څ�o�BV��4x��]�`�1W�$�w�	Q��Ν�"��_����'ʊ&�~^��\N��k��mX�Ly�#}���EY��'�h�w�	�#"���{�Y�bI���84�~�[[״P�5��%��#)U�Q��� ��[��ݺ)�n�b���A�&��
�$��`� ������B�j�Q;]2&���aÁ�����$�s42:L�,�vv����o�~��~�mYZYd��A@���!�zi�@Xo�?�|��'
z��;$oH��Ǖ�N;oMT������	#��j����T���@M\�h���)g��i�u7A=�9�{�u]J�&e]�긠f�]\�G�D9|�e�k {��S���p��9e���9�|boCl����3R���~�)=;M
f�m ��<ν�j\������\�N�}�Y�__��&���Ok��?	V8���=��i_1�>����g�LT�A����㜌���|�vyN�#���1�5��tj6rB
"&ܙ�L2q���S�`GcJRt}vH	$׮]�æi��o���X+H�2�j"p~Em��]Æ�fB��Jf�t���՟R�������z�l���`�盤���q�¹��z���A��@e�m-�F�F�	���b��  `v� �#Pcb>gDjSq_90�23\#�a�I�Eg�J�L�L8�af�Έ�L�h �Q
N"-�ψ^�p]�%Y� ��;y����ݷ�mU��y�6+V�:C�Y�{݁t�:(�&C��C��t\[}v��8��D9w��������0,cC =rV�TOɑ� �0�����C_>`��X�D�A�)MB�Ν;r��,>{Y.���䠫f6�,��������po�j55h�n=i���^+�l��'��i�jdj�#W��Tj��[�j��پ �7�(������L	NUL8���d�@_MAP�6M��Z�	����8�<p	W�~����4�~j�`8k0�����K*b�¤j�q/G��nmc[���b�^k����ru�� V+�E��G�8�y�]@tiw�A�_T>S'&a�N�ٓ�Gv��3I	ف���<���]�d��z5��;C1,M���H�9K;V�L���a���xVj3$� 8�l|/�%p��@���ݕ#���ۯ*T���������Yj�~�Ht��۩5�q.xO�L�l�M=��FC����2��c6Τ��
�Wd��@v�Ԃ�C"�#1�&{1�����O�BH�>#��W��45��`ڒ`�,��(g�M�oj\�!x�=A�6�C��}x�K�7���:���?�[��p�H�#����~�|��_�h��9�C�+��|��kf�p�|�2��y\Ltz]�֞,�\��V~�'?f��9�3�b��p�������o?�2q������<���b�`�G�.��CΈ
�Dg���n窺���zPOD��@[��p8h&l�?���Ac�:2��Ap���nk2�AGp�b^�S��0� �[[�?dP��|��I�Y�@�A����u��,"`F�$�(�4�7D��T�4-ED�$�J	�ޏ.���^t0�����W�ߔ%�+˚(b��֦��=n��8?��[�u������L�no?a��צ���h�z]3�7���)��S���W�,X[�u��g����3m�1;B����	��p"��3QB�=������T�1M[���C�:Bc�	��4�s$����c�, kb��S>7.b����l;��~��<X �4O=�x���d1I��Ɲ�ϛP�3�Sje��i�LuƠ�s�:�d�j����-)��dAmL���+�o���G���Q��+"� ���y���+N� ��]�MR�u|������O����7��h��j�bVY�����9�غ	NЂq�����i�����!�PiT#�� �a�C2`�4��|�� ~؃'�H�Y�$%1�qf���9	�F�w��oK�ɍˬ~|�˻�0t�������'�~��4������=���jā@�<��i��u@$t���̮��h*�O����:��E:��l�0��L��af����Z[�*v�����N�ؗ=5z}u�F��b.פ�+�ǀ�ru�i9�qC����[�4aL誟�j��+��>ո�#7�:XYD�+A�1�P �Q6n�")��!Sա#�c��t����G�^�j��a�׌�2Ϥc�&l�,�9�KEZ�����T��l�<$��r|��<��؁Hm�L_��P�DuBx�Hoo4y�U�X�K؝�0+�C:FGFw+��!�o� -�d}��V�[�&9G�!K��Ab(����'6Y��������Y����8C��{<�0�����a�;�YA���e�m �Lc{[6�ߕ�q(s,b�X��<������{g�v�Q�$�D� ��L>dY@�Ό�&�4zb47ԆU��"������Lo`sS=}9h#u��	8�اh�=XW� ��wߕ��}�d�h��H��{p ��ם�U����a�ip9(��8�F 'VA��a��"�@��s�'z{$��k\���
�tP�S�T�h �����h2q�qM�B��&|ǜ�G��	�v!H��͞���`��L�"��CSZF"���x�CS�7��lV�E�W5Pb�JG̎i���P-40�04�$��`��P�.������Y�5t�H��9�;b�$є)���z<�9��'������S��u��h.w��7ݳ��F���S$J��,U�����j$�1�.�V|��Kq��|2�m0���/�;�%�s�.��5j�u$��22S������-�b���۱��&���7͞����1��y�m��2L��?�w�'�g�3@�ob�J@���d��:ɩ+����%an�������$&H�l_&���ܰ�]wB�⁌3:|����kB��*X��w�����١f��V??[õ&�8[���y¾vv����C��l;;�����f�������$���MR�G���������w?�� ���������0�Y��1� �!��P�0��Y���>p���?�8(���!�Jq�Qz���s�B�@B�2�h�*!�$Z�?�C�����;d$���i@���'ҿsG��p����z��鬀bT���rowG��0<n��tͱ����&	Q���G�)�kD�=��L-��"^f<L/cPQv46*��3��V��jf��ge�4{��9YYZ��jA�zm�� 7��6(���& ��f�sg��K�ʽ^WһՉ��^~ft6&�Ժj0��3S>��� ��N^��WD���dC+�!'ӆi:�����x#<A<��M��}��b��M>��g������w�1��`>���~Ȕ{y� ~~ntK@cz�MlA7+�~t-��x��,��M��	\�6�$�E�#^rL��X�煉Vh�8�W�e/�k��?�p�%t����>@����@�������;�6at�>�!F��M��&xc'4�
=)Q�������uw�'	�3�!^h,��r�C�9Y�=���F_]��*��|�����I�j�O�禦T�`44A૘Y0�up�Kc���u�� g�=1�ȏR�=lH�s��q��}t�P�FבM��=��$ҭjP��/����y�2GpV,����r���o��v3R�� $ �?h�Io�@jz���J�7�@m �C%q�^�V�EL4����#�4��-T;�f�P�v�d$͎1�hr��)YW�>`n!v{k����� *�?n�2�g}a ��_\#:}@� SCȢ��/�VKU��N+'%�
���*rش`�
H�Ç���g=�S�Sʚ��@3���v��P�*�ܢ�Ы��~n,j�ڒ��}�$@,,1���:��vLۀ���u�{��������O4y]P?k�R�{\v�=�K�.F��}�D�U���@w�i/\R`c2��x���_h��#Bc�*ꙛ�b�%0�qT�q�+hD���:�����o��W��?��;޽�N�}ۉc����h4p���P!��E�*��h�z�g.�� P��z��5���ڵ2�d*ΐdG�BWf�R9��R+>�}������Ⱇcb�{�,�1'��LM-�&�H�I�%��}ݳ==���	�cs�k�c� 5�8g�iTt��V 	&6M\���O��P�٤����7I���?���;����+��w�����6 6�*�m��Y��h��ٸ�4}('�
�ё�ba
1)��f�ǈ�y��]�BJ�,"x�����é��@�����K��j$� `�b��-��Σ�l���4_Q'��W�J 	���;E�D\��(m>`��+^��4��t��ț2�v~�h��A�ӡ��Z-�����<��3�Z�&��@�[avA��%��@g]%T�f�]���32s�f�d> �68���A���[�`h�VܬB���,�dE�3���Z�&��n�Ap����ǫ�O
*��S��ٴ��q��q�k_� �d�U17\걔V�w�;#Ec��.cNR2d�Y9Gbݕ���2�o\����6;O[o#�0>~jY�X��4�x�߾�?_f��ޥƓm��.��ܐ*�N;$5ls�M���̎�������5#�;��u>ȝ�˯����������M�Al��C����������˄.������̧%�����o7�Ep�P��ϒ	�*��$)��m���&��R����v�6��}}^�;����1Ȥ�Y��u(R��R����AC�p�X]]�����������৯�fe{��PO��Y��m�HxJM��v��p�ryeMr#�.��V�e"!(�F��q����!�Ϯ��Z����!�{��ygc��)^xF5.:���~a!�Y}�@-.ɩ������֎��i�? &��$L���s9���}K:�y!��Ƽ��t8o��5C�0��@wDQA݃]���4QRS�!g����vYV.^��eݺ%IS/�9�W��!O���lO�XC�:$�zPDƼ�a��/��1�+�ZT3#ah�5��Y�뱠�.e����r	�����:��%��N���}v`��f�D��NF2t��ȳИz/���g��ލGϮ�kec&��������Ƨ��'�<����q~ ]�2�3`!�V�lV�je�(d�GS��4@��Ѕ���(����_��#��s���h8Jn��0��5Ĝ⃜&�E�$,����)n���P?�'�r,E��%�&�Z�@���A��uD�=����Q�i�L���<�h0{��]O|���������y���V��.|��GK���I�vb@!3܈�y�P�*��#pB�%]�2�X@{���a��\)yq����~�DD��D�v$����hG68�D���g��
 �?�V�4�`]PcWV "8|i�ϋ��"0�J1 ;�;�NN�J@Y���H�J��`�8zPΐ}j:���I�&��#5���D܄����ef|-�z�	q SE�)���R޺'8�iiNz���=��,?��Tt���R]^����ˤk���y����� �"l+!6�= u�:�,o\�Q�㣎� $60v���N��3D���t<����A�������#����aB8Z0i��E�j9u���� �bt:	��L(�Id)��;��B�`q�
�}5�=w�1��]Ǯ3Zah5K��w]�1S$�Z�e.%0#�����Z�j�Å��W�H4[B�:(H>�hXYx��{��9*6ʎ���f��e�P������;��Iݸc1�̧�d�/I�x/]�.3enR�;�����Iq(�H����<b��� �k�ق�)����J(�<�{�?�k,�b`��F��ʲ�Ԇ�	p�h&�����ˢ��m��JsOr���� X�;gp�9a�6d��c��{��~HH�;*���A�٥�����ֆu)5X-��Af8�bY-�YaF�߁^�쌜�z�Uͭm��@�Έ*˦�`�/��:^���&�|n���o�{�Է�ڃz׌��*Q������}��ڦ�>x�u.Uǰ_�U��9h�z���]����)�ܸ+���?���}����C^��..���-1�=���݃H`�׉d�^�S��,΢%�M����0|�F_�|;c��&�$$rVN����~�����;28��Y�vQ�����%���������j�iZp�{�U�����N�Ęa�g0���_��
�Q�yά������V;s�H1A�̆��F��Z�T��|��#1ּ�?�m<e�q�!�����P<,���I��9�k�������u���q��H��4w<IxR���FH����e�K��:T�Ŝb߱�QQx�;n�,�C� {�w�W�cw�M�w�=�h��7������m������<�mɨ��
s=$�6�#>�uG=z��6ӄA�k���o#��V�&6
2rz/��Θ��!7�d_���a�c׋���o���������/��������������#l��d�a�36BWQg�G[~�R��5�|8�/�X`�3c}�C���]ˏU���O��|�g>C�->�3DbJȐ����%�\ʀ	8�8@��X�?�a3�BR���9�|P!����O�;r��l8r���UY�luXBC��x���%���Ϟff���Kǋ�d����~Kv{(^�� 2Q��g.ʙ�ޔ��O�ő��K't5Ա�����Z����0��0g.���J3�9T7G�r� � -@ҿ���F)K%�Y�Ϡ�%j��ۊ����}��_1��O��di�G2�x�k�����\����W`�C���c��ƙU�2�{������Az벚�}�KR��3��)0�M;UKKt@W������\��(cCqP�l�%gA8�p���w;b	\RbCwx.�c�M�ΙFn��3���#�p���S7f)��Ԙr�1��h?:{R�8�D���{A��};w�`�B�N����s�y��F�����|hI���@�AA���p�p`�sluR���K�R&}B[�܂g����51Y����}�YIN��������e���p��'ցm�ՙ#p �9`#� �; ]!h?��&�t0!:T�1�tbE^}�M9q����j���a4�8W#tGC)`�	���\}V���y��7�Z����}W��B
P}v��d�T4��
����k�1D����������iP3'�rM�LT����b����c�:ܷ~�sr��3�f���r�ݔÍM��rE��`�g�C�j#���;Q��9 ��S�N��~�=9�&F����+��bsh�N�+S�_1�(5P����W��� ���xrE��E}[��9���P;�ֵҤpI�����(t�3���%Xy��cF�Y1�	l(V�����}6��(˚�|�2Y���:�L��o���"s�70A �N�������h�"+NL4&sdc�q1(��N6�@���;8�*���97ִ��)m��j�q(�8>85�>q��OJ���u۶){8.@�8���8�CMԻ쇘iΠq�����ݤN6M8'sD�$��C�;�K�"��u#�y�r,`�������'�<��=3�֐�B�nS6=������۲��.�v�3F�-zԓb,�I2ʗ�F�> �0�\%G��(���I�����E9BA3�����MR�5y,�y�޵k�������{�%qa�5��%Z���Rpڑ'C'�4�9���
N%5��Rt�-i����8�\!*3=�hV��������� XE��/��_�����s
�^�l��'�ԑ���i碔s r +���.���j��P�t�*�\��0Vhx��!���,����S�����\�(���eMp򕺔f����Aq6����\A*��I���2[�I}	���#��2_�Hb*�S�q���e3ܘ� ~��Y
v��,�%^t��*���Y�)tA�E�*�i�{<�y>I�*��%��xBu�}Y�vcx�X��HIll.�&0�)+ڽp4E[��-��'q|�6��A�{$����:�Rf@�O��Ag�nP>�jq� |�㐱Kl��6�,.8��˔4�qrGe�����6>���ž�ᘀ|�ʼ�����ڃ��~��bo_1t�(A�a[p?����I��t�q�c_�����-e����+���i�U .��c� Α�R�/543?�K浑%�QΨ9�T�A�D�b?>���,� W� �O=�m}�Ip���������ݗ���r���R���mo˰ՒbZ	h⠖��*g~Q�����\������s������\}�:u*6VW%���T�v���љ8}��<�����+��jp��F�ے��$X�X�Ap��C�$6=0!�������6�R 4�j�������W�g�%ͽ��>|l�ۜ�Ԝ����V��j��˒�w
�R?_������+����
 ����g�v{�D`�y�[��3�_g0�����5�kN�B8���k0X���iO߹��2��e��Ԇ(ND�2��Ò��sn$v̀&.�B0��/�=�i9
ȥlT��E4�7�Y����܌\�}���c�NΛ����kN�#c�	m��?W�׉�ەsxS�{���E�LgvV�I�=�)HIE����>��L��3+�"�u%�qR�$��4\q�X����t���ⴿ���.�  ԭo��T�޹-�[[Ff�A�H�=�م�wG�L�-6{����V������1bGt10( �(D,���($bV�V-��ʒ��U�=�+�K�g�O�Y䘋
����(V���JEK��=���K�;9�փ2쎦`C~?L�}8!���턩�7I������~�����/��v�Y.A�bNq��S��ÓC�9��"�96u��b�ɖgO�"x]We�ۖ�&�æ������1˨#�n��Ąq��(5؈�iu ��e�0j`hl`H�a#�jE������ΰ�h�6 �Ü��q�&b|�����l���n��AQ�a!#
I��U���+�߅qp���L!0�r��aT����:3#+�'4��Kkg[
��,]8+g_|IʧA`�_Trm�#���X������l���a�hP�����@�		����c���7Q����o�YSFL9b�WMU�3�$�`�3��9A����P��,e��/_܀�P��k�YKwz�b�p���n�;(��ibp��]�����|�Ă�([1G�� >�/�;�7�k� ���0��� ��͜�28fP5��	C��Fn�9p�i�(��D�]XR�~��<0������LX�A��+�L��ӑ�e�.��t�VYs���Q��Ç����M�ܟ%&y�	T��ق��31��q�03�_�����'�1�������`E�1.U���oܔ��_����K�וx�c�xd�5�f��i�b@h�Y~=�pQ}�P.��	�Y��֔8\�)�	t����H�jV)���a�����R����| "F�)-%�?�ZE>�O�3}r��O~"�/�G�����٨�����f��O���n�g�¥	Ș�]0MF�����f��١v5ֽ?d�3R�{3�P[��7���g>��2�0/\��L�Q�f������~[N�8'��w����{Z����5��P��h�V��X�kD��ە�h��5�J��$_���P���[���	�-�N�:��R���4?�ܖ��i4,��9�]Y���l����ߓ�5�!4hr���(�����Yl���Az\���"�P��a�ۗp.�)��{+�6��A�
��^��v���SoK�?q��J���؟�� zֻ�4G��uA�l 3�8�0�q���l���`%�,�8s���E�����s�7� ?��5[�n�K*��Ɓ�_K};R�4Q4̉��������I�؏{?�
)��5)�t����{��7��o?�-`��ohA��1���I{�� '��"5/�Ρ��Y�w��hx돮���0ᖒ��O���I�ߺ�u?6t��,Fa��V��ġ@�q>o�e�6��5?;��HkZ�i�x�h�Yhh� ���%�����4����z|�|��Z�����o5vd��x̞g�^�@aN���G�Y���~?r��V�3B��� X�^��F�`C����MfM|�X��S9�xC���p��q4m�����`V�l`k���5�.��B�&���:RǓ 8/��~T_f2i�}��&Jh�#�G��CY<\�d)�R���&�'X� ���ؒ�T�gd"eɠ�/�;�������;D��-u�ϼ��\�~U_����E���ȝߓ{������3^�☤�;����u*����o7�Y��dL*L�X�XhKנ���jPA���ڷ�DD�\8� 6�I�G\?�Bpp	���A��xv*b�#vep{��|��{5͉����n50v0nG��$�^b���3�;Lb�EO���5����"FH>QsI�O��y*p�s��a��?�8�� ]�d�����rA��И*/u��,����Mw���l#�fc���O�C+���xp�P�F��m������,�kݾ��d�W�q�.��xh8�4��
Z	�b刅621�O�!�!0��	Du4�¾@���1�	�E�r@LU�6�`3�o0���� ��J�������1�א��̌zR #�*a_�&�f��)sKR���*�u7"^�HlO�2��G��1���h ��Ѡ�P��֣<�ruN����n�� "���傴���S}|�^cU�Z����~g.��������7�i$K��D�Y�e��U��˚4��})i2��ez:Rυ6Ӥ�<�}������|��IIE��Z�T1�[8�����z�
��Q��~�t���������瞗��e(`n�јB�unfP�cV���Dj'ڭ�̂���?/�R���ȹ��,U��7<�z�*��$�h2[�a[�LA_3_�~�+�n��^��ِ߼�����JU����
���:�Y_ߔ/����vT��03��]��ZU:�
m`��~ӃfCwX�C����V)�P��y(=�������:>QNm�Ƞ����8f}����;�6��q؎��?������ڐ�����LH^�>1��R�nc�z�vB�Y8"�5IT�Y���e�:F"��Q0/�|[S��1mG8�Ep����դ��h㩩� ��B��u�U�S�q��.��}Y!%�cW�ɕٿ��U��$7<lxy+�A=���\��(��;;��`uK��{LaM�D!���x��)���u�RD{
[a�[7Q��.���Lh���tlC9�6�����b����w�U����3�/m8X����`�*"�Ȥ\/1Y�uA���X! �px�5���f���vw�63 s�g�K-I�BO�E�}����N	�I
�V�|��W�c�K9Je��?��-���kٹ~^<���8�� ���yT#E�ٵ�}U�ZYV��IB�mٸA/�Ъ�5
x�`s�õ�=@*(}z����?z0��4lJ�N��A2 �rh�� �Y@cK�M��i��9UK�����<h�RK���c=Gd���-6Ę�ztȠ�c�~x	���1�BP<����{we��	�]�,��E����v6�O>����?���ߒKW.���oJi��ڍ������EДE���t�K��Aw���J:*�#K����-V2�D#V�P� ��팕J�V7#�+8�F�b��d0�G����52�h�3�qp���	��oJ��C���7��E�#}��7�Vf���&i�� *X�L*�nS����QA�7\40�PhՔ�~����wM��ȺM�鈙��T�51��z�>+A�|퀄���#xY̛���s� $�>�*ż�H'&DX���N�k�� <�A�3���{sp�k8e$���֖������A��y�N+��li��3�w�.q�{W��^��>;?'3��Vl�PP0���hH������P��*��Ca��_��w�������4�~E�S���2�t�����	zG�sM�\c�N����C@�K,y",���B7 șR� ���%#����5G�Q	���3�پ
l�A�I�.@Y����{Vk5i�m�>nK�t��ċ�r�g��i2�@���.��;���/�����<��@�7wt��X������|��g���B�lJ�^��rQN֊��g{I���n��r�I� ��5]X�����I�U�H�'Oʲ��<�"0������k-,,ș3�dF�5f���A��C��-'�WȘ����:Ԥ��ɒڜ��yY)�P�����Y�캙���)kp�����z.������!)��a�e���,6�7��<�W.��m�;�ʁ�-(�#���ͅ��/^�(e����\ ��	tc	�[�L��t�	�l �G�ŕc7�LeV}w�G�)w��#�9���V����ΗR��gk�U.��g���`9��)��3k	|!"�-;�bԤ���	��d����u	��/\y9pI���!�������,�/�X*Ɖ��cyL�1#�W0�`s�����x����o���"	�i췸_�$33�.H��Y9�:����iP���An@���abb�Sm� �t3�S��|S4ImV1�A�f{�ghW�v7	�,&T)2�(������x�H�}u��:�ϲ��`�(TB�,F򐯲��}1���n�3���v�v	��*�Go��$_��:���hX��Gŏ"&�\��M�U�*�&3�-0y��+�0��Cƪ��^EP��� ��;C:4E`�#�G���f�LA.�웬pt���wr���Ҳ�{�9�|�,i`F�ή&{ے>�'A�Pr���\)�C�-�`�����Q�G��B���=��q���4&��5���������đ�ڠ�>2Iub�a��T @�`���8No|���2�YN�X��9��s��M�͇�o�;�?hJqX�;�{R��r��g���/�(�DF�%���("k�'BPN�TFp������oՉ���"�E��^�!}�|T�7 ��и�m����t-�fϠ�!��i@��B�DK�*�ܱ���ǣ��S�Q*A굖��������A��D4Yu�� lC���= �#���;��f�d
QD�0���� 335:�|j�7tE��N��~���� ��B�7��jb���h�:4�eVcc
<�� �R ȇ�M0J!�A݌Ô�F���"��teg{S�CC��@{nA����ST%|�A�A�P:�-�eq�/�p�1� �Y��`oOv�6��T��U4p��fXE/�AD/�ji@��]�p,�,��2���������y�j�[����Y©pP$8<���X�w�ѭ@-�{5J2x�q���<���m9�k��	�<f4��S��;���#2ep>���}����zj_�0�3_�3RD�$��+�h�{�s�9�X蚏�~��AϘ:z|��vu_�u?�~��3�X[ga�m @�S{�{�;Y�ߓ��;k����V2"���ggf�.7��.׮\�������` [��^Z�gO/�	Mf ���ٰ�3�R�=~��9��&W_U���ݽ�ܸ���
BI��iȽ;����Y��wG~������f��"�_�V�+O]��W����	��'T*S[P��U[�"�z15@Q��8%��^W�}�hb#�=r��3UvP���%��-������A�;�D�߲{�-) �J���& �#c"���<u�llJ�3$����(�gt�׍�]7���U�Ǭ�ޛ��~ �����?zNKC��7���1`G##�C�M�4�#�L�(  8O}L�3MV9��=��{��X�|�����ž��c�
<�3˦*ߡ�*�Пd-L.��g��q2�`?���2OCj�(���%�L4��4�$*�^Q����j8s/mK|�4���%l�H,iq�d�hx������K�ѩ���G	Գ3ҡ�MLl@WB��1<�N�g���g<����D��Kq]1eb�u��[W����y*�<�H�z�@$�'N,K��"馿��+��hC�;�W���,��}\�E
�1e�WU�:O2N�l���X��ĉ�$_�G��Z����<�l�gw�tPa��`ٶQ{aqtt�E-��lՔ48�7��K�	�{��9L,����t$~�51�1�f_<��	�7C.�^N��R]��.�ko�!?�������x��(���� ������Gk��@,��:�Q�m0(�j�z�K�5]pÌ��o[N�&�K��I�HY�a4r{���#8��*j��w��ဆ��G���f�dhQ�C|x�si�~)w>���#H���Y]�`��ɳ��=#�?���?�"�֚�<��!ڐ\�3��!���1J"hC��}�>�;5(q����e��21���r�nh�y��G��5��:{Ffհ�-�|u��l�e��C���0�-��{Vi �9$���C�n(��=�k��W��"���̵�9��5��}�{���h�ҬA�-T��F��_ |���:<ؕdД͍��ʭ���,��u��v=�U"�xY�6��:ZD<*3s���R(V�ӥ{�I�5�FsW�^�	o_�k�\c�q��In<8��a����Z��58�~.����~�'��ݐNs_���q����&4g�.��ʊ�!�'������ll�,�Ȇ�����}�C�%TX�L�޿����D�|���N�&��T)���mm�ƣUi�s@�
Q���N�������CIZW�������};w��,�<a��ޓA[�۠#mM���Qf;�IO��=k��J5>�3��8��[t)��\;ĤxfR�#��L�g�
�+��@��@׭� �-��M�w�az�U0��:,0!'�]�¡\$ѸS���m����ۚ|�)�˼&o8{���w����J����5��hb���-[` �Ҥ�X/��Ҷb�ww����sv$Ϝ:�dxFv(��^\�9@1�\�z�^��:��<�RQZ��
sEY�$���32x�#w5H	�[XX��ʹ��^Ӎ���ȗP5���+�~�ە9����%��+/�\j�.j�5����_jj��{"U{�j�af����դw��%Y�)�jAj�J�*������|D��&��iJ:Z@1X���\h��I��$��NC}X�JΥ�&sR��j��<���Ä	���	Y:yJ�4�H��{�IxGh,x�k#����[an��7��.p�"�#�B�Q�y"b�3aB�H[�� �j};!�����.�\�/F���܂.�ƐJ���Ax���\1w�����A� �!���E�OgwfT��8wIb���M+z�����+�X�����Ȫ���r]� ��~��Y��`j� ��D��&�Y,${��իr��e� ��D���Y�̱q�)��h<c���<2	�yܑ���5��l�{�f��{k�[�$�?l-��;ۇ�huMj�"�l��.���7
]Uݯ E@���/����^D��2� ���÷��3Ez���F��Y��?�|�|M;Isv������ݛY_�РIA5��p�8<<�y@1��e���w�c��A� u�)�1�~BpK"H�j98��Xn�(���:�EV	�4�#�k=��WN��.W_{Y^x�[���3lS�:��ݓ`�,���/\��j�<x��nC>���oI��00��F�1U���U0�8@;��nh���jpnk�ᐲK���QE��x
3�p��:Gc��Y�A9	���8q��׋IC_������~�פ'����Ғ\�zM���w��_����D��Ňr�_ɗ���3���#C?��Y�&	��� �u����U]��^����3M���$� ���=�[L^j���/�95R�r��������JccM�r�θ>�(�O��������"yA��m��7�`G���C��YW����mY9{Z�sUҸ!��Y{$#T>�@�TlWȿ_�tI��+\̺� ���-���L�ݾ��v�35�g5 ��k�3 �ΐC��>�D�ܗ֎&�=���;sV�z�-�k��s������?р�!����$���������r�٧%.���AZ�y(���J���!I�7Gh��g������b�����ko��4t������?������LS�\��|q�39� ��g�1Y�i�y��Yy��䤮�O60����K�����ے~�kI���/� W�QB��E���Z[���My����p���<�����Re��&��;K�?�?�}]s���\�~U^���r�$?�t� �Z���&l;���q� X�C��\E�t.N8GP�`��
���9tFR�s���&��������7{e[$`�R��NGr��фfJ�c=IZ]YȊrR�_��\�D>�)�����i��d�CڭC���y��P�N�|�
���Pt����k����\����I����7���&�p��j����Py^?��u=_H��67%9ܓ�z�f*	7�f��B�"�4;���@�N<W��P�@�B��_�K��R��1���R��R2JT��W�l��2:Y`8�|M��ث���0�k���&]��~E�oI���y���3Ék�e[���/��P�M��^:#åyiJr��)����{�Ch����lX�u�)�1��Y�����M]�C���P�Ҥ � ��(�O�]��w�Yev�_�@�q���-l�PC�00|H���!����x	��c��/t��tNހ���loKK_�w���������i-�~�>Xq��%Nd�����	u�O���+q[�"Y6�5�5{0��DA �zم�V�ʜ&
a6�O��Xf�hB�!"���}+c̴�td�]�Yס��I��L�2�e]2n��� 6�j��U�G���+�g�/H����F"�p�|ҽE��	�Q,1��&��q�(��ў=�`�!a�$����� ��P-tia�XHS�|Fr:�ga�>9�9!ҠP����	A]j�������Ue��	��48��t�`&q��u1H�b�Y4U�t$A�[
��MR�5x�������?���|���`*��+��g��؈�p����ҍ��R�̵�}&�Yl�DC�� �!9�zB�ĝ�p ��t�H�����g�����I��u5@}i>^���&1�{��4���ș׾%�_8)�'�%�}$���CL}.�П����K�d҇�F��J$��@��1˂k�?�ϔ��F�3��}��McCI�`	.�5	�	�%�*%�ʜ`8y検<ZNh�t�\�|A.]�(�:f��2\{,����M�pV�@P:P���F�9��Y�<�Ac_T^N�,�w�|S^����F�v����4�ɗ7>��A��u���� ��s�qȻ���dW���κ�޺)�޺�C9�&/<���H~��gb�Z��'f䞾�L���X�>uI~���;����5���G�v����O�s��E�eV�'��_}M���±Bi�H����w~�	Ƕ��Ԗ��s�ʏ~�#� ��e��F�&!*�����j��}L��+W�?���W���ؓ���Ś<�{SV�� &;.��4��^Ѥ�B�AgY��{�ݔ۟|"��������[�ί�.E�����StK��o��7���!+�'O��k���FG�j�^��{_����~M�ɢ�ݧ4��sWN��k@�Z�}��)����rG؃N�%�S�+���^�4��b_^:sF�6��?���I��3�����'/|�e�:��@�ϲ:��+���s?�\�~M^z�[2��, P���2�gm���r�]=���^(�,�����gd��z�+��z�H6�-й(憀.��'����"��dIr�?�{��
��������Me�T����c�@!�a�a$�,��*�2����G�/n�? -#�����x�����RQ�_�"�.^���.$�=aQ8��N�4�"ADp�R���Җ�l���d�{(�G_�!��i�Ҥk�a����#��T1 <q&z��K-CE���eM`�r��o��sl R�aߍMAԸ�T��	'
�Q,���C�\=%�z-4Y_��s	;Cv)J��=G�T������=��B�v@��p�{꺞��4��}�y�=�g7`�����S��)�Y�$������H�Ȯ�R�K�^m6!�p8����%%�ӕ�>�D��S`��?K]-94q?t�l�7��m022	�= v��v �z���~�(�0&�D Y�)z�����`	���u&�cۭ���I�չ�����`RW���?�����I�T�R�N�2�r�p2:A�HG\4fN�&�N�IA�پw�,�':a��y��sp#b �>�e2�0����ׯ�^أ_�{�ə��V�#�f�cj��L�&O�)��"^�`lR���j8��E<�E�b�v����T�U8σ�!�BY09�0L�L�E+�,�C"��Ϊ]���&�1��a�d� k��d#p	@��: ,uQ��of
�y�����O��_����ޯ߻�����ƁO�h��E5�,�7Hy�D3(�K�p�	y�7�D��Љ�箅��
�+�x.%&�@� <flY�����;Ӡ(���,��(��� A� ۟~"����d����H��Ai�.g�yVN$�W.J�`[v�H��%u��Q��`��Kvt��cH���Qླ�v�U
E��J�0&/q�����	9{�,a/�*�2q�8qP�B��}ؖ���^kU�Ԅ���O[��ԩi@��Uy���+�=%��:�ɝ?�P��5���߻-�>�H��B�����k�z��Q�������l���X&��Dj�]�9���%�]�ԥ���pE�0�	Ac�5tk�^c��C.����g4`�����������~�Y��
ԍP�(D��&�R����T"U5��z%}TE1`�����L�3�RG������ xny	%)��%�T-��KR-�s����޳�K���5;LVd�d2[/30t�֙��n�Zc�#�"�����.h�W$~��6�_��%��s�eQ����9)#��vE��ųH�Θ��).E�t�x��A� +X/�Z[��ؕF�)D���-r��,�y];b�{{qiA*��"��t����J&��Ba��!قz.ß��"���u��G���W�0�u����d�\T-��E%�7r�	��~ւ�ߚ�w^�P�^l��ѳ>��tB�k.�l=�T�F������A<pf�Ea�L��ľ��7��v��N
���(1��1$(b"�ᩉ�\�= �Q���8cĔ'�(���p��a&�JU
���G��p^Nkb�=��t ��1��<q���`/�n�}H�yN��j~^��5��5�H� [�Y�z�t1�	2�D�FM�J��|lA�̋%=;z��>/-,0���~v;�� �f���'b���13[�}�"��	7�$Q[�C�� ţ�6�0�'<��a]��4���`��4��Z�?��?��ɐI8��Z��d���`���4@��P�K�Z�Gk����C1������ds��J�BV:�o�+�Nb����Ad�]=pF?D�z����4P ^I�5��	�l�Fb�a��tb
��,�m���h��k�q ?�	��9q��.�p���U��M_��t�����h�g�$)�I�q�c?4;=�K�-�O
<�'��_������ ����5�|�IΦ1ĥ�?t���`������.��,����:�W�����=v�/؅x�0W��m6-=R�N
���u*�+|?�S����P~���PP�n�Q8��E0v������>�z�G~���K����� <Q$B���9G��G8I�D��i������7I���w���̿������;�|gww/FƊ�"�t}�;�x����
��cL��*'����!:�d|F�sP)!�6`I������35�P����� �ٳ:�a(�/^�+�?à�����?�������eN�^.��%%i�w��o� ������|({[;�w���)����R��K��d�.�vA�U��9�(�8�b1/�O��KO]&�\ڀ&�ga���.�<�ek}K�����w��-�3�S�3P5]��+�����"���wd��)ѽ~K�ܾ)�>�L=�݇e{������<�+�_�d�����Y$c�Z�K�8m�4�k��s00N|�������D�}���:D1�H��+x��R����N�VԀR�>��zy��21��I!���`!C��XK�*G6�u,PG��m�����S��b������^{Q-���E�:�lS	�Ƭ�<�6tL
�Y�L�X๙����Uw(�Z��� s�����sF�-v5RM�*P��=��� M���5_	�tp �`3��l}��Å%E��ֽ���O��Ռ�GTU+�gh�3��R�
�E$�!X���G�o��V�)��]�얮u�`���U�Bѭ��vz���>W�lv΂�dS�"R���CЈ����;��{b�C��%@U�����B���c�]5q�:)���C�O��t`l �ƅ�pߠ*+z4!]72vql+�Ę��/������]��AGD�P�E�*;��`��
l?��~_���M�?���hC&Q��L[�<���Br�X��0y��>�|��	�<G���{�{�dͮ,����ȹ��׷ʧ�د����A!�g�AҰ�w��� )��o�yП깁FAW?��lKkw_F�j�;��މ���l�[B���v��?hJ{�Pr�%�פ��	FP�X\�IK��|ny�(�fGp�e¨�1[��������Z���?R{�%��q�b���*�Ģ�!Ԏ���IF 	B���c䉘�4��>�B7���Ͻkd17r�ɚ�L	`���ޣɲ4={���ڼi+3�Ww���`NR@0�Zh����Zh��В���R(�A	�B$A�I��f����fUzs�;N���9��"�6Ø�ۓ������<F�S�kb�ߗx��e�Ke1е`%�!�w���g�N͙�'�5��z�B�0�"���S�"ں�B�0�g�P�`�����R�"d��v�"p]ɯ��M;���d�GA���[�G�7��[�Ai�Qq��[��f��򊷻a���.ӢxB�3qn�c�K�����Q��Dt� ��s�����N
�kU%U�P����!$���i*�}E�\�����^m h�W>�;T��a�IQ�V�A�0W��|C��i�8V3��o|ĕ#��bmnۖ�$5�e�젉�R���<�M
~�?�ӿ�������?�G��O�����T�ڽ5�,mp���,[$<�ן�n�/�l��HG���QM
���Z&�4tqG�!n3EV�6)[�P�iR^�R:�>�K����K)�tS�Sg�~�%�����{,;�8x&_|�#��]�i�C�5�KZ���D>~u*�}�L�RN�dQB��+�<Ѐ	J��6$֍���L�/-�µ/�V(]�o����f0Զ�kk벷�N�5)X�X�C!&��2��_Bu �<] W�X����_�5��PX[���_��k?�U���k�Q'���',�g,��|.���$Ҁ����^{��z���2�{6�p�ך�X�P���Q6��	t�Q�ˀ��Es���4�C�A�*�l���]�m]�75���P��OH�
]�ҹ��y%����w��Z0�IG ��8$K����%���/���^%��f-oJ5�rJ�4���5)+����i�6���L���&�xz-O�c(�g粘j����S[2`D.{u~ƅ��@�ɗ.�89#�%�5屬*��L�@�D����)&#E�e���A���w�����FS�Q�L�t��0���$a6��t8�`�i0QU*��^��2�6�J]k=�"愁�FR9���b���Aʞ�M..�����]]��ё��/�
D���J�yM��r��(S>�ɏ�ۀq�l���!�jv{�ݰz�����9y�R׋\_�sBc����- �>���c�0�C�� ��ɷ��m8�V�H� �"Fj4#�4�{L9eg�4�kJ7� B�S����|�#�[��͍���@�,k�]͇u�޿���F�k����0l�;�}yp��ֻ&�H*�&r�İ��3�p�Lt�
�����z�W�d`�wt�̿�~��ZW��]"���΋�K� ��X��3� ||5e����$_c}M�R�����g:Gu� GUu���}��7]�g*���\�x�\��!�����Tbm�� ��� ��̃+u"������I!�
2>Bf��e�F,� ՟s�1,O�@�! ��{���vH��Ϡ�"�]d�E��)��ËSY���� g0烉\��M�g6�Xd�[��E�P�T($�����Q��"A���SP<C%�ݐ��<��ߐ��X��?���������tݱdv2\��`��;=	t]�{k^�GC�X�#Q��Ǽ�M�$^ܷ��!�X�b�xf0f����
Sx�M���1��1�B���L6i��
W��*��8�������I��mM�r�S�'�ɱ�\�K��s |�����lP?�8�n�Rh@��D�͵J���]gV�ss.r�3p	a���6T�W�ѲD�7U5��U�E��Ҋa����UNI���u�c޼'�8IԼ(�\P�Į�ە�#?'4�Z�I��9�s�RN�8�9o�?�d+c�i���+�&����o�m�� @�����w���������nB\H(F$*̣q<�a�+������L7A�T;*b	�ah^NC�K,� Ѳ}��!�
 ����G>�����|^�G$T��ic*w�o��ֽ]I:M'���i|^U{�f�\-3������S#���Nm �~���� �NAV����վ���e���F�yF�
��d�6�~���dkgO�7w��=کg��[�A�T㧙a�/c�<�a��ʈ�|��4HR��m�mtI�n�˭�����c��s�z2<8��ɩ�ޜI6-ֵ����\0]P)�(��`"��˹X嬨s�aՓ�P��J�hW��`�Z��y�Ҡ�KH�#T�JWm�z�l<���G�FhA�.r��og����I6�˕�+M:@T�qƴ��j7߂�9�-�t�t�vp��g�A�$���pa�X==??��>�{ӥDǸG�]�2d˺���Td&`{�y�$��dE�hP8�c�au���]U�eB��F�l	�ؐ2��<����T�p|�Uj���R���P.0��G7s��i��ҲP���=��@�����F�1�䤨Zͩ�;8�x����ǯ�1����2��0d�!���a	�jfu_GԬj���a�
�/H��G௮d��$�����s��8-9W�,��(�$�P�X�������ǳJ~�"a��*6i� P�~]���{�$���@��*T���!t�!�����'L�='݈N���VK6ַ��� N�(j��G?��f�Wz�[�;��gY�R�0Xd�.��

�G��'\>��ZK�`8c�꘹���Wz�����|�2�]��`��iR�c2#��IGs��A��P�:9�ْ���У
s_���KFq�|��+��J�'���ڱ��\G�Q�*/�𴀭l@� ��P�%�!��,g������]I��#�N���P	��J�a����k$�}ɑ̠��s
�yqb$P&�c{���:��V��VF$��ER�����U!*��Z��f>�)R����Wxf�U�T,��<�*z�K纰t�7}��ۛ�/���\�N�e6��a�SB��:�9~(���[XB����6���ׁ��7�)(�A������CE\�m�����sa��&�VL!����9����6�9�sv�71 �1w]���_��BH5�\R�{�=X��?�z��,�.x!o{4TR�Un�1��E���T�Lv�:�o]��96�X�d��_�\J�������>�b����ƶ\�bj��A)I#g�Y�՚%)�O�S3��fX�o튍��KzuL���N�]d?/v�6)�%}����������ų�����ژ3��4+�m~-�yC��%�J��1�YՁ_`-lhHr8@t&��,8G\����6[&=�Ao9�i{�]�+̚W�$�\����Pz{}y�1�M~W^����Ԥ+[�۲�����}�������	N�+:.�BT��@���!��+&'6Hd����i0K�F���D@�)[���wؖC��Җ��#����(ۈ@�?�X>9w�w](1-'��է�J��	1��^�:�?����������*��3���O��D�߼���+��|Y,��4�("������sQ�Ѝ0�[��'�vS�XW&�p�t~�
��+H�lcϧS�>�lY��kӁ�0m���]�P9�b��������5p��+$���P�-M.��M�f㑜�X�,$�*�z��ts�&�པ�>�L�O_,����a�@��Ҡv�P��NǼ/���e���h�����6_���<�� y�wr�6�
���R8����R_ș&ox1�8,�����X}G����<>|-�^R��j�I�m8�y��-�}�p��݀�-�'���6*pX(�؞Χ��7��Si6YF�|���P�q���Y���&��%��`-��ƺ�y��ǽEEtxr���B��h��:8Q4 +��9z�Z��|�=V���{�j�Kԯ|7�|�x����<��p!�+�4T�a�G7�ܺP�s'�7�&�ј����.���c�fZT��a��7�U��jQ_A�*��ۏW֙������ؽ��jC.t<��+�s��3���ð�4�m���L�(i�M�ºN����%������E�b��4��O�^tW��"Y��K��+?vtcs�a��h`PI[�C���]ۥ�u\�FT28��g�wD������|��Խ���$�17[ ��E���^_�8�e�N��d���!���Tz�da�M|S{Yi�n��z���qV2Q�Bǃ�Σ��U��G��83CK3W̘ه��<6��f ��[�.�E@y�L:�A,2 /�:�6����F�a;O��4(d�/d�Z�Á}����-�N5�J�pc�gcYk̀>�*��SHQ����-R�U���yR�Ţo�UbQ�wB�`�� �z�7��
jc<`�v�5��i�sr����U�ﳳ���Z��|3	�c�����7���p~#՞nFi� �ޯϩ����Gi~u�0�����#�H�
���1{^]�x���T���?���X��]�r'�T�M�d��+XE։�M}�w]΋��'^g�J�,����7�ﯱ��y|���>N������#3	ۭh��/n��������@De����og�r�>D����4�7-��\������i��vif��j*ǯ��hd|�9'D.���C���cy��}پ}G~�w���\�����'�K9���.�~����?�%xg_�?�'���Df�^J1^��R��ł�� U��}�WkxW_��Lƫ�˜6 �ѝ6I�N�����C����צa2}$�>�����>������?�{��ӿ�G�ˣw���{�]�vWD"�/��ߑ��+���B�|�C9��K����F��Bk�삘�L�%��,� �2��,Α��T�(�8���	+� 6NFVy�_Oc�j�t�C(�\tEHHčJ�ۏ*Ǻ$�j���j"ã#����TtLp��8��C�ӟ�|]P��H7z�?*������ ��p��?䫡\�S�_��%9-��1��B�n���z��������RM͕�DPE�)5�#�V�_\�kl�F2�9f_.���Kb>1�/O��駟�ӧ_�p2d���H
./2�B��_ȓ'�����5`�	��UYi��&���=�g��T�`J��g�4� ���'��O>���&�`"T�CS��f�9%���L�� ��t�.�:�A�C�����޿y�L^�xAؒ�mXV��ɈL^�{��W��>w4aA�3
]���X��\a٬�ruI�FrWUV�H؋PM�������i��j�X�1m*)eĕC"_=JW���Ǎ�:�T��R��E��1��CI����m��'za@U18�Br�I��K8vg���wT�+c'�L�/��
YG@ �m�?�h����MBq]$O���k<s�nir��ܠ٘��j��d"Y:O#�5��2�j��Y�`��z��!ۭ����o��tM� �6$��K����1!��R�nue�ۖ�����0$����A�aSjc�3K�̦�̒�4�5%��ʔ�Ѝ�/��][���}L��.y���΃N�$tA׽Q��(s�h��Z��ݩݔ�8���p�$�c��k�9��R�d�{�O��'�ɩ���[�+~�C�Z�ukK׆���<�$d*ggg�D�QG��@����C���['���Ua����7����랟�q|�s�:Qy��oA_
'p>U�qIEݶC�ks�{��Y�lmC��{z7
��8.xe��dN�������^Vz�`F�E��^�7��y@�M�y��g��&e�Eŵz�)1:BhƔdU���S.c��I����G��nSQٍ|��86KdM~%��)v�� U1�#�[��:9����E�Փ��~�y�S�9�o��_�G:_����v��=K��GF4��u��B�>��B=��A����z�U<T�3�q���a2!م���)̲��6�e�`�:[������g{�o�i`��?�s���>�ǿ�벩�7ci���K�w3�h���G�����#i�Z���-y}�F�.�����AP�X@Ǟ���a�O��n,���z1@0���NX0�>h8��������F$k�����5J��o�H�\JK���2��g�ş�%}����>�����-���"�������|�]��!'��{�G����ɿ�KYM�$�B��6����"��ru�s'+�u6yu��7�@'(^�K�jx� �zvt���nV��75Yz��K9|�8��f��_�"=bu�K�/���y�L��1�-i-6��yh��r1��չ<}�!D4s�|^3,~P4f�PK9;~.�����^X��m$E	ݗ������`<Ҥ`$#��i����K�[T������s o"��Imk�'/��g�|������|ᘻX-dp5b������W���P��W�;�=��x=Nu�G����h���?aqtzL~7T�ѩ�s0����t���R>��'r��-s��D҅d�X�u5�	�&r�����?�����b�A��rS�qL��(-z~qJ�<�-zzo�����Grl4i[�1�������$΃�y��4 ����H�z�1�N�d��[ǳͪ�׀DZ�FY����E�u���t��9u�K�����{�?H���up�
�@��[���Jbǆ���5!��u�.I#����d��.׶7���!w�>�	�ՙ/ܣ�Tp�J8������nd�?r�M�3k��������fC��L����I��|���4�c@�Զ$z��SMV�n���l렋t\�	�y�X!�9�d�	RnB��`,���z���<�{�Aw�q��AoH�F2 �Z�p��O�y�$�F`�`B���@�����%�u�(W��c��̩8~V�)EYJG�˕��|�9f���+�4��᱑1!����(�u��$����Ѐu������|#<P�Gv�qC(��y�d8����E2��3��#��C-n��b:�����:�E=�olɃ����Ǝ�onS1���������f�|���7��;`�H��be�Pr�
��Fd-k�@KprSk�ڝ�ΊvN�ӻ��W����Me"<n&�z�װ#�[Ϸ$�:%��H�u�4t7��B1>
�{�,�q�}�\:n�!���s�h��:AG7��bn�Yq��yo%Q�/���r�_��M�����uEj���.>p�+�3~����a��$6Q��Abq������R�R�H�p�	#������-���`���n�e��D��ڍ�ӿ.v�6)�%|�埆���?�?W2�F���Vm��j�U��ZU�}�}M��T��ި*��9�"�3��,�'^ܤ�@�B��0M-����,���v����<��H�|��N����11�e9g��/�R�3ѨVù��a�C+A���Z �;���{��TU��3�@�sJ `�g��xv�0��X|V.3nRy`�9)��.fS�糉S/�xa�ѣ2VR�	��Q�:�b�kP5� �/����~�|��g�۽%�֚|��~]>����
�ֽ}�� ��mS��PCO�����I�0�ZjaxX� 	@"�����s�����s������W$�&��C�o�
�&pO�K�e(�tJ=��Ϟ��j@8�D������Hз_h@y*_~%O~�9a&l���i! �3���Jf��28z�A�O�����$:��P_��;���Yq!�5p��O��K8��b��F7�%�5�E�kr2^�=�437bY�c���P�>�-���~@����q��^��=}k�bs��;��Lƃ�&ϩ�as�͵;�[�#��h�Uʥ&�_��3=?�0	#{J�k\�&.���P����_;��k�Hn���]L&:�.���Ħ�1����5�*�G���89=��>7�k:G�u2��� �gz����Ȫ�AX�_����{�h���Q � ���G�u��6�x�0 cG<����# ,���ɀ"�̫�Ζ�Jm�9dRA�3��Ü�K[�t��)k�� \3�g&J��ؽD�^�ղ�H���/�y�>��7�9v����I,{w��;� #$���2դ����Z�/��5%�2��_���[����8\hb�&���|Q2����+�
��o��\l5�kln�J]s(�$�^��f�%�&��Ր�_3��M�*߻V�!�*��O��x_cH;����G���z. ="�u1���,Oބ�+�1��H�!/,y��������#$a NIN�Nذ�)!�H�B�dc>5%it)��n��׀izx)o�WF�]+=��Ɔll��_�}��L����d"�7|7��s���Uz�s�q��d	� �!J�3�T�7F�-�����v6�L��v�d��-���4�[sk�����J��?s5BgD�I��2�b�PP����+�K�դ����<%�b�A�X�v����|3c��F��w�oT�o&AYyn�fv|51�����I���%�u(�����I���P\�)�:�������#������9�I��L�E���SB�1�������9��@�y�+��Vu=�P,:�3<���|��b�ߐ`똅X�Q�4�NX��9(�8z��c�pw©c�VX-��Nv��w�бYG�W~��^��w�{g��<�M
~	�^mvuP��A1��w� a`%�RV)�T1��a�&��S����7��U�,N�(�jQ�fKB0૎��L��J�߰�Pj�?��Gtr�`L�M�B�?u��3:��g�O�8=��^G��3)޼�n��Q����������r����'rzu"1��O���ܨ�$�p����n{)G֡Da�&he�"u����dtEhH��6�Ɠ�%��gG�f#(�$�Sl���!�)4�)gfR�M}��饲:������.��zG/��ٓ�FoM��/\�[ d�t��6yo#�1��� �}rch�B�����8��`6X���� �� Tj����n���]��r��b��ό�8�f$�!V>��rDf`��I�&w|9�R7�،���X�k��^[�U:�h5��ׅ\�������D�F�?��4�
���;��4��L|PQ�5�����=����T�כ�_:L����������QҲ�KgMF'G�EQ��az��~> ��ݣ%�::��c�Cr���HE�㝶�{p_�m�	��ˉua
�E��Ӓݨ���r��ӯ��>�`�%Ԍ
Ýs����Y����Ç���͒H���Υ�'4�]�{�%���˽G�4��q�\�7	$[�`H78M��o�Ȼ�=���6�}_�apx,Ͽ��%ρ�z�0���ݥ*`u�dz�^��;����	�oW�}��"3���P�>�XCJ �ZdpHG!0����gd�$�S��X��do���<x�N�����-tU�İ��q��B*>�m ����1�c~�&�f[�<<7�I�ml�e���šL��4�fj8f^�2��Ry�̸6�t�� s���a�'���R�sMV(=��Y�ZW��A0�;=�l/_I��`.���)�UM%Q4���Q�)��7gg�a�/	$��9��/P�z���XҼ��TX0;~u S]��|�Z[�{�����A{S&����T�М��\�j�-��G����:��:���t�����2��䥎WH���4��%�u��k�:�1�ڦ99.0JyU(���i�c��Jy���2v��)�	���zEP�X���LI[��:�!�c�NCǅ�A�}i��X�Y�9�H5]����$"����y�%}z(�A�xi>R��q��)��_�tr����XGG]����!2�WQ���U�J �
2\{<��r�-ov�8��F��5+?�R�M툪i��$��~�>7 �!�H���٥c�{5�oX�ߑ�����ǝt
�y�:���t���q=M�0(�����]��<�	!F9w��:tk�r��W�N�vϒ$~l8CXKJ<x�����2$
���>L��S����[��TO�ga���V�O����7��M
~	��I7]��t�����؀� �.��N�k���5���۟����*&�\q����l�M�9w�3�����h*�ݍ����4	G�ߛ<�t�ȇ��%t�C���t��@V<��xs =�Hv��]�dF` $��\�z!����r!�鐲�	�@n��,*M7b����F�f�����e1����@��V�g�b�� � r\t������R�������f��O���rW �=Ś� ��zula�BWd$O��r��g����_Er��I�lB�=ɗ9�`�4��v{F�L�w������]���پ���B�#��JW�ȥ�����xpE����u��Њ�}��%j������f�&����{�?�N���[�C���g�4@��X�*�8Ⱦ6u�l����;��ݑ��J2�@W�⡗ء�>AW7ם[rG��4)�5���L�|���ݦ�G���Q���{�#w!�k98=���O,�E.��)��x�{�} -��>鵜\���-����Y�X�]�=~W�ˆ��C��&�:ΠS��	�.�%J�٠�X\ n3�k��hŁ����Dȷ��a�ly��ɊA��td"!��դ��G�>��D���Ʀ��>`'c�#T��5!��P���e��as�[�ۄ�!�E���k0��s��jr��*V>|5�]Kx ��n���?���1#@�Ak������h��X"�Q�[b�&����1]B��9�z���A$� ����}v��I4"�m��UORs�*���
�m�6G�}b�foj
+��;)C24G�pځc#/���S�n�%��7L� k���7_꺶I%�����|1 ���K�3�Z�.*�~;/�;1� b>�K�rL��h2���~Dצ�IA���3����JP�*`�4l�P��4[�Ĺ��l�WH҈gUk}.xH�[3��z�E9Ŝ���zx�.��oN���T��B����@<�ڔ���d:&"(s-ڄ�B	E�`�l�Y G�
ET�Ѥ$2N��V���fW�
�������s\�T�1�|��I�ח�~v<�q�Dg�7��+\9�r�D;��G"sK�0��Ypt ����n����r,�ZSB��Pk�44�!_����NQ&ruq�"Ӛ(X(
�
��r�Ǳ08J`�0$x���VqwP��\�"���C�9�z��tN�?�&c�#���������1P:�\��IA�:@`~y�KYc�K�_��!臺�R!=�"Ϋп��p�t)/�$�9�v���"y��ãȵ^w����6T,J�T��ρ�s�I����Z�l�̔V���~X'�gX���I� Q���Yh���1�&��N��.�¼�l+���@���a�<������S�^�)�����e%z�-ߋZz.��i
�+H��?�c����eQ�w����{����I�/�cR.{y^t)wg�uJd�	�84~G�#�>ڑ���J�(�QLA�&*I%]&�u�bS�ڦO0������]u�Y�ʣ_���n�M]|W$��ɨ����l�`ʊ�T��yF��ߔu����2Ǧ��4oh���W���7R�Ҡ�R�F[`@�K��؈8̞];���=᪊ss�A,��Xj`�J70�L�/0�H��C���%��+���a�������1�� |���
[����1�{)G6+=�ɫS槢O'�������ۭ�H�L�V��/�р�
o&-݌��ݓ{�$�F��IC��nIS�^�X��<�
H�������v�� 5��Ѥ���VuSߣ�����H7¾l�ܖ��ޕP��d3ѝX����\�eq(-��q�S޴�ߒ[{w�[��ߓt�ȣw3��������¿s������Jc}͂�t*���$bn�6y]@�k��_�Ҡ��lhp���j�,RV�n�{`���P�zO�oscWBMj<�3M������k����M��D��;｣�r[��m�]��o��Ј	�_/i�B7@�Xܾ�H���t4��Μ��3z�
'�P���~/��P���-��ە����n����Cg��X9N 5ܒMM�>~O��_�<����֎4��-��z��MHt}������Ksm�$̳v�	��1i����Y[۔Fg]�K���g[��S[:��ʑt���������A�(�F	t����)	�'��W(8Kh�)0-��	��"��U�5,� �E~a��T�)V�WUJ̓�֙<�]��xR!yU:Q��fE�1�\fn��V&h�l��[p�n�a8.P;x�d�����90����t�57��#AO���� Q����3<�\+���u��Z�����-&֙���)�s�!m�r	h# ;2��:gr�X���)�-?ffT��s��77t��#y)�n��gt2AzzX q�uLhͱ0�׍�}'nl�N�p�k2k@�����-C~W���pg�z����lR�:�U�u]��A,=BF�~�̺�u梭�J�+=s(�!`�B�&hg:��e�nʵ��c6ڄc$P���D�#6?*�2�%��1�8�]�9bJ�#tZ4ʂ���p(��
M��e�c���+�ں�}t6L�ap��݊��TuT�{:wM�?b�8l1��R�+t>`���5��'I���Vlθ�#�B��g>���͑�_龒�sR�<iн�R0�8s�C�^�'B��*(.�@��07���X-�"S�x����ͻ�u*������'RIh	b�F g����)�ˮ�	�t� Dh�n��K��]y�{�3�'Q��t��Ӱ��cx�,�՘#09`kP�0
�����8�Һ�t�\���Y�_���7t˙�6�p$���� Etg�+�z-�Ź$����B�� �k���m����ۯdc��vwv�^ks�%�"�s�'�K�e�,[0$б?�3_��p���K_�b}Z�%�Js�f��q�����Ə�&�d��<�����ŭf3�t{�`�+.�e`@W6�l��J۴w�"�z�S#�����`��D�8�H�m$f�LQ�):$��&�J��B�ʚ_�1��7�JW��`�dR]�F ��l�^�4�y&�ـ-�R'��;�Ȇ.Zg����ⱒ��L�s�BG�4b�g�542Vm�RU6 %񝖸aX�!QZ�;w����aK��	+�)�W"6�����9�|��}�LMjO?�[�f",F�WWb 3�]�g�#6�܈M!1��%��]G&bmTTS�;t��T�/�3¢!�G�IM�5��oH�n��M�a�9#��w�r�k��`�.�	�^9,���Bt�*)���h���7i򆖱��\������-���m�޾E 6*�������a65��h��� �k��Ze9B����"N�r3��ܻ�@��nM�2=���)$�.� �ba0����L�*И7PV�#=ބ�a�8s�J7D�8�}Z�:����`T��p�$�e$M�����8�Ibrkw�	 6��x���{� �������>%Q!d�s2H����M�>���;�S�m����
 �a���l�mH_�(�Y:�Iy�3CR@�l�:z�:�:��Sm*X���|C��o"X<��a\���!��L����)%\�����m��PTw5+��el�_a+_�n�T��Ҝ����<ϩ����=J����zX� H `.�����3L�=C���	����;.7� �P2)�	��	S���֥��Uf â	�Z=ھ&Ͻ�u*� ~.O���4��p�������7Z��Z�%���{�{��ϼ\Mg�(��W+ѱ�s3��/��Ǝ΅���D�%�^����Z�����z�4�F(g�" )�掛�J-��T��Ω����I7���x@�!,"��
�;c�UBu-�+5�Thtgx�&���B\B�*>�^�f'ѽȗ�έ��\i�7O8�VS��{��豴um+5�(p���cY���]�+s�+�XS#g�I��0?r!����W�C;�G�7u��������=�_���BF��^��Ab��j3��oz po�!``��Rծ[��R�%�;�����L�Ng�h�%%�C�5/2K
X���ɘ�5��#}�"E��B���مΉ��ܧg�o���rޚ��ҽu��}�Հ��{:9X#,�.��UJ>��ìL)1pk�#KG�� 1��¥{%�i�{���z���? �#3|GPlK�]M�tϊuMG���\�'Oe�䩬F�:Eueh������G�{��[�?�m���{�����ߟ�/��mR�x����˯�NN��=�Y�WZ��`�	#���.��7�����|d��}utt������{�ְ�@���� ��AT�b�'>7Y�V-@"Zq0)�J��UѨ?L�!�lρ׆v�M94�0��M��,9@��!u��46��'��2O%L�0PW��5�����@�X=��T򫁄�请���$���#���+������_~,O^=����̳���u!���&1�z�@��A9�'L�N��W�T@��LT('��YN)�g�yMFL!2_�0^�$Ǻ}��A���NP��#,Py���'/�!k�+.Ft�kI�[<Kڸ�2�	�F�d>��5��E�v��1*�$�3)3WH�d��Nq�t1��`��H�ݲ���ǆ/]T��ӅS��9ݾ��=	*ȅ�.M�U7m�8���`hg��l�sP�0��<��,��um1��;���2$�N�6`��ϙ�ߠcc{g����$6v�Jvf��x�Z�?ߺ�-���w�	F�4�_�`z$)H쮆cٽ����6�\�"Q��J��$h\���k���������x��i����΢�|L���qhR�l2�oj�>��&���ZR�O�4Hy]������eF2��m��L@�\��!��a�������.I���|S&��Q=���}�����+�lX��� ��X��=�9-?l�G�'�$� ��
	� ��g���n^8�u���5��
�f�\���,����z]��/5����w�^�K�9W�cM����4q[�utDg�N3�n3$���W��"�~h�shk���0Hgkg�9M��:&�AՂ׵t�*$��k� �Kh��F���+Y͖��u���#�]{�� 8����s	w��!1�	�M-Q�AB�j0`,��E����w�P�ʸ����!���=��[�k�1�,5���(�~�y�ò�-K�jS�*�q�I	UD]r��f��'A��~��Z2��ڈ�m��D��X\�?w]���8[7�k�Gb4$gO'c9\�H_?��lYCW�%�G:����&���Ģq����撶������w��p���������驼9:�C�3��s�{o�����t)�٥�ݿ.G�'�m �9g!.�y4����c�-� qE'�0"��y�h&&!�&R�1W���{�37���0bg0h"Aׄ�"3�=%������b�H݇!S}��G�Zmy4�m�$M�`Ը\ѩ{\���0	`zp��0��:�1��ݙ�	�\��)����W7Q*��񒒦w���Y�lib���fܒf��K��,�4��(~:fbY�&rrv��E�*�I����<�'%��|�I�z��J�����4���y\o�b}�������������Kw<IY"�n�0*��������}�˱��*�W�b�-}��<�����2��|.��e:���G
h/](5���H���5x�ו/�Bg��-�f�������,�H�H:�Ա�;1��R_Y�V�>';e|]�i^t�4�e��ʕ�}}v��u������w����۷�K�̸aWzӢ�j�x<����>ԠuI��U��@�]$A�{��UƉ��o�xݸ߸���l�M'��	����T
]0�E΀X��x%������ߐ���_�?��!�X�M"�G�z����f���bsK:�ޥ߽�C	��\M����L�@>���T��EUm.�����q魰XRA�X�"���B&CS]�5â��,�Ɋ��JB��P���t&Lh#c��sEР�xP��H�e5�鲞m�xT���^�g_sD\u�Q�*"1�]�"�9%��
	�������"@9	�p�n�\4��>f�]D���B�Odww��x�ƺ����xu��A����k1P^�
Y�UzT��z��zPT9�%�2������r6
W�^G�5����s(��T/Z�&96��6ci�{$�ƀ��G�NN��o�
TV�ƈ�B�j�$;Ǜ�۪��� +��<4��Fv�,C��mF��=�J3*r�k������.Jh��$�; �(b�` 9�����9J���{���ni0���r���H�s�
�<�ljn�S#�A��3'!Ԃ7
@"��XX^Z�P��P!"�
�f��t��G\a����d����,p��uU�O\��
��\���#0��j���HuT���]4��z�k�����u�.��O	���x&��;f��X,�.cq���6�)}�L�G!��^S�R�En��P'
P�Gd晩Q�����t�I�ip�����'T��#;..�D�r���L���Q�jE@�����3���
 ����<�u�m,���@������{O����M5�˃���w�5o��N#���S�
���TmBh�p0�����X\������D9;G�������X��B�Z`T\v���w�*~MfS9׵�|2���S]����c�?��L��tOk��{k��յ$����+$9�[�um����ʣ�נt%��2ֹ�����x>#�Gv]�6w�������]�>��/O_���,�r8�vVTC���9p�J]2�C�I�<%l�&b�n��ݕSX��X� (*z���`�5-,ٷ��4wg�[�^.�OY�,4�6��Z��w��+��?-Y�o��֮��]B'���o��{/�X,Y���'��FQ�r�H>bd
�I�B]0�~��_-�'�N��p.K�������c�4e�5��c��dy�r%�E��lԊ����?�ڤ@oP<���yЍ4�Jo[W���7/��>��,Z�1`��Q����^Zp.9Ɉ���t�
2^&��J7�zZL�jyYXUs��zY�����p�,M��!r�@�h��Igh}���Y9�3�;�R�@7�2Пu�Ƀh��&�F��A뛁�Ć��������������A�q)���p�mЄ�KPM�r/(��%�0t���ӟ�R���F���������|�x�����-Y����@�Ј*��c�ܥTA����������E�**O�b�?LL�V��h �鄸w|��C���$2eܘ�aO'3��s.�2�l|�[�W,~���"w3�V,��6CKMe� M�<MT�ts�©�h�"zC��ߝ-������?�w6�d�ߤ�����t�wEg,����)�wo�§T����/M8ٱ�5xSv-pF�+`�Z���%�b]8� � ���Z��L�^�k�P�	�0��Ď � �n�X�6 2!̫2�`C��t�R�r�}C�,�
y��R��\�|�_y\��Q�b�O�\ JU`����QP�L���M��#�5�o��C���*�6:��i�;�!���;$ؙ?��!���Xk:�y|T9A�I7h3<�`��g��I�M�ٚ-4�XPm�A��0���B�@vkk�ݫK���0�H���A�~��7����z�F�1�����+A���@������TU���ǃ*k�*��7S�z%47���r$����>e�J�f��8o*� ���hB�ګ��A�sE���k7B����8�4�sG������ƺ�b�Nä��H���딸��H���#G�r�OU2�İJ=`~|�s��!.�3���`!H�K���	� ����5K��n?q�Ǿ�&��י�3Y
�D�6�+�k��:�4B!�CCI���>"�4��&˧t�Y�(`%?㸋��0ӫ`f�Rb�͝�y���JV��TD[nױ���5M�Ei�m�|�P�@�<����Z����t���z��!t�u @�Y��u!�[�88iI�Ǉo�\�
@h��UxM
$ �aY�zl���d���M�eM��.��*S�^�*�f�e9��������<�0V�fY0�+t�J?�����ZB��1�r�����u?�;f�x?e����r��m�� �`������)�t$�7�����Oa�TP��`vUPJq�Rt�έ+���S�+Zz�A$��Z�HN�����9@7� ���&�>a�;�V>x籬on�y��-�RF?�\fӥt=H�z��&��8	�@���R��n��	�
r�@�.3�C�-���c��-1���J�ԑCs���y[%�b	�F��	�3!�O�9Ѥ(�+������my��}��C�'-���|���n�R)M�R��5�ĭ�����/�3��%\�7���=�v���VH�v��15�	
סl8^D��@4��t4�H�z���Ju�^��H��"qm�_��L
�H��8z�����K��W��m��z�::����6�bD�~#򩽬ax�^尖#�7��|�{�pi��G�@ � �f����Q�K�[;��{�͞��7��yEU٫1;o![�������U�l���Qp�=9el��TF���b�J�
J���6%ˌ܄��70�%�����4R
k���V���n!�L�!0�Js�l7́Kڴ��$`�*-���d��h��
�aQ9G"ptt�ԩ�����I��v����-޺�UW��U%T���B��z�b5g������l1�Wo^ʳ�Od���MP(��|t)W/_��#�ޮ$z}�z=b������L�Ϥ�Fv�������B'~B�����w�C��0ӱ%��)	`���u�2��`��:��;	Bs7K�¥I4�
7^Bb��@��N/�Tb�$^9"K� 	��0np��ߞ�����g�9(�
Q�Bd[�Ďz��%�����t`�C���T7V	�ʺ��~��[���d\�Vٻ���D�Z�H��~h�c�kA�P�JL-ٍ�M]T=�ۺ�$��u�K/�{�H��/�	�+&�_����o�at,���%�d����͎Oh8z<���ޑba�l��]H�x�E�i�Xҕ��7s~�A�2W6�q�������b(3�
�Qљ ��4�)}E2W������;w]s6��5L�%����]n�/@}��q�H����:-w-}�/����kO�tn��߆�/H�7]�y��w�<X����/�j�O,9;!\�#&�6�JY�i���@��0�^��p�4�*�+��C�e�=�T��:�HH|�A���5��7 >��.F�G���T�J	5��r2�"��X�� 	���|�������Q����$m\�8�t��'Ì/
��`���\��G�Pڛ۲_'�4�+��X`���;[��[\�f��ȘP+�st%��:����t�n����T� �Y��]�4� a�1U��%�(��	3C⻪1�u;�6ֲ�0w{,a��K1�3k2�.т��!:�1�S�m(t��4�C���c��ܥ���d �T�~�c�E0@� �����ӡ�����ޑ��we����}�10!��zP&�p��>�P�U�����$HyO
#}�FCv+�!����b���t�"X�D��ߔ�����+$l�7w�7=��&J[��6uΥ��4yjU%��EΝ=w���+4�j��&�	��5F\��5�-�
�4x��:w��r"���5<�|�a�\w����2͌#���6���$�N9���7�y�6���)E4ڑ5�4*�L�5<k1��l�bIE�ΜIk����z!)�G�4�Me<Z�����D�_��2%G�R�td�/��;��9Nt.��� :ׄ���U����E���+�����׋t���F�{�r�����J��t��\���Êڰ���G��E�* ��ݻ�ʺ	A�f`3?0�ґ�\�U^��(��Ъ��ͤ�b�߫���U�*��A(Gw��������}�_����� ���. uVw_��b�gUׂ+����j,]��#c@#1������K�Yp7tr ҃�P����Q��dK/�BY!��0�[V��f+�A3.lؓ�1��|>��0�X-�"��r��$��j{�Ee�}��]�i=�+�Aض�8ք�_rK�!-C9>x*��G>��?�I�Jnz�"�r��5�\�Ɲ���o�����0�������D���x:�A���*�1*��,���p�ْ$��Vl.�ؔ`��i5�^�Di�`S���VC�����1�8�ά��m���_&�`6�Qr�|R4��$z^�U ��Ce����yn��*.����զn�9&b���N0|�B��&�L�Y�u��ۜ�26��H���ۑ��ڴ���y��*e�Q%/x�@$�[�6��� q��dssS�{�2�.�W��Y8��}��ʓh���K$n�ǫϙ��s��t:&�eC7�F��5Jv��Z�,���tl������ǜ�kW�P4� ƪ�����cM
���h�w�e{��u� J��H̠ԑ`B��uhl�߾������]�=�E켃��I&f��f�*H︦I;`bg���cU�R#����&�?��}��^29��9[u�Lg#��KS�q�X0�x�5p5��w�}qAD�[ ��Z;�4��2�X�܄����:��#``��m���EU1�+\���P�d.�]���3�G51���'\�*yfy�0�	�B��UJ,%�`��B��L����^W��/����=K|Vy�\q�B���q 9WB��g�����ȒnV���O]�`� ;���l�%�D�o%����G�o?���MP�
u}]H4������0��Ԃn����9�.����^���ȫO�����,�C~��ǒ��I=�TU��{�5��ݒ������>0��{�v_�����/���ES"l���\i�g�L�P�e��N
T� (`������2�^�h�?@��.ᇀ��P�c���I�O���0�vL7�(�`⎪/dbQ�ñn޿+w������������v�E��d�{�:�q��2si��g斥u�@��;;�(A5y��K��ݾCo���&9,S�KiA2jX	T��e4
��\���,fL�����
E�cY�i��f[�E*vJ]2���J޳tp\�Wr�w�p(��E踇�{-Xr�1�f�`�9	��9RzL�Wa�=[�' ��NnR���&+�4$�5��4���q�]�#�ۋ�A����fx%;�̼9C����������T�[�q�s)�L�SFc���4��0���i���ڤ�,'����?�?�@h��`�����X��Oƀ*���;\Y5y<b%�[���NQ�t�}�D W��q�����]Avb��-�h�P��3\�9SY�/|AL�=�lS�]5�2�`h^Tm4Ørs�D�#��e�Ë�D!曆7{HMe�<����X�m�)�܅�6	���;_�6eX��`bb��wȴ�x=
������E7l8�z��|�<�XD�W��9t��)]�i?~���z^�9��@VWx���y���:A�^w�K�����}���I�`J�m�k������L.~r"��;���n�������7�Ś�_�j8���}�?�}a�{ъF8ȋ:x�?�3��EUq4�-"d���7dR�bh��b��ޣī�_7����N�)k�1�I�%��h:�wԙ��#� �έDw�`и�NǙK
⮾��q9ts�wA1�PY�M�fm�q�^�0EO�Gp��6e�Ȩ*�L[}��U��h�0|6�Ȩ�L.R���7���ʨ�Y��,��x*�6T�UI�z0#�޳V�aQ-V���a�������-�[�<_�Q�^+�5*0���:��8:z�C�L�Х�Jz�	\��_�_��Om#�`����g[ۚH�2{H2�:6C�Ļj��k���;8Ht��D���2#���������@1��K�����O�o �J�@:���#�c,Ṅ?T�J蘝N�t`�����i�p�^��!?%�|2��\�%q~��^���9x.p�5���nC��FQƫ#�ja4mu��W֚��V��}�&�R1
c 
8%9-�J��^��� �YXq'7���:��ֺ2�U���K���a��/�9�{�{�9b�� ����?��߲�Drvu!��c���"^W^�ܽ_��&���bF�X0tݞ��4��c�q�aFz�<ǃ�g2^^J��iRe)vAt��2RCߪ��T����,����zS��i0��r6�ڲLs�:��X1hukK�ݞ��˳�_ɱ&9�_���S}﫻'���\N���%��k��ABqdc����O�k2Nr��kF�<ҽp�m�}�Q"]�!}���屰cC�l������ѡ|���R���ք�^��:�����C�	=����:�o��x��.��Pl�đe-�p�#ߑΫ.�!!�Wa�V	8�&{��˯��o���K���#:@+"�U�9�:s,���Aޔ�*]�T�!��0e"�q_zW	hu{���#]M`�Ꭓʰ���hrѰB�?� M��hKϢ�1�l���6�G�9���Q�+p]H����rE�4�dq7�n��a�ؽF� �ꢼ��։���|��^��+�7�8��M���q�`i���T�a}ߥOƏ�OY��Y'���+3�|��/`Dm�k$��|@ei�qʒb�\0�����0:Rza|����Mb�_���N]�Yf.�(4�Q��~�Jc����S�,zz߾�7q�Z,��]I��UT�!C���u��]����~�j�DQ�	�ӂ��d݄���=��9��ӢN
*%
B��\�Øz<���I��nS���[��zTA-�Ǫ��{�������+�Fn{��wk�t��78��T�r�t�u�Zk���A��M�9��\L9�VT�!|(G5PtRt�Q�Lէ��F��#�	�~ђ\7*���R��>�ͭH�Vň#��A(ͤI�Iʤ�%��__W\�ժx�cp3q@��i̶�8���>e�|n��6?x�@޽�'���,�z.�-~�f��ݕ��{�|�H���G���96�B�\G�>wj!�9B36�Y�*��*@��Ԡ$�7�$g�K �c;f�>�qb�l��Y� iO3y1������|N���t�(F{�A����j�����������:�N��"�g�p�E�V7l��/��T`8���o��s��:����Txq|i���Va�q�5P�D{~5�π��\P����#Y���Φc9<x-Q��@��VX�ў�@|Ɩc�d�J�ֱ�e���L�AĘ	Us�ߺ*�Ձ�..	V��ɶ�P��5y <bDB]���#�/IC��b.o^ʩ~�o�_��=ܖs�lpF��o���}��mO2�Mf�Aͣ��(��@�u����-0g�P�V����\̱̪��0� ^^��\Ϲ��*|��e��~zz�`	���=�=�ySV�X�X��B�ֹ��qr5H��g���4ie0fDL��V;8'8��ᥜ_�i22���$�.f��;|��;�@zz=���,,��j[$ă�[I��JX!K��v-&x.Q��v�u�.�A~���Äp��w�ꏱ7*�"��9�.���d!sP��I�! !��~���z��ݑ�����Fz�H�|��f}P��<�c�24ԑ�͜2�\�k��&s�KI5�/5q�g$�B���.q:���̂T����屼�:���sټw_B�W��L���k~4�x��7蚣�5+6���4!�8;%�A�D?s��<��Ty(��~��}p4�(��ҟi�N��������@^������<=|)��L8/M2<�Z��·ߕ�~���b"d�W(O�&��NC2���'�ɧ�/e��
��+�O�$^�tNt�3S���5H�>?���c�6��Y�7�0e�*?��l.�DU�6T3�������w��Ǐd�݇4қ�J]o���,�y.�2��M�|v�|�`�� 4���E,|o����a��������6����,�Σ�ؚU])WL#3t�!:b�5�&�T	=+�cܛ��#�g����Zs�������ևk)󠎧8+蜞O\�Y��f�
�>?			�b]��:>)�E�F`�
'R�ӳ#��3�Z���L�p*�x������r>:�X� m�s�Qb*t˱�N�3i��@"�C�hi��<��$�qS�Mw�U�������ҫ�F(b�Y`�L=�0�[���'�p��T0ސ{���;Ek����L��*�I���;KH��y��j묋��<�
��Z���/�1�V`D;g�]���u�D5�r���c�9\X�PW�S:g:x�]����F\��Ƌ%t�E\U:	��k
`��)�0Ƹqd�B�+冻$?��HX�)��<���UzX�#xD�F_�҂�9i��{+�h���	�.��l�`Mc��w��9$�2%�����b�q��=uI\��g8��媇%v�%��d'��\����YĬ�w������%����\~��������~%�<��wߕ���H�~��y�P��D#i��F�D�H���P�?���_�lac{]$X�<����*��R��
��f�U�R�n,\�`v���ǆJr���X(G .AC����`۩����e��y�V�F�U� ����hUR$?�8�5ǇG���s��ί�G՝�P\l��^�3���ɛC:dr���tҋ���~�8����X޼y#[�=���W��,�֘��T�FW^�ql�G�~GǴ}Z���ϼz�B�\Ne��������9���B���'T�Aք���_-��|)��oi���	r�吁2!�z=��Lj�NN��W_Jwg��a��z,K�+�}�{ϝo���sVNŪbqI5[���6���_?0�G��������mHݖ�M�U,Y̬ʱ2232"c�<��{���Q%���$�u���y�3|��{���Ԣ7��ѡlomi�p,����8����l|�\޼ْ������&I�������Cy�䉼~�Z�/_e���Sl4�Zpp�����r4Ll��c�8��������
n}�P�
��� �1(����I�1�PP�
�e��G�������<�G���j����FFG��uԟ𵠏��=�������]��*�id0ImJ��
��=�I�Ni�����~@'��d�(j�"��jftkڕ�����x�n��q��m���5��-�h yoH��Ne����Pvr�3|�yތK�fע�$��+�~���vZ2�Ϳ�k
�}�}��'�!�[R�L����F��R�A���5�c��h`�s��5(յ�T����G�����P��MT-��%8�C�1�~�����Ϗ	��8`p��)f��Gp��%5�g�^��ݹ'�:�>2�^Jfa
z4����yW��tQ��!�H;�~ ?��r����^X�z��A7.��as����I]��uR`F�P����r�p^�5`�~�X^llp�cL�WD���LC�m]F����1�ZS��5���ukP](��*˖��	Pv�s=}�>�c���L:��Q��BS����@��u��d��C�	=t,��}Y�a0�խ}d��sd���) $��g�eV�Q�NJK��S�g�u�CV!� �%5��	�1�w��@�'�ζg�~2K�f��IR��B�ѱS����yd��ʳ*����k�ꁥ��V��g�k�L�1�х�ܐ-p������c��ݱ�Ï�s�����{)b|C�Tڌ�$q���N��`�9�@ N��1���*�l��i��w�;� �{/��4�����H����B�o��i��q�7�8b�W���˹�@�6�>?Q���=��=�,��h��T"����;e<��1n�TҔ���5�OY-���4�` =�w�	�>���,�{��$}�V��&�]k����^贩�+��<zF�0���XE*�1���#0p�z���AWF�;��tcoi@З�I�@%6���h�ќY`i�%�Y�䛩���mN}d�&������jAL�݄ ��h
x5��i(5fC* ﴢ�AEٰ�
�8Z��}"�P
�DAa�#OF
.p}��@� ��°z�+��w�@�oܓ �����od��{_�=���}[�;7D�`+̂ �W��2��� ��1�l#�"�2�wc�A�Y(��Y�ȳ���k���K�:*���O�;�|1�&~p���c,��2.H5�\Ĥk��g��%y�w�3�+��4!;����fs�A�v�]CUF�%�4�����_�Znߓ���*e����
����ޑ���<��k���7�|�;P[P�AU��k �X~��������wdfe��"���RЁ9��)�<m4�ݺ'K���DGÉ^�P���x{�|z�w��<V �|���]��f��_�����Y�:�ps���m�.ʱ~��<�O`�:�V�_oɧ�������`c�
��:m93�b���k�
���U���t9>��ڽ7����ul�x�B�ÒT��(���S�7�8�qb��t���Ȍ���<7L�s�U*z��)�KPQy�bCn��U:G�e�TpxfB����縧�E(��|� `H)jJ�4#�ֱn^�o
(:-TC�ev�C�?�+*���z$� ��sc{� +FPI������$FS �o��u.
�/�it���$��Pg(uљ�ҳ��F��FB+��$`=K���M֙QD�:�YT;�)���FN?�`ͫ��#S�y(����Α^��~�kH�H��ֆ�k�=�P=!56�}�@��K=G��B��q�K4�<LI��~�j�
�Ɠ�
��Ć{E�u�4�ck�	��2�[ohk8�0qB�C�P�@C6�X��P!�Cf��L�0τ���S�Kl�6&��K����A�<A��˞,��2�š�'�����t\Ֆ�ȧ�fc3�
!��]Q�\�P��ӧ��O`e��0S�D	�:��&�&�?��lsI�͞���} 0��+@�bGI�{Au鲔��B�08�cb����8�(�&�>��Hn	��(���*���|�{J�Z���-�>{$(���	�*ܡ���-�Ȋ�UzqOS�;���=�@T~MD$�
��L�~"�2�c��O!	K32"}o
��g�+����	Z�,9��MxZţ��7}��}�N���L��;�`�ɦ
f�)�_˩��	F$�ŷ뉤*ծ�͖MTk�p�&Ϩ�����{3żg�q�	��CWʾÂ)�M1�̛J&���XqY��4�
���ze�;�+"(����Ƌ���Rzwӟ�I��8N.��˒�Ù�6�����sQ�L9�|:P!��Rg���< DI�5�f~l�4��8�|jC��3I��l�>o�����ܠ��XI�FW��x���5��yUPt��0��c<�y�'��x�:L2M�z�OkM������/����ID$���<pҬ�P�ZfZ��	3ޑ.���$(D���d4O�l0�����h��jM��t�UW��R�U��2�L�4P�W�j��]IE�ɥL;�o��� �.1K̃ј\d��P��4�˦�,1zg���J��PE4>�� &��tA�尠`�e�Vlz�P�E�2�(k�nKia��[:ю�p����]���oIx���G/_K8Ӑze��ҕU��C4:"� lB�J�O � p���L����"��.��b	u�����,d֜�S�2k�)Ȍz�rF�>dّr͑�F}�{Ϋ��}?����|�٫���+��Ɛ���cv~͜f�vK�:�jz�`�#��7o�4����t�z�
�7_��H�}sɬb ���;��@ ��&j�P �٥9fwP�B ���&{�i@h�Ԫ~�+_�"�,�D?�͛7�g�7p$�FPip��FF�t_\�$�P�s�m�j2�c((�Sf� ���r��-ټ�P�^|�>���ǅ|}U�	��Q����r��z��t5(����+�֍k��סQ�Z������U6$oh@���� ���"�5��2���Q���q-�x����fE(W)}�͆:NA�Z��.���hO�m,��e�t�����Wd}uM�c��#����˲����&	P�Y�����&�"�8�\��Y��*�4?V�S�9�O��34(T�f�;�\���=*x��5��U� W��׊��������/���R����T��Ql�=#�#��Cp�
�b��|��������x�#,�$3����0{2�w:�&��y9I'[�y��r�4���k!� �)i���Odc�P�Č�*aX1^8�y�>)eФ��#7�3Âίr*jUR��qJ*!@x��AA�gFq�94��*��&��>�����.��5�S�)T傮�o��?��} �n�`���\,� Kx|�rM�t`�����h4g��2Vmԩ���[��s{�rèj����C=���0�p�s���&W�~_�l�����׾&3��(��A�g<��������,=�F%�kU���C9�����.;�<6_vڇ��`v���r��;r��[������UT���҂���|��ܯ\�*+��)�5(h�wUI�B�k�G�5�]����>�����3;?�k��/�Fr۱�2Q8aC8�>4���]:6ڛ�pG>6! ��xLas6�>�Z  YM}�h< [`80��r�U1�^3����o����������>�g���TgG�W-�e�Z7}�9��
J�-��i;�*�-�����L��T��%����* )��\��F�ʰ_�m��.��.�ySf ���%�'�1i�9�A@Al�{b��UB��2�W��b� u}�vyN>�c"s殸o��%�����)RjR��<��X���L�<ϛo���m���q��3��z!�z��3x}���cޓ`� �)���Ȋ��/��׋���}f�2jo� r �SLqV4%/cG���iRC�P�v�E�$�S K� �#b��Y����=�џSW���i��弄x/�'8p�HO?�?�e��m�f�๊��G����B}�2}��]B��L?��ev���K��e�Q�B<0,�AX��Ka� �3=��I��L�Q�����q�$'q:���ec��f�i9�'}]�+�����������6+R��F�Ho|#�R���&A
��^w ����x0b�9�h Cq��JGA��2j��Q�9'�����ڜ*Ȧ��/ !%)v*%X|&X0u��..K0��I�w,��3s#ڔ��}Y�/]��٠},O_����CX��ڝ�Ҹz��r[O_��O��5yw}���
R�gjR+BL':�9n�v<�irR'5�ZIS���(ͩ��͕��ֱ�%�GB�Q$o��r��m5��8y� ��y����b��|
��a�'b��f�y��~�z����X�c6�^l��P��uq]����_�B���P ��
O�`U X�q]��O�X�޾e}�𔺀����[t@˽�w���S���F.��ug#���	�M[��4�f�[�nѝjXt+0z��6rE#�_.���W��U��K�Q �I�*�α<�@a �HX���9y���ʽ��.sK�
|hPP�M��M�~��֖tC:�^W0�50 ��;��f����\���$��o�uC��]
xS��Ʋ^�z��>�~���o��E��w�+7n��ģYo�W{aeU�
�H1�e~qI��ܸz��+�p�^^�H���=���+�r(ׯ\��|�2���s���^\�Ź9��������k�䭛7d�T13��굫./ʺ= e{z�
��g5�,��t,A���؝�W���u�(*�D�@Vf�6gz~ ���}N�����6��-�F�ʁ���2�c)�2�.�W���C9���D�e,�Y�2�dA{�}3$��\s��!���9m�
}S����ZLa��x��X@%�X P���W��
�ƭ}��Vt|�g�k C5]�j��E����������
�uM�� ��8 �ïNנ��]\�9�8^eV��x�)%`���������^BQ���W.��7��rr�/��P�vM�{�c	�f�ԍ�,+J/7�����3T�Ҁ�Zc@�9�b�)h8'��Z�()�����X�u+w4�ė<���H����xzܕ��CR�P�@%���%���,�o��Pׇ���B�{�r����.Ӊ���ŷޒ[��'R���;�G�B?��5���  ���t@w��}&Kk�kE�']�*4�L4�2��&z�\�)f���ΤS-1c4��\���k��2�����a} �D E
�l�Git5z��I�aƉ3|�X���b!b�ɠҸ�]~�v���бrsI�21�L��ӄ%m�\��o�?R۳���T]�%>m^��@!�y�W$;PL��.�;����g}��n��|,2����'T�C�_�Xp�d�4o����R�{C��?�-99��mP�k�����=:nFtYB��THPQQUF�K��<��1��3vL�1u=oJ�*�c4��q���S�����v���^��ߌ&�;q_�'��a0\�{�|j�a5�$���D�8D���@1V2A�43���b)�K���1B]���X����0��x�7��t��b��C��8cY�w�4@��~�@\,'$�)��3fH��,�̀�3�X?#	 �_w<��.�B���	�&���i�����Y�[U�$��Bf�6�2ر���3�~���gR�RRbC��'�I8�������I�I��nD�4��R؝�����(�ܽ{w�ygyc�
���������}��X��>D�c��ޑt����X<38��I����T��A�ቾ�,��5n`^!ɩ3��Cr�
�e��CianiQJz';��2:�Ѡ �`��f�H��\\�!��>�ޗ'[/d!jJaF�2��	)O?���˩����R�)�Z��rE���JR39%%ؚ�L�L�ё	ڴ�Pʹ��$v���~Z�@ʓ�����O{r��|��>stJ���mQa3���Ҿ�w�)�-��4$������>gjZg�pO�30�>VW�|��6�L��-Def
����'�)�.]"�5nzK�@�u�;8�
�H?��A[}f�U�3x|�1Ѐ��V����Է����\�kdi;m�r�|-͠�mA���9B�k 0���8����K
�C�<p�i���[��2���dpt��MEl3&�������V.,K
� ��5�)𖲩X���@��*#0T�F�]d��h�vx�[U7O஠��:/�w޺��Œ����� �FAZA�� 1Y�
�\l�f�C�7�Yh��B���h���?�{t���*��ΐ��s�QO{~F���xx-��6��D����N�9֖al���`}bh���*$%�A����a�<ᑂ�v�>���B�7/B�ml�4/�;�?��	�i�h~ᙙ��V��A�|��8Ò���͆�K#
��}�̶5p��&o�cl��u��BC�EW��dpYQI�r�I8t����r��cA����&�pބsO4��ݩCy�J.���^��{w%�`��x����� 6:�.�=�pc�6�O0���P�B?�8���\^�{KL���z����t~��^��5�=���Ü�`+�9��)���2��4`Z0�-�~��vy�ք�*��&�̤��<rp"�ֱ�>�ʤ�աZ�+/��;w���{�i�H�f�rљ���\rխ���17g��-}a�d�� ��b��x���bc���Aa�ەe�D@�M���@�4�2� 0R��
b1
��n�)�V��H���K1�IʆakFW�0�2aU<=&�6�����#L����D�Ѹ�j<�}��-�ԥyJ�v)�$7�n02Ua�=qw�e���o��@��&��^�3��2�+���U/\�E�Tr�\$�'*�f����)
M�c��He�U?�T��S�S���v$�Z���NZP3̝��E�`B�m�+��iV���g�N��	��&��q�%E� �C�f�@��E�](����F�"���$���A�[Nʃ�^3N'M\�,��3�wE�AG�!f�
z��c����8�;����
�>�H��3j6�l��L�����8�x�BS���m��_�M��yG�ybEv0�����<>|��Փ����^�Z�8��'T�`�Q�݁e����Tś0(@�-W��� �'���5����h��&�7��g�ĩ�����������	+��MQvK5���f�IԢ�Z�M�<����I'����T�F�@��4/*�*�2<ޒ��g��ٖ9*�+���7��ڝ��,sYKe������t��i�˂޴�l
��Q�2ρ�Խ�#6v%Wɻ�A��u�]ƀY�u~�Y�XhN���@L݊�gjH#�s��Ϗw8�\6��,�x&S�%o�q�g��zcԶ��X��6��nbSS`&�  `�����MMa�J[��@ ��h���k1Lɕ�Fp�n��d`�Ӿ���{��Y�H��L�釡�?4"B��G<�������x���Rxt�ȭ0 *@:&�m�됂�c���0	���!��b�(){'
�z���3�����
L�X?�#h/HEA&��P�"EJ7�ǋ��m�y��<��46�aE���mܧc9$p�
��$�[ � ��J�?��ru�����Ҩ��~q��p�>=ٖ�����`�WP� �ŋ'z�ERaq��h[�'��)|$�ʅ�t����T��"a��5�#�NW]#����Elĩ^��b8��G3���~�&ސ��������.�ܜ��WjlY�R�9���ǈ��hou,��!�>}wH��}(_T�W�ϳ�����k��74�g�E��6gQQ��~��7ά
�h�.��eL��-&�}>��5L�f��zڧN	�r�c^[�j��q���.��3e}c�~e��0��y�|%C1π!���n�m� ���X����0H��VT�@����^�ag�[�l�g��}�5�=���|-�*ȃ|h �ڜ4�iྤ�<l3)$��5��Q%0 ����!�wa�_���Cӏ��	�h?��fZ?����nkZ�;b�F�&���L<2Ŵ4_#����f� �����]���k��׭ׯds��#��st!Fr��,@�.��OH=B�+��(����F�:��w�� (𺖹�33�K��ѹ`zڻ3�N[�d�g ���Dg�X�}�ǵ��� ��D�(N���܌��)�H5L2��a�b���d��4؞�`�PV�������~JP�Я�rU�Hĵ�u>�:5�tM��RD�j\T��0�XA���Cc?�c5��bs՞�^%b,ܥ��<&B��z���33�E05�F�i�D�P�R�K�~�7	KE�=���o�c!�I=�t��<��"��]�mh���������6�l���DX츀N���  ��IDAT� ܉5ՠDo�bn��L��*���*�L���;#c�:��taAٴ��E!K`��z�1��17#�ߺ!ua��~CnݹFS��_?����ѿaa����ίNWv���s�_'v13��+�T�����8���Q�����<��D�m�dey_��<7I�������)����eH�J^8��T}��~�)�6�&K]��7�Ud�(F�*ໟd��Up�2n����nA��j�&a�I����kjg�X�	�1{ �Н*6�a�J �M���.Γ���v�]�Ӗt��Lz=�u��vNuQ��׈x�d�4�띶y�!�׃"�W�J�dHJ����+���ɄM]�v��5��cf����]x�AG";DhT�t�>>ܕ�=����������;�Ų��){/^H����g����y#/~��C�-�������J_O��_*�_Nx��4��5V�\��S��@Pw��7��|�o�ۂi��
PC�EeP��n<����?���
�}J�tve��3V6�J7��W/���P.�ڐ� @�ou��ǲ��g�>x-af`nkC~񣿑Ã=�w����SQ����#Y��Ը�D��^}r����g�&��������/>���c3�4��=ŢϦJ� �S���9%c��M֏s�p��@��f��	�9-	�^��3���|��z*���!�r6c��5�ft!��:6��]�{�T`>���R���te␌h(�֘8�"���4u]*����c��?>2P�8���Gs
��!H^K�4O6+*i��'�o^�/�;����r��fE��.�=*�%
��:V��C�y1�׆�hG�
�K��r������@�z��#]_��]����@;��G�-�J�a��ґ�^�R�� M��X��*��u�9�����Lv��������<��
�q9y�%�$~�RZz��3�4��3車4��mɜ�KU��Y)ӰF�=�L�{�ٗ&s��,#��g:Z���]&�%��$^D�����w@�K��hܡ��M�0�u~��ʫ�y������K�^4�C�J��5��%���M�en���>��sAW5��tj���F�	�=h��z��EX������������i�����y��c 3y�=�3ު䭝��.;����u.�C��L)��r�?{�P��^�dN�)��� ��*�(����Jʆ��֪Rkԍ651?�A�UTW^�Y��$��X 	& �Z�}�v�܁�Y�q�N��a4���w��/2��$��}
���o��[Q�������	�>|������i�tr�B]jA2�ެJ���bRhh�:�s���.`�-7����}�Wt=EjwcZ�$	�l�iDv&qz�A`	�	h�NS:�_Gr��#I�̍�&(�";��.�Aet"��ɎWeeqM���	tC��2kC7ddC����RӀ��{��VEz'r�����Y�<#9E����q���ޔMe�� ��p�����$S����'������BȆ0��H���ɗ&=`bՄ�h���O�eG����9��cڪ�j<0�x(l��ו�o�ؓ{�N����J���7(��X��oߑƼ�0����~oO�z+%)(���F8n��2tp+����O$�HC�BiFj�ڹ�L����b��*@�u�^F�U7�>G
�[
Hn��*�D�9�q��8T���y����u�U�M_��
"ِ�c%;z�hv[jC(���R@�~��@z@��tA�sH3?,���o���&�}y���=�4(|#x�|�n��I� '��S��m���#y����B��f̷�-}�H��Dj���T7��WϤ/�*�L��Q�@dkW�`_�Ͳ��{��d��J��9�1��w���Hf�m�k�JE7��γ����ǟ�Q�'v�|Po��Q��r�D�P$>�O�l�C.��{dp�������֠g��6�[5&�JL�Zr�@(y��?��
�	����5�g"��Ę�5��1��'4��0��4���&	0=}��4z���w��E)2gF�~������@<A�f��˨n� ��AC3<�$1Oc��r��M���É%I�{z���uN��w�������(i9���u��m*��Q��VW��{��w���.���2���L���[
��`!4fgdny��=���ۻ:]��=#88=>��'K��r�����䐮�3}R`��O�ٔ�������N�~ld�[��x�Ӏ�.���V�ӱ�c�*	�)^�Fc4�/��p�ky���̊��j]...S;?�8d�8��D��u���\m$�03	�T,d�Q���aM���F1&ъk[�ޫ��=�B9��/���e�̒��t[f���ף��`maY���1����ّ$Z��.�4	D��Xxej�b��֥�A[(I��o����5�Y�5D�(''z���.!��*�xҡ`�@׭��My���n�~��	QP���@4F�8�6g(-L�r��qT������[�>�	����*���2/�Y�[A�K�le�!妞��絎�x���K��5�O�L���LJs����;3�*J�g�g�ܾ�˛[�nRF��%uJw�u�
̶1cN�@��_��ޓ���=v�.�$�"]��-9��pfa^JhD�*�I�^w���B�����ˁ*��4��BdE�H^�z�f"H��Mw���$�P�D����T$M�޵J�4�\��!{�$j3j�q�))LF��<�
~�z2���H�d� �@!mB��"]茎tAE6�x�s?�|k��$�ɤf��;�x�3=9O�����Yc�s�E�����f땜*`>=:dY7p@&+����x&�>�H�|��\�pU���tG��'d����b�t�\��F�����@	2���L �rbn�y��l�s�.��W� �ê��P����H͓���"�td2�ݞ�^el�̘U2�68x��T�#.�0@C�,6�89���1�|S|��/��?��+df�a�Sx�h-���\Y��
�F-��Ep�5�i�u�:��t���S W�/+ �C�+m�w@���o6���`Pk�Up2��Q0;� �h�T�'��x��.�1xD̔c�Q�*h�_����c���;��tl�JqБ:(h��\dcU��7� E���KI�%k�t�k��g���R�6�,�p�hݺ�|K�I4���ͧ���cVG<��+�f��l��D"@�DAuo�1<��4)%6|d4A��LMw�CI�_���}ݜfه ��nZ�>��^�%�OC�<(X;|��_�!l<�
7�I�X��=�P���d}�N���*�p��xX��̪1�'�(=&����pH3>b��1p�U�B�ߌ%�ͧ��j����ې��oc� :
�ąe�2j��TO7�Dֈ
Ffկ��|�T�����w,	�U}�8���B �d��h "���Z���q�! i�Al-+�0�P�-C�k���/�����{���}z"�0��#�_����_3PA����W��蓦��b�A�� ?pYhćh..Cu����נ��f�e}�t,��A������8i0<�H^��	�w�L�퍝��. ԁޗ�Z�jK���F���%���M�?�ܐ�j��`PQ�{)��, ���s�T�[��.8�%�B[C!��>�̓]������Q�)t|Vu\��������w��h�^O]��\�CJ�����y��Fn����8_׫�X���\���@��2�^וR@��ԥ���=F��+�(:���)1(��\:,�ܽ�?Ե(,V�ވ�ҔQ�p,o�����r��/o�}O��槞0h��{te�ʭ[w�����j1��3��
I��T�sհ��t&S�G�W`���� ��3$Ɛ~F����6U%'�.�����O:�¦�e�M�iE�%
HA<W�9~�Ok&��S���۹�,�O�������yP���8>W�H��w��e8��
M��[�o(����f�Q�+�	�!���;FEu�qINN��Ս�	�f&q�=s�Ǻe�	�����O�~�gC��m꼆q<tn����eP���t�X<��$��Tg1%hg�a�L��O��I����"��G����ȷ,�k0Ό�2Uh���J8VvM������/�����L7���7bS��{�������,�A*_�|O.�uU)�ܶv���C���ǲ��ĺ �#��@d��|�����gOe�i��3�>tS�x����� X��6]����}��&����gfh�,(}�$u�����C�/1�3��(w��;�rPb����7ntwJ���2,��T�(�eǚM���̚���d�V��:B�4��޷�^$k��D��"��+X�UASZ���<�۟K��5��nXo�J�t1�La��2�}!�-)�J��Qp�'���>���耛�A��m=Qpߖ�0U��YG��K��`z~����qK���|�Ff4(eC�R�J��}9���r0����%�<~B��`�*�.�z}�z\;O7��X������Ah<�Ҕ�wX���V����qW�?\��.�ʞ��%�h�M�Q�H���cb�O��q_M���!>䉼�˿���E:#�
����zmOe^7���Es�o$%=�����}��I�ߕU��:]=�aB�}��Hc�R�cfj$
����� K�� ���.f�� ،1�I+������JSB��F$��}�e��wO'(\ڿ�9� _	iH�Az��2��aHI�䄘�iN�p�<i>�t̀�8�ey����k��#¼,"[� V�����t�Ae�T��)����|�w���T�4xE��KoD��b�*��
��p{�H�;��V���h�-��Լ� �t ]� )�V�5���ܿT�g7=��oqz��M�s���v�2<�q�+���k[��^W��	]Zqk
�  �jP����i9+�ԣQ׼&&�.��H�5Aq�"��m:�^d�!ܠ�O�s�T�eV�q&��@��f\�;���������:҆�5��k�
����'=c�:��Ċ����P���=hk`�u����B3OS����P�P�?�A��:z�5$�/�4"�A����e�m����*���tyyo�o�Mi�ǄTL	�bQ�V:��PF`����w��`���zS�Q��]�1�(	����L��z�x���zܠ�a��"V8|��M��%��񉟨 ��F��X����w�hw�@Ϡbl-��=�y���=g����[[�^�K�fY�Y�hZn������YK�P	�\TI�z,u}mU?�ס:7+�0�vլ���1�A}#-ճ�}��|��5A'�Eb�m�`�psa7��V��_5���i���{n|�1��b��:��*��S�t�c����nAiѵ�f�||�>��7G����߽����q�Du��	��m��bF��n}q��bM{�Qλ��M���y8���|!�lEȲ y�b�h�p��n�tU$'�d�4�a�+�Q��-�'���+�;;r��23[���t�~&ǯ_ˠݗD7���K��'�|sC>��Ϥ��I:�T�i/�ɁE��.aՄ �)�&s?s� �)��g��X�)�z��Y[�)%0z^�Kt�{ �:+2 �=,K�9 -�c�k6#3�� #B&�� ��(!�=`9�]8?�?��	���3ҕ��!
R֍���D�((�UB*�Ds^��IOv^n���)�39��j6�����H�>z*s3������ѩ���=i���Y�T�����RV ��a��o�l��yrr$��m���d
�~k�����������c�΃N_j��T���"ۃυ.ܝ'�ʋ�m�$#�2VU^�r���1�`v��\�v�<w�h�t��xg�1�E�2֠����>�rw�,q9��vB�eХd�k�24�f�ѨW�1`P&S7]!F!4�C4k������/~!��2A��遌���(0��}G��� fJ�@<��}�n���cH'N�f�)���W���c3��hP�\�(ef����%=�2h�A�o����4�f�TH;�Kg�)q�=kv���� +J��%�L8>�
F#���:�Z� 0�-˖f��^�Y�>�V�n�%����A�.�b4)��7)GxT@�,EoG�����D���XW`93#�ׯȅ�uY.�u�z
�����Z��g:�_J�n��q5%�ڃ���P�lo̍�TrN����K��[�z4Ǟт�%O�(	�� ��*�}�*��hq�)�)�!��!OS{#�I-Ě��$�6I;Ѕ@$��x)�JL �A��$`����':ӟ6���:!b ^��[�ӷ��@�(8a�i08��@u�|o]�06�����m�ِ!Tp�R��K�	�n���Ա��X�0����K���~)�����*y�WE���:�c�P��,i 
���Qg� u��盳ܚ�yg{����LseV�
x�3*{�H���S�Jw�5��dw��=��9��]�v��(�|y�D��7&<����"k���y�R�ޖ˗/���E��}`Yh��>��S��
6~7;m�`:.:�FO�]vS���s��AϹ
���?���w��<sN�qL�F_�G�S�'.ɘ� ��/�ύ�_�d"��s�N�r:iI�w,���^Bo���'A{2���-�,oI3J4��>��a��:�@��� ��>`��h�j&/�''���L
�4�AŐh��o��b]NP]�}�&˹֋���ˠ�w���~�/����Nok�ߑ"LO��Hf�<R���e3�8L� 0C#9��/6xL��G���p���
	��I0�~]���B#*�?X<!�Nr	`W'O��21�@���
���@7o��7��A�-O�][��n�kK�ru}Y��c��������G�<�����#����5�����TvT\������qI+g�_L�(�r�����Ō�&��f�����C -��(-�=����i�.KX�ɬ.XP�98ؓ��W�M�)����4+C:|[�߽y%��{8�4�2c.�5{{�� �&�����2d��usFٵ��s�m���v9�Y�L��`,���$=�r��딼l�^��)p���42Op%��>�qR[�J�)���ZH#�Rc#F�SP.��������iL%A_b����h$�p��3�E�s�
��ސ�:��s$%�؆d�C���hgu���-Y���e��2{�*���Ո �j*P,�H��/e��Z�?y&����@���q!�I�,�S���M�,5zE�9!�1�n��@C�RMx}_Q���s��>ձ_��k��(���T�
���x$?��|vԒkKKRQ S��u���tL $��-7�|6x��5���7�Q�6ޮO-tN�ׇ�2�`�S�Y}��r`6`�S� p8�3�(��tJ���=�	-��;du(��E��;�fwuJ��W���C��#{�d0	�7Aj%1�YO�����9�%$=����lR𥧃��v��%Y�=Y�y[��Ň�n�����c����է��ٯH��K	�d\�"h!}z�$:����X�sh�D�  `�ܛP��� ��{ Td�=�r/p|�\���y�*�ȹ��7
2G7��e6m'�Π �1�s���5J���6��4���L��L3��x��;n��9�"yZ� � �)$N��>9d�a��������EVj!p��ܨ*pN�҂R�oT0��ơ5���uO���k �<�����H�5r���N�Zž.�;A5��ZMVt^-B�����µ��?����N�<�� +c17yq2�XwQAE�&�r�~.j�E�~�k��¬�ɘ���]y��A�ǵK��\�Q� Yx���Ot���G���;;;���Kp������s9�q���������d R�^�씂�*Y|��;Y�UHH�27-8���! {���������?����ӊD����^d"����҃���wf{8�������G[[�����mi^�G�����-,�I�F�NP�����M�<�@��*�pa�o.Z���m�t��I
0�`йk��A�I���
:V	��y��>�M��O3�/�����;�����������j�>}��	�:ر�Ys^�T�ڂ����{6Q��'3�RPN�:����*9F?@�] �P��L��*8�RL�j�2�F��CFY˒nXe�����ʭ�����n���N֐
,��҂��~���H�ޗ�O>�B��z�p��Q#�P+�<�`�9�ʭl�L]@jM��p�^ �����$�{��s�4)ĉnV#��	�$����+��?�cy�{�O���.X�ޛ�����ˍY:=C���P�9y�B��������hl����N�Y�=L���h
aB�#�\�5U�\s=�qJ��ݶ$��OG�=��-� f�.���r�;�'��y)�q�� i��}I��u���Q7�b�*l������'��|.��zH��``����5�j'�,�j%=&P�D��O�Ҝ)	Z��G�o	ԑJ���N��bH�t������i�u��r������ �3�� �<:ܕ�g��𳧒�o�T�����:>5���1B1nݾ���b�o(�ӝ���6@�A3bF`>�;&rz����� <ZAp����,���[޻+���D���������`΃,\�Y����𓏥�Ⱥ�cR�b�����>�Q9���y
y�̩���CZo��m�4�qT�P̹���	Z���[���1z@�:���}>�+�d������0�+������A}I�9 �	�t?�� �;Ȭ2��?B/�����4�Հ���E.�Y�?���W��ܚ�yI�ί��˷���39����3���
��Ln@e���II7u=�B1���)¤�=5 f���Q�@�� v�. i^jN�(r�]=�1��gr]���gSIArM� -�����p[f���3���Ϸ��[	E=�Sv�T���~��UT�O�d"��.!� l�t/d#�@�f$��#%��RUj�6�V�:p�e9eS�b���u�*�zP�DF!B�{�
�~O���e<a^�s������d&x����45��nhS�|j�%����vT���4�:������)`�y�\�g���}�Օm>y,Ϟ�����*u��"C��D�}�|��߭���~��<|����]��F�
9�����#qԠ'�F��֝�S|f`�F�����%�\�H�����=�L�/���=���{l��6_���N��g����*�j�&�����9�'�� ��})]�,5>���*���hb,	$E3�+�='�:�|��iIqTdb��T^��	�>�j��B���J�5��g�'��z�Թ�<��V��__>�q������O�7^�T+F��n<u�	6�6���}s�F�ܴ�-��e ˜��q��3����g�3u�maʛy���4q
$Bp_�y�����?��>���u^���}'��
6X��U
e�������@���oIaeVOҘ3Т�dA*~In-_�YX�.,�f-��O�������Puj%�8d��8�������9�sS�}>�)�Cd�|F����Х�w�Zb\f2$)���9Ӕ��ɍo}[f��M�2�66�V/�˅�ש.��s��L�]邽�yQ����IopL�J)������&;��a�e,���zN�:2��N"�L^A������璎�������|����'�݉,���5���� �>%P�z]��\zaO���ӓ��P�c��C|YQAw&]4��emPF%A�*�s5 ���j���!d���We�h.��Íte�k�S�1��U	f����Ml�d��F��J��}��J	�@���H��60�J�]�O#�K���8� 8��kU"JY���;6VT@7Ɍ2�B��3�-L/��c�@�ś��!�K�Dn�%��eYD�����4Ț8#0�n)�i��ޕ�ɉL6��w� PQw�eP�0gA�2c!ט�uT�<'Y��=Ex��A|s?-���P��3��<�hz�� !���PВ�,�
ꍙ��:��6f=g�dFHg�A̦�Ԃ�,h����8���`��o�XN����T�~Kf�����2��F��c�	%9�g��va]¹�"KWD�uY�Rip�iIp�k2� ��h.�5B�\��(5E���\V��IE���Xb��?
�G�g��I��ȦӚR� ����ӭ��ف`;�϶t(�etHO�ZR&dA���I���0�s/����V+�t{��`�����k4F�2���w[]6_M�*��q�s	6Ro����D�03/G�>��Qu@0�z���1�|����2:���]cx�0H��^��P���*z�#ςN#q<Rɥ����'F2�u�sXv��2�/�8ŋ�Xo���PDC������tΗ��a[�2+[��jsS�iP8�>#%]��9�4�z���3�e�d5tAP���/�\���uy��B>Ӏ�7�����,��ͺ��b^� �yP���ʆ|���,�>���9���3�o��}��,��L�t�����鋁C�+�}!��� ��ܸ��=0cЌKc�{o�{Ԭ���(t�R��2p�ƋQ=-QJ4��.؝��}x��>0����d2�U���Ľ6�d��ȫM�9�VӤRQE�w��a�?gS�&�4��՝Y~Ï/�����ҽ�w�=��_�G��4���t|ܾ4����.J.�^�I|V�;o>e]��+��l�iy�UR��8ET	���-PY W�⬛@:I�;�h��v��L��n�$�}P�>�i�>�y�ko�׾�)\�M�}$���ْD�?���5�Ss��-���4�%i�N����p���Fbw.��`
��M���<��S����.�S���gena�M��;;��.H2]{� �~�|o؝<�z���.ɍwߕ���i@4�H[��D�/��� J�w���i�rQ�/]���¬��Y)4K��}6=�943@e��[� �ƃ�-(���`Y-T	�0*I?r���}�ە�~"C��b� E���J����;
��LE�pho#Hh�L�_�&�z��YZ_�.\�����	8�.P���q7BA"�� -Yղ��B*.�z��o���)�7�Yp<)�3��:؄4n$���RAu|���R8�1�o㔜jd�:�:W�b�>Y6��:pk G����Y^+�d�,FZ���	���i�2�1qF�mJ�ՠ�ltl
#�����0����k�4�J r�a�A�2�Y!�O���3�_ͳ���%�L�$1�=ה��;I�qH/6����M���@�y�@�����R�@�X���,�"dnku��'&X �O��~O����f�>",�a�R<��`�:����ќ�Ʌ��ܫMy��G�9z-~�X��s�^�%�tsY�e}߼� 	����q�> /�=��@�9>�x��o����9�z�9�8��-2'[3�x�{��
L�?��*=(df
�����ű3��D�BFS*T���;qQ!�@�c%�k_�@z�)�UL $��	��0Z�N����MĘ2���x�ɑ2��C��[#���8���A��ta�I��\@ A��zS��Pz�ak�@�X47iT�@��<$�-h�A3{^Qal��(�LѠ8����ТĊ�uzP�b9Xxh4����~SlK�sx����w�[�YS/�x�fPu���v�o��=����K)̯��*�ɀT륵��0��9R,U��ϳ�"^���������ܢ�Z��W.����+���17f�5�P���H���.�1#d�����Yv�?]Pp�gv���ڤ�����x�r�����ϩ�ѹ�"��������.	䬪����@�|���5Vbº][P}��C7���;w����|�=�,�{;`_�>��Kp��yL�+>��� �~R�Jv����5R{�n�Wj}��Y�����_�㏛7�?����Y�yo��o~�/N�I��P���K�A%"�]t�&w^n��x�&e�:�<_��i�eDB�2s��$ÄΎ ̡O �z�n��.C��@��ԡ����n��B"���t�.^�����7��L����=~,O~�ٽ�H���fQ��k2�λ���=�z[J�/��oM�^=��gO%>1�j6����4�f&��sJ�&�����
<D��<�g|���������?��?�Q�C�aQR'Q*@X�� �IQϿ��=�H�~������_���>|$���.Øf�;�#}�����_���4޾�F�=�Փ�w��< s�f�6)�,$	K�<ϗ+�-�+�����u�5��۲��ˉ.~c�BAT��(���|���L�7�r�kߑ���I5P��7Ň��nV��KO�s��4�KLw��͆9��t�TD��pm�G(��+�@��q�8Y)�mM�&r����2�m*�&";��d
e����X���c�|X���ے6�|M)^]����m/ܹ#O���wt,�D�a_�,��~z��c@��(��*y��#XK��-��5 ���<A����0Ҡs����8��@�r���N�؋������	��w�IE�K��§?�n �u<,�^d�H4Se�0����� 2�=�p�ļM�Ck��V��~ޜ�X5�P޳ dWm��S�I���m� �ߜ����2�x�x��O�iR!vk��֕��+�z��R�w2��=SP� �$M���������%{T���#@Bp������z�TJ��D�);<��lO��K8�*�׮S�5TP�ԫ��c���4#hΜJ�SJ���sG�	WNt�;[O���J�{�bL���p�G� ���%d�3Z�l����V���*���z�y�x?I�H-�P���&����d@pc+Ft2��K��H�2��l2ֱ�^W^{���+��Rd��W�jw0�����X�qt7џ¦L�f��:GՂj�^{��:����6���k���z���s���1�jV�l���C�Up����L��U��ɚ���s�<!��eG���u^nw�^�@��H�%	�y���J�ӗq4�ܐ��U�v�����ӭ�T�K�Z�R�n.�ЦרVu^9
фk�k7���Dph��tJ��/�y����G�ꂤU�<���E��#������*��Z_ٴ����?�*���R�S ��}*������?G�1<������?�M9����v�IF�H�.�/H���,�U���ri��S�o���
��~HE0+�B�0��)�Y�$M,�ƀ~Jy�(��]��pZ�U���>�l��,�`��9_V
�|��?��/�����nu�}�����T�����E�f��oRlgQ{>�éԙ��z.f��M���f�q	��
�OL���T�u�cӀ�2d}QC=�"d;A9Z^�@&�S�=ߐ���_��O&�#Z�G��<{�R&�_��Ζ|{��CM
 Ns5�+gÅ0��B'S�C.v��";��:�$51O�"���鍤���ߖ��џ��WnK��R_���ɱmT� �2��.(>���(Ejp���^����{���<�կ���>��QG�P��r�@���n��?ؑ��e�:���=�u:T�(����`�{i����g�,��������	*�n*=����m݇[�T��5]ù��à���)h�W`u�zW��e)_�,����eE79��㧏���_�J�������˻��4L��M�~<fF�� &�J ��:���s��lL�"�Q0�>�8�C��qA�P�
�?
J:~'î�={$ۭ]��R�rU*7ޒ�KW�:;/��,��e)\�.�k7,Kp(��<��$'����c��鞕����[����LRR�
���c��'@2�qjn�ୂ{�L~�l)���RU�T�m��ȧ��e�3���Dv�Z}�_��\��"�[ϟʿ�W����|#�������O$l�( �y�q�fH��Lz�_r
ew�f�̉	�܌2��~#����:����s�s�{�II��m��z����e/�
�TӅ���ut�T>�1�3�p�K���j���L ߲��rD�S~�`$��N��\�{닒�l��'���-9����Cճ����g��U�2@�)�����t���S��*�I���`\ReȌ�p����Q]ֵh�scw���d�?M4Fef��P�7b��{�
�9�B6��NĚ5��9�����N�^'-k��e����+E�kjM�"�l]C5����~gWA|YF�GT�b��T!21��[�� 1+V���-�MT�f楬�q���P�<��dV��U���)"$�P�D���IM/���G����(d�O�B����*f�y�#3���Z]�5Ei�+�:3����w@.��ں\�qGf�~Od��WT�����q�^�T��y��K�e(��\��s�\�*��s|G�H
��������Le�+�����H��+#yF��<�O_s����s�A�X�7����/�M�K�(烅i/����93I��\��^���
��Ѐ������YUn�����P,I�G��w&c3DRT� �F8T�t�+��ZW�� T��S(h�W4�3�)�낰W7��/+_>��:���϶����`�+��nb6�6�����n��N
�	�Y�S��I{q/��`����]�'�1�22�kL�t�@9��2S_@&���Yt`1��R�M��ڪT����h��X���YoȺ���;DP���k����'����k�8wEªn�5]("R)�g�"�W��RRܠ@T�h�B%�ޠo:�� h�	:��@y���+~�k"�M)�,Je~��(���Hiv���lك��6{�i�[0�Qt���HY�HCbQk��y�kp�M|f���?���#��|���Vq��Tn���+lڞ���ͨ��B ��	��{���~ G}X�Ǥ4���h��0����u�CfO��RQV/������%�v�hoW676�ߕ;�ޖ{�w$���xk��%��r����nfP��㡔*5.��?R!|I�ׄU�}�"dW[���c s�+(��p��p4H�����y�R���d���r��o��7���,��
�?���Ty�-ǻ;R�k�����f�8��>HM7?D�&�'�x3�bu�dx��37�Ĕ&0w�a$�ҠqY?��F�����5�gu�/]Z���ݖ{��=�)��~�D����dg���ٹ�j0��7�!ք}�B���Af�|�Z�4��h:����3��5fg�B�I-ͩuH^��;�'�I�2���c�R�R?�	�6�s)��l`9�����j��̮��1׻��2��G���hK6��NGң����Q(�!�&��R����h�Pޛ��׻c���߹�@szPOG��du��{�w>���k�5UCRE�PbLiɯ�)Յ��#e��͕��h�^"�=@Y�;]��.=��ŕ9��k���&�$h�% h[F}iZ�u����Ж9�&�Wţ) dE��>�:��4���T�p�TШ&��>���0�G��НVe�٫�����Qa��w�-[�ڨ�}n�d&p=#�{"6���5р�WN�� ��}�B�7C�����P�9l��E��P��>M�`�bz�)%X#������MzT$�sSj�	R�X)�4���?�3jՑU���Fif���ٜ�P�O�SU��J>Tu�"xyƐ�����y��)��YY_����i��iFמ١��^��9zk���^�m�$+zo�T�%(H1Hr��B^�\2�� ��7�.�U?��Qql我����=Nb%��T&����H��P\X h��D�\�U�!3���_��h�Χo����J������W�7� N��M���w�4����&�"�j��d2�A�/_�@u���g�M���ZV8�����+���F�4ƺW~�^�_�9�����OD-���}�;�sОm���H��o��mP��䕫��N�];sj�{���f�=R��:���o4�d�;\l���үE�8��[�2�M�%2Jq��,K�j�8�R1�U6�12UJ�)�D�|�ϥ#`��p�@K���'q��s�"��чa��CL#YSS�a0~4�x�[����XA�
H�ё��v�\V�࣍�
7ff�0�1Qi4e��ZN��&�Yy��PUHx�*ciY��@-�O�S��������� i��3sX\?����>�@�}#WDE>��3���⪜|�V���q�����}*����φn�\	M9x��edrK%H�~_ �A����.�%�����&ٔr~��4��w�y��*J�ǰ"�j��x�
B6pR
�QC�YG�\��Xfi������'OЕ���I�VRgӌkiGo�@KY7<�'�eS΍��~��m��T�+-�9�yԍ���L���΍z2�1Q������i�`4� ��MV�59!�?��w�}���qc���,�c��ZI
��Ч�cRWR��}Ս�W�?�$f�&Q
F�(G����cp��[����.^X��/��k��~j�3T�CYƸ�j� @�ajF2��G�IP�����rQ4�{u��+�4Xp�^��j =b.D����ٺơ�ݕG��u�H��G�@�&��&cm����l_GApF;�� ��� ���sH�9̠f{�i�C��X���=*�{��dm�km�N]�L����u�x~���3�%<�����6N͝ù��Ѽx��@q��͍��}�:Z���@*���J��j9:�Zq=Ǔ����|���F�1�FF���
��Xd�k���*���u��Ҫl�8�?E��U��C�JDk��I��;=����f3.��k��d8���E����{j�ȹ��^+`�K��4X�eNWX/$��c�8֊u�ɂBٗ{���{u����D&����h��V�=�<kU"���j���>h�����	���SGJ���k߷�@�F�"����tH��g(���c�*���J��dB���سJcD���g�ӑ��|������ׅ�����笚�UL9g���ˠ����`J]G������0M����A���oBg{e����h��?(��VE�,�`��Q|�M�s�l�:�-��OVl�w�Bl� �ʇVߘg��M]���/�w��dZ9�]v_�1����tB�	.��9q3�
��x0��A�HSB�i��o��mP���U�U�Z��W�eٰ�
P[ݑX�<�C�hC_<�3�Nی��S���@K5��t����rB}��k�z�F�d@ِ��@i�qD�J�툒�4��Cf���{=̝kb��办�)�\� �⾀��^sgN�ԛo`��q|U��t1�����r��~t���,�:��~��x����O�wd�-�>;�`��^�U%���D��׫�wW�B%f^�4�K��U��S%�����w�ݻ�� ����+������|�6�=V0������'���`��I=��{�z����\I]a��������QeHn6��h��`�+�T*q�@�v�(�n
ڐ.$�&GyO� CH���lV_y�$ *��!X\0�!Md��/.��K/aW�o��	hz7�[3�x��M��s�p,�z(s"�"+J#ve�aIa{�p��I�{���������p�>ؑq �XB��P���0BG>?\<���z�wniY$��|�h������l:;��p�zݶ6cS�ʟ��+�*%�6v�):���}�_7!�)1�w 0S�o4�
�� ���}��bJ��*r��p��K�=��g�	8��0()�sϼ�]x�w��i"d�����{�/�B��H\��*�H��R�˅j��w>#\�I<�!4�Ax��i����c|(���
|����^pT�8kR�ה6v��x4(Ȃ�L;��o�sz�����W�)�Ĳ�y���1лy�Ǐp��Y��!e���}{�3�u63�
�|~^>\������w�}�t{��5����ׁ���l'�~~�5p�{4P�L�G��i5>l���O�N�!h�E/9�����/����CJFf&Ğ���5�3q�s��ܣ��n�.��j.][�(�j�'��оJXf��L59Ѳ����2p4�dV�	RZ؇Y�?�=?�}\������Q�<�~��	�mY� 哕*�U9���:�o��!Rk0�2�`��d{t�# �U���=�4���l�.u<�L�J�A�>xkR��.1gnO�kN��]�$+�����R�в �gCjnʙb�w8/T�68"�I6��'΄?<�����m.@�>�t��Xf�e���r��ZXּm�as0K8�������B�4'�~�oA�?]�]��$�әڡ)��Ezf�GIo_rf30��ʙj����]�ǌ�����#�� >�Ҫ��Km6>�L��e	 ��t3ח�ܳ�u�hs�a���0UP<��zE��^��\^�!y-�˥|�Q+ap�7M�ĔMT)���7�����6�$���Ny��ɏDh�X��f�Ps�U�01.�.N�l(���H>)�����'8��ǧ�}�ŋ�b��p��e,���I��0�x��F��E<��b����3����_���ϯ���MF42�?�T����4�W�z?��� �O�.����)���J���i�dU���)7�w��_i.�2�B�@%N�QN}T�)�R���>z�m����f]��B^}�O�����В�3[W�i`f�����|�>��������T�MW�����C�+�s�Dd'�I�9����p/�ЗQ�����V��>B=Ob+�31�ך(O~(�c������b��׀�'L�T6���G���y�O��韢-�f�ѐ�*�Ž�<�k򜘜	�U����08`@`� Φ@�"���Y3�
{�CyYߊ|�/c��k�q�~5���D��_BC,,�}Ʋ�A�\�m������ѓ�H���&�@�S�#�Wd�c�j�<3�̎�MU{SX��R�>���i�3G��J��L�w����7�����l�Ke~I����॒Wy����WZ�?!�, W��{wn���Pu0S-aF�Լhb�+��ЋD�VQ
�)�g��/u�M�I�|G�_W�o���R7�T�u�ǚ�=
�����k2���55Mom��ٻ�<uS�D��uR��Q���i�ڒ��	����9-�!���oFDZ��'�1��'io+�]�^kEd��d��]���+/�y��Jܺ���|}�.�O����Qk�V�DjJN
jr<�#Y@�J��*����[���4�O��J�t��ޡ�
s�� �0`�{�2��,{�Y�ɜ��&�<���d�u�1����z�|���i���gy��O5!�]��h\p�|�2�S֛,DA�`�|͚Ӽ�R�Q���h)KEs&P�/��,G����6V����W�W���LmȦ)2z�D&Ӫ��XgN-<6Z�fs'�o��u�E|>Ӧ�$��8�o��Ձ�K�����A�4��$��{r��6�hE������{&��5��)�h�~zˏ}فB|3���= ��z-tO=RE����+X _bRD��U��\&}
���V�y�3-��� ��4��@������a8lP>�:lg�7�^&��ӾC��oUJ$�v�O��D�R���hϰ��?��JA*��:����Y�	)h��#�jp���Z��O5�1�����'��^�Ȥ�:���׷A�?��(�4�$=])�l|�,�����J��	Y$LU��i�>�����-��lI�K�Q_�ۨGal.��rg#18����.��Z��T,�3��Cl=���~���^��s�6��r���r�g��h.�) �r���'�q��ctڪ⨽���g�4�47�!��u�*���eC��~o��%���GL�TrÛ3(/�c��A{k��}�EUSޗCޓ�4���L��ݍ7��k��_~�E���[�Ū ���n��ٗ����\���q��0�>QPFID.�<��U��&:94�j�u�X8e�@ h��u��� O%��V%�H��8�n�.ʪ���<*�Y?y��\�:'�#���!:ۛ����D���a��9TN���0�����kױ'�C<l�x���%*�"���u���k¥jLr���Yua��YJ/VzP>)n�9uЖ;�5SVV�r�8�>#�G�����h{��>��ь'sh�ٓZ�/�͢rI���.zw�c�t_��g�̶� 7���|��`w����	�&��VV������������z�� @>l�s��JS掄l�o��������
ν�`u����`���_��G�Ⓩ�Vs4�fFl��L��(�H��&P"�)c*5.5���zV�"��!�9k��>�*J肆	���݇�Y�2�P�O�O�`�\U/ݳ�Ws`�i�Z�=���[a���;ͦ9,G ��ʙ�V��D��Ν�W-�����'�cW�)�(|��<^���d.�q��K(,�hm�-kb����X%�}�9��0�)c�
P�e��$�#�烎�3C
ܟԁ?e�q��-���2�+��<3���cU%qj%�D�a���g�����T$W�q�o�֒���g(�k~FMb�=`Г(�!�g!c�z=bR�>v=�=5�Z��2[��,�BQχ��^�a~��:��}�B�a��4�H0��&�� �8��B�jόTQ&7H?r�U��"
�g��K�Fsb��=u:�Z�u��i����2Q{������XPg\�x%�<p~M�93�BF����1Ub���3��yѩ8ȫl-ߊX\��h���R�r>]C�}$��=���u�٤s��5Q�f�Z<|S�a����؟�u���:	��?R%���z(t=��2�G}��T ��}�}��oЅ�~�벨��LC6�R���L(����XOz�i���G�3��k��o�%S*U껂����G�7V�Knr^X5"e��<V&�i����G?
�?��
�}��_2)�nΌǣ5|�~_7z��z ��M˗���*e(�2Wj:Ua��:�y�������9+2#��ƣ<b �U �?{
�0E��Čg|����3jPd+�Z�< +�"z�}<|t��E4r��i"a	k/�*?3�p�P��F���^K�$���BK�2|9h�+�K{,k���Utw����ԑS��t5��(�$fA��D����?{/��-�����_�Hu� U�nՙ
b �^��TG[Ʋ��w���=��^Gsv�������$�ٓ�bF�`g��W���A��=�ȡ�
��@`Y��M=�=����au"���wG��9�
���'O�wL(���6�:+AY�&,a�� ��j�B����΃�x�ݟ��obr�������2b9���;8��ۺy�N���$:F=DT�`F���p�Z�^����I�\��0�����9ϛj�S��T~�������28̔��T, �<~��Ͼ����o�o��NM�{vK�_Ƴo� ՕY�8��d��I�e�cm����۟�	P�k�<�Xt#~f��|���A[�)$�p�M�0ľ ,f��"��1��e5����W8��s|u�w�b|�$�Q��?���)��2�%��w1�d��1W��41������M���"X��%�B'?L�?���v{T)��&��$c��pUB�<Z@�s�t��T��4{m2=���:C�uU�ٌ����PRӋ�V:=w���H1:E�*�<JG�)]����/\���(�PUd���s�Z�w���h�,k�/J8u�4*��e�ؒOھ�� �����"_ҜB<��p�"��@RG#Pe'Gu��'4EJ���
j���ԈH� �Q�h0��l'��UTr����I����dW�q`��u*�ʹw�rE̾�	U��R�ѕ���O� �X��2���I�I�d�'{�(���#��y̖�'56��Cϐ�ZD(��@���T����q�AŰ:�H����4�	���5�b/@H3�H@�y�^���43Lڔ�)�C�H0�q(�J��g
��dU'��h���%.����gZh����k��\�b&-��0Ha�H�i�g7i�B�bU�ؚ_���5��c���bG�s�>�s�=�R&
�]C9{X�VWlW�5��;N���ϙv%�_��C�c!(j߆���A��>�Qq����{9�@p�w�iC���AfSrAA��Z�����;��qY%,� �	�!�$�oKL�Lˌ��E(����St:�� �˦�ї�${�~��K�0B�dMI�K�W�ed�[�Qj�C�:�	�Լ#����`��"�ⴀ~��C��o��mP���-�q���wO7�p��#3=�`9N�n"���mF��m�MA��P�C*A�F��㠀�6GJ���F�ȝA^ �ܐ����㐥?��xE]�yu���x8~�.�p^�:�g�>3�O���%�|c�R��r��i�TB�9����Ytd,u�Չ�e���{R�`�5@;�2R/x�%X�%8�I�1��@���\�n���8�/�&f��[B1-��"���=�Gi�>��43���QO60:~V��o`�aO��5�f43�r�6P�G�kw�I�y1W�{gN�@O ���'(�vQ���X�}��%�����</�jDE�|9.�m<l�cS�~3�cšLyP>�q�����JuzXȳ�ð�����Q��'��I�p��]C6���΍�q��ečYK�
�1s�2<Rߗò+ �/mI��n�4n��F
�&����%y�6�`Rc������V&Od�[2W�rP�A,׵oKP|�>ￏP��Ʈ�Z��9<.�����qn�u���mC��OZ]���2V2d�T�&	��d�T��o����À&[�
������3�aD����;�1s�תDq� �"by6�����oa���o���6v�����˘�t�k�_^�b$s��no=�ߥ!��`G#�):^��|����l13���8J��_j|q��M�ǜnYP��4�Jj��9Ϊ<dl��Kr�,�C3��J�j!e��#s�����yL��$81m�S�tϕفiF�"��R�2��;QD_�Scyg�P�U%��[3yL��<�P�s�Wg��F8ɣ2��SC4����+�+�m�	��3��{�?�UF�kF�0��Ǜ	V��8�\Hd������7Ǳ�S�6��e5�*Wd̺v'��<��	!�r����R�ݼ��|]@t�4��=Y*���/-����#-WTԇ��l4�
+��yl�#SQR<U��}Q}�(������A47���<z�	lgd4ٓ2 �j�Q�/�_Mѽs�{;�vQ	�����ߥ-��1�걳�/"Z\�'{դ-�h�)
�[2��9?��s'P������YH

^��pH=1U�6)����6�'�C�L��{f���zF�`�d�2��9>td��Z��Y��}g/���l�V9K�f31`냓t(ASW;�������UY��ƨ`z�f4��9�y7ʌyL8}^�O��Fz_�:��He����J�7pA(��	��@浽?=��G���0P�z��cs
�m����e�a�̡���56b��햶��k>���Uc2CC���4������
\�,`	��'p�V��}׳F�0������P�ʔ/N=��L������r��%�iN4�u�j��<�b�*N��s	T:ڳ݃ϝ�Ӊ��*����Hh�+�g��r��o+߾�[���p0���w��]�~w��L˗1J}�)}��L��'N>.���앂�8�+��oOlS�j`�1T�aV�b5�I|+k�$:Jl�i�fN���Gy��Μ����:^z�$B;}ٲ���	(5���ڨ:N�i��8W���u��,��?��KEt����pS��9�`}�\��G��}�X��
��lJ�hS�A@WS@o���x�V��l�%����3�!���s<h���ʋqT#�Г�I@\���[�l�؅ek�I(T�Mо^}���>�9x�@��}�PQz��|�s�̜Y�W�z}����<n�c{Ї���l��C�	0�X	ey�JX��S=}�"�����>�`龀�����}e� ���m��_!�[��7����ɿ©�4W��� �ږC�c�V�	b� H�Xy�m��h+��b���3s:O=�43�Ǎ�P��Bd�俗f���K����H�6<���}������XԠ+�g�������#�h��I�񨇧��
�&�5k5�K����@/nрM@Y��D��G�{&�I�qUPʩ>�D~ �$JPi��x�3�p��gq��A�z2I/�Ӎ'tP� ��l��\@n�Po��{��y���&EI�NzXL�E�)$�
U�ߪ�@vM�SP"�3�wUm#�i�� %��=�"��f&�Y3J��h�)3��n�kco�����!L%H��i���̣�Z���4��&�AUF�Go���<ݻd���-�#b̓ab��M��2�3�;��z�m�X�U0�����%9NtYW��M���q�KrS/f�Y`vp ߛ�=c(�x�Zٌ�>f���(W
�L&T�����jP�oQ��j�K�"�I�i����Dk<D�� -��<��t�T߈P��Js'N�:)b��Stw�U�8���ͬ;�1G�f�쁠p�N��'PY\��ٳ������M��eΗ䦺������N��Y�����ɺ�-�P.c��S|����{�J�{ {$e�C�ETd?~�{?��o|���U��>����ut?��;���n�߆����Ysq0m=d����F5�]��?�ڹŹ������e�0ȢK5�����2�I�h�*8�^�Y֬��Z!�Z��8V����g_���e����!i�No�w1m�u��/�ևk�v�I\���F]"rf��Λ鷡e���3h3�C��@�6{+m�s�H_��{��=��h1��c��|�e�l�2	a�ɿ��z=R�0Ȍ�T�ɽ�Q��N�9� �W
����S�� �s���d;{�4(5�c�ܼ?��a�(���by��;�Je�?�\�Aۃ<s5�`=c��P�����ѧ Z)�J�>�T�-�0&�T~�g_M��d
y���uh0�[|}��"+L�׿���������;7�a4��.��r~]F"�k&�/�Ɓ�%/�de��-VO7嬼��Nf�Gf��g~N���d��$��송|��L��Q*��p���r�D��p����:���#�U}����s�
JO�Q]B6cY�r�?Auq���l�U9s.��b�/�����u�ܾ��_\����0��.Ǉ\S��)�|�8���(�8�|��?a�ݣM�6����ҫ���nc��{�����h`FQ�:l��^U�U��!�3hը����Y9���5}�\o�#cF�>�\�%pRG"k���e�����v�)��N����*��RjjMjql*�49���q�)�Ʌl�-�/�̲�ng��� ���aNM�":5S2��)|r���Ob��%`n��LuB�j�3��0 �R=�o�7���i4���8�~�h(�͙r|-�-�߃�ed�e�A[*�jf8�lY,j���)�x�ɵ�W�����`A5�% �z��xHJ���	�r���T5�K2���U�E#��� @-r�����k�h���
�l�w����
{� ���".�6�w�.�ܼl=��̵�����/��Ԁ�m���1#s�A9ǅf�Ȥ8�J���˓���l��(
h<m�TB��<u�u^fU���i��o�s�ʹ��#�����SY��!�-c��I���:3ڣ�@�T0�_�[V�*j3����w\�/+M��c�Y!�]�_����)+=����^��E��y	�+�-�}	 �s�n�AE�r�"�<Ԇ�L'�K���D�]��&Z!%h�S��2�t4�q�{��Q��C��"�OiOL�X����1�_E��':�k���3�h��ۜ��O��������8�D��	,�.`,s��ga�Ț�XCe}/���׊1����vQ��� wS�����\r��k%\��q��ױx�j5ɒ�e]�1Wk`�O��X��?��Be�/���v�SǑ_^­?�ֽ��u1�~
�_�N��G(?��l:%8��eqF�kf%p��#A�����.k�}yE�U� ���p�k��~���������_Ө8R�f��T2��[��k�3i���w0���D�3:5�Y��z�Zc�Q�b"��>!��.�M}��Z�Ɍ�#I�R��q�d�3@�s�+���V�S	pΫ��M���b%��>Lq��e�C盐s ; Uo��dE	��r����zV�`U#�	�-SOKgL{a,���o��`d~�]�2���IL��<m�>��һ,�80���5s{�A�T)��Q� /V5C_�,5=��ߡr��e2Q�>�h�`�zNkd��j4v-�q��I�K@�¤X�.��1�^L� �W�W�U�΃z�@��\XQ���+Xw�[�A�]B5���V}���o�5�z���w������K�|��w�<[Wz	]m�Y?v�M�u4K�Q�ag�n�I��l�"�Ċu�
�5��{+��T� �]6�	A��r,��S$T	�ey6�R���>�x���P+qR6j2�{cl޹�����o��ƚ�[Y���38����,�#9_eJ�ZH�}�������#t���w� �&Z�P~��ʡ׵�,eW�1�����S�]�w���;��$AǢ��^�w|�H��&���j�r`j*p��Ī�B����P��#r����4gUk��'/�3,��]��ڏ�c��scF��F�I�S�m>�S	�X��!1��&Me����p�����k����%���-�T�3cH�"UP�9�3�K���Y,�Y0b0�Tj5(�T�4�h@.��ԥ��kU�ޡ����-�f�ٞj�6�h��F�wi.K�ͧ�,��g9�Y�BQp�H�v�*q��e(6¶�w��?��K����-�M��t	��=f>:�J �FZ-b��*μ��� �ZQ�Q[��~g���T��n�fJ>*̴���z�R�<�JU�#Y�D+o�RWd\s�߶�7���ڀ����G����-�	(9�̳X:y��f�N�,׽��G}e�S��A��޽�{�|���S$w��B�o��D���3lM�Y��2l�v<`�{�9C2m�3��o.�����_Ѓ2J�e���ڵOU1���a7`�AAhT�1+OA#)Y���� >�����9�����+u9��e���X6�؄�o`t��%��*�+h�:���QZX��]���.�{кv#[<�B��A^�� 1���X��*�<6|�52���D�9�������s8&{G��	`^��|E�P�u���$��z~f^��̫�y�r�UL�DG@�ñ�"�W�c���ӗϡX�b��]��o�>FO�p��Q�@�̡cg�����}���c8�B�즯��
0{�,�%0]�?
2{]�(ȵ��@{83����޵��� ]�i�E���V�ܕ+���_C��W�7�������W��c���LzH�m�x��k���pa	�7��P�{��k(o��e��*�t�O9��4�]6_�v�fe<��l����ژCAn����H�y�N��k،H,��U�Ly������kW�����G�]��H�*��P6X�m�M��%�U���{R����צ��9e�x6��9��)�6�V�`"�	��������ԇ����L1_�+ �K�#�Þ��Z�[�F 8�I��.,�"�e�W�]�����@<����V���+�����r�qA{�rǉ�V�%(�)$)ʁR��c���2� �>O�W� M�����J�>��(�7�o�=��L'w�3Z=@xo��?H�LC=�,�a�ewFǠ�����o_��W�nU?��_�������~�N��R�i��i������� �bU����A�/h��x�f6��	��M����9��4�Aʐq����!�r,����%�kT���TUY��,#�4�lˆ�������{��-���Ê�"��zqq��#yx;���]	�'��P"��|��̱�j恣a;��߸�	��6\X�����q���`a�O�� �Mm�<����}�o�C�٥J5nFv��O�����?4~/���g�8w3� i�S����N�����ZFZ�w���̷l�VK�w�|j��^ِH��>
̐�m�u�F�����|޹�R��t���lC�zN��ДgC�~3����}9��s3��=��3gp^�� ɱ$�x��rɌ�����K5v�k2e�#�A�΄}]�vGJ13�N��S�\/U59�qj�����|}V��[��@��6�Q-ַ&�"�e�|����/�-���Ybg0O0��hwG�Wϟ���x����Fe����M�3�H��΀n4@0�+��ቝQ޷���|nRL�����R���F���-`Bʜ�~�%�iE���.�{\��X� A���Kk8�r>��O7�a���'��S��^r�H!vCX$u�B��Ϯ�4+�'�f��If��0��եK�G9Y�@X +Z�&u�Ë��a?�8����D�� }y�Qn�aޔ�b��������N/����]��%if4�(�r�;�̡�A�L(本���r�Á5��KǱ|���.+�\����H����/ѽqY[2���Fi,����Z��-;j��2n�S��>����>QP劘	�/#���k��dM�}(s]@c3D��i�nʫ��[ac�?�do��-�k��R�,Č �'�w%H_�#W�Â������O���>��ұSC�tn�%�`�O�O{��h2Խ���S��2������B_�#��9�������p�^yU>��NZ�AS����qCx��v��1� �`m�U�����I�������!�9��{�>n���|�'N�vB�^n T#*7��ʭg2)�@�c�Dj>u��n�d��pԲ���y[=3���������q0N���d���ޒ�ɜ��̠��eg�q�XC�
vl)���z��&J`H
����U�1F �G���88��Ol�ss����k#�$'{+�BQ`M��
L���J�g�fD�2I���P�@'������Y�2���Lrٮ�e�0W�#��Y�_�U�ZP�D���zPOjh��)�ђ��M�R�f`�=��|�7�$��V[������"	��Iֆ��wmD#�vDwi�T@®�z��S�J}j�'H]U2�t5#��5*H���5�����@��Vh�GQ�O����Y��j�s��ʪM�_���_���.�����O����'����@G��\��&NNF�I8m��t��Im˲�moj��9�6�$�s�Y%�@7Ir�!JX]�l�ƖM�ݐ��( =N���{���P)1��v=��Ȃ�ª���³����_��7_��ꊑ�=����x��{�޽�pe�,@�h'���!��y���������h���BI@CМ�����W_F��B�Xj�����������A��6�Ȝ3Pf�y��(2���( h��S.c��,}�G�3/X�cP0�|6�i�!�:h{*_#�zw�����Bf��f˕�=03���@@wm�o��i���},`q�cҲ��<�<9�1���:>�9���wZ�X<}
ge,@YR�{(��!��|q"{f�s&aK�Tr��n�����hSl�����'JqJ�WYRu*����M�01���X+O5�h4���c<��g�O�Tv���-�߾���}��N	�o
�XZ���w�J�:VWN �Oj��J/=z�m��k���iC+Yߚ�C����w���d�M�<�%�� �raj�ee~���1��D{"\��_�S���"�����1�ZZ���K�f�c��]:A<J���kw�CzK��y����$M�=��t���b�����4���*5̂�9g~����8�9Me�t>�����(�^è^�~/���=E�E�뤣k%�X�?���0��F��=�
�*���UzH���V)�i5����3P�-�J9F�ׅ�n���f6�&��5�7P^;����TOK������mtw�л�ݧ[jX��W��U�|���������)0��g���(�T��Y2�c���~	�����^�@o^>;��dw��z�xz�c���ȘH���� �5���O>��7���Esf�\����e<�~�G�-k�ŉg^D�^G}yQ��N����2.]~E���K/�g$�ە�T��NX}����Đy��~��E����{���߾�����P���O~�3�'��̠P�`vyY ��E�;mLn����)��q�7$��]<��D�Ξ�=b���~�.~���%��������&,k3ט�}Y��U�&���h�2I�fc�}��e��b-�{��է��gc�һ��z�h���T�ȼS �R[˖�N5��5bҚ�z�򝞽�?��8�JP�1I�:W�BӤ���t=
�
�=u��L��L	ɌC�w�{��m[�3%Û..���h{��>���^Ro�dk%A�^����2����g�L�l�<s�v�.�-.8�����d�7���T��+�U]��4�6��l_�x_SH2���&1�� ���o=4Pޘ�,2rB4���D���'}4%x��{Pқ1|�^*g��;�W߷Fh��Y�G�]�2�j<����̿�3� �1d����Ƀ�	�e��J{�o%HI��j�yXC�m��
�����O������������/_j����Iu/�K2os������X�A�YD��s�����+�gA�V2�q8qus-��f��]�ŪR;Phf8! �NN_3�\��ڌ��xˍZ3��2f���̋/���!.��r+sH�C��x��G����xr�#x�9�c��Aە�*�,)q�=�Q�w�JE�w����������k/a��Wq��E�U�;�������&���66�s�O�b�+�'�V	H��vˢ����B"u�̑�h/@e �GG �֞l���̌�6��h�P��OT6��e��z��ob8h�&���~��(R7�:�$(�k��'Ǐ�r H8�j��� �FTD�MNlT.�O��PRCt��4��a!��`h��N?1Ы5�0p�YhN�2�� ����]t��$ڮ�[Vz4R�廳����'����Q6s��^G����BQ��Z�D�V,X�Uh���>�J=�ΛＣ��sgOj�j#�9?���\۸�,�p��ݧ��0�~��w0�Փ�,	 �\�P�Gl�d��	V����ǔY�&U�j�6�v��^ʿ��&:�曚�̕|�T�\���X;qZ]���é)ER�$��_>���3�w����B���O��l�%��G�J=�e]#!)��m�J%at&'{��C���.9��u�/����(.͡H�J挬��̗J"�A� 1�k��h�E!��0
Y���Sϵ%g�q����HR8���DךA�k�8�e�%��P�t͋� �֌�/��/ {�7�y�GErlY�	r�M�jI���ܟ�d�VȜ}S��82�׆W��N�>�@�t�.����1������7���;���{o��������:�IY����ƶ��	n�9��!�޺�� �����"?�%�U+>����R�y�;�?q
'_xCƣ,�P�ʬ�c�|����`(�3�S��	�,��<@ɟc�T@����_���Euc_�$svW�Ljo����J�z|�H t�������Er�;�螘E��2p�"Αni�T@�C|�����_�����X>������d���V�X!�s,��.G��B0��4i�i�p4����x����6yFF��c���ٗБ���?�xi���J5�o*�QE��ʂ�L�CKi��L���H~n[Βk�Qd?�Ӽ�T�x�.X�3�>�Ukb����G�y��gs�SZ��*��IK#��I���^1\и���t0�qak_��H�hLn� S�g�^B&�\o��e�ͪ2�[�2��)�Ů�ܾ����ֻ�aS22q���T�
�� ��@$��\�%�K��b_���&z�ǈ�����p(���]�7���1�#�=+��73p>�T!ϋ-�"h�@Y�ЁEwҤP2��q�����i��H��$Lt���c��]��P1��xVp8&e٧�T���o��o_�����w���|��ΙwߘѬ)W�/��Y��e�����Yi6{e%��u�s��A8-}�&�f���	�2������&j�j��epC��h6Gu�KU�pW~�xQ�yzQ ��,ށ����-���bD���99���C�N��������f)٤J]n-;�elt<��-�V
�y�j@�'=�*�{��0��6�=��~c���M�ӧ@��f�(�3�FK2��	�F�23*�?�����mt��k�CCJ���U��R�T�.��%�Z�WQ��~ږ��9/��U��o��r6�'��GLu��� �MV���Lf�E,���ߩ*�3�	h��/�?������}9(��_EW6�����\L:=[]�,./I��,�����N��ڥ�D��8d�{�o���Τi��<Xx���(�W�T��C��\���pt3���51zwZ6{M��&��̯}�	~q�β���0)Tq�����
f%�d����{ػs��o���)o�@�A;tVyQy_��D�}y -@ҿ��hΖs�@�h42�� ��� g*�p�S?;1���?h#,T�H�s��gNc�7p��?��w^%�O�YO��S��l��eu॒���6�~������|��6`jK״�XQ?>1�7ucu�!�.E��fv5P�@9�G��L�q�Or�w	�v�l<���yYK���BO�RM�YҌ�s�^��{��²�2�$�ے5R�:��J C�À�jf���D���fV�2p�oUQё�^��9��J��|�Q�pa+�
�N�N��k�	@��i�L+��j����%=K����.�|(���}�zW�I݈����
#�U�+1]��ϱ�'5#�,0Y����er�����������o~���y�>y��2.���Զ�Ĥ���� ���̧;Kװ����2R��r(�9Ľ�W�ٙ��z�<ϝÏ�u�N�����0�?����k��>/�4�pN����G���e�1ӭ	�%vZx��W>�BI�6�'�*���Qj��ɸ��;��ӿ�%��Շ8- ����c�=����Y���7�p�F�mm�Wo����%�իh�3k��UǷ�W:"�SJMu�O�J�%�t��y1夨� �k�W��a��1W���s�������O"ϷY����j���,�ƚ�J�/!���*�U�8��*����l���=ET��8�嬱�O�l)����]53��J��:�Vig��/���y�љ�C�7t���E^{Aױ��!-U2��$�pZ�}�)@�Pp��D�Q�}u�cZQQ�s��9�r�z1(b�]�x͔�^�H� ��<[�~�f�pJ�p��Y���v!�Sf`��n�12
�����Xྷs��#�^rV�#�2~[^�۲֯�6QZ���˗eKh`�����I�/�d��;
&ߚ:��t�~ļV'�R ��iz p�J���.YQ�F(ș���I���l����W��ԭ�Yc�o��mP�O�5��|.�Tl��%5�?��@&�����LR�R���wg�L���9ajrط��49��$�V3�)'p�!�:O�w:q
4��"�DQ~��T(���FE�ѐ�(�y��[����W�ƿ�Wx�_�1<Y�c��l�tNf�����k���+��(��ऩ� �]�?������[������(V�߱l(�A�2���_;u
����ܫ�cf�����c9`�����~��6�
����ϰ{�K0�V+X���-;O���X�����(�U�}$�F�1�r��"�-ƂS摯��{x��	Fݾ�j��f>iF�����}����H�0�X����05�,X�l�VM`&K��|�)�>#�7�ɛ�	�-T���\�+`h��E�Y3rno�Ý	�*9}�E�]��Mtfgp{��NQ6�j�AO���'��}	p��9�R+Fa����ڰN	U��WI�|�G��3��{��1�|��4�^W��a>b�G��W$_g�F�����ǹ_� e����jE@�m������"weN<x��`G>+��|],=u��>�6��n�ӍQI����)^��ό�gZ��kޓ91  �L�jKy*qi&/�¥+x���XK���9͖v�p��g��;��ݽ=��pϾ�.��oqx�e,�9��������	@��A�|f�;h�͚��(���\�p����~T(̤�s�,Lk�S����}G�n����6��/�}&����Kؗh����^Ǳ�Ǖ�������w�	ߔ@�3a���[�]�e�9B�AE����RƮ���S�9ԁeb������I@�p��nϤ���N��*�%P� g����Du�
��sV1a�U���u���&���ng�,72�5�����*m �U+X�L��ͻj�&@�ݑ@����2F�'d-08x���_]œ�wPu��
�1!�;'�<jw�c���\�ҳ2g38��4۸�ŗ���ULdN��J�8�
�8X���l��y4�����&�Y�5�����&{�����T�j�O���	}V�gh4�o��S1�d���?I>SVY��
�6aw=F���噿\�{��� �R��;���GV`FX����r�3��
���GE�M�WJ��g��xz��Y9լy&���ip��3�+�U����4��i�4� BM���&�Y�}�&[��Lu��Q��\�/�P+�:������L�w�EV�ұ-r^r��3Q�������R�L�>1���%_Ɖ2����z�8�!/��yD��d���D4�}��BU�s�ld�]O������DIY�{�(kueԝ��@e��i���`���e���d�3��� M)Yݖ�7j'G��X?+�kʱ�:d�D�@�Q>խ�5'RU�$�����������B6����oYv6n���f9�J#�u�q��܌�c�7ѕ��v�4���������Շ�V��Y�^���3���	T�U�D�R>d��X��(�1�86�d[ �W��Ƒ5�1��2R���d�����X�"��f�R�G�ɷA�����_iz��o��?���[J��b��m��D���93�O�¤!L��M訄���q3(��R����h��ff2��Y'_�rr,�ժ(q����(	�܇��Tfp��eY�W୬j�q��1���P��3�n�T:a։F-� ⥏1��@~>�61[��5M� X<q�_y�_z��|hT���������d����q�+XX��_|	K�*f*|Y}��!���T%����gJ�,��Ų�G�N5�8��E�=s	s�m:����q������Ҁ���<��&�-(�j��}�T��Q����x��M��{�^�'A�٬�2ֳ��r0��:V�|��)0�эa��}	:L���:����9�
������
eR��$��r(����-aN~&���ĪJ[��Nq��$������$����Yi1#}{ط�D5��f��>��e]����b,���k��<����㟢�������d�����u�2��q^�o��޺���#��m���%@�|i��Aa�?U�� }>��2�Y&��7�L^3�M͠y#��X��%�|ᐺ�
�<���=uR@� �o\ǭ�>��?�~���n|��o�ď���o� �cK��2dnl���Z��Q�3/�ˑv��A3R\A�z
<k8gՀ �k��i�4(����P!��X�Nw�`'y�%���Q��y���xS�d���h����k�|�Ǎ�x��ה[�����O7�bN�� �1��d�FC3o
&2�B�2
�2�Uih�Y[<\�M[�7����b�/X�LmU���΃\`���_�y�� �����>�K�-,b 㟛�=Xd���J��>����$qM�����	��M�T��g�4�c�:-��ϟ8���.]��&t�֏!�����u�XYT�ݵ��q�³���?�-��.<�2�3Mr�3s���5�êH$��o�����ﵔ6K 8�$�u&l���F����\�|E�*�U����I�=�8G��$H�u7����{%���L�g�e˞�xPā��TuS�h����,�2��z-�%�+�鱠�/￻�������m�ϲʱ�ћ��ʿ���K`i����0t�X�*�/=,��Gڌ�X�z$��,`�$��g�W��}Y��&��)	���C݆|k���{�V�ؓ%�X�)5(MJ��03�j�z�S-�	������G�Q=���0��9?��V�\}����[^��G_�.�4,��$�H���F�ZB�b_׽���fP �2��
�@��\�/��'6)��h?���(J@d�(���خ�@ǒ~A^2�@6gp[������bh����JY��Ƒ	���Q�g^>5z/P.VCH�����f*�I����H�� }I�nI�@�����Y� �1��&��g�7�����2�\���Z�6� 5�b=�K`$�8�
'+��B�f#�48�� ϋ�-��
�)���T�|�7��&����	�Sv:�~��=mR�,���f�h�@��Lj|CkH
]��[���O9��6�ꠚ�D6��S#HT:.Ԍ['���P�:i6��r``����,��x$���n�/4�h0P��}��94A�^�_��F��b"?�p�[���@�Ӥ�6��Ͻ����_�r�\��n]�'~�/>��o��ƣ9�Ͻx�	({��h�z�\�����[>ꨆ6�VJ�!DޡO�*M�A��\i��������U�5'AQ����aL�}�?r�+�(��Y-"���k<����ڂ�r�˸�p��N₭�Irp����r�5d#j
x`�nƲ�(?$�m��#����w��LF3���s8}�����K�]Dn��Ͻ����<���+8���Q9\�6	^$�
j��e#ޗ��u�G0L���܋�y_z��.�oBO�E�W���<ˆ��\����s�l�**��Jpue��KO�޵g_��G�d��]���;����!������[����W��Y�O, �y������Q�yD��.|o��x_�=s�Jr=4h���}�m�D�,_z�OM�xe>ӹ90��t<���*G2�2f�C9{�"�O���w�����v�5�`u��r��	��<g'���b���3ؚ`�M�O���Vj`��C��z�9?�0	&S�g�$���'j藫p��	�>y
5��ǀ`@��~k s,/�Y�f�Z���9���"�:�U�|P�i%�yU8�1׎*�yM���j�8ґf �J��8��q�Z��MQ%a}s^�Ha��P�1*�=����ͯ���ꔜMj��%�d���{�����e~�yY�����j��˲_,.̣ɀn���<� ����y��l὿��2.]:�K��곳�N��9�(s�8���a���l=������U�'࿽�X�]���*+F�wS���?���Z�cOAs�ڔ���|��9�4IR$ի,�AZ@c��=5�]_aT@�I43��`[O�j��97������re��Ĳ_��2�2O;2���j ����V���nc	�� �^��^�t��E�x�&�t��ӽ�JԎ���(�S�G���X�}\3o�:�3.zb�\�5������L��&5�L���L�Bj) ���wn�v�
0�����tFJ��sZ�L]�L.��SUۧI�	��}/5��` _�-(�3�S�!�ˈu^Z9��>����yz��o��������E�I|�n�r�i�$�%3 ݫ�Ne#�`!���\ߗ�'m�/�5�Dz�4&,��e3(�rK���OQ��.����$V�u,�i�3P�;�_��'��- H5 45�U�Y�aCCQ�I䩊"�1��?����7�G��.JssX.U��=w�|�%�����;u{R��	&>3�4_��>Y�K��CJ4}+4�UW<�bŪ
����a�`�-}���o�u�+���pUVت�9���0
F�*�E�Y��@l�9��Sա��L�45n�h42���L+>Qڐ��R�T@�E�p�N��Dr��p��}5��!"�U�J���VnlbA���`V 2�XY���j!(��5k�+]7C9����+��S�DF��2\��d��e�ɡEzj�yܿw�߼���;�:u�<�t�mu��w��}9���	^����-�ë�|�P-��e�syO �x�6I��D��#-�c��`s��3�FE7j̴�����H��.T��T�?�W�di��W�������j��g�gk���.�4�Q��|�3��D��HЈ%��;3;;�j����EU�V�3#C_�s��UH3�4 "̲��23���~��q���(#jX'U�xC�����場2g��6l�ݶEȦ��s�Yr氱~6��ۓ�m�����ԟo�ɽ���������@?޲�?�|{b	�Ņ������\A�Azo�\r�����I)�]��7P̈́�g�-�F���x��]�t�<�� �.!XP`�b[p2�k'�c˯��f�o~���/���}��6�����������m\��W���ן���g��s��{(Y���je�u����@?�������@:Bs'�ƞ�[jw�4OM����]H�þ��̦����:��]�~ծ�9	p�f����j$e�@X���7m�E��lׇP)sH�$N�f�Л�F�	�ٍ�5<� ��O/e���.���îh�jO�k��)��~�akg�ۅ�ޱ7�����i��tnre��[�\���nO�;�w �8�\R.��(��ِ����c9q�����501:��iI��}��k)E�Ď�:a�gOY��<�Q5K���<L�Yk^a�Op4������vs�C۸w�N.���`K���&J7����J^S�v�@�S�S�x��`�&�����ۜ��j��e{��&�����>�d����ll�����a��ܶ����[o���׬{��٩Sv�غ�g�X,���ܲ��?�����c[ƞ8��Kv�G؉�CU(����G �TJ��d�νa�������;sA����y|��p�����pj��������]�p�vl��<�3�bo-�����[|���1Q<��Y.t���k���e{��GV[[�9�g�q�����jX��I?>�W� �I?T�Ny�C��
��tl>�9V�k����iR�f{5�T��>xʳ�N��CU���)��}�,Q�,�1ؗn��>xQUb��᪗�}�VeH��S�Z���9��y.�.�(L%�	<�Ey�lc��gy�M)��6c�U>4��>��(P!�NK��,00P�n.���vy4�����L՚�Y8kL��w���5�R0@@p8� �,��iSI�E�|붌�k	���B�����9h�'�a�*=Q*���s�g�9�����|���("���W
�*iLfV65�/�8�{�뻶{�eñ]�R&�R�}@���ʊ
Fc
J�h�E�@�e�=iJ��Fd�(4�c��~����{6)@b&&D��ѶkS��_�!(���Ԓ�� ��|�`I��l�o^�La{�g t�	���ˊl�������;e6<Ѹ\���!n��R�8���K���-5�E�x����5*��F�.jʹgm��
&;3�ԙ��q �nw��F���(���8z��BK\X��ְ�cO�ʁ?T�`����q{�7�ʵ����2������Y�n- såY& �iea褫*��OÝ��o�-ğ���ND`s�7�"i�>��>�6��~��O���j��#���m��|�o��3��j�eJIOa~���)̂A#g���mD5[�1\jtuASt�6Ԫi���xfOG���$I'V~�������+�J#�F6y�`gl��%;���웯Ў;��C��-�>@����2�K�F Ě6ʊ{/�jj�����"M��-�Z�}�`�lVDb<ǜ%|�\,y��+m,�l�`� Ʒ�@��K��1\��~a�~��U���������m~�i���,Z���n��N X8a�NX��=.+�1��g���u>\_N��>��a#y�g�So�Ǡ��a�+��[���¢����� Nx���r��ʢ&�$�%k��H�6[��C�P�W�J+�-.��Wm���}J��FA�A��2����q&u�������
_$S�+=LD�&�Y���Nq�k�K�;}ή�����w���+�q�)hMHG�^�tɮ"P�`�<����OU��ت���q�}�^+t��P�6@����|6y�5� �XU�u�N�@LR	��33IjA�C�z+��:}��cӽ�M(QL��X�jf�5u�kmv]����" ���A��[�ͫ�F3c����|�ڬ<
�8g���m��l�Ɲ��<)_x�+ǎ�I�ϭ��,X9y�%[8s�p8���ڟ�����v�-?8��-{møi����Y*0*��Hݶ��m��k�n~e8���#%MUfN�X��X��F��B�惖���3�~,a;w����W�N�k�.�lk�����ߺ���\�:����I�N]:o�/]���~�&j6��m��
1��V�\���.]��ݺu��|���}�][C�q���aK���)�4/_>oQoIԌ�RϖؐD��{]f>m\�`���v*���p�(���fMesSe��o� ������uf��N�k��8#Я�ӧ%��!�~�!d�ѕ�����3��<T��̹�5��꜠\��VQ�J�hM
T*j�<�7���&ޘt�Ӣ��C�VÞ!����Ɯ�i���$z�ވ3T�	lK�'q�	e�I_��ge(Є��L&�L}��&� T�sZ��"��>��6�ݶN���3��+�.��V�F�#��vﾕ�}[��l���.�e�ٯq�ۑHG=�Ü"�銪��,�VOT���a��N�z$��U��U�ҦV�3Ld�k=������@��t�f'�?�5L���G�����.WSbrdX*0@7o�VE+	.�AR�6��
�����j����CQ�8c����l�������A���/�����Wr�5f�j�S��4��)��eP>���&.����K*N�7(F*�U�S��������/Aʝ���"=�1&o����恈4�)�H�	D�]Nd���s�Ʌ�88
���ܳpn�u �Ѿ��[0�8���0r�1y#^c�_ ���>w���-6G �h��4��J=��tlC����g�)n���y͌�L|�1��EM�@jM�6�M`<hH�0Ē*V�(^�6���X4 `}���������Ma����]{���������m�'��Q�m�S�׎/�)� _�4��9��E�+�0`��P����RO��@�፻0�Tb�3Cno���.�il[�f��'�X]}�M���>��p߾!��C;y�4 ���| 6d��3[>�j�g��[d5d��kx�U���>v�Zbϕ�� ��JT�����f��l����ab�9Ĵ�p�8��x��x�؝ʦ����M�՜�l�'�o\ڐ4��=�|�%�M񄻋vl��=)�I����S �T��+kUc�`�ٲ�P�i��0r&��N�&7�@`���R�6�!��j>�V����گ����l0q�W*�`�4C�Y4���7~rM�T����܉S6��Ȧ4)��Ӝ=�%PK� ��̩E��c�ʀ�d�:��(�O#H�����N^y�5�
`w��ҵ�-(��={l�
ė��h/]�?����o`{������k`�Z,�c��2<��;t�I$z�j����!��W��k�Z�t�Y>��UC=Tt�ފTk��<<�_`�~���DT#�3��X����-^�l?��?����WmA�vk6	���,�z� ����:UMe��#���׏pD������_"�[�����ŋ�ÿ���G�Z@Pw��v �)��+?�C�r�e+�m����68�KⷵΙ ��U%iYy����Ap��Ol+�����*��]-um���&�� `

F�Y��:zM���cK����mv����Ȯ^�d"N��9�Z�^�t �`ʗ�:a͓�������52���A��������7_~ h����ŧW��~`�^�(���9sB ��6��Ȝ�Ϭ}U�$���
�Uk�I�5�1�,k�L %c5@��C�x�R�����mz���u�s?#� I��%I�,P�@�/ͺZ�c��5�gc���뉃��!!)�8��f$���h�d����.�Ig��}k?�*�V	q�� ���=�=��c�tΞ�����|LA0+slp��
؀�
���	&�����d���Ή�T��0��}*~n6���>���A���^ηi���C�y��n~��}�ч����� �r�ɝ�+ ��� �i�bH�1��fd5�vτ;��T�{�%�@&�
��Jc>w'	M��f����]���sKK�U�9M��ʂ-�p?�����+����[�J���ޑ��Y���x�-uV}G�PR{m[��SL��%&@��=�AVHN��mQU1\����A��g����ç���j���/i���$<\�-T��T^�MK5A��^@GC�J?�89�z9�Rs����'2�ׂ�P��d[�B˰y
"9d�d��ю�@l�YJ�X���#�毇��`|����	�͆����m���-N�V�9p��M;���Kv�w�����8��Ifqˆ�"5�9��uL����&7*pD�4����S�y���\�^o�� ��d��,��)�F:��q�2��*�����M�$�Vl�WO_��_��gO7�η�T�lnX0�I��J�t�N�L3�J�X3k�0�������Y�م�Kk���:� (������߷]�C�fc�_��u�:a�%���% lf:q�{{{��7_��`ˎ_�`�X�U��޷�>��N]=k�k?½�,o��S�x�U�Y!�JBv�c��U��D��73�M�����}��3M���+�sK�W� �V�T�y֗,�^�'�l���$VS�t���3gl V���>��l���+�U�q��"��-?��b߼��cz9�fط))l�cbtX�L �Ӗ�b��<�Rz˖����
 Q�g��i��ݰ�ooZ�o��4i�gٰ���g��E=k�z Y=�3,ʱ6�����B;��KA��īW��I�q��O����.���ܽ��U���[_�k�k�?�@C����Ǐ��� �I�N�>k=�W���Ko\s�� ������綿�ȖL�@ X��R'���Y]ч�S�~0(��&>�Ѕ�FA}HSkS	�y����m5�Nѥr�� ��v~����?�&��d���/�5��6�>�cK~�N]���v϶p�.P���`5&�;�lmX=�^�iZhO�d�CMI�)#�Zem�]ئї_�õS؛ lg/ٙ?��-����I���N��}�)��,^=e��.�*��f�,���T	�`:=w�	��;�`o�Gd��?��dyO_��d���� ��@&.gZg�Ii6c1dUu��o�_���v���-�_=cW#UAR�A���ӧ69ط+.Z�Ա�.�|�Y��+_��;��_��=��o��޵���-�*���΋K�z�*s�Vt �����D��4]~��&�J\���2��"`%�N[r�����{����� V�J=<̀ۜ��a��=p�x*YngE��q��gՓ�U�=@ /�9@q ���ڻ]�m&�O�����6�ش� %O�@}R5 H]VQ�J&��sC�,��}���]<z��JW�;DP؂m>��[�y�f'��z�
�ՠy�-fu�~������>��5��ne.T��b��ɥƱ9�?�J��7�s�`O���x}l�'���ށm�l[�}s<�����ۇÑ���\Y�c6���aQs�?+��"Iv�S����z��_sĤ���i�Ƚ�8��������-[�64��i�~/Lh��v��>95;�s��m�"��O�gX�e���Ğ�y�)��\I[��X�a�A�3�3=����f�,�YQĭ,�w���r�h�����vA�^f�?��?��}���v��k��|���;�V�����JB��~K����g�Y�m�ݝE�ʱ���|�?H^y��w�HA(�F�6�Fm:�d4�C��� g�d���Z���-z
�R��	������0��)�G2j�����Lny|�@ ��9皙�:i9�hRd8<�ᠯf۽�O�_��m|���|�k|���lô�e8��;V[���+���#q�c/��\J��R�7)�� Ki��c��������Ɔ�ɘi�����=u����O�إ7ң�K�=���f ��^�;�b3"��SM:��)c�� J���G����^����=qҫ���>{�����ݝ���������"9�0�|�jZ)( ����dVe@"�@kʜi��y+�9ۓ>�5�uQb-d_9d�Ƹ��a!`fS���QA���Y=f��֢�&��7�ް���?$�{r@y6Q6LJ3Iȸ�O�d���C�I2g�U�O��*�����Ԃ�����Y�@��5��ἣ���/�ښ8��[�Z~�=�r�7��	��N�w�ޟ�O�����$e����n��#;�}6>T�h�grɔG��H��hgzι(a|F 
�HV�#��7��'��^J]�ej�kz�$�x���zç���������X��U��޲��xi��ƾ�~��h#ć|�lL/*���l�41������CT	�^Ω.<Ħ�YV����!*�xWT�j���� 0 �BS������=���ɵ�v�n�3��/���2�;��!@A
�����
�U���QA�<���sS�y�ü:?��޲�E��J%�!@� ��c��9�}ק&4�\��fϡ��۰,��!��c�"�<u��p��Rڪ���T"F%5�:/�d����Dl~����к��*�� ԧө��o�]��`
��uRœ ��)�>+x3��;��`5e����kO�y�F λ������{�Y�ؙ��m	6�?�xb�^G�&{�<��<�������^$����;bFvx��M%������_�c���m����X}mY`X����
�<{bw�e�!�����O�Ȗ�x�A�x���C��_��������z���/���&��}[�x�z�. xG@|�k=�=�5�c��L� ����S��;��{����S�z�k���u�̅E5R�P�����g`̛���n�n��n���BL�FYU�Z��}��tU�Ϟ���/<|dɇڽ�>�퇏m��_r��Q�:i���� ��D���F�i._�B%ڪ@�g�*k�	U����~Ǘ�*C]xe��f���\��iyN����ż�_���a��zN~6rA��5S�Wꓛp0Q2Tzm[Gp�8�n�S� ��a?��.+��lv{���5���[��Y�^W򲃳�3M\҇�c A������L�՛`w9����y���4�����؃�tD5�U=W�B`�DD������W�+�V;��`�̂`�Nvp����Sb�6c�EM٩��l�=Az堹��H��Ė��h�쮖;��e���
�A��dy���PU�m��V��Fٙ��G�b�2�u�4m�8���O"��0c�Km�U�6kXU��e�r��Z�b�]��Z�^�Σ[��p5��1���3��UUf[Гg.	�e:Hx?W�g�Qy�1��lT���ӬU�k�3-_�iz����ޒ�������}���l�w��
^���on?��B�)��n���"��Xi;,S�T��J��9uG͟���_̒*F�d��)2qoȦ6���Y�D�[��>�'�n4~�8�뇇�?��ŏN��ԛߎʦ8d-$<V(7�� ���!�2��i���<ɏQS��?@tG�`��p���8$�J�MU&�+JQqj/,�2�������R�K%Z8�Y"�;#G��)��rjܳ�A����/o���}[*�q���k����#;���z~]򥤗4Ӯ�2l�}lY!G���Nص�_��p`w��7����d?������Fq�kV�Z�é�?]��pƋ��{le�ng� �x�ѪkbagG�]��08 /0fvu,���g��~�^��Ƕx��IΰbV��u ���z�0J]+�vm���}��z\Y�$6��0��M�=���6�"�˰�t��z-a?����c[�{j�UP������ P������M���� �k ���x�%�S;�Ə-^=#����޷_���c���3�gU۟��7�+�}k�^��3���u�?�#Q$��	��ӮWdG��� �s��d�$o��Lҡ�ޖm����_\�O�Ο�����O�`�Ye������ᶭ�9fW��~��גS���.ܱ�7~e{;�m�*R�T\дH$�X�K ���w}�v!`5�e�9�il�v׬Ŧ;�f��f#��_X�f�S0k�#� I��Xn��Ң� �Z�Ϋ��PSM$Osk��}Zu�'�8��k�xF����� ��jr��2R��5���7���>�m�q�p7��Gڇ1�:s���lZ��U��̝)y���c{��wia�7R�I�Ns/�Z-���;�}��}������v�Ӱ؛L����Vj���Dyc1+{j����#�zʚ�`P@�ӣ�pI*���'v�)�Ó������l���� j�I��+p�W�_���{�kF
L���ެ��u���H*�}"�'XJ�(L]���qf�a�7�/u�6�o��_�_�޻m���Ҹ� >����>�j�v��y�];w��KzN f�U�ް��|a�o}i;�O$��bo����9yNυ�a��c��ܒ���#d����2��+�U�ĕu�D�Z�W�t���3�Ox��'��[o(i��x��}ɻ>�ߪ��Y{~6$z������i�=f���c�w��2�Z�Q*C^=��C��o|jg�]�����]�򺩤{P��&��"�yh��.);���*�p�80(�}�����;f�.a/Hn��8�T��:!�^��r��E��ι��p�%$�0���7����i����;���2{͠��:�l����{�-�H��6W#�����noj��9�P<z�K�M��!ȦG���w���j��6p?����عs��������/���;}����_��L��0��貯�I��W+2<Kb�=ئ�c�V��?�������6�<���>���]��
���f�k^�������?�7��};��l�ZK0���~l�ا��m�����������5w�����5���Z2����:�����0����X�&�� ��"�����c��ɯ5�$f�Z9�(G4K4��}aV$���ʥ�ֽv��/�>�T���r�Ae?�J����/L�t�b>؍{��K���'�����SRI����v��j5Z�u��_��A�����I����i����Tfť"��آ��ZC��
=�]T�J��*`��+��"��VU��]�Wey4�\ǅ���T�(d��դ;~�T*AG��2���8�G�D*J㍀Do�?��GJe��y�F��(�F+�y#��f��ٱts�mA��"��B$�ג:[h���?�$b��BBO�,A����t�%�UGM�bRHX��B!� �**�jcQ�:^RK�v�0�Ƣ���!_�!\��.�{��Ά͸��$�!��� H((Pa:c�+��������=۰8�}R���2�h������r:z�AנF���+yd���q�_��8$8�}�����[^@��u�pk��]N%LK��w{��Rv�)����J���3�g��,��\�������� ���J95^+���S:��T����9��8=��R�ݥ�/XM:��t���KW��?�s{�~b�S�����n�&3Kص�_}�����3�ۛ��,����S��*���HSs[�{l.m�"	XW�Mb�qo��"�Y=��١=lg��2,5���<�ds�j�8��}�Z����j�����ߎ]��"{���a�\�p���5k�����m�?z���[<S���@#�rRdG���
A�-e���\�H힊2+q0ה��S��hgS+8EC��_�����؏5)�m	��g`��q��9{��o[���|p������c�1�%8��>)�[mu
RYɂ٤��
�]۩��
Ƅ��,MG��`���"�13M��d��Y3��{_iW.��d��=;{���� 76��4��Ti�����e���A�ֆ�=y��_������$=�dPC� Y��	�U��,�`S�IT�<
h�X4C�0�a��'�ܴ���I�{Ͽѭ
A�t��L��A��- H�|�۵eJS( ���+�S�@��i>,IM�܏���6f�#��08q���Re� �Ο�;  �׹�-_���c�8���pO4�v��e[�^{ s	�� �b癥���c�K<����٥ҳ��b)��y��I,&�����d�k��b�hh;Omp�7�����  ��c{B���lqq�:[�,���ςN�}��3����<������_����<���*:��,:�#E���)Y��8�-�EK��^��=iP1}����.���/~!�?�F1����̖`�(���,{�����XQG0�{��Tz5������ć�m������&i�x�5݂�Np~i��
o ��`՘@��h��1�U��[dg�3Ȓ�^�fr�\݃=����j>ڛ ��!`j�Ⱁ�6��g<�SN�Dh���:4H��v�l�f]�7[ 
@��Ol��]{p�+۸����T�	B�SYPC
}���F!�5U����w�rg���`������S{���7�jO��L��,ۣ�'l�=)�XC��N�g_�ͤ^q��1\?�mG����m���5�/��hc=YA���CP�7�p3�O��֏��v�5k_�g� �勰o'���Ng�� xh�+��T���IJ�;������is�����P	;qܙL�4B�h{��q����h��?=�.u�t��7j�(�-,9�D������>[ƽ"�����4'^��P=!�
Q�^�8��\��(�����s�
zB�E������Ŵ�]����o
^6���p�_�f�0$��,�ՙ�2zУ��z�弫ގ2�Ҵu���a��&�L���/�h�_X���_+�E/r�^�V����8 g�~���r�~/����7�_��I��Ux��:+��2��:�����.�4�1�A\��:���k�C6�R��� 8gm~�ʆ塍E�`Mt�R���9�t�l6Ie!B%��9<a�$�?a�ۭ�����5�򋺾j$&��A��!�!ULd�	��#��X�`�+��#�6����)���KA!QrG���Ia��q�` �N*`����n�� �?n���uI�a�m��V�w��E;�֫v�M��ls�v�<�a��1' V� Iu�v��}�r�Zv|u��]�h�G�l��w&f��;��� �׭�ܥ��<{d�;��l�06|�9�Q�8ڞ{kX�p����p�[ֺ|Ƭ۰��C���M{tﾭ��7�����O������S츇��o���C�`�;�Ț�bǹd0;���V�Vj-[���J�%BRv�0N��%q4���4�+��8v�4�	{v�<��{6�WLm�eW_��J���]������7 �c{��;s��(��Ol��]�X�T���I?r��	���s�s]���0mӧf�� I����5��*Mp�����/~i+������EO�v�pl��ph�Om��� j#��Ƨ��'����{�{�l4� ������5�w*���#�w��ә�q�y-`(pSD8K�LU�l!��f1� ?8����ۯ�����|�W�%�c'�!P8}����ܕ�`/�
i�(;��{ۛ���،].�t7q�q]S����"���x�,�	��)%KIb����<� ��P��A�rl>����U���6�e͹]�+}La���5��=0YǺ<��[˰W��y斀�����Ϯ�aO��+��!Fn�]u�Pq�y\܀%k6G�ئ������*���9[_�cm�ȎHUhu���p/&{b�s���!�k�ʧjZ"���SK���[53�#�R��|aqО�Eqh@�m[{� H�"�&g��g�?�uxF����ij%g��cu<�޴oU3�b�tk�6��ɔ���+�x&���+l֜R<#��R��|^���� "��pw� �R6<͒Em��V�6�ӨPF������VK�a�n��N�I߁�8���T'��$����F9�6x����	2���\-N*>9�*�Ϯ�B���ɿ����ݷlM�Uʘc�u�ijP�6P�H��3Z�Ac+���[e��\��}���9%�-�?�<R���MHS����m�֔zN�w���B�$)+����;u��7�+/`�4��fT"�0�P��1g�����I���z�:�P�@���>Zʹ���e>LO��WA��ue�m�T��`#�d
=x"�!�8|��Y�^�����س�m[}��/_2;�n��"\k��:KF��J�Qud�}��t!���ZO�pw�>RY�Zi���^�I0���!S_)�G�#:�)&6 ���|��%�9��hR����P�Jdl�WU�}�v���MW{�:��A�,�_�?;���&���h�ρko�'�`=�E�;�C���A6��qh��v�v1�2��Yv��BR����D��K��`�FȅK\���\�B`�4f��.sT�IoQ_k2�*��9xN�o��}��X���k^~����y����w�9?'W�w�z�@Ј)��+4Pk�MH�/��À����;�P�$B��%��F�?�P��y��~�<�e��i:)K��d8���6��|��_�����!�@��n��/a���r�W<=[���p�r'�P����T\j7H��hs\�(�2!�9�8�!I���>\و���Y��B�t�<ߙ3aֺ��Q�f{`�v>��Ʀ�/�U����s���w�l��p"� O�3�jĴ��ml=��{[����kL|���&K�n��ȖO��K��v��e�#�����������}��={�e�Ƃ����}��d/���N���]�������"P| �<،�����[��WJ\M��o��n~����

N�:k�������y��gD����'ٍ�Om?�M����f�h�{�u�v|qQz�:�ڴp�)O�3�ҥ �^~�왮���}���R�)Á�:(3p�-�8q����ݏ>��9���i��.lY�� ۏ����w��Z���K��ѝ;v���!��	 �8P��,+]� �E�D�b��!�R����NBo�^S�a��I��e<�ѽ���/��8�wwl��[`�A���#�����n����ho�F��0�c5�rzk�h�Ip�>]��� /U�N*5�d�h6%�7�����b�fo��&�����Ǳm��Xm�kg���6�sx/������fo�����1_�( @4n�nݴ��ʲ{w��Ҭi���� "�~�ֳttM;V�8R��<|�Zcr��B{���Zlz�2����ݹm��m+�X����}���#Y�)WȤ�����s��c���V�:u|���?�*]��+��vH~1v����7��HȤ�/�++w +�����<��b��U�p�8�t�3v�Mn}n��c����sW6I®��~^c-|�@�~J�"yazd��F���l!8h�|9XN� S�+�\���{loo���?�2�.w�YnR٪kY��a��H�a��J�{��"��B��4ޏ�`�`qʘ��z!3U���P�P�� �S:�{�쨏�����T_6�w*NKǿa_u���"	�
d7*�yN�d��Dqk�-7�1�J5N���v�(��j���t���((�TGI?�GOoܴ?��57��� ����@0n�A~;R�AYȹ�u�l��/���c�' ؤ��);��T�0���-�aWIE��)�	lb��iN�,j
�ǵ��V��h�7��Y��l�"�'4��ɿ�-���ќ��ϋ��b���<WnG5w��*X1��lfVRq�S�G�!AJ�?�K�0!YJe!) 9�l6�3�ء��b�,Lg��q��{��J$e�΃�6z��F���/]���V��`Q�>��GVA�� �s�/1~>�JO�ɤ3������GA��b�i�K��]��7c�<��������O��ݒ�[���lp�M���K��5ۉ&v����8�Ei6��,"�o�y����V�N'�dH�3D�3�Ft��b������*�A�d<T�+�m������������AA'g�(�cl��Rk��)�Zs ���|?��l�+�L�K9�*P�u�l���V���'t�:P����A�\�s�L�A��A�g��W^|yQ⥢�jC�����{���4<��Nrj�������cF���G�ˬ���>�K2*�x�z���%��q��V�J�N��u�8�g��<�3���a�r~TO��� Ǉ�J�r ��-�}�L�Z�!���Sq��i�$�(J>MN/TU�+U
��o	�+	.H��bB��P�x��$����9@���`<>%yx-YPb���d83])ւ���w��3��O����%������ۮ4ط�Ӈv�ӏm�I�Mx��O=nH8Q����X�hZ��I[���v��wl��I����m�~h�����+v��y;��5v��=��{Ӿ����4�*��y�ٔK0E��*�2��������_�ܖ�|���������3n����� [��[����mR���?�ǟ~��/��&iIp^M|���J�e]*��>):�SOZ6B@�3��#?[Ӂ��5^8b�f�����jt�g���I���a�ؘ��������������$%����ɷ�v�����͓o>��N����_����>�:@f�,]��CH���}U��w�}枴
{3�"F�+U�Jf^RR�`O��Ӵ&���{jF���"�$�� 2������
:	DH-K�u���ɳq���*���V-|^���J����G��=d��@J�1�JG1����$�����v��a��N6�ΩU�ݕ��{�{	�x�Y�c�wP��x`����_���|i{Z#8�{�Fe$.i�\j::<��P�/�u�!�X� ��Z�%vz,�#��"ޤ��EX��A��A�y6�Lm{� �6���9�Y�G�b�p "���i {;�܇Z[�>Q��av�Q�H����SY��T~��`c��
���iY�_���]���/�{�m�u��+����Q�Z<��g�s�S�,F$��=%0Ҩ!�����L��	(�"ϼs��l��E�F�qdS1�N_R�봰�V�L5c�-�V	^�*�y<S��ͩt�	���B ���������r�#�Rkh��0i���Mn���.q���pg��µT>�	!��z�Մ��8^]�E+�@A�τ��l�;�+g���*���R�~��~~0=�d�o	�`��Qb����\5?A��a`Xd�gJ�i=�]�?������llZ��  ZJ	j�&�s�0���S��߱N ����"����{�;��4�hH:��Ce~;���ᡥ
ڸ86��$��nEN�O�=�8u�2��C���#��<�����̇汱�xJՈ�{��f�3)�E�yr���~=����F+�B%k���2v����� �C���=���u|o��w��h� t8���&�o������Om�R�f��>�m�I5�vq?�^A09acqk�k��ְ�R�B}�p߶�����q!��^ϖ�X�:G6`�`n��l���#K�k�a�	�M��D�jo����F�?�R��u�}J>��B�n��cͺ5��������^�$]�8��k�=dCxL\<s���:��0��OWm��W�w�b�Ƌ�}ϯ�Ԣ�I""��ˊ�]Ԥ�l�s�_A��$��t���uR�աa��D���T���=��;,۳��l�������u~���0��躩��B%'��@ga�2d*u���K�I�R���h�O��U!�~h�#�1jȗ�)%Ň�!I����&�g"s)j��&f�Q����m �����
c�`F�������/��	'f6����j�eM��(�KUI|"�_��d<ց��^D�"ʌFQ�܁󥩣I�mP�k�����yD�J��^*<Ғ�61�L�R����#���3��|l��~��k����!�C��jh�߱��~e�~��(j��W��G9q�=mN�a���/퓿�K{�[��W_�Ɖ5[Ľ� Dp��������ʾ����������-ia͙&@%؊�f
�s%I5�b0�������|@���{}[ſw�����n�o =��gj��kjis00U/�����]�G�
#��jy�J�W��f�	�s�Գ���� N�)��6 X� e�
��X���T�3D�L�������� ���z6��V����O���x� P,��gړ�R�p����@��Z���3���[��UhV�Y�g�#��j�l4�jx��5d�w�3�ôn�5���f�#U���0cV���F�j�7��ә��RA�8��  ��s�"5d�Y���JP�)39ج�	�C*U��'઎��ߢ������5��t�N]{��+K�-�m���Sooj��ӯ��Z{�gN�Ӣ��'MH�#�"�J�@j%�+=��+B����h+��K�6AFR��d��v)I>^<
SҸ���ϗq����R	v��M-��/I��8�u�J���(�\М�B�`��2���CR�r
Q80��8W~�s�H��.����v�޲��6����g�Z�zܢ� �(P;D����A���I�6���è��WJ�2l9-�sΛ�ǜ
���\�%��n��LM5�I�p�45d�8e�	'��"Ń�X�|�}� 4���S�8N�+��$Z,�cq���&.K�a��		:�f��s*Mx��3�O�5��bY1%���.�9j���s��z<j޼<ce���LlqM�ćUf f���W�P�h��9ך����9)�o_�+҅��ӂ�i�j~��A��/Wq�8����N���VNPC�C�V,��ܕ�4 -w
@�G+�Ŧ��4�� �% �Y�L�.*�ܨ��l5D�#�#T���wq��k�D�2��|��+.q��+Zr���V�+��W�1'��"U�G�3�|5�^֜�$lT֏|2��\�8
�p�@!�ϖ^���4���Zj+��E�W���c �A���7�Z�0��hW�[q0������կ-��b�ڬ���S(�eu�U��XXZ������I�IUV���~���vJzM�G8�P�J��\�@/K�����ė5�\�����=�����;s|qM{�ם=�k��JI�r�o������A�C�R<)_Ly[��I>�'ٞ��m�ĺ�N/R���~�������W �/OF��y�腩Oh�$��:�sZ�^�ߤ��$6�[U�A�g���W��9�No�+�(�����@�9�
�W�R�h��v�^���&�s��[_Q���P��,d�LT�3�����9QP�zq���� �z�<�ҷ�w<H�OZԠ V2磋Qο<�C�!��F���j��8 ���x�)�&���t�N;&aSM�4Z��L���e��D#��r�gGA��"�)qc�~�L.����r�BJO�6���̃������) ��͵�V�Zĩ���&�>}d���=��_��/��sg���x��lo�����u`��r�x��85����$:QY�J"4;[�ſ��6 {k�'v���H�!�-k�m��?�xf�o}a�?�ض��Ң�1@���^+���g�m/5N&�J���I��t�J�ԤpN+��=4N�o�� &��p�z#r�O���{/u[�խC}z��Tԕo"(�����# ���J�zM����B�w�%o��)��
�44,��o�����P�����3���N����6�l6��sd������LV*MG��vD/���ۼ�^�ʴg|ș�]�  R=�����Rgj����K55/��9�ŵ$����5�X
'�FZ�a�����\��׌����"��B՘���a��v�%�툚x֕v~�,�M(6�j�k"��~�>���{���vú��E��_���e������~"M���f�m�z�����ZȂ�z|�ĥ����
�q=��xNK����_��%���{�1ld�J���?�%�/�:zp�ɈӹGʬ�z!%�oĞ�����SQ,��wK��E;�!����2T\-�����g��P&9��J�x�J�������~���6l�`8Ip�KO�436<Op�2[��O1�DTV_���wI2�՘" tל���L����B�낸N�f0և�#� ���I.�#Q����@j;����&�r�yQ㏷T����E�)D���4�0+I{կ�B���4�Z���ɿk��͛^p1�J����wic��|���9��Xז���;�d��T��׎~7A���2p9菬Dp9��&�����n员Ai�g�^�0A�áͲ>��A~������{���=l�ܧ3KA��R�
��Z��Ed���P%1�j-ML�NT=/��`��d9M������y�˼�1r��ټ���@�'<#�KNZ��9�7��03>���G��>;��+��*�_�]�AIF��ҩ^�ea�0�@�qU$[�hB���g}Z�r�AlU6�1q8������ �L\·_�l��];�왥� �����/�9��  ���*�i�!p�^��{=�+ ���e&Ok��UڻT".�fN[�Jg�$�T����PP*8��Q*E�~���`�U�$q�m�&I���L�q���J��Q�9݈~�v���@�ȃ�(
Bs8����^�����C�Ғ��m��&V�)�QEm�Q����
�������8�VG����i�
���D?6U�('G���s����9�GR��aԫʱ�	�8�^&��b�J�5Q��XvDKq#��s�������!x�^�.U
�W,��Hc\g���*N5�+G��Ѹ�`�쿠���3����Drv�<
�L�A� Q<q�{ƥ�qN��Z3�L�#�) ��z\˛ɤ��T�v3m5[i�nIt9��٪k_\�����E�P�}
��}������jj�����Pr�!WNP�w�̣p��J#��SD��2�/
�Ň3�=�G��|㼲"�D:#��l��i)~%��eX��XM���M�+�p
�t��������];vj]�>�5�	���3��D��0��)�W'�4dt�4�i��������al�W���NӠ ��[���h6�r23�E���¹Z�s줕-58P�+%�#xI &i���)��]r�I��o/��gҍ�r֒�0Y�\�^��X$�����"�c�S��#M��Zx�S��C��~Δ��\Ґ-������H{^gz.k�����$�IU*+���0�q�睮s���ܟ��Z��Væ�Tv�<e>{M�ℎ�'+���t6�n#Up����^��jN}"o��s���5�	|�R��‵ޟM4��"��~�����{Y:c�2��do��<����FNn<�Nd��&A����㱡�F���;t�F�?K�R�LT%��5$~l+UE:�<s��}��	)G��~��s��^K\A���tz��ΆK�l�Z{� A�2�꫊��Nc`�`Y���h��\eě�B�Ꜩ�	��(;���ʘ�V�<PQ�� ����@���RR5{��U���$s=�-���+�2 �*��P=��F�)���N5=��إ�q]��;����b��&V�dz)ƗS8W@��o-,ڴ���T¥����}vpߪ�i��ج�g��!��z3�kNW��fM�3����Q��	�(�+��W�q�i^�77�DA���%�
��� ��!%%�ٳ��� ��6�}����0g�qS��)-eV��Y����i�>)y+}����y(<O0>����)`�n��nb3�ӱ��5<(*K�z����4ESJބ�A�ʷ\��e	A}] {R1@�ԥO�A�ԊAA ��J�s��Fql���
/l<���*�U���h���1I����Zy��u�88+�k[���T�SѺ��WBbN�,C򓀺	XϺ+����`�����`A����^��� 	@|8���\*�uZ�N����d���u����;b�(Nq�'G�����Xأ�:��UeڃI�s����6�W���+J�lb�9�(YT��y�w��P&�{e��&�K�Lz6�bV�HYb�o4:<����>Z�b^�1U 4BX
X�L���WH���%2	8�>�D@�>i�
4h��v���~oP�͒Uխ�������?�ڽST�ZZŽ�^�sjP��!�TĚ6�	����JFʯ�uT���Ń��C�	�_����r�����+�FT����aQ���;���PБ�ں�*�ʲ�����0��N��iW��]Go��i�^
ţåk��vX!�Z���*�ȫsBUUqc�z"*l@\.I�)e��}n�Z=F�QVi�gѬ�VK���Y����Z(�!K��9��`��������w<��H�x�f^�^��c�+�xvz]��x��Y2:ޒ��};�X��<��h�>���R;��bBs�TC^D�i�7��K���j���l<ef��(
�/��%�ďkt(� �t4�n%�U����?��B�f����BG�\'L$iX3\:��[�mhp���K�qT���2�T�I x�'��P6R�p��?gI%��6�fI��\WKT j(�
/����(R�ĝ��$��q�SQxM�&��' �5��@�H�"�����*�g��0�A�-3-��%� ����֦�d��iy�\�3��9^=�i�{bfz~4�^�t�Ik�t
����/s�'��X�&���z��3u��fu%�<�+�J�N7�x�����wN��w,d�K��ug���ф�Ol�0�S���a��:��?8�ޢ&����F�������ׅ���;토���g��a>�sl��L^D^��j/�Y��i�pI^��C:g����#�WH�-�����)��L�.g�{�G�R��X[�O���f%C�l6TmH+���.G6<TS ���a��ȔQh��<i5� S���	ث�ܳ����x0V�Egn{o����v0�d[$+ة0�vHz��ϭ� �U�č���h��f�r޲�Z����kzӴ�,�ϡ����W�s��\t�{��d�V�[�����@Aڜ! "+\�� v8�<7��7?�.��b<î��$�M�@hx%�UV@�3�=�������&�|\��@u���[6"�?;�9cE��X�=��xH�7��-������I����6ƚ�gC{4����`�4S�z6ZM�)��d��b��tW�n+-��4A2�$W=�G�`��Ux}���9/}x�!�q�fX�'��αc�<}�z�� �h�����>ٰ���MU0ͼ�{ձ�ج�JEhF�n����o��9`?T]��D�I3Q02�Ǣ�p�q �" �m�6��r�v�YLe

8w���Eꓨi�iL�Y,P�.|���G�5N���>�{�)$����}�RW����p��'�k�F*�GG�b��Tn�d�J�8��iK�@��<R��d����Sz�,�W�T���3G>?$f������zB��ώ��7D�a���"M� ��s9�2 �0���Z�H�I��a]5��2��8�t�g��w�v}�G}�o��h��>��U��m�43�Y����m��x�z�VQ�u����A>��8�z�Ք�i��(`���֋F�g*�¤o��4�%q尬R�o�#"��3q� {��M)2��=g%L�#��E]���0��1r�����p|E����,8�p�q��R"7�0�u��9���{�%I��*�U?~���K�py4-�p�ݴ�I��*c
���G+�I�>��"/�(�\�2f�P�)c����+�Sc.?P�j����|���G�F����/�N�(;���FE���߭=/� j�s����*���#�]���?�Ls\+5Q,�'�߿�?��4�dR�9���(r��\���Y���(�N���эĉ�uQ��&N$7C�ke&k�5�/�vЂ@%�L��%Lo���7l�{�2��E�� 
�rV��<[M����~4j�d)����$�r|��#}^�E�Q�s����Ԥ���IX6��x�f�Y2Q��:U��Q�_��6WU�W��s�aDN���Xs�}��H���!㳩��eU��������:��<*�/dE4�&�'�9��L@OU�&��̚�رr�� ��yv̞.��h�F�����xx����R�(KC��5㩨�<�D�
�&Y��e��
:n������`� cD�"���u��?�i�q���:�$�W��`�nWǝ��m��xL\�%���r���lG�(�l2���A����y�(�������Ulrg;��X?f/�X;�1��-����g@�Ѐa�%���(�({^A�C[*s<OWA�N�&rZ��Rsav�UN��� ]X0;��Zg��tĸ����i�px`{�؆���r��W�K��F!�|V�z='���f�S&I�T�z�]Щ�_J J�R�C���Y�Bi��i�i䒍��R݋٭1 �:y��5�S�+<�1W�2~V��x��Ғzü��.v
�F(U!�=߱����Ý�4��+�)26�Gx��o++��-�l��v��@����m��<�R������qv� ����=-���{3U�H�j2s�D{�����2��J0�VH�h�#	?Dp�p��zqCc�[{��]^T�4��:����(�@�}G�9�}��ڸ�{q�P����,��i���R�tJ͇�*����KSC�x��&�e͇���Mf3<�	���b`'O_�3 ���U[;q�N�:g+�����w�9���=5�l<����W�@�;S��6Bo����wo�mްͿ����?�Dk]V>�ޙQ�*_%�� ��������ĕkv���r��[�9x
�"�)��+�"0ళ�w����{�EiL�5����? 7q�&���G#k¶p���r��!c�^��hC"0�}�E�`\F]�d;���]��U�8u>7� 
� ��5P�``����W�(~!��@��|A�2y��C�������O��ꮳ2�ly=�b1o�԰[)yQ�N�bn�Fġʨ��t�e��T�g6*�do��O���93�Fyq<�Ң�9���p����ym��v[��,a`o��\�RyPP���4>yj����,/���
�T� ENa����{��K���k֬w�-���5��{�"��ph��D`US�bJ�TN�m�_�y��I����ƕ��%�X����3�Sf�N��*xT8}�VӀ'%�$�C�,<&���4}�O}�kqAMj}Vqs��:X��)�-Ѫz���Z�wj�}�	qC�*_��Kꐡ�	���o�ps�*�R̤�r��}ϯ�׉�gϞŉ1~=y�߫���2O�����l=���t��y-ϋ�v:���S�Q}�i�D	9 ��r�TY`S1����|���a�iR`0�!b��C͹μ3pcop��Ϣ঑��}�ũ�έ��!�aƂM���\=̼;ht�$�U�$U�SJi2��Rr��	��^���fM��G���-�%3rϬ\j�Ba)�XHv$��M�����c&�������g=�MҫL6zP�Lf�ʦ�I ��j��=3�������Fd{$3��9֬�%�d�{�Ͽ���ω���e�67�T>Y��X�����sW�"�H��F6Z��15�'�#8\J��8�\8�2��9+4^�BA���C�J�M ��IZ��:���\?��i�r:dF=.!y��Rԝ��ײ�Q��?�N�L����X����}9<>��?��(n�2��zAJ�]c����7oPE&P�C7H��|4b����BG��TZ��@�����T���l�V����HM��7YO�zl���uGi��67�B@�,��\�47����T&�kF~>�gn��ܕvKJkK2�X�ï�!UЀƃ�=��VF�i�V�>@���e=Itʐk�.U
��̆�A#�a��f�M�j�yz�b���\��my�{%C��f�Pg����.Ԥ��%��BQ���"��,���!e=��'��g;�4�	Y���w���ޢ�^-W�PJ̵��<���gn�y��B�|X�Sx�OJ<�Q���5.�HuiY6._�K��9�n��T�ۧIV��@�fwz.�����8cbg�dUK�V����u243���%��a�bI9{�YQT�VQ�Bj�$�=��:�JMF��Lu�F�k.�IM�m{{W��;%�����#��p����}�P&��J���J����(�rHHF�7$h&ϳ,���l(Lh7�{]]$Ct&��j���̮��o��6�e��5�v�Mٺ��D�E���{6�Ҥ�
[~w^M�z���������B���t�Itt>|�2G����0�o6��}�b:js3�"�	7; 9�������Ϥ�m�&[7nʛ�'����DK[�e�z�,�D1�kE�G]����r˿��?��O>��ᩌ��k�Z��̦��C��Jb:տS ���d�Y��}ZJ�I]�y 8�vu��l\�$Ѣ��U]�%&h��C5�h[�3���(Lzz���|j���z���^�Sz��o��67T���	A��%����w��[�������xATA܅�Ĕ���Yd�I�c�Z�2OzL2)`?��b/���ߓ��s��/PSa���eY^ݑ���dqe��e����c/�jB��caQ��vdQ�HM��P�2�Ż��b+�w�����?��~!e}v�A,Py��F01����>��	/��kW�����/�֮��Dڭe����]G{��zeG�k������)5�lT��b�0�u�g���416A��@?���o���6��&��9e�nL8�)�c�����ȟ��cN��q����T4��cV��k�����hs�5����5M�}<�?��q�\$��z=�^c�1KKAC�ܗ*���GQ�G�~;�?�����'�|���Ο���O���޻���-�3�vT�X[�ԟ��YE ����C�oz�C�d&���.�&2�1#��a'� Eߊ�f:���&�ݕ9�=���+sH�L34*\`~"��)$2>�w�X\�^����55c���t��5x��)�B�;�|�]��2�nDG�b�=���}���'	��g�G��g�� �m	�,&<�YYA��6��!%�(��%zZ���T�M��.K �8��+Mļ��#9=�ꁕ�Z�,�r&K
`�ТFe�w$�Pa(�m��������_��f��i{��n�a`: w*��s����~a�tdgc�U�5 5}���<{����&?
�J5�xe����#��|-�g�'4�r�}`�Qn\m�9,fV�:�E~<�y`�!U���z�)P�,�I�� ˬ��HA�Ӕ�K�/��𑜝�IiuC�vv����#�����jZ<�m�t���p�������X+���1+BH����"�)G�	�����UR��z�NTL:˲��!W�������*qT����l����@�����X��->��>~(=P"2-؂+�mrPCB�I��{م�]����i�sY�øaG<#?��:Z�iT���E�ۯߕo�+��)�^�(@BL��k6'��Re�Z�-=������W��X���S�q�k\�b��scv�d�k��M9�JE4�S�� %���u1)O�:x������b }kM�*��/���o���[,.�������/\Z�
 �pW4�X__������
���B��L��Z�t�T5��e��X�}<�p ��Υ��|����H?ϙ&���F���[�H�=M&
zj[���]��λ����tV����L5Z��Jpz�Rj)�=��׾}�\�z[~��)>�D����#c��2�����ʳ		00+�2y�sy����R� ����  �pIDAT����e�o�t�����[r���d�Ϋ"� ��ӵ@`�f*F��UoGP_[_�ΥMY�zY�(�_�"���C]�HWc�=k�F2�b��9�+��ÂH/�Ifi�Ԙ`	�Y��H�?ޗ�q����,��mM�D�+�t�3�^�ˠ�]�)%�W�3o����{��`�V���VC*����_��D�}D5��^@b:�>��Sy���z�����0��Ut>�|�ll�|�	���qVD��B�t�w�1m� w8@�"7o��7u-)��l�[�&߇���?~��uM�'���&T�r���ԓ�jD��JdU����.�_~$MM�[׫\��L�*�FW�֥�g[�We�W���o�¶��&U���u?.�ۺ���Ɣ�?xK*;�,1�F��ϏJu{��v��������gO������4�9������"6!��z.�O`w0a� �GX?ah3?���ЕeIgJK��䵺�	g$��e���R�tz����%]]�xs]x&���ٚ����N�����QL/9<��/ے��Y]#O]���n^�������_�� �ۿ��͟����h�?�V�����*U�M(Фƹ3����Їb�ڤA��P� ^���` �Q3���,k蔗���Njդ� @�X���%WC8�g��SqՕ|�
��(�
e���Rh¤-}=l�\������嵦�����A�*�=5���'������@��hϣ� �$%�2�+�<|�
�������8�Vfd����v�P�G;��ԁ��-����&�Վ�U��&y��@��4�cI����T��?��7�=�zxUH;:Mq</\?+�S9Ԡy��sMg� �Ie�b��8dr�01��x�@&���K�.ɞ�����dM�{C�Pa�Q��ptp$���@z�͖\~�M�^���_���_Kzp(�٩��Ϸ��]l�΀mީ�C�JkPL �q��Y��z�)z�~J-M� �7��=ٺ���޾�J,�E18�k�٭8���H�/�7�;K����@N�>�_(h��KM�z��iTu���Z$ޅ!A�{�& ���l���d�*�hs�a�r����W��&x
.^�}���۲peO4s��󥫇��\�����ﳺ}E�r*�"W_у������>��>����B���u\ð%��S��K&͚Ë.��
:�gq4�F���>�����K��C�xuEn��]���?�Ϋ��W�N�I�o��fSʨ2�s㇁g�+��?�s��,��X>]����G
���Hu:Q��Ɍ~a����^�9�8�j�e�q\��)MY�0y(������voO�WoJ��mi]EB]����tW���x�{szړ��S�n�T%���Y�K�R��YceE|/cM��}$�G_����SEcH�~*>��
bR���	�}-`��\�ܹ&Š@f:줽�>8����k��O�\���~�2Un��I�b�jiQt�*����)nP��]^�la]�w峿���g'�_|Ǝ�j�J����ά�C���B��Pf����� �֟�_U����r��Y]g�۝p��K""p�}��L��,=�O��jT�y玬lh����7�k��_��r������.���5���5���j�TQ	�M������� R�"w�c���y�T��iR(K�D��{0p��)�]\��W�d�[P@�q��D������8RrZ+�f]��iܸ)��-T�A��"��\h�����c ��65�L��D����!f�:�����(�F1�368�"2��H1�Y��ѱ`G+ȅk3�M��5ګ�v��,闏.	��ҪD����^ַ��.���!�U\����b�fRoP�����"7�}S��{a}S��+r�@?��
|�u}�(s"�&e�k+�������P��7�9�	9�h�*Xn4z;�^���j\�gue�hga�y��%�.��Ҡ'rt(���G2Գ������\�5��v�Y\�_�lI�:`#=�i�<;z(e*5҇bK
�B����ҳ%�uM�aEB��L����i[��M=����e|6���s�<Z��3,i�ڪ�IeE�B1��8<�8���J��CS
07���ˈ4�����2)�g�������{P���F#"��e͂�9�N=	@���ب5��'�Cb:3��x�1e�t�����|�xRx����Lpm6ȏ���&q:�X�9�Ȯ�`hn����[���#���vK�k��/�E�-WȇG%�ӣ}��ɓ��ͯ>�GzpN�V�S/��ehMHs vv�B�T����:e��[� �a$P[�e�}:KA"*�W������\�����U�X�y�_�a�GE8�Qq�`*���}�+�>�,�^Pџ���q�'
�z
Bh�$�L�)�)L>�� qILX�Kꗤ� x���ҍ�Ə,���}���1�z�	�W_|���w���ٕ���|��,�����;�����W_�/��/��/?���?ӳ��ԈP�F<6��3^( �)t�N}�#�/+B��0Z�^P��p"g�8��������X~�/���
Dњ���O�K��Tӷ������*���l��U9Wnܑ+�ޕ���eT��(��,�MZD� 
>��F��M�ڷ�%��iJiH�6���aUꬺ�@��ݑͷߑ���i����T�jw ǺNϺ
:�|O$�ZS��T�~.}������k������HK���ן������X���е�P�\�zX>���n���
x@� �Gg��{�����"����\��yW�W�Q��LHG&QE�mO�@߃�fwDj!����UY^^�ÿ�{�!w��( �T�{�W2���^�s!c�+|�=���3�)�݀��)�f�G��Mu=T{�w]�٥mY~����wE6v9��?VP�`�)�L�R�� �Sݣ�<l�d�$��z�4ɩ�:R����%]�Uy������4�ˡ���[9�eA��] І��[0B�\����t5D���v��Ο��r�?Vй�kzڃR��c�B	��$KQ�G�T�uh'��8UnH��yS�KI��#~�!+�+�XB}.09hvvs~�Դ�\�O��뛱�4�c��X���k�Ƃ�}�W���c&A��WhF�V`գ�ؙA�������uJ[[rU�rg�ø������?=�|�v�ԧi:e���/$��:��|vI�MM
�(�Bܷ�$�Aa6
�K����<v�#rI�J������c��r_�U_?����iC��&$^[ϨE�Z��e��q��!4�B
�t('�z��w&�+m�A)%=b(�4�Mx$�ƶY:Z�[�X��Lf�8��>Kh~E�.F�h0�r�X�Aa��k�	�1|��2D=�mYЄ�����(�U!�Q3�+�u����C���	3bFV��i��������������	���XY#?w�s-"*M�V�{VL�-7	�i�Q�,Tl�bZ	���u/5��;ҳ���<�?���c��!�g6�ݐ���_�ֵ��3����zԕ�o>����Z�QWc�&Y�H��"U90O��!�Q"�3rO?���ٻ��b�]][�Z���@�=z,�|!)֊�Չދ�S� �5{�iybH%7x8G�J<K�|ų%���Y1[p���_/�������hue�QT.'q:)Q��S���8D���7���B"Z^%s8���mڠ"~|SV\�����!s�ԻwF4⪪�3j+��Һ
�$0EPl�����I)	�ńK4���Qtư׍�ٻ*���|�5�,yr�e�ip��0��rU�eb�F�C,_�*K�we/����^��~�����>���|D���i�����)Dqh���\���`�T��(�@��P�+ �0��]\������?�3y�O~�� N��N�I�`��?�GG�h���B�)[����Ր��u�0�w.IOA�<|��u�R���xv~"磡�Øf�Vح�c���A:�	��Tb��!}�X�naYn}�m������7�[^��?�G���7�}%��ZgUW.���4����u&"ߜ��u>���=y�Gi���I��=�<{��l`�$P9��9�8�Zd^	㕺n��ԛ��\���bc����⿔��'�����|����oPqkgwKA�/�jC��,KgyO��*'�3�{F㨲(��y_��my��������|Е*� d�+D՛��3W�ǽ��6HN��˥��A��H�����Қ���%ڻ,�5����/9����kv�7�4�=&�
nʵ*����s�g��߽+7�ޖ��׉<��#�?=�
�tp�	��	p�ĞsM-@	^�(��7�{8dV햶w��{?��?�d�l����ן��5���g�0_1��r��u��Qф��fK�3�脯^���������Ӟ������YT���i&
�bЗ ���"�H�nb��ũu}�b({gKں^���!�	^_���ɹ�z�^m#.v��̍��9ӆ�i6�& �I�bG����oM�c�U$��L��ʂ&�5���xjT�(��x�M�J�w����{8�"���>����oސ����Ot�5�h�?�Kn�z��`t4P$9x�UX�FA�d�����Nmo����	�?h6���K��X�f*��f�u�8�[g q6t2q���Fu�Kr���ɍ�}W�fKzoO�)+�P��p�W65!M�H�Uκ����VM��u�b ��@{�W�N�G�ӄ�i�i�B����	P�֦�������O1}L��)�jeJfh�����ƚ؆LHiJ�@����Д����5!8~�P���J�=�'ݳ}�/Cv�&ބ�ZS�G�L��4OH�J��t�#(9��@?�R�����N&�&2��g�>8Oѵ�\Pt����D�ɗ˅s�%��cs~$&/l�=gz�L0"J���l��� �P/C������:�X����dt#�Z��@VXc<^��=����h���&��Y_��H��Xc��]xaO�e$4�#]���yU�j�hB��M�9\��#�u��l$��Prz|T��t���4	[�/5)�C�ߕ��$��
�{t2�5UP��8]Ap$PTx�L�"h A&�!,W8_�g�nfVMĠ��{6e�dr����^F�6A�ߺ���A,|���-�x3R�ˤ����ߗ�6:����}]]5�.���G���I�e�F�$�;�?�d�g!7��܉��a�ȥ��$έ��J�A����*�2K
�¡	JH��j ��^�j2�xob��8�Vz�6.�+��P��я%	��_JU��רՎ 7�"��������~Q�U]��W5�@���^�/������h
Ξ��)Qf�p�1�^����41x�y
�D�Q$��+�r��ț���~M��"�w�c�s؟c�h����Ր�Q@�Z��X�3H_*8���.��Y�rM��R����?��8��^�3P�H�,:.���dc�Q���S��}�gé�Q1����w��?�O�s�����>�/���yG����'-�m�*�l֗:r���9{����|�s��ޔ;Ww��#rV?���M��2�?�f[�g����#�U��PH*��~�1�T˺�A}����Gr���%_ݔO=�����_�H���.��ƒ�
A���dݫʂ&Z�Dē�� ���MYX^�H�.�E���p����F��>W�e8�V�1��*�)����<y̾�'�چ��Z}v|��㌟ea
)~ui*�.�Ȯݡu��dU,w�fzM}T���ц����*OFI`�3��59[t�`��$,7C%)��h9t|�L��b=��;����������\��Gǧrt:�ݮ�dq�C�<�5��V�ޭ��W�T�^��}M*�q_�VZrU��M�O�ʗ�]���d@l�.���(��N�N<��dR��Щ�$	*b;��Є`�wD����?>�m�������T5�
9�4%։�\k���:�i��h��j��H˯K{QA��+����o*���'yo���N��d`g��Њ�������R�=H�,�����m�~�-r�x��j�1r��D���`!��!���Xf\e$N]\ow(u���U��GD������L�ŲWbM��-�����b�F��(�E&���z-�7oɭw����<�4!J��.�ڂ؜Z@�2v �q��e��>I����ys�B��QnՖ�o�+���FN<��_��ߩ���x��-���(.Q	���!���d�ũ��y"V��h8	ͫ��x��<º�'�轛h�쟝r�sE�F�edH��4�+��8_��� =�Rz�� B���MG���ș���7��-3#�LP3��}E�������ϩ�e��,$`i89=�8J���L؅# ��^P���YRh���+v�n>o�\"�r����?��Il%�RN��8���EE�R���'G-r���H��D�sfk�gr�^��P�TAy�ٺ��� faH���s���5E40����c���(+�U�I�Ƃ��w�q��`<�A}������k���)]�,��|��؆�݂��J_�8�Fi�W5fO'=��`]��11S��!d��&=�R�auN]q���7�P�ݽ^&�L_�/�p�������.��}|~���Ǌ�}�� Q��eC��O0��o�P��4�&���*5��R�MO���%E?0�@���۹�6���r.eh�{�y@0:�d��������[�1�Ç�d"1l*Ȟ�2
kR۹.����\z����+g�cu�uE
�1�_k��`Ź9���ԫ5�zrtpHP�����{�IueI�r(~�39r_��0�F%�PYߙP�8�DLY4|����z|'i(=Z��-o|����g��ƛ��m�=�/
L�Y�J�B:IeqS�
L���e�OGȉPq<�J��d,�뫊�
Jz2�*��@��]W &�Щ�&Ee��0�PF��Ǡ4*�^��T?�@��QE^�λ��O~"��m���yrړ��c=�e�RG.m�����5 ��J�T��,�.q���/����ˁ&*�^_����(�=M5y�C�|$��tB�=}�,���9Ws��grj2� ��4�V5(IO׃�|I�����;�ɾ���|�{`���,��6���&�
�E\U��K�]�J.�ژ�89�dܖ\�5��a.��3�i26}���2J�/���9hH�8��A>v@��D�iJY�q�#K{7d��+�tc}�S G��%Y��qs}C��;
@�@��κ8$���H�B�� ������;�IG}����U� l��N����^6��M������c���ج��+���'�7S?�Н�^o��zKښ�T+!�<��_�@D�%�c ���@� �$K��o�J9�=��ek������?��_}(��S��)����r�H/)�p-L��Q��@b �]�A�	bcQ2�P����v��#:���Z��2��\��Ȕ�:�LP��yXǚ��&��š�ϲ�����Һԯߑ��'r����e4��@a�����	 ���#_���%�#P�t��4�
�ci//����,�^1@���*��F�bW���y�u`J]
h�����OE5��ި/=Mx��7�6��w�/�����Ne�?ׄ�O��Sx\S�&c���-RS&�L�������ڕ�;oҀ�HcvXm�Oc&�a`�*唋n�U��z��S"��,ș��p@IL����ݷ���@>;;s�q�4�%?P����W�gH��L4�'�Q2`$�5�@�
@k/�Ӹ��#o�ZF�3��F�'�����@��J���,��䅶�=��jҌ�����.�F?A���7�5p��JD���FC��t�~1i�v�����,��N�o`�*'݅�{�%�gsI��� ������L�߄�+�ԧoeJ��a6��3)Nm���τt���QN��U���ҿ)֩G�?���O1X���V.HH���B2ѿMKT�:|�H&���Г�F/}�Ӂ�w(���4�pP8��<%�ߓ��#9?;�\ �Ē��n'�O�ª^G�$����<35��g	���T��V����sLlx	H�doq��S�S�f·��S$0ΰ=E��޹�猊U�H��?�OK�B�=V<�Y�2(�YH�dA��O�8G���ߩW�ˤ�����������w����?.��{o`c�P�W �.�:*�xF���| C��
@A�)rӊF C���9& %�����`)3��B���N>����jNb�PnK@?C��Sd*`P�S7���5���?��;o�=ܿ9<� ewY�r�N͋���� )@�v�z-M����&\��z�
�n����L2�">�C�LZ�Q�lpR�w�����jA��&L�tS}�;�EÃ�\�-{o�+�z�OG��QMD�O�j���e�����B|/��2M��!M�N�l@czoO*O��7�g�V�5>C��Y�ɒ����&(00ykЃ����@�ӑ�}#�N�����wdc{�T�z�r�pS�3�԰��v�����[���-]=��==��aM^ݻ,�^�K���^�g���P,1��v���33�qy�ui�󉿂��Wj�z]�������)�޻/g�4���Ȧ���n�s�հ�bx��*C�G!�Ԁ��{9=;@�>���;�1��������IPh��I����fv�s�?��5��b�tZ߼zU�>����ੜ�3X�\��KW5X�5Mbh'�!�n�3{�\����%(*-vd8�RI��	/8��7_���W5�Rm	�1�gH�\xI}�w���@-�&IՅ�lhR��ٕ��X��0��Jk�-M�H�a�:�>��?����b���Yϧ=����ټ����ޱ��ۥ"Q>1����b��ޏ��JW���b|6���,����W���]:T�+e�����hj�p~-�D��Cf�G�آ�pfEܫs��c�˦�JkA[;2\�\��䌤U/��Id�g��F�L�O2��L[��r��7dE�EL3�@Ah�=���MRB3p7�e�Ԋ�+��!�
W�r��$)�����/���w�@���3*k�V��e^b��u�@wtY#���!@�{ieW�&,I���-��$��H�ff�ws�7Z]�f�|�Ǥ0�#��=cR�R��;r��o�c�i�o�ف�@���g���1��p��s0�IL`>/�m �M��aޅ~�i��2�������D�NO	ܛ��LK�'M6��J&�t0M9�j�TF��o',�&�!����"��b�(�.>���8ŵ���Ly���Q���L����
��@�4r�@��4w��3)4�7Vi������e���`
��#�3g8`�x�`1�Yѧ�T�tUJ�*�bN�:Mu�'']��i��a�z6ğ�q� 5�����(@<3j.޺�IoK�a2���H�U��OU�&�y�ٽ�M�/����u��t ������^$��:�	ǔ&��Σ`
��XJ��f���Ȳ0��rࡀ.Mjs��I���,.f��f֭���I�N����eR�����[o��|��ɸY�����?xz��fM5��J��,#�:�i��5�p=��}��L�4�~�Q�a�
�q~Cϟ1�r�%�$L���zP֠���~6������ 4G4���AY_Y��Ҳt��<9?�<����Kr��uY\�ЂxQ����:�J�(�,-ʸ?Пӗ�nO�zUv�ܖ��S9��J~�+V' �
��d������ϒ&��t-���������H6�ߐgg]9�!�2*#5��h����I�H4�o����4�1�6�wv"'��lU/+h�}�59��9}|�����i��*vGT:�RY�w��y���5���[���-�4`?8������ζ\�v�m���N'V�beѸ�80qVW�j�������O���P>��F޸�+{��&��|��$>K�<JFN9Ĝ��!^1ll����QHy��ƪ���ߕ�7��9�[}��x"k벱�ik��8��n�;H;L��] �*��U���#L�JCAf]�㯾��#�y��ٵ��d�Ĵ��a9�4Y�ʗ[5n�~�TŠ/�������۲���	b]ʵ�6 #�b{��$�*�;�"�E2���3���������5a�����O}G50Z#A�L�x��1T���\�2ӥ���N=���҃�-8��F�"�6v	 D0{F��;�J��ޮ<��j�{�D���Ŷ��λrx�K���Kv5�ܤ]94���$�1��V��<	I����k�IAE��Q���D��~S�L��.!K���/�Xu�|眝�s6���V1U���X1��b�$@_�,IM��Ɖ���E5�Q2��W��)�9��
�]�/�3��]�����]Y����4&+�̠Л'�:L}��MS��<��U����s ܪ&>������������'�t]��_/1�5�"> Y��+�[���(���Z@��wkM���"���R���܅�ܐ/��M�4T���K�sb�1��۝��a��;k�ͽ_J�I�،전��+i�L���u�'�� U�L�j%V��'�<`�z>�f�Z׹H�^`���1���MP�a�դTfF��.:���> !�1�R~�/�[.h?s��0;��"[�␸�Y$��l� �g�����9���g��zc��O\L0�B���c�����%���9�����B=��7K�5Q���=�a���"&��H�R��<��"Q�ʼ&.qd!��[('�9x��f�Ip��l���h�S��CRJ�S��(��S�8��S������l�-�܃�oF:�|��k2��ew�
�}A��e$�ｰ�4_F��2)x��w�Z�s������kk�W������EA!��TW����%��^	f1Ng[�DV��d�����)Q�����S_���ʷ`�
 ̯8l��w8�K+��+R���hP���*�sSmaqk[��?���}�ڋr��kr��uY��&1Yf�����4τ�<QY��R��A����)%<W�o޺%�Oߔ��dO���j(�Ā�8��B��7V���Ʊ/=�)��޻*7����m��LJK�So*XA�F��`�yf�E� Ȯ��j��,�u�����ī沴�){oܕ�_|"��}I&	|���s3����gN�H0�@�C�����	���ߗ_�?O��W_���MA��e"ZQ9���`�6�l���5���2�i��?{$'ñlv�eRy����'c�w��&l�X����@v�,�`e��P�J`E�C^qksSv�(��1�ۺ���s�5�e�l́�P�[Eԇj�e���Y��pu"��]�>��9� �\��=3�1U�t�,�}�y�k��n5H�@x[�AY��M����4Q Wу^� 5`+�烅�B�1C�"�����&6Kr��+��������E��|��ی{�4��+R =�}߅�>�뷤���T�>�i���Uh�W��@R�nG�68h7��0�t}T��n�~�������k��`~��-9���2��8�d�씨@c7��u?j1�_E%�2�����H�>9��Պ��g��G�΁j��ߣ3E��Fo����9Q{n���sG��v��*ʘKUR(�o]�d�s���+��9t,^�$j�Ytyf�R�!bI���kmi�G��Uv�
�ȼ�~�r��ū ���.��i��0�v��*;7�Kr�+���T�B�6O��d]���c2VYY��LM��ս=�//I_��4�\y(q�H�q�'�*�w�����3��]��j��JجJ}}Y�jd�}(��*<��n?N��4�����2���u�d�b�X̨��ڇ��|f�י��8���l�P��d��{�Lm7г���sv�3H��ر�E���3aQ�w�F�͜�L���=�<����=�W���P�STٱXT(d�C���إ�d����"�پGo~�i�|88K�9�(r���s��|Xg��{#���+2��UB3_c�")�jd�4��%cZ�8H�(4yu���ϱ>1TI�/s��*~f	��s���d� �f��rJ���0�B)f��Tf�0q�b&�Bah�!'��R�>��s׽���+�d�~G��I�����ͷ�����K��g��|=�S=��''2: �TAT�@G���j�� ��8f��-c� �NH�ݝd6F�V9(hD�4�� ���/A2T c���/�	J��]��_Oxi]ڕhyM�5������ի�\h� ��[d�?��c+��E���!��d8��>�Q��c8WAouaQ6nܔ�����y_?k��Q��yD��U�f��Yn<N�Q�#յu�j09�ćJ�r��L���!����td�Vt�peJ�&;��
��`����P��Ɗ,\�*�K����+���h|�!�\��{g��0 �nA�Քu}�_hR�y��W�����SP/F�Ǹ��I1\���Pq���#��J9�M���usc���Tu��ݺ�+��{O>:=���=ɧ�T��
Ս��iv�`�=&G� &�RK:H�~�t���x*M77�A�z�:�4p���}.��L"<��L$VZ��n�@�{����������숉�l��RD�G� �U�ό�0�=V�TU���:Mu�7VW��{���#�G%��,隁���A>T�r���DM�X�K�>v_�+G��?x*��qT������QY���^�7)��Y灬mnibq[�zK�
���2Aq��X*���l�lcX�3Xˁ�xQ�N�n��QĠ)�����`��eMd��ttl�F��`�Fp����w������6�����`u�(,8������*͇�IKfU�"F/K�@�3�,ĵTA+��ARf=Sp�b�\ޑH����	5��%s�mҺ��
�:����5��5��u$�Ѓ�R5���+������ͫ�b!��q��XR6�u[�w�š)j�	�]����g�x#>��g Ш�@?�H`�SĶ&�%q�(��f�<h8���i�L�~��Y�	�+������ܴ��=��]�U}}I���LO���%,��!�:s�HK�yR/�MJY��R���=�f�����yK�}�-YZ�$��	�G�O�i�(�%a2�T�{���胹K�B��,�H!#�\�	�J�����م.�E���ffA*w�U�bxs=a�Q��OΊ��'�o�,���9p&!M�37�q˯�D��EL:6�}A5#�-�DEt��S��\�.�4�_�K�9O%s��Q��U^�R�c	>*^�]4	��"V�39הtN�3yW>��b���5[0#���{k������e�ϒB�	���$�sjS�9�p+J��c5K���#e)�������2)�=y-�m�޼�;�?�J)�I�(�ׇ�$����ֶ��@N.p�7Q-=�Cې� _�&���E��gV� ����hR�aW���_��^��SS�aJEQ��T׷���&S}�M��r[:��"���2y/x.�٦8ol��'���6齡&$����l/�d��I���{����������)b�1s�[pafqkK������3��۲���+T���.���t>�N1��������Y��H���C�׫huV4Q�J㢍��{ѽ���w(	xb�媉�J��	+_E5-����[7oʽ�T�~�L�&��Yݙr ]�W�-����9SS��_N��HJ��7�����+�^�KmkSn��<��C9<��H]��xҳ��9�y�3w(�Lm0<Xi���Z�s��D�I�Xj�� ��"qR�~Q�{�0-:Jl	Oǚ�`H\��T���yc������L*��v��Q8�{	3�9AU &�s�&+U$�
3�� `��w*��3�W\/�_��VV,S���y�@e�`p�3�{��dyk[��פ����3�*O� Q�u^$t��@}�*���Z��a�|��*]y�5PS��o�����;��������^��$�� �aP��8��;�8�niB]�_M����eAhn��`��֔�Ɩ�.�H�^$eIeL�9!M ��5�=�>�g`�s�n^>'
%.�a��L]�'-i2�$�8��$YgA���d�ꉮs�Ɍ�``%�c_�W��`Q�@my�k#O|��c��ʜw(Q��]�K �T��	]ѭ"�4�R��Aft�?U�$%���]�t�@��ٟB� e��{�P�*��ozL�T�R��X�b�2�f��37P�[xx>��Yρ?��8���Fe�X\��ZgLD2�$!�(��@&���(:�,�pFa� f&S�iٽI2�'+�^.s�Y�����r��Nϫ�:5��8��y8l���=o$�Af�=�;��a���"��<b2G�y�u�ڊ� /�g�h� �,�j؜�Q?�JX��B��v��y|��[c��r1�5�~t�Q8���0�o[�n���뗚Դ_�SP:55/�ΔL�ͩ1yN�Ϝ�H�u�D���T��g��$������3�$�y��L�����{u�Pǎ�s��� I_��0;�au|� #��ݚGB��S�[�g�����e !p����|N#ʲ���L
^��	^І�Da�^�/��4�Fe�b� g�KX��TI7*�h�\ȺQb�huف�*\q㌴�B��՚����w-���&���<B�ǡ+2�&�*��둳.-Ȓ����h �/�ʥ[7ec��I(���� �*�'u�bx���&�	����/�^�A
�!8�RD��m�v�[������Q��f>�U�<ǐ0y?��;���^�ђ���^�+��U�i��(��cV'P�P=��S���.��ک ��@�lLi�J�)Q�,0���!�u��<�����|.�Ȥ�8�+*�ur�\�?�h����5����i�I]w��f�C.��KP/����
��TT�,~��k���n�L��#�)*%>�~��ڐ��<���;J�L��(=�Ui��\�Y�iF*�4��DrzҕaM>S�Gwk	�H�qݳY!.{�5��Uv}V���LdeO�z/6�djݮqP���3"z�;��zL��F�XS���1�?ԃ�y���	:�ǹ��r�qui��[ܞK�+���H��gLd�AM�aE��>��,�����M��L���jY�h�U�'K�HO�@.��5$8�h�g�t%P)�j �\Ll KcF�h�����P��� �訏���Y.�j�δ��M�y�� CL�� �H@Hm�䰹�'��=9�.�$�wC�b�od-(��+�Q�{5Gf u�9�ؽ�lc�Le��p(qɓ��/ZZQ�?����'թ�p+�0��/,� ��}��*��5ːX�~R���@t�7���T
Z��VW�,� Y��l�@���QA���.�&�Pfc��=�n*�\�V��Ll,��jHëj�͹&e�����Q�\���gq�z���g�K�)+�1�dT�7�5��a���.�ل�9���ޡ^(���u_i�X�d�XA���=s2��X�r*��ޚчr�����=i(iAPz��b3>��ieN��:J��� ��{R����.������}�.^O��)�=����E��?��w�ϋ�Ν?���=GO�W���$MHB��c+���)��}f�Q��[��fE^w�����	��<��rAH�^�]�d���>a�!�Yl&(�q���(yL~�v}��A^����\�� ^�o���bO}ƶ�Bw�;��'�X���t�m~�Wt�@U�I�%
���ˤ�����+O�DϴiKA���"�I�6\2�L�	�:b�qN�\�<(x��;�\\���L�Mb�)�l����3#������䆪 �3k�O�3�d���\ �P[Z������K�6e��5r��JD~�����Ϯ>pj�6r�d 5!��P�\���gþL
�Z�@VQR��\_ȭ�⒛�I�[Eѻ@�%	.����W����7�lT֟��&cUn��� .�˔r�qY@�dn.��Ҩ�e�������&�PAa?�8L��Vp��$^%�3 ��h�^9$�;e3c��
�J���'i�}���.e��w�x�T�Y�L�t��i�\I� ���rE������D����/��i��]\[O����u]������q!�)�
SK��*��RC���6;�J����8A�#b�����A�b��Td����s��t�T)u�{��*��ي��MvPAƎ��{hv��.�}v�H=�����Nb����2�����g6�$���Z4�gU��k4TL���j�X��� ������Y��r�6ru��WҴ{���%9>�)�J�Su�x�J��>�T��ȭaTT߭��QA��r+t���TH���iݓ	|m�]����q	��[�10�-��U:���Hλ&9��{�q�K*%�Ѡ}ST=�go�Avp�80(�k�#�lT�#���|'�T���>��_HN�y ��B�!5�Y�5r~&5|�M~v8Jf���T�\�}q��_yρo�S���1q=g=�J�l�J���bu����%��f���}�>fbBP42܏��L�uY$SY�����}s���Ͷ��[�
,��(�S�դ�4i��bv ����Y�/�g��^_[�`c�
7rv&�G�2�������1��p���X�����İ��ְ�%xnAP!��UHc���epx�ݾ��g�4�0P�FL:?.I�������p�s��ǿ�uq���1�����/������*8� �w��2�[�%�g��·$���,sBb4��e��%_����'* �6 �R& +@Կ�1�#��t��1�-;c�ϩ��.3�ޭ�C�/7 2KΊ
���&�:�b8>�64O����Q�_ތ�`�y����g���f	rG]�/$9�g'E�)��w�{�7�����2)�}yU�� ��ఘN$HǺ�`x4��g�.>�@˙"����j@�W���v��3���^K ��d����U�q��@�52�1���!����%�5�w�6[RQ���W�zC*�>��b�<oۜE�]��v���NS� �SM*:�?�����=U�݌dG߾Ԫ�ЙU ���P��X�Ί Eb���z�J ܐ^DE��%�}�Q��	�%*e���.�إ{��w�!���IBcL���k���fmsCt�{p��Y��Q݃4$j��yH������v{2l����-�;��oP0Bs�
y38b�$w��C	��e�sl/4%����Grrx(eM
���4� �P2���W0��S��R�Ԓ/\������I8����t$�)�F<��C�������vg��3�Y\�K��3E�z�Y1�5@е��H�F�ox���*�$�^j�8��B����h�CUg���%)�� .�c�T6]�C~8ڨ��Be	�{��c���p��攕\tkJ��ul*%�BK{���J*F�"��U~߳j)~hcM\"��QQ�6*䃳���S�����~�{]�؏��F2՝�1���]{��@��{T��@p������V�ٮ ��7
ǧ�����#
%Ě����H��[�U�Y�Yur.h����I�K����U���}դ��k"W�ϡT�G�%�2��M���
W�aO�I+lijX	37���C��y3��|�|6UOlh2e�)M�9˅����<s���g�P��Ō�B���"���M&3E��%݃����B����`|��r<���  ���O��c}փ��}�PpA���l̫1n�^(��!�	k
�ۺ&<sQ�&�<�<}D"���^�G-���c�>E��e���B�Vf���7q�Qt��o����0�
�c�T��.�[��Xw"�A�֝�����=�!y�����>��&�Yj�t�q90]�V�X�t(�,Y����ln�Š�h2Ht�2�d��e���9�6fQH�><EWԵ�����`�J���%�8�[5gx��=b� IA��g�xo�S�+M�3�~Vfb�&�>ϔ.۹���Q��wםZ����=tNr���k�H��d��n�^��Mb�92ic�ep�*���J!Es<
��Lup&5����^҇^��)^z�#BkC�a`"oeW))y6e*%9g
BRg&P�+���>�������C� P�&�=A���<��M��1Zp.���� aC��J=|���r�*�ଈ�>��K1�� �O[
�A���zD���e�,��Wī��Q �wTX#7AW�`�d`1� k��R
.��!*(6�mT������ݞͽx�����gz���DN&8d����#�jSV���3���6��4�3�S���B4q-o4���?�2$�bt�U�����6���x-�q ��G�z0�dt��GI��ֲ,,�88�<r��ܪ$ź!�pkI8Z��5�J����g�P�	��=W�d;�����A\*�4E���Ǽ�a` =ȜzO��@C2�C�����sV���D���D��-J�K��ԋ[ֳ���C�s�����C]���C����޼�8����F��Q�@�*�&����sO]�n�����X�,+��1�8�Z,���m�NTU�R�xX���*�~>�p+�Q@�H����0��h�����ީ���d�K�&�A�9�:��Qsx������� a������i�.���ß�$�%=�s|ntytT��
@����WP�\r�byFt����sh@��:��t�{I��ފ!��
�<YL��^�t�0�@C7w<��2$
���J5`ˉ�b�s���s�����?K�}ĶNڸF<�ĸ�X������]=�=��cL/�P'�g���d��m�k���=��\bť����q�l�/�o��+���f�8��?V�(:	.����+����b*6��Z��љ8a<�B�b��.~-��AM�at	�H뀙L�Q�
����{���^T`�Tn�{ �9���{��Nt�Ƭ�� Σ�0�Q�(W�ؾ�u�m�!PkBP����?�f2�pgs��5�8(�>���QAb�y����Rb�.Pa���6I0G٠�g��:�
�ptuSMrzt��.��8[dl�4��-F��f����b�w�R�{�N�,ɒ"ْ���"a������O�z���� ���y�j�)���}�<$r���32c�������xӌ,F�X��g��;�T����@F��X�R�[��d"�@^q<c���Wi5(�Y�C���]SЍ
-^�r�J�y�B�����g���0f�P.�!9։;T!��J6v��� )��j@̞J���Ԉ���.
.4�GO������h����%^�J)|#G���@د����ɮ!�V��\o�bM�VA54���
?S� �>σ�\�w���*�yu�C�����%�j���.1wm�R�s `�{Q0Nب�|�]@��*����.�_�>B�&�W���u`ʐ�S��\1�g�4$��S�I[9 0g�.��D�h����×b���啾�zt��H��
iO�qJ=�);YE)�u��a�� �> HQ���*�~�&���뿉��r���s�ً0�uf �����'C�p�����r:��r�1y��߂�o����Gs���!P�P�Q��_�X2F��m$�3�]��(����W�\���fK�EF�6��<���̇�i���%�,��w>�1�iJX��~Ȃ�_�g����i��n��9��\K�m�漿�ދx�����)A�����N̨H"Y4�@c�E�ߌ�;����h��5+n񋃧�����F<��X����)����(f�#��gB՘�fj����6���CG��9�-��u���:�f�*s񜋂�<�A6�\f�b���_�y0x%���v�K����[��9 ��Hk^����ԏ��No?e�ȋ���b4�Ϋ��s�=�� 1u/b;�F��Xjj&&�Y��{'Vyg巘��i��FϿ %[���腸�"*�|1�%��B�������a���g���|����3���%0���]��y��@����1�a $z1*����$����K��s!�1r�4�e�F�
��pPϊ�xV,c��m�
E;h b�_�p����Ɵ�C��S�NXNY��]1��g�N�Ιb���H[����܈��L�S��S&޹7b&�� -��/��,(��N����Z�*����2)�}y�˙�	���@�I�#�e�f.�-��U� m�0}N�!t��������q�cݣR�ja���|����q}Нo�[�Q��ʦ�1���tǥ��<�:�W�?U�>��ت
ŐO��Б���^z��-���,0��3�^ЇN-Ya�Ԇ��7S�pQr&=���i��,2�`Z�`�d'.4H6�i��/ݙ�	9v��#�[���z�~�Ӆ�	�b���L}��f*Z6@;�lG�*���9Z���pq)(;l��_�Y��x�F��b :��0���:���*yěd��F	)�k��C���
�ȼ[��ie�y��Qs�����	�3	�-i
|��b�������:�^��0�.���aM�OT�P-Τ�����%�}�ܒo�c��+���<WMx��p��AS^#��d4"8����%�	����{��Wŗ!~�D?�x("�7�RѤ8�O��h�
]Pr�����,q�U��{�~C�<�P�u
U3k����c^?���ۿ8�K����Θ�@�!ɠh��)m��T
MK>tz8���9N�7~1�(�J�{��"���t�����H:�zĹ��8�\�i] �ʩ^c����H���4�P�I3f` @��ph���6<�@c{;$%�*(�{��zG�2>?5�����t1Jgo2s��4���O%�OI��	��S4-�b2KZ/r��¯�LA�p�PlR�N�P6���a�*�}w�p�S���g��;~�T�K����j54��{}Y�Ae���lH��A݌Z��S��h<�N)�9S�T������`���:�ή慟s��W��qa����c�U�̑Դ�3Z�w�P8���.;�;��{x�Z�,�����Qt!�?}Sֲ�s�� ��\���HH/�I�T��@�fJS[H2�k�!@��[(�]����>��<���¤ ׄ}2н�%PI��<�iz�5U�m~.#R$*�8ㆮ-fo"���s�#/4ӼY�JC?&t�ys�)����c[�����\���%ě�9�w�?G�9�3Y˲�i�O�z�����r�0��b6X���o�s15��VO
�A[ԙk�{�kr;Ly<����{����E��5UdJ����r�� ��%vׁí\	�٨Hm��H��yWZ��x�9��r�oUQ�p��o��M�x`��	0�i�����ڎ�f_&���@���\7E�t���^0ӑG �NF<����I���ŵY�-��Vg�������~�3RrI��(?�ۆ��-�&3�����t8'@��I�Ք��P��?��Y�h��A��y�oV�E���< U�MXV��� ���� ��Լ �*Ʉ��b���Y�R�NP�Y]�x;R��~���*b��|��`7��]2���wԻ5�*2�h��T�A��b�3)��֥[y�Z�HK9.�͔E4�NP�:S �c�8�8��M��n�Ӷ�XY���$q��S��Zp�؋UMh+P
�I�Xyz@����X�:sM'�#a�����]
8'�5�M'Ҍ<&Ch����E<���r�.�ɮ��x�l��`�#?���~��鰯?2��F}��+x��1e$&Δr�Xr�{�x���iv�u��V��4C��0㐷X�y,�W��)�b�#�4O�,6�eXq�4x�$���ϛ@<�u
:�����V��j�Y����qȐ��a&���+�ʼ�qh�ʍ�*�2]����@C��B}��O����L(�Ab(����؞��W:���y�k��ׁDk�y��J�pE�KD��W��'76\)�.�A�0��g!�W�p��]�Ώ$��
�M>�/�E��w��X�u; 5��ɯB�j��n��z$K��0���=��3k�j�93�(� ��_@����'H�8Ӝ5����<|��W�]�̚��'NQH��^���]���ٱc2<:��2��6��� ��T��7��6c{j�jMU�O�����gM��[+�i�����l{�w o�p� �����	X ��:@_7w�=tއ�����.�(�0�MS��zk:��ik���g�r�o�����w�6�J������l��V�l�����TelX����]m�И�0Lf���H����c&���L|�}��c·a�xxx�I��j���h���j�4�g�Y���\d	V�7��G�ܨ����p����x�|�m�x���U�0�v[?!l���L\[w3X�;Z��R|��@�w54�0��j����;>�A�Gr�����Ϙ;n��r�X�)��-+c:���]V�NO:n����ݤF�;*�N�\9¾M*f�Fkx~J�e0���=�$�qV���Xj�.W��C��Y)s[�Ǟf9�y?ʭy���J�iG���i��L	�c�1�f辰rsà2g�vV|��S�yBK�f�}�m�T�Q��)��S��qL��J�V
�@ʝY����\[y��R����͙u�,����)�񱽻�k���D��;96�̓O����3�X/d��A����/%�[Y��@ݵ{�9��Zq�.&�e/dC�aS������1ο�a�������x�ݭ/���˜�G![���E9[�����kw|$�����gE�p������=���U���虌�rx  �G?�3�����q�y��@�-	S�vw̵MgR+��Y;�e��e��˔�����h��ƻ�v��s��9�]@�,�":W6�֋�l�si�Y#5D��P�VkM�F?�i�v4I�]\fRo���6LTE#5հ��	�IG����.����,ik�6 �T8��;�J{�ߓ�h����n�����.ۮ��5]s�������/��X�J��3
���b|�z2FX��05�yG#sw�����&�%��%G[��Fmg�4��d�%�\Ju;W�������'A�Ϡ�a���� LT�%��XT��p5�k��ڣ����*Y?^;=t�J��W+�h3�`?7���dvq.Η��5v�j��{~(F@>8�f�}���׏`-���r9��'��CYVV��ݷ��p_�R����'MB�"���b � ����i"!���5��P�8`¨�jmX�A�*ّ{��\AbH��e ���wm.���K����Į�nBũ��|���vC��]���S����V�(�o�`����|ޮ�b/wWY�>x��o�������U���șo��Tt��He��"���?�I�>���*eގO�ڬ��T�.����Q�!���{]�tc�u�'c��=C ���:ߩ�E��h@��o����wA*�=�OX����:�~`u���z�b��Tm�&�Gx�!S|���+?_��Z��e�?�])�����#ܻL�I�UK��=R��!)�����|Τh�����8�Iw��j�V�w�,�Qllʱ�7T��
���A��}O����9MYc/����{)G�kV�
��q��!Nβ�4J�K�;�d@��vͭ�_XV�$?45�P�+6+��Y�����{��S�-�_��(��cCO��lW�ͬٶ�C�E:d���z|�!��W��,nG̔,�#]� �KS���L&�SS��F_`2;l����Ҩ�go�җ*ZUE3�@�6V�xk�Q%�'#�J견wj"ڣ�#�����J8��g�0�!Ñ�g������J�����훲�nRnG��sS\���D��B�߾� �'�ף�@|+	��%�<�dw�+;�o�zf�m<���"0`f��iȁ6
�|�./a�����]��lbW+�;�H��4[K��m�@��H!#RGb�XMP�'^G5���TwO��Jg�\�lS5�w0�{G����͹,����@6q�﬷6Iz�;Aw�5]�J{ ����`-S���r6��>�|���N$������x`�����ԍ���m)��s�9� ̬R�Y����Mh�n�Z��Y-��{xn����ă��B0N��'|���}%���H��d�Nљ2�׹�sg����>�`�A(�g���oTMK����^����Z�lw?����\�rz%�����K�m& ω�Wit����"�e�>m�w����Q?�g�T:�Gv�A�QH@�MgRb�&x������*��[f�6��v�||܇��L����;��J`����J�0eW��Lۏ2Ɣ�dկ�԰ �i����������M	 #��J[�Zcg���}:�U#����k~u%'��$�}ێAUS�	��+��$�����X�!VInT=���:S*�<���sz�vs)���ܾz�}�᜘��
��T����l�wC�0��R�ǊN/Q��j�׻��Y6m8�~!* 1�Y;�\�Q��{�wA?��h��~#S$z_��4�U�T)3�r��k��|m�>���ѱ>�ڇǏ�.��[��F�7z�N|�}��Yoޏ 6
���e�w�d{�艪�� ��m℉#\�&7
'+ܮ����{����(�L�y�~��O	[R����B6�_�ç�?~���Yy�I�
�1��u��S��:[��.��9�nJ4��*��Ѽ�k3J
�*W�D���]���v����BMt�kӼ{/3J[�u��))II��w�/�݀�]ٛ��ٓ�*�e���ݥk�'<�A�Gr4�P�~TQ��`�!���6� ��t��R�y�EyXMG��p��Дv��P*����W���`4�'`yѫ�bl
�[e�}��8�	��� �?���*��b#C�)���x�\-���5��:�R%9�,9n����[(v@8��+8��֬(A�m�jIW_Q'�EA6Ĺ�����
�v9e��u�Rf�U��2!b��3û�N����"�N3�1���f��Ž�\_���R��Z��������4OFN�~�(=C�������0�l��q߹�s�]����=-�g�Bb6�j"��BUw�t�'Ww�
N�"�0��{c�u=)�Y�\#����Μj�{�mV��&Ck������&�8A s���Ƀ��\ �%�Z��*M`�v;��~�:�۹����Ze�5џ�7�$�S�dЙ-g �[��A�
�m�z��S]���{>�>+�GK>+�[ @�!�|�"G0�j�nIi`��!]�hf�wM�;�`���!��/-m����kVs����
AW� &�Z�o�y궾L�T���2�������]�a� �/�9g2T�
��|�81�v��}���w���e��8U
+*�Z�������[��7��hT;�sg4X�r��m�N���|*��?S"8(e�J3p"�*�03��~V��d�v
`��h��`� NƳ������a�b �!!�k�	�ㄕ.���#��R�D�@X��v���'��v����xy�{�KAa&O`_����'�P��r�?����&����F8�׸����Y_�IL:���B[C��P�!��h;I��Ke��jGr��̦r��;����Lz��}I�H��U� >[����eKw�]ݰ�;�G��l�=�(������Y��.d}�Z�}�Y�{%��#O���i�q�	���o�F���Q����8JT^�J�z�w���p�Zrpu1�E�TG��;P�5$s�P�ɤ����>�jS�ͺR������A�-L}�]��F�3���h�K���]�^��|v�	n���A�ͳ�;@{�@	v�AU�8�Ta��M'��%�&lB{Y֨ǭ(PV,��Nsؘ�S<���`�V���������m)�e��~kϠ�\j���L��Wr;���������O���ݒ�uiI�iՏ����Th��k��`"O=�%|v�7�,f2;}��A���,��kj}s%�f%u���VJlaC3o�S�i<v��4��d�Iq�l�:��h�ېz�j@���gE�~YR�&(B*�R=P�w�.er7� ��x��s��-����5����O~����8:����6�}��~6�e�8]�T��ˀR�4i`T��N�e����x�Q⩱g�Ч�uQK��Ó{���������d{�Sߒ�AU ���{��3p�f~��L��0���l�>�O?���6���� ��� ���|5�AGsv�C�ңw�Ā�bz+�۹ X7pH5���h"��ק )ӥ��Z&���r�u�P3t���* F�t03�sNN��9 ���rx| ��(H���qăN�1��+zڤ���}"�V���r�Y�{-�1}��ڻ����fU1��:4�u��&�`Y΅`6�DP��\~�;~�<{p(on� D L��� ?��BC�M�4���N�JH1�dI�5�=�TƸ�Ó�<$\�ȷ��Q�rO�����%�+��Hu�L�X�}�UѢ���#��Ͼ�%�XO2\����j3_kF�O)��)H�鿳b��z�����g��zk<� N��R�a��3���A�:��z�d7\B{Ip��^"_��O�t|���jy��A'E�Q_����s���/�QgA�Z�`�fg�Fz	���6���}�w�.:fZ�����$~jJ8�����H{=���s �3�Z�dRߪ~ڗa1�5�I����!�b�a/�3����\>{zO.3Or�tа9l��]ZQ�NP�5�7��=0��9�+���~��X�����d� ������#��[�;.w���co��oA��q��U�zJ'�����;�?ӀC�I l]��p͕j�Y�
��e�t��^Zs4���g|&�h��'cP:�஘ͥ���;?��#ܮ���T+ ��'G�Yh:��&��p������R��s�#>��-1u���4pq�6�f?I-��RI��a=���D���8�[*�=���C<�L.�#�DxdE�Uj�UR���%�p�Gf�=�+"�]&��/���sڈ�ȳ��Hf�{A��:�^/R��L���uH�4� A����龜ơL��b}���T^��ey��JI[�|а�U����>	�[��{ѧ8��ø��F��QR7i�X��Xr>3�|~�K�m�9��Ym�J�\��cT�>�t�qb�V��'
C�e��7Z	#�l�����<ꨟ���lk)������y֠�$]����� �=�L��u�U+f,��UY�|&�zi(9���U������i��3}�D	S��X���0 ���󘀘pP({1����T��T{��23e���%�I-���!�ZwE�}��l$�7��[|��?4l.��B��q��J<STC�N�R��k4S�h��t+�N��8e�b%o��L�)�Q����Ȭ���Ky���Z!c��	�	���CKm�\Cb���ɣ.t��O�d�  n��j#��J��t�*��8�隤`?�t�$Jm�2@~�l�R��ӹ)�	�ג��5+ܬ8��5lz�����C���訜��R�uL�ɧi���6g���sV���FLyM���l�8�30V�lth��vwJM�Z�d��)���\-N��(�q�B2�M�!V��'x4��[-e�����e��\..O���P˼��\R5#�N���r13x^x�̆����jC7����;~��)�
��>�Y�z��d�n�q��f±ڬ� ��r��r}���K���J3��Z�Y;�C��������b�<��G�r��9 �p1g�(��頣�L�VrH1n
��ε�K�[^76���Z]�.��ҍ�Y��S��x
����#��'� �0���+r��ݥK��*.ϯ�L�oj*\���c0W7̜��[�����Pz�_\J=�@03�ώZSJr���~@֠�������cY��^�q�s�&6n�zkH�/a�fش��(�>� �kY6S%� T�M_��B��kDpn�-��ϥ�/$�������n��]n��TiE�6.9�!�.�'��l�_Ks�N&�}*��HΗk���(?�}gv;�+����ZK�씨�Q�̏�Y�d6�J�B�=;�A�{�Z�g�n�㖈�}�ғR��.Ӹ�۱!ո�ʣǳ)�fy�}{�?{"/�gR؏p�9�-��+W)Ma '[�Vt�� ��H���-���x�� 1~f<���>[�13�;���A��5�_���k�����R�6R����b��Ř��ͪ77���;Iq/����ٰi��� 9�t�.e�!o��h��X�Û�*9��A�I%�QaD'�,�={�`���R�;��3��V� :P�Ͷl0�hPM5Vv� �����)�xFg��������+���>f��Ű��j$����	X���B�D�Z%[�dܗ1�[�L_� ����${�F"�;T�G��I���]�N7&h��ж����a�F�{|���2:�'��r8|(Yʶp:G �[%��J�;P.�̻��*e�V�k�8�7l*��0�|������s�N~�����,IbmJRc@�I�X'�������A�-��ZV�B�IjUB�K2h��U_ߌ7����������~�?���3#�
�"�T��ǉ��Ʉ�#M���	�/��nz䜛�2��F���p�"9�
M4�� FUG
P��z;>gkC9@�Zio�RmC��?8��Y�kP@�&���a%��&��$��V�H��MɈ���*�S��Кt��hpZ���1]��>(-d���'	�#+��Q[#��x��vG��l*ҿH�5E�>�k�u��]�lV��zo��Ma�5�i�&�1h,$1���]���+$'���|��_�n7���o����h#��")y�B�V%�c���I"=���c ��F���S�F��r��@c}�C`�(4�T�M̪X'��|���I�#1c�g�P�IT�c2��8�����CpP���pr�����*� �� BB�T5Z�)��Ӱf-�����(u����NT�A!�/��n�_��YR��ľ5�Q��Ɩ��w&}I:����K��������c)>}*_�.� pVظ��4�{,Z�ڂ_:IF\Kʌ�
{��Q�j�%��ess��� *�!�wy%7���ju�� t�yfu<��oZ����jJ8��`w~)��L����''��+��:������P��f��~7k���]_�vd�
Cz ��c�~nH�^I�mEf72=}���
�l)޶R�{�#AI����+(��Q�������M��B��J���2>~(�y#+�l ������&~O�{J ���	S������2��,�s8�Q����sY��F����W +p�0��[j���Ô\�Y��2S
_���p
����޾��M����M�sB�Pɫ,*8��A�=�F0@����t.ޛ��P��Ñ�IE�S�����ϥ8�D����|� ��mM�)�s��9��+���Z�ݵE+3��9`�J������a(כFf��dg���h<�A�5�(%���[L�6��y�X��E� �^�Nl��t��\�<�go�ƳK�Z��y;��QQ��V5���yԤ����R\cm�~.�o>�	���QOVxRF�`��j��I�^7���@����1�eۅ6��̎(�������*-esu&�v-CVH�Df��������PY���rP���(x�n�Z�������q}�=B�(*����8ٮVu0�t�#s�6>3xa��n\#%+��U���)>��D �������r�ð��s�_��s�) �u�k��6��?����d~q.S���o�3����L:B`Y�<P��O9�$�z
{U\@A���k%���d��N\!hY�������͋\����<93����O����G
��]���0�՚�%�2�湜���&��b ��H�$�I�E�j �4�!��>�3��f���;�=#�ܞ�ʫ������^�3ؠ��7d�>Ezn��N9F �J *K����7�l�a-,j�x7�ۛ��Pm�U� Q�둺�+�HgUtt�V��=�S��GXs�,a�'�' �k�o��j�^*?�$���7-~^g����z`J�ƓA���k��Q��A��V�Z��C܁�Q'e͠`GR.�g���껦�Y�P+q��\<V��,h	N�g� %\��7��t��H�$UE1&OTdC+���i�@Z�
D�::V�i]k�`/q�w�@[g$�JZ�6�[�O)��
B;9���������">���$ĺ�
�E#�P�;3�L�� �YɪZ�מ�R�=x��K������J�Z����j�^<��Ja|��{O�&x9x%�!��Q������u��fX�ڱ���dp��ʼ\i�f�ʁ�f�*,�IV�8��-�g��^k�'��V8���6W3Y��e��ҁ}gr�0H����>(�h��kx&A�k���a�����5�9�6�2�
|'U�i�@bf Z��R��G�4���Q�H6�І�t�c)K��5әj��	 W~u)_-��}&�ů������Z���Ҹ��P��H�I����h�RQ�e�\�,����ֲٮd�O�O�X�����w��<��n�"��
��Tv�g��`2��#��WSi/a,�r��O�O����Kys����i��ƄS|����r�I�bФ�C}/D!UV*_~p8�" w�:
fg����������g�u'�L�����o�MY|�akԑ�7C�>Qk�f��%��r��_�W����s��.uR�c��Vϰ����l�S�Nd�Xㆤ*�V�������˓�9��˯d��o�:%���\�1S�R�����s�Yɷ�p3�]�w毿���O����RKR��5��|�60�K�0�zuuc�jT�"����ʇ����X�s8�Z&x�jz+�/_H~z�y%�f`%���[�67 �n]j�-�a�ZUR��0����?��\�䓃��>�B~����b&� n} �΋�L"�u�w�.�n8U�m/��vv����/��oe��ײx���F����tn������Pv�*ʏ�!j�$
����ne��y9���g��/���V�,Vk��I7�<Tڡ�>QY�.���L]耱a?�1�K5��R[��5�m�� �o5����u7�"0p�#9��3^8�y�N�ɱo���R�_���O�Jt8��Ү2��F6֔�� � �x�C����4��P�����V?	�FI�`�����؋��%"�L��(��:�Z�u�}��1d&M�	��a%�7�Ɇ�L8��/�v�	�'��(�K#8�k�:e� W���8蜾T6)�{�sVn�� �L��F6/�K8�ɀ�K ���׌�� ��!T�N9-�L�R۬�n�%�z�'�t-�w/�?���}��6}
@q��:dJ��Z�3)U���g� �Y���~����a�"���/��V�w�`]�:ܲ�
,�9�G�R�L&� � _ұ��G��6	es���n��>�,��Q�t�H�$�
e�s�/��pkS�=D^ �����8յG:ē�N�ߨ`/��������������n���:�c@�-�� ��m�{���w$8�A �ï:��*�]�r�� �FZ�+�l�7{�Ϥź�P�V� ̾� U�\�ͤ��k�K]K���3_��ae�Ɍ��g�k-�DP��K�5¦�T��nՎR]��E�o��h(��t)Ғ�}>o�T�3�X�ᡌ|*k����������۫����8]��
�SWiw���n01k���M*�[Ӌ��OX��,"&���Q����P�.�z�����A"n��{q�π��d#祐�F۾�eu=���o��
�QQ�����'	���\1��j��'��&:�U�1��p�G����/��R.�J�#��C<���^a �;�A�Gt�Ax���k3�j�S��p����{fVU�"VЯ�T�u��g�ƂE3�Nw�^'P��[A���O��4�����(�$R�x�͑��M&���4�9��[��y<}����#�)���g%��Q G�W���ӹ�)�N�y��Vʉј�.�evs����'�`*yw}.�/��_K�oT��Ƨ�NTh��gY&�����S=_�Jv�F������T~�d<:�+ ��w�rَ 9�]3fPvkf#?�Y�` ��z�%�C��	����~@��,��V�����5�"�o�P֐ם���!M����X:��m6���d���<89�{?���rv~+9����W�=�  �����}�lq%�
k�yf�
M aq��*�,~�J�7ߋL�)m�  L%�l�eW'�TB�N�_+α('UՒ���/��ky�����ny�_�W��@��Bn�zWY#p,�,�p��C@�s�$:쫒jS��/d����'#�?Dȅ�e��p��7�}�R�I��2�CsB:��τ���6���g���Q9�p+8� |�g~`b����O?�L������~#zqx$GG�J�⻕�걢�2��RY�M8�������_~/��oE.�$�J>��@�=+hz�^����m����S"����qW�d���� ������K������%�#)7�8�_����H0��M�6/"�Z�#3��}X!ؚ���x�7������&p�k�ф���@#m����#h�C,9�ꫯ��s@w���Rf�ƪcm�OA�3@=	C��(ZS;{/�'&{�a�0&��ؓ�+��[���⢣����� g-0� �����+)����d�ɏ���Xɐ���ޜ�e��l����%x� (=���Ke�x�w�`��Z������1�.p^�$�:���W������<׬�`+h��٨䤯*W�3�B�`e��:_%nc�"Ϛ���I%y%s�r+��k��L��	|Ǳ5+�$i[���IɪH�ʚ���WSܯe��\nߜJ�ꅄפc�P�Vيt҃H#�jt�!�U�ǳ��d��"�7&Wt�E�I�]|EXP�e74��5��[Bp�������ݡ��www�n/�������nU�E-�Ω���~̒>tPI�n�p B�7yD��e7"�(�P[
#�nAA� ��Kz�^�;H�'�J8�f3�Q1Q����&�#\�FHg��(,�%��骤.	.��V:vT�!%9�6����_���H����~��
le`s�p=�U�榛���?���r��3,��C�=L�k��Hc֘�r��xF {�{���Z6�/'o��a�� 6hONz�r��\�2�s�JBLχ%��kQIܑgs�f@]��C��6\�T���ۻh�6���C�0OD���Ȍ%�K^��7.ppxc�Eo�}uv���j?�v�k*��=��-�C�L*�ӑ#�I=pb{՘?;��Y�#er�ͳ�%®"�U��})�ދ��ˠM{̤s�'��|yˎ�A�M|����^㚽���3"�!!��?:�p�o�Ȟ+t���N=0z_nݏY�ʫ����Oʔ9K��]�7Q��;�`f��QIK����7��˹{<�sG
u)�a�� M�s$�0+f��n������Pxߛ�r@�y�aQ���uP>��^d )G��>�j?�aO�yG�g�ؒ�2D)�P��'҅��N3q�3�����'�qo�*6T2�����D9�F[|�bߥ|r�ݽ���R����Τ�뵖�+	zHN��:��L~�7�i}��mLi�e>��:qe2����OlJx�k���į���?=��XW����o��s4���Mty�)�P�qO����r�x�d�����Cc��U{͊l��?-f��/��u�Z�"����h�/�-����bӋ����$�pS%�b��$�هG^vl�n�p�\���v�T8� �]��b}]�r�Ϛ`���U�$�]^L���� 0hZ���B����s�U� �"�e���O龒,k��K�l��}�>-�3�J�@O)@���G�f���Q*�(��B�}9+U���(5.?�"���[�|���?"}�k�$YQ6/��tw6J�]�{NLt�̆I�kG5�������B<W;�'����g�Ph��I�:��:w���+�Q��'TH���N�:z�h��ӆ39�?���K	� �������Y.S{�ȳ�C"@T	o-W�����Y�Z���/�VE3��_G|�\��R-5�����s�+��8>V��^%G౑��ڔ�u��>�ݖASޏ
��x~�V�,3'ɸ&���[�l�o�)�&Z�q��Q����*�KI4� ���i��~Izg�PV_���~�v�:+2�[��Lo#��Q��S�� ��7R���u���WЇ�o�+O8<#��[p���)����^�ڈ�xeޑƆ���߅A�Ӻɒ_Z�üB��a�e���p&��d��<ɇ����ާ˦��o�#�wd�H|܆}�.���i��w�ʥlH
i-�Gv��<�2�M�M;ڣly�`-XC����2)���}���Ya�Z��Y��#�y���?-�ut&�������f�_��%�'Y���&Q^4��&����3��A��
��Pc�S��S��Ӭ�-�O��Vj�E�,n�� �om�A��w&@;m�o�5�	�Ŀ�Ԗ�υ09ݩ�Zo�*��U(;�]Ta�\o0���#6f$B4�
|&%�� $��&�j"��	�0ph��)�l�>\�2�a]�X����¼�/���A}RW�2���0��oud�ɘ�o*���1��v̍(P}�J_?�}��V*�v]�F,])XGb J�Ө�1}Ǹ��`���y�p@��D��/)	�a��5�-ex�I��#(��˨���!�	6��b�ot��0�/u�x]t��m&�y���&�.�!�9Z�ꊪ�/�ATϾ��g�ѽ��Xì���~.>kˑ8��̐h��r�?��j��%o��GߣuZ���7�Ɜ�����}t��:OqFͶW�����ݤ˾gc�8Ы �������2����[kP&�[�x�x�i(��)��3&}*�y�/�Y�B��7_�?Z��һ��˜tF�#�i%zo��,�.#���m6%����Z��ω�����H>�m�}�M���^��
*�r����.x�����ҏ�/� y	�_�g��x�.��D��WGM)`��)"��zT�?t(�"�ڳW!n��f�&�LJWV%b�H�?�8��|�u%��VS��I0��)=ƩKK(\(�A�m��wN0)L��'�x��/Ѯ�j����߆~Ǎ���6[K��W*���E$9[k���H��B�^����|�7.N_�]��-&tyG[�I6X��Ya�D�d�+��ܥ�UE��^t����KL�;p8� �t����_�S1v�.Q�������	���C0?3������z �ƃLM�-��)�+�]wq=jt~��sE+Kǈ�T�nW���_F#L^W͚���٠��V���ˀ��ߏ��������3}������!��~J���x@r���q�����Ӭ�����QBGw���aX�����g�`3.�!�B��?��O�I
�}��2�nN�O�%;�O(G"��2�/�oc�%Q?i�Y�9�M{�o|9k3GWY�RE��L215H�����ɵ���TJ�a�0��%v����<�eYo�K��R��.�.�)���Ѷ�M?�>������y��<�7K�}&��x�j��<�ȑ�����W9������[���2��ʖ���N҇�(��GG�*%��/B˺���N&�H����(ӌ����qҏ�@r�Iu�z�<��^�}�SF��*���;��WxҼYf;��6��js�#6��?�` �P�^�_rU�"-8`�[�^�4�?9�������M^�UpVz�A�<_R��2�hJj����o�*!��ٟ��&-2�"�)S�w�p>~�]c��������n���K'Ի�A�7�tW�O�Ih��d"�
1��^_�q.��b��h6Ջ1���lJ_y�^]	���6��݊}j�4��V�O(�2X�cU_�H8�ݴ��j�� o_	�{1���I
�k(-P�4(���<�e���c�f	�⣷��C��+�v+��a���O�*H����=��+��t�* ��Y/Ō��NNY�w�)L�T3��U��v@Ft�.>l�ǩ��Ͳ��3?<u5t�H����,�&@D|�y޸S��%��_U_��ޜN���i�,��!k�6�h�V�a���n�.����?�+M[Gqe?��#DҖs6�;Fw�(����|ە3K$h�`*���yc��2�1wbh����_�O>�H�BOXȏ�٧��pb�ej�ae�D�9m�Lr	�<�iT�=FO�ϝ�5?�%�v4��������o�V��_%�����cè�,�-����h��h�oVA�vE���E�)*��2�ڈN#�E@J������h0�Y��`qoՙ�D��,��[F��4}?����D�,�d)8v��u꽓�8�x6�8�1+z��y�[������h��R}���6my��V�>�ʇt��Cs��B���}�,��U/6.
g�q1��,֧؈��/��؍{�W�"ȧE&��|Ȋd���e���e��;L�M�sa(�)N�;C�ri`(^a=���?����H8;r,��Bw���*�ae#�pfY���?$1[�n��i�d#���(Z����h����P�9��(
�J4��C�;�̓������}d
a�V�0��I���Mzv�V��o�I!8lV�ِ�LN� ����t��춎���O�a�=���T�#uW��c���a����vL&�7�ZC��TB��e�9�6���`>8��!�U66X�r]oj�'t�����<	l����O�4<�bB��S�hO�ȣ!���oN:~{P@'eX��n6�;����x~od?gx�/.:U9e�*E�֌xێ|?�F3-A,_꼟`���_5I��f�Ӭm��8?2�v���>t�Ħ�9z�ی�qG2n@�|Pv�)�Wl�V)-�<����!����7�y�˅ґ"l�=��:l�eV:�hoΏ���&�����l�����[��8<��:-T2w*=m�v\9'���K���V��!�j���wk����O_OdS�8`��s��el��x�o�
�P�߂���� e@�Nt�X���~5���Y���awUw�>D�r짦���=�>���{5�׸�c�D��[�7���o�J�,�?M�a��:��z�+Az �=	.Ҷu;��oM7�I�ʠ��D��݂�&��r)D�¯hN�zqq��+;u����M/����й;㺂kv�@�3ǁ�:����R�^W��w5��s$̹i�6P��ƒ�oׅ���m!"�E��є�l5PŪ�n��T�.Of9��P���i��c�#	N�p�sY�=��MES��V}\%8�^�%� �{߻�%}��#�
꒡���v�3�Y�w <]ry�O6��$�R��B�ŧe�Qa�~΀���v�h���=����/lg����󕗝��nQ�N��_���~Kb�N��,�P-h35���ּQo������<LL7��� M�E�*z[���z�b�-�r����	�&#�en�#}��E�g2z7h
�툃1dY�%���Kb',�&o��ı,>W�^�7'گ��/�n���=��>y��q�dOLY����B[��f�ٶ?5FԂ\�`����9'̊�J�Ԇ�`E���i�o�����{̐X�i$�����4���)����Y�=���=/�u����6%��di%�s�#��i������&�P���h=�n]�~4�&��^c�c��<��7��u�A�ߘlޖ������[9����sf��ѴB{�{�D�Ϝ�A}^5<#�����l|�p�9�L��9tWQ��*��+s��Ëg:ڡfE� kz"�ʦP��.a�n����R�g�5�������ӆ�GF���E�~��L��V6�ztո��g�׋�d?z��M$c���˙bb@�w���}�Q+�;�J��R`�e����y[�e��:�Fڴ�������L�ܟV�N7j��9[���W3޸`���A��|�׶G��PqzE�҈# 
X��mm�]������[¤�ȸā�4�r.��ʚ��b�}��i\���W$5��U�@���y=U^�"#_�l�������8΀�ҿ�I��z�����,��Xn��w��:�����Րq�8E�Wrf�p���%��S�V�Ɍ)�"f����ґ
it���i�$��F2��K}�F~�T��us.�;��,��wa�8�@#�T�}��K�S[p"͝O�:��,-�n!���ٟH#���z*@�0߄��Q�	=x~�q�h"��6��b�\mo�`��k�)'�����%��?[�.�[-�Lg���������}4�]��������L9�1<]Y�&���~/F�$��e��o�I�s'����W�'�#p��W�/15ө�aӅ��h�����c'�q&E )�2�,�gn�iS����m�R�z�}tW�SØ�I�al��,�|�+I.�K�^蛪���|`��ұ��e�>�]�����i��	+Z��p`T�n1�*^2�/b ?HV"�p��=��h�3��f�51���)�[%���~.�R��-�~ʶ�8[��g�LLAn�>�R������k��@K�R ��U;O�c�ھ����4��DL�ط�T�Z�>]����.��G�O���B�j�2���tP�/���ǅ@+w��c���RO�c���j�6
�Ϸ/�5,�[���}^��#����:�Ը��,��r����o�5��-�C���j�8 ����g`+��:%x��7[�p.�l?��?�9��g7��T�@.^����z����Ȧr;H|�ʼ����5���ORzg��|'�������Kձ�Ї ��ǘ��!��:?F�C��+�#>�j��-̀��>*��ff��		b2ݶ���綋�beF���:�=z�������,��`�@�|;�����opOgw�w�ke�ijӦ����CA�ߓ1MJ~zAy51��`��FCn���]2�k��W��v���a���R���SW�}�M�
$�˅V�*���.����a��q����܎֔�}�����N&m�G��~F��Uۿn�������mh��A����}Wyd�m�i��Y��B���3h�iA���{6��]"�g�7	��sCP}\h��jQ����k�vQͷ̓p�`áM�{0�kx��R�Ǎ�����D��#Q��|��TWIʛxh�1�Cv��,�r�'b��yl+�%�����]8���ϱ�tRlu�>6P�&�d�ӑ�� 	>� �P��R�S_s��9%�pb�6A�XG&�s�Xc+��3�k�P���Y��ԓ�sLr�Ѷ)넴4F!�4q���-��B���ѓ?�:�_f,a��M��˗��z+�9P��F5U�c��ѡ�a� �0v�$->rضS�
�׊���O7�G��es��V���j�%��Yz2Bc�OrGO��?�oF>/��c�K] k�rG$�EFm�.�@Y�HHy�ߙ��Qҗ��R�p Ux����I'���D�� *&Y��Ґ9v&{Y�M���x�g�%�&/G�su�l���JА8Ʈ4�E6�وU��7�f�������$S��7o_��s����8��Zi?k�S����X�Q���D}��5����\]|\�̩Sϫ��j"
H��E�(`R�Փb>��}S��_��1Qy!�a�׃�S+5�a*>w7g`� ��q���e=�Sp�t�qB�*�c���C7�*h��6�Q��b�6I��w�{��Fny��>�2�Zu$X-?6��ZXx/�0Χ��l�k��xU���*�����z���,Z�%57H%Gmp!$�Q�-�Y�nT$x�
Z�W��෪�D��Gnvu��
�T�	�"����t�݁_*3��܃��D=�)��]U�VW�����\�I� #e�Y�����S���'��%�b�y���/j���� a� �PU�A�iq�&����$R�[����ջ@�p��~�9��=�	��t��x�.?\?�p{�R�\z�m+�U���c�k�۴i��bp���vaT�'nzEƐw��~fɇ]�|����R����\��0���.�V��k̶n�f���W@l�%l���\klެq0%�]�}������Ă1[+K-���
WE�i����)���=D�|�p��6��<��{b��P��Zt������ӕ�x�T_��p:�<���T�(��r[�+H���T��+,��c"��6�/JI��[���l5��c��S��/U��8E��F'���vJ[��XZ�5U�au
9�嵧���eMʻ���b16��,iW8\���nN��	p��`LlЃ�;���FW1!�l�O0
��l�z��Хv�8��#��S��s;����3�^g��ԄJbYx�����2&1U�V2�'�wnWr�#Ȣ&���V�����hS�J����A���Q��zZE��'�IX�BO ��j�&ve,�3Ki�
t����*}���k2�9�-�A[mT�<�ДN�ήv덩"�n��܆��X���/�$��OK�aq����E}_�D�Z�hqǅU�S�J�
  ��"M�l����c`�g��,">�˭�J{�j�`��W&��> �~F�1f�p��j�R먤�s�� L�n���9�"[+8@Nɰ�Z��J��4�]�Bq�
��ᨧ�����$�=� _�1HY�%�	���>�UC-Aa���-��z�I��)�x���`h`^[k7I�"z�q��R �.@���$��_R�ٞ�|�7��IxU{�S(������&s�k�˲m�}�d��NMU�1�0�Q�X4��a������v���tN
e�|��Ep*0A���j��:��;�lr�j�g�䛘/�^��]�*�}ϰ�n0)$IN�]`k_�Z\`gw\��EĤ4�U7f�$7��h9�/�� + t�MxU��t+���;6��!��Sz/#3�҃�e��.�,��� M������?�L��x�X ?�Gy�j:�G����8(�w+��\Z�x)�g����l�h9�X�T*q?��:8��6�m�"���d���/ί���/�ړ&U�d��y����jq6���K����	�T��.ˮ�Z�-��:�u�OH�h�U�e�o�O�:��'��	E�n�Y%ܑ+�7%��>z�X���{�-T��N鄆�&��j ;��E��'q~a��-"��Jy7I��,���$p�R���K2 �pa��A08 K�y����bta�-CY����o���dD��,��,������]�(���[r@k /�;�;�ұZ7	��W��.�_H	<ָ��2K�pʟ�ɚs�� ':���I���y�b?�jCk5�Hy�(�k�/�����
��I�W��O�E��I�E�D>c㯾�Ύ��
�%��ל�����?O��,�U�s�J��+ E�i����9d��zv�`�3g&��'5N+��r��[�v �������K%
j�T�&�+S3hϣC8�C��a�nwC�)�TC+�̆��S�"蚜Cs�~��������+�Ew��f8t��?���u�P�@�F�}	�۹���ޢ�#���ɂ���b��X,���i3я�l��g�)�?Úν�WX;x!�n�a'�,r[�����6ȸ�B��v``Rli��#~�傔�k]?�s��P����1�^�=�kC�M�6N��Oκ�s��T�-�K�Q�ǈ�!��(���K��i���7����dK��#�-��0���C�?����z�d�c����!���z�L���f0��<ݩ��\����b����j�]���>�X|���{Ӕ{�"�.&���Q��"R�k�>��;����Q
��Ѭ-�jC��}�R#�b�K�|�ˣFƙ>����L�C������c�Y��j����^(��Y�Z3Y����:�'?�xYCJ�g?�vBB&0��Ȣ��K�޾�q����z	�٬��uEBy>�{j���� ���<��I�.��Az߬)�Es? ��W��ayӊ����`����2_y���S��7��{j �ߴ���l�)?Ol#W�13��)\���lf���I�@P:��82-�L2���a���X���cR�������:�u�\/-�<�ۦ���cW�r*3y;m
�><gai�΁�T<�����X?V�`���_+����'>낾r���d2I$��Ӌ��D+��c��Ġ��:]�W����.|%0C;6�F3.m�ǝzd�o\�m��W'M�~�;��|�!f��H� .:� �g��	S�<�X	��,�� ���	�Z�̣��E��]�q���#'U��c������
Ui�	߷=��eE$��jp��E�ܹ(�x(�����c [w!
햹S��V�(���#њ�Fp#b%͚���]�K��2�)�f�?�>��(�`X���5��2�؃& �`P؇���R��}�K9�e(?����Ʀ �����hK%;DDOv����,Ρ �فU+��{?Σ!a�Eu��L��}L*��O���Ѧ���j�����#���3	�j>���z�ނD�09�.[,���"����W�.��=��a�vT?���a���'�{it���^z\Ӿ"N)m1���Կ\� ��Ncs���L;���V�@y� $��L�n|Bci�P(,��a2R�p`!�_�7Ŗ�v�m�Ө�q�5�xuS+�e&�Mޡ|�x��L�%~g(\��q�?:�4��m��|��R&9��]����y�w9��i��0��Ěs��gE��mut �uTؙ��uc�qG��6W��5���w�xs�w��Z��� }��vj�����u��(��D�o�M�o������o�L�ױ�L���N�?%I&�vj�n쨤�
�$p�-���O��$� �o}Q�� )���\��38�N�h� Ų�^<%s��d$�����&��sYK�]�L� 0���m2��Q��p����j�'�
�*��9��|���k�e�6r��,�����z���;\b�"ڱ�Q)���墉��ě���Ŧ	Ƞ�hv�x�O�!EΆ��K]�f��@#��<n2HUgad�� �?�;O1�3I�Vҍ���`9�b/�����G̭a93n�}�ٔ����d�����_�w��(�vG)�ꙶ�u]�z奴�]�$�o�|q��a����q�v����{���]<k俕>� �H��ػ��z��	uN�����ЁXH��"Sח��d]��sv���b�B̸��\��$�L��E���{�xmQ�X7?.��2��d�!صxR�{;���3&n�����d�p��k��v����c���s����q�7Z�?c��40 ����=�=��u�oQ�c���~�^�Ӑ����B����������㑗���0��m�ݦ-Np`6-Of��v��0\�3J m���l��$3�F���% p����術��e�/q�ɹB�+�X����m,���1d�Ͻ�<^��?�-�c�[M��61{f����i�����B�]�a�mɸ�^���4���_�K��7�afwo�^/$_vO4w���_�_�+����'$�lH��&ž]��k}���}]����w���������S�(�K �;�?�D����PK   F�X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   F�X'�Y��  �  /   images/df4f81ad-bfea-4377-beb9-28b9cf54631d.png�9��PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK   '��X��*�  �  /   images/e8e17911-f8b6-4995-a3a7-245093d5e388.png 0@Ͽ�PNG

   IHDR   �   �   ��o�   sRGB ���    IDATx^��^�q%x_�S�n�F$2� 0�IIT�Z�q��=k�3��^���ڲ5����-�}���ؖ�#��HV���@��ht�?���V}���%0(y�<8M4���{�Uݺu��_o^�9W�z�j�y�^�7�M{x�x� �4�7�Mx�+�x�:���!����'@8��-9�lvh��ڰ#[�L��(����#@��VhY�������C����V�Y�A�q\��c��FW�16��j��QTγ�o�Q9G��m[�e�vj�^�3�
����R�z���s���k�.��>�a��p��5oC������1�|h���d3�5'Gz�+Z��q��geiO�55И��o4]iV�4�r+s�,s�<��4��;�ae����+a�V�W*�k�jm�/UǢ4������x�ࢳ�S���M��:eYV��l ���_�S�_;_�Z�����vkzs�j������ߘ�r�d!�4�$��(�͇�L��3lۅeY���b��>,�I-Ǎ,ǋ��=�C柂�)�;v����78���S�����a|OD~�+]WG�{�Wo��c�'�/m�ry����@������m!AGpm�L����v��ZM��U\
��;��K�a#M!�i I��u}�j�T�4b�ׯw��?<o�����������Z7�k�{�0��b��?���/��?�����5Ƈ�M�Y�Yw���������c8y&���-8o#�@�7�� �4�c�m�����"���w�F��aؖ�v� �4������4if��ԚJ,��޾�K�}�o��CK�]�m��Q˲�-}}O����x��«�����`ޚ�d%�%v�8q���c�w2�����c��X�
�A�ix��(����9���3K�q����v=�y��H�Q
�y�R� ��V��f�[��w,��������_[�l�Ѳ���_��5��j�>�H�ʩ�S���N^<����mA<����n+iۈ�(��#�Q�V
d4�6O��p�xs��-k�d�7���BCr�B�H��wYJ�`S Is䎏(ː&lǃ��b�8E�h���]�����cޢ/�.�׽h���;���w����4���!�О��K�V]=w�h\�3���
�遚�+���@�!di,��w	V�"MB�Y׵�2��m�2��6�9�,՟�a0 X�].��r���d�A��p� ��!�#X^	Q�"�yN/(#�l4�an!�|4R-�4nW�/�]����~eђ�J��^Z����M��]g�|�g�䱥�z�������p]	a͊�2B���<�o��Ln� E�F�a[��ii?�`+�$7Vn�����)3rQ�=h,��/�1Aeŀ�DZa���s���#����Gi��v�Js4 rJH�rZ���0u�w�[�d���Z�~�a����W?~7�w�A�L:������<|��Ɠ��kn����V����iN�x$l��/N7oOv��TO��\}\�^f��<��Z�|@����1��h|1=�<?���,6C�>���ϑ�;X6Za��*ɟ0�Ў�ȲKײR�p�o��:�/}lպu����#�1��K��g�-;}x�{�Cg�QNZ7z�d�׭��4+�t�� فe�M��!`h�V

n(n�K�"Eð��|Df���|���I#�h�R���D�|��@nKf"F� ��3�UB��bi� v��د^��w-[���+6�]T^4d�w�>�w��;n����#W���r���O�{����u�i%H��UW��#@�"I)	"yh� lON.	f`��Ro�\c�1
1[�Ij\�d�Yhh��?��>�4���d�aFB"g(�q�KdhG�XVq�"N,�3Ӊ�'~y���{�{��_����6�8ӷ󇦾� ��;�繽�68r��͍k~(nL��F�����
n�c�Å�H�<�C�	��ˍ$(����0��w(>d�;e�"����M�]$	EÙsihTBn��!�M�+/�FaBw�II;�E�L��f6"�G�N#�j��Z���+V���m;^\uǏ�o�w� h�?�G�.}������o);��<�F)o�+����X	d��%���8Z��lϕ��8B��.^ݼf��h��[*n���8�� �T��0}�IU�4������wyFb�v�I����B��8F\��R~���&���B#��F��՞=K�o��u[w�~����4�o�A<������}0��n}hC9k��|^I:Yq�Y��G�0�zCsQ7R�Yoj�	��ğ\
� �G��!&ȁ̢q���!�)�ĜǺ��5�C�D�!a��)��Pw�!CB�)�J���Lf@��z����!�{H��a6�w�Y���^�y�׽o�������D��O9��������C���g���F5k���٨;�7��!*%�zE( H�X^x���ieqs�X�&H�
8$2=�@�����O9��,�"A%f	�£𻦯�yrGq����p`�
K� �waJ��(i,��ip�4�
b���f��Ě΃��KW����M�߱v�Yk�O~���6��gx�_<t�����?�#iszew���N�˚(��,B�d���2�� ��rA�Zx�a��T�H�M�Z�Tj�I ��!Ă%c�;)&��/�%�3}3�%�Hh��xw3���ňh\FVp�1hr�C2U(�(L`�Zq.`�
��HmL�rDZ��q�k��tͦ��v���j���D�����3Xu����ԯ���rm,[i`�u�����e���93�������� H�p�8�<��ӒM��g�@a#r�F»Gp8&iPɌAq_��p�s��&��pr16�	9�s�	=�\`kRWI�8�%|$LC�"�K򧑸�+�b��x�3=KVz��u�u���6| �V�o�A��G�����&/��Q�9����+]�����N۰,�3d�gz��3�g<Y$�|�d�v!�+-Y�T4ś�G��]��h<t���LȠ��g���`*-y��Vq#�e
����oLSV83���O���PXA5�4I���)ưA�-�}���vd��[F=u���8ݹh�_.X���w���q�[%���������ɣϿo������VR��,�� �YB
;K@���J�2���|>�^C�:3r8�x��Lxњ�z1�=2���d9�V`I�/us��Q���c�5�����Qy}M_i4}��Ij��:m��C�h9�'[�����h�@�8�� Sa�F��ξ#n��'�m���[���^�Vx�o�A����?}p׽c����d���n7��1������2���!�+5�`P>�|Sd�mjbg�q�z� "aC�fq�!^F��O��ErU7x����K���D�B���!������Z,c(bmC�
�#=�dƛ0l�#Iz�,$gmF�E�	Q�0qPO,�S�[�����jן���;����?y�6�o�A\x�S�ǟ}�����.m�t��� o"Hۨ�:<�K�@ǵ���I��L�an�t;z�Y�0Y����JP)ajb ���;����˿
L�Գ^�"�5[�K���䑚mں#2^j46-,�����@uB�1�����8��_�%��0M�21��ܲ���[���]ot�[b��/U��{әC��t{��[�lz��Q�#HQ�v!�P�<��%`2Ϣ9@Pek�s�A�:o��ԍb��(n�\j�|)��KQ��/7%�l��H�9�w�)D�e��"��s)n)�B2 z��S*�4�EN���,Q\A����&J�&yf#��T�h=Ahh�4���{�?�h͆?�x�]�z���nT/���'V�9��'��?���;G�j��f(!A`�`�؁7��@�d*u
Q����E��pr[m����=��	s���g�����9����^�qs��������@jXRcUy��ܔn '�P�U��5��Ȩ��2Ik�Dg��[B��#�;Ѐ��T�D3��t-�������Mw���7D�����#�\pr���^>y�?yc��7]��({	�*.�,A6����@"�)$�b	5�"��>6�0�½;J]��8���?�1��xcn���E
D��UP����*	.�8JR� ���x����A��&aءn#��x��H�%9	�9E�Dxf�6��[E;s1��h�C=����:��������_[���G�<����y��s���;�s���;|4j��BN;�8�,�m#�c�2uA�O�6B��Z�������3� ����I�d�������6���J�[��
��~Z��q�jJ4&%-�����9p�UrsM�ɎChjKc�v#C��p��\�MI�,I������y���F��y��Hu��?]�y��X��^~�F�D�?�������lr�mI}��I�*{Ȳ6���o6.y�Z��=5�\Jے>J�/��YC��C���$47�(�8��}h�:c�Q@�؂
*i��ڄ9�R8#�%��q_ho�X�=u4���-&ʟ��؀Nz~Mo����s�
�%�0IM���wzIK>rWȫ0��N-�S��=�=�������|z���~=F�ą��rѩ=���ԙ��k%����p�&*>?:�5��4�)�5�c�Ju��he#�
^hr�͍�����+����K5��1��1�k#������1��*��|���n�+���4Q
�:bE%� _�3H<�6K�H�D~L��K=EΌg�'����D��Nm43ͼ�����[��շ���[�G_O!�1��_�<��c�M\8�+���m�t�T�[��������ħ��d��4SD����&�0'�*��S`.N��(��B鹘%�^��䢫o7Y��uMA�6��?�q��V�������j-4wF�+�1CQ5`��g�#�Д��M���$�Y��PM3e���K��/�n���C5���4���\�G7l������9t�!q������_� ���]
��U��Y��h,u�Zy��@� (�����i�!EB�����n�)�kNo� G�3�����77��[�)i�a��Z�(��,���ץg+b�r�>lW�3��J���	�)���Ak#Ze��:f>��V�IJ��G"&1�(��"��#4~D%w�h��f^�ʪ���_��w�l{뮾��&���6����9���w�>��Cv�چ���vy1*yvކ�ѽk��B0��kbs�ט��U5��,F�2�=1춒ԍE-�y�f.���t�?/�����K��֗�Ss
aE]"U�ZN�u�ųoC\{�g4X���"�I*-�AK��Ρ�"XR�{���y��Bh�9�4AB�����+�-R��h�>�c�Ry኿�t�[�h�;�ݱ_���e�N>��'w=���K�r��}y=	��4��䚞�*� @S�Ԗ:�b��1"�7z�3L3�
e)��zS�V�"�������זmd��.�P�C+�����7���.��b)l����L��А�Kr㰲)�>����娨��{t��Z��ٰ���[�'Gdyh�ld~7�v��˽�����#7�q�ݯ���u{-O�{���|�Wky{]%kڕ�.�R8�N����:r����"&�ь���M)�5s�� ���p�t��#���� ����A��`f ��^�A�I��*�P���N2�"c1&Wp|}�~i�1� |ޤ�UN�J��C��`�TL�nA�R*�4���_\9fTv9R7�k�{#���HT�'��H�
"���4�x����Ǜn{�c���o�� g���B�x
^N><��¾��S�ʉw�q���M����ّ��q{
�G��Ffbs�0β�����( �*~Q����I
1>Kl6�_~�q�����a`�fBݸ����I� M�&��4 � |����^������� E)�;ג�1��,��bo/��i4�+�H�j�;���݆eg�Mva�i�6C�V���9�d\�a�6a䠕�H�&cm�+�+��ݰ������/u/��Uu��v�8�H��������=�pc������)��,�0@LPD�j�$=��wQ}T���bf��$�O�`���39�x1����!GN>�?��ބ}Z�֮.�Z��4�5%&	�2��;��� }1���1Rz�4�K�IGU�ôёv?�=L�	�-Ua�Z��wu2���%5�3Kb}/`��Њ,d^��C4쎉��k?���w�Ƣ;�Ua��l��_��>�K�K��E)�-��v� i�������!e�Y#��&��~��(f(e� c3����1�Z�2i爭��U�.\��x- �"���\UjӪh Ev!����R7��O6Qt��T��V*�l�,����z�/W�Z��b�q� �c��FU\KHL�P�AHWJ��5��Rג���c,j�I�3K<4B6WЂ����h���Y|�Ɲ|���?e�p���F��d��GJ��޶��/~,9���jٔ�W����V��\	�( J!�\0�b'��� $QĴ�!���������^�Έa�)AkKH�!���#�N6ԗF�%IM�b��k�7�h�,�t�
,m�p� �C��O�ȼ�s���N@��I
J�@7#U۴��C㊄dp(]&�+�L����1H�[C�']���x,F����ъ�Y���lc,����篹�o7����n~��o�A�\�����c���h��`���b����u䌆�RI������HKӅj8��g�g
��ϕI-�����98х��*���r��J*DE`���hq�#"�#@>@N��}�LEiEn!�B��z�"q$�K~�DZN �D�@rVY�]N� ��C�H�!�n�jåA04Iu�� �`��߷�M��6Q���t�C�5�A�n�M�)�UVڹ��*���L^ˬ΅����_\�q�sւ�5��(^��8�����g��������X��U�`Gv��C!M"��'�r�+ѕ�M���k�E!46��d�n�������e�l��)K	�x���Y#	�\�����L���QF;u��	�sJF���-�8}�
ᰙ8c�õSXi��^i-MO������yN�jb���%V�������t�PO7e�r=<yc��.�H(pUڋ��M��7o�)��cx�T��j�Ȉ[r ���e�����dZ�����w�������o�.uի6����������h�ܖ�rbW�6�<��)c�n����z��d�T&V2�� ��i&��Ff��8��
��D���j$��5h��6z:tWnY<+kI�4pʰ<�����k���B�����V���UBW�%'���>GN.E��8f��gb�.g@ذJ��'h4�sm�t������}��8~���V�J���e�hK�Ǆ1e��v}�����6ډ�d)���!���#��v���]����n�u���� �/~v�����s�v���/�ZS([��y<�f�v�y�/�tL�J�D-�4��As	�R�4�A�c��h&%�W��8yn�.N`�>��X����tc��ʫ�,4Y�'�Woz�8���s8s���i���dU���~7,�����h����J�a�m�
qxBi�~P,1���:]��p��y���ҩ�X��kW�c�+G�R�`�O�����x R�'�|�P+
*3�JyN#ϋu����p%$��m��Ch��BSy���{7�z�//�t��ւ��4l�j�y�O����~�o�=XJ&:J��t���;�S�]i��483��]�{��t6�Q4A����&�"L+�H0<�7�C'.�����C$�� �:��/Ă�Y4!Ɩ�.ZY�vZ��p�]{N��X�k��D��
���İp X��wn_���
'X4�T�>]w��B��#�s�:t��Mab�S`�|���q�̓��rRRqz	�.V�Ա������Mau9�0�����[
[�R>�Z��s� �qif�29���D���D�q�-w~t�]�}�����_\X�    IDATxU����O<u���������r2���$ܴ׊�y)|�����-_S�V�r�;�n�'H���h
���Y�[j�N��S��q��ƚ@��Vfx��Ÿs�b,�L��c�|�_C=���H��.��1Y�W���h�)�\���z��n`�B��[W`��z�6�l��#b�pJ��*r���΍�x��5�99�+W��T ,������o�@O%k嬩�$����	3�5 �v�NDoI"	,�J�V�wc�%[a����Q(��dX���A/��Zc����t�;>ܵ��'�P��>��yC��|ϡg��+������Qɚp�l+��)/BLJ���Ѽض�sMc��H�3|�Wm�"؈����DVU��#�q�X��0Bcȁ� ̈́�����v.ŝ��bQw��=.������C'��'^ę�2l=}5�\��׬A+l�����!Iu����N�u�R,�P��Qq8����؃Y��'c�x��|�<�^&&�^�Av;����티h~� G)�F�GD��#t��@R���C���&�fS�_�J��h�4�XrM�%�)�v�vN�L�׃�����[[w�?�p��=��|^������W�;��t�����qW)�DI0N}��0��"c��ͷ���&���jJʽ�l1��f[e�v�O^��C��< ����.O'��C,��ܹ
�oX�%�|�:�EhWpq���G�૏�d�����l޼+V.E��x�����i\�& �R��w��M�*�_j!�B���$g�]ӑ�3�aבx�D��@3��Z��>஛����U��^��gc�D4
���X��=:L�k�hBh9�&�B���r���>�@Sy)��lJE�KѶJhڝ�˨,\wtŶ�a��͏Zw~CE�u%r�ٻ�̾'>Z�r�>/��:8ᅌ��t�s�j���5=TX���CSL,`J������5��خ����p|'/^WV�b�^/N]Å���-,��u%v�����\'������!<���	��]��u�q�M�0�h�Nq��%<��i�?r
������Ÿ���XXj�m�Xe8~�Y'Ώ��k�Q<sh�@R��>�`��}�ݶwn[�]Mx��l�L�d]�(�Ef�Ny8��S)����L�d]�>�(����-�ߥ��.�y�Z��]��a*+a��ճ������;���ڊ��~��q�1����w�u��SI��l�bw�������RݤwH�ga���X�蔒�نQ4��pA4ozS���W�q~��ku������0��}�<
/iۗ`�yX�G�/B�����³�.bρ	���p���7�������K7��~�4�uD@f���<�}1�vİ�S����DX��S���s�q�|���k ��#�`�)� oٶ��<�%)�l�lAJNB�p�(!�/zʜB�*�%�I��� i���%�?C32�d-3a/Y]%'�b:�1�xhy݈*�}ko��M���C=��y�1��i�������]?��KK��$�Iq���O�OZ�!�L\��U���T`(l����J"k2��"�`d��z� �j�b,���h��v�s.I�1����A�~�|,�?�Fh{�;5�99���:���)�V.*c�-+�u� z�}� �|x�|���B��k��^�}�<���P�r���x����m<w��?>��,X�(w���5\�|	V����6�߱wnY��j��*���	ר�b�!R�]���9��eI=��fn��~�,��p�Rk��br �3�T@��A�t�]�:W����;����������!�<���WO=���S/|����[���[va�l��,���n�j�kBx��b)�#�d����
%���,s�_����.$� �L ��[x慓�}𚜴�2b9�ٴ�;C��8��E��������e��YR���������G�j��pO쾆Ǟ=�4p���U�eM'�-�a^G7gN��ƮC����S�2Ic���oA+�p��	�;u��4Ԁ�l_���.ü�6�E%���6ኾ�B�Db��r1zL���L�%�@�T[����X���=b�����$�����C��Bu��gn���{���X�+O��n�8���m�rd�o5.�x�[�\��b��J��}����28jr77AU����NP���BYд��(t�R���R�!�"rz1u���1<���k�� ]�mv�����%?D��1�xx|�0�9p'�I� ��p�-˱��.�+	��8w���v_Ó��H#C��-��b��. ��g�?���=��Lw��=܏%��`xr�<�SǏ��Z�W�q���x��k��;F���m]E���R0˃�x�v�V� k#�����'#� du��X���L+�6A�\�M�L�Xy�dʝ����D�_��������w���oDP]�A�'NgN}n���'?��o��.�Y��Q+��N!;T�Q%�!wYȧ��U("]��	!'��h.:JX�m��F�b����n<3�Gwþ��m]��w�Zܺ��hA��Sc��^�cϝ���:Wj�ܺe�n�CW7ۇl\I��cx~�yLL4�{m��a���X�|�����c���99;	�V��5K�c�N,Y�'Ϟ���<�cG���%=.n�i%�۾}�6:�I�����8aK��+B��h��!x��Cؤ��l��ŐA�[�������d��"Ҿ�K'�J�`��d��_zi��m��w��o�p��ĵ';N?���?��Ĺ��h]N��c�%2_(n�L?#���S�"��;�(�M�dS�~4pD�� t�����l�m�cI^<;�����ǯ�ey�,{x�m�cm/�v��&b7�t���}W��'�`��:Vvc�͋���t�hDFƁg����{O�Պŋm��a��5X�z	�O_}����i�q�-�l�TJe�<{�_܇�g/�5��]6��Y�[�.�@g����d�^�
�rGO���EqS��!X$�����&�KZ�i)y>�^+��Y#W�3�Pv���2��:��|�c�xu馿��������W�lw}qqW߱g?��ˇ���R���Z2�]�Ҥ̅g��FC(�YD6��V��Ґ}�r� ��3n�h`�=D{I� �;�r�0��c��i<������0w�Uv�;��u�X�݆���	���]/��+���ի:n�`�m]��7u��� JJ�����c���3*.�y��ܲ�,�G#���!=5������~�\��ZI�xã#8?z�u��+ V-��ʅ]X2���k���M�ê�ÉdF7��9o��T�V�؅2fH�C��)��W��3�� X����7J�]�0��o�����H+�v����|��ZiͻN�>q���܏��3�x��M HR��܊d.��c�QA��P"�ӑE��A��S�Ӕɓ��a�Ի�@X��kh;�0��a���{�O\B��e�wl���a��U�qDv$�̋Ǜx�s8uh���y%�u6n�A�� �LL9x���x�٣�kje`�M=غm�z|\�㑧����c���=�Ƕ1٨c2����?��Y�*�x�ޕX��F�P��(Q
�a��*"��Y'��ލ�̸d�P�������5/*���%�MO�yVBE#C�C\�k�K���?�˥�xEY�uy�����Ȟ/����~��v��q�Ӧp�Y�)
$����B$g�f��#</D�"M3���p�*�|Ko����H����W�t0�����&�{�!N���{�ⶍ���+���ma;O^J�������m�`A���V`���!l�8n�>{�e�U�k��yǍ������x�8q���1�Ц��<�^B�ݳ��I�R>:)l�Y� �W�^�m�;��ê_EOI�"�8�:�����AP�GwO-e��&K'�RxW��2-צ%�.��BD�(��$���f�Ȱ�8��e_�������8��<�����s_�ϭ������!C��YH�*X�A	&l��"e$��a;%���P�}��l���͓�C4�3*kK�EI?,z�#i/��k�ѽg��	�!]4��W㶛����cH��S���2v��׾v	a��V�8[v.ƊUњN�o�i��s�OK�i����5ؾe9�tW��a���6�b|�3�	I�5L�cL$Te��΁� @O�Bg�ƃw�Ħ�;BT�q�YqëtH݁��*�Í�(BF��R)��C�}Ba�hȫL��b�N����P�.�f+V5��{}+_���}��=����S�����|8�r�}��H�c"����AU�h�³�hE��i�ЫƢM*����F��L�d
,9�v���K|ᢝ�Ѷ�1����sm<��,^<>)սN��Y���*��Q�^�����ƁCc���N Im4�}Jؼ}6ܴ�Sm<�����	��
�^VŽ����EU��i���	d��٦Z�F�e~u����XG/\����7:��ݰ�V.���nX`��+��&�a5dZ��+,yhI�?�JΠ��� ,����Z�QF-�%�饙�%]q� �a��gX��1�Y���I�yk�]��m�0�-�,������u���_��ڱ���v|���kɄ�T:zc۶+)&��b�Έ'���yJ�Z��\��PD3��kF�ee5��<�)G�p�ߑ�m���;��x��n�=q�Ę|����jܼ���IԌ�Vs�j����<��,������=����֠�Hq��9L\��3���Bl�i�ne�����4{^�3^�������x�8x��V
����e�:ܱc-�D([#����c�Yդ<$9�v�T��Ljs���M�|%/��cvt0G!0eaP5f�Q�#O,��1�BVe!��{n��K��B%v��y��2����#G��^x��[jɄC^�z��J��,�t�;-l�+#|OQt"	��A��r(A�A0�$�p�
�&�!Êỹ�7�!"{Ɠ>��S{/��1�J��o��M�r��je�z¤�OM`8}���:�3@g����S�9ʞ
[�-/c��X��^6-"Yd�hD9��O�L�
ZY	�΍�=�p�t$���aÍ+p��U���F)E,p5d��qGFg���\GzO!�L_'���5�i�a�R��#�{8.z	�C+|P����B���ğt-�7x����l�M��������~{���ؾ|��l�.�S(����חA �"&e�i%"xa*4Ӽ*-j�y��x}u��vi���aܘaX9�KZZ�q�UFd�`<���3M<��E;J��7o���7���[��Q+!
9��'X��� GO_����S�V���b�38`c��A���K��U&]<�,�2B[�E]F�T�Ъ�ę����9�>��Lg�~�rl۲
ݵ�|LTS^ޒ�N=`�L�͙�C�f���.ZEW(�v�itU#��2Q�r�bb8��@�bm�Qm���<��+�������>�y���O�W��ޙMZe���#�"���ɤ��Be+�0#��KGG&��LAn^.��b�k�@S��@,�}6wo�̮-1����Љ؝�����q�{�������X���0�hߒ�h�׃�����2F�\��d3ߘj��ZEO�����pPr)�'�l"O�E��#�4ajxk�R�n��#�X����&1j5��;P�i��Ti�jA��Q��Tj<�m�t�d�[1S��Fdet� Dz��SZi�*ڭSm-� ��[u�C��r������������[F�����Փ;��)��:J.Og"�8�8���)
�(-��~�q��g4�	�R5�r�Z�Јm(����p���Xb�v���6D�F3����\�b|�2z;st���\_�!ŭ�b��ׅ0+��8A��F9(��RFɥ&�ms>�)�+�Sa��Ż��4�$������B���n #�[,tvx��	�h�w`j���H�T�,K:�8'�M�f*�6���p���R�����>QzQ��afeQG����љ��%{���_Z�yۓ�C����2zl�d�N��̧l{�\���iWTP^�M�:���26��Y�dl8;A$�&2'� bNM�)��9�U
=��Ӵ��"�F��GB��JPF�1��O�}� M���)�y�Yc��Ȝ����S�Tg6��ʥ@&�K�}�>e��#қ�;\����,�:�������+(B��=�&���)ǥ�LHh>��	3	�j��[,lQe������ *&�B�mi4��� ��&"1�M��� �+E���6��_|`�W�x^��x�~��C�>���wtc�u�1���Ԧ��1Ċ���{`�t�&v���7�=���tQX0+a	PZ4D2�;��B�7lZ�-_�Q2u�^F��gx��P<7�ĭl?w=8���H�D�r���F;JP-��X��N���)�a\-�6�X~&��<����.Zt�<�TR�~Q�U%�&��\H'���Q嬈�!f2�d�L�+�ThvX49�F�*��u��n	df�A�%���G�;���?�����ʼ{���������p����u&/�וO�N8"�,l���%��{3SY� �yE�LȠ�تƋ,��9!��S^٩d�������y
��`�Ú��82%���@$da�	�����z^��4�F���!5���}���v�)��|.6Ӓ�q�5}��Wcy�b��ݠe�q�{88R��%����L�^F��Q��<2�L���t2��"d�+5?׹zu����~� �o 8U�J��r���S��Th^F��5K�|v�[����m?z�u��/���#{?_=�P9+W-�O�p�J�=�f�T�h�R� g�!R9�Pc���g�P��/�dl�I�j9��,U�L���ǙK�6G��yt2n��� Vr��?��wPb��4 ��&a$7��<�cqaȕ�x�����l�2E����DgL���k��^��%d讹,eK琉�뱌=��FC�Q��ʇb́���2r�k��%3�j��G\��he>��2"����ƿ�v�C����_�}]q��[>rd���N}_9�V��M؜#�i&�P�TKI��8[A�/:X�I�#���!PEM���u��΂��B��:k�X~&�^xperK���n)�,�g��T�#R�a"s�e�f�s+���{�����[f���Y�$CF�LL�����|ι�{g:ot�3���� Э���B.1;3�_D���G������(,DQqG�>��p�\�Hꠝ�n����0��\r�'����߫���W�Rw]��s��⾧~�u���k]U0k��iV��c�ub<����-V���9�m�(G'���2��V�_�O�p/����Bx1����Hd��{V��Ƴ�US32(�ZH���"�"���eׇ�riQ�RC�:ҸkfM骅b�,?$�%l���|)[�K%#u2o��G�4�r� F� S�2Τ�j E_W����kS��i�q�U3�L��������*�J���m������E�-���<��O-���?8u��/x͡ye48� �� L$,9]��dc�'�I���x&�b��&T\� Q �}i	iVB��*��5F�8�-8���h1���% /��@f����,��V�E�P���e��7CxN�j!c����&A���U�H����X�Ib�2gSddқ�l��D�ّNo�{ʥ͑d3 ��o��ʌF�!~v�tm(Ab��5�r�l�)B�N��}\O.�"���iqe���+o�/k���Ş-���\��?��+��z���{˭_YR��ܶ{:��}.L���.����&\~�5�b�2-��A�������:i�� GU�t�m���L�8(������깋���J}��N��d��֛�io�Md�>3Q'���i�!�'��VșO���oB`���jZ��Q&��A@K��4�r4YPn ps���ңa��A2N"%�!��T�*o�� a@���d��/�r��9���er��s    IDAT� v�u!�b�3f�S�TV�d^A޵d���~�;�?c�����2����*���u��#���=yym�OSIc��d���2l�sP����,N7.�T:C�T4���ٲ�D�t�6�c�hy�Ճ��Z8wq��C�
8�3��a��1C���k��m��K�Ba&�ҥ�z �Y4ЇJ��f����	��(&щ�4�ٌ ��e��Y	��� efD���J�z@G��xa7z�(̡��3����;IeТ��)��mAH��2����4)����*^�S2���T��A������z�W���^)\��}��W���������&.ne�/±#x�A"ē'�R?�x�K�T8~X�A��x�{�\�n�����wXӯ"�{p�\GN��ęHF����wby<;G��HW��*���]X�0Slxs�/�E�����:�\� ���ZHmV1��f��8��'b891�cE�������U0�����If(�\m$v]�1��x#Ep��/��Id�5�&�MR�j��PP�z2�.�0aU��k?�ᶇ>�`Ǐ�y��'��oo<������q�q�L%��7��1d��ά%A��"J'���v�B8u�_��q�� u~�I%IKH�.\����I\��7蔸�.B��n�i	6�]��Q�g��Q�̀\���DL� �q�������N4-]�J>��%.��P#5\��!�R�=u�.r-&���ep��R����tQ�;maQe��^��j��p������Lw��A�cE�]��4�P�A��hEJ�q�_�`4���ALZ#��b��o��چ|Ñ ��!x��>�G+���ѩ�*[SU�j³CM;9·�
vQ��Y���V��n��rYP&r3��g!�f<%g���(A��̪ar�B�e��C�jd񈹿�y�HuK�3&d���S��d��d�H\;����IZ�nX$S6� ̬l��f�J1$��E2I� ���K�ԙ"�`$~�j�8��%1��`r�LSB1�N3
A�Sf���ers���8K����z�/C��0E��܇�<�D��-���ַ��L��n�y�/���s#g������yN]\��x,D%`��F�s�(�a{�[�/d5�y;�%=D�`���.QR}�k˗,#I|D�/���I�J�:�=KUf����QQL��M��WB���\x��F���rt���s	1E-��qݦ��(:	�dH3_�Y�f�蘢!�3<Yf��!i����4dS����ҁi�~���h(mɖI�����[D1q�e��p:0�u��[���;q�ʍ�Y��/���u�Ԟ����~��W���Ŭ~iy�m��IC��� ��]k��M���c�aZ�(�q�$��vp񔐿W]6���p�����,�YϬ��C����g�>�����y�jvY˔��1�5��M���u�6;S��������B���µ(����nd��\"��t�쨮uTa��-��U.S��f1�N���V��ln�U4\�ka������;}ٝ?����B�� �=���q����9uKͣ��z^�CS���ɠoV1����BX@J�=1��EF'��2x����IS,�A��Jp�HΊ�$UA^PRŮ��1�Ɣ���bi��3xn]�ԡ���fhz7�q���EH(�s�j�ْU16Y��K���i:[K���܂뗌�V=�(L�0�ٽb�����&�$�'�8�p�<@�����92�~ǟ,�r��m���ؠ��"�U{���M��=���Z�#�#��#�t�2�;A�:��Ι$?A�]}���4�b���ڪ���$��y�S�O_����3�N
8Ji��a��h�=KL��p
2|Ԗ�~2L�}������Dg�K]�N�}�bI�)�ڨ��gp�Q8����l�5�)7�7�MG4э�}`��,n)��:ǃ�I�~�˕���bP��c�c	����G�o��?�ڲ�akٻ������|����́'~���?V���n�RB�`��9P��vN���=��t����x�(�
zS9>��,	�3$M�x"A��c\2����.��A~ͬm,��0}C�P�W,p�z&��Oa �P=n��xv��f6�[2�jh1<�����,D������m|�<�K���,��=�'�Bx����3�� ���m�Y%�a�c˷����Z����ֳ��:y��7��'�Ϟ:x��}��ѵ�,��lw� �#�X֒�B<I>|�Q��Bق��T��Dt$��� $iD�)/=�,&@�hs֒���gf��|����2�P��J�豊��/ۙA�@����<��C�ZzW�icV<�{Y��v�Z�O%;�ϥ��r�0�t�!fB��l�Rf��k���V�nU1mUF�n���r��ٽ���:d�E��'ޕѫ7~��ߏ'���eǨ�uT����S;�S�RV*!��M���:D������1�-P��lӂ�C�������f ���v�nTA_��w��vS��ͪ)	������J�g��:I�>k̪tr��t�MW��E�JV;�M:rM*)�i��C-�G���pZT��b�b���%d8WE��c����M����[����6n�J����	^��_U���\}��V�����Dc�^k�ԝ��'T=�.,�`��(�%��n!��1�ݓ�`�3hZ��+-��!<}���8EŊe^\YT�_r�f��ߋ�aq,0{��M4Xc��,f+<�̚g�afz(�gR�0Kߌ�B��YC0�Y����pS��b�e����45C�Q�;��?d>'�5�򼇷���_��|�ڶMY�o���b��O.8���?}��O��J4� �F- ���]�MZHS7#	�TrҌv/�J���j"s9���,n��L�:�s�Es@������U���e&��)�Q�J&���9Feb��j'c E�i�����0_"�������f�tr�;H�E���!i�]oI��if���Ŧ>Q_��Nȳ<�!�����Beњ?�r���r��k
rR}�v�ԁ{Ox���hꦠ5� �B-`Aƴ��,n��Tʼf�T4�"]�&�Pq������ll��X�dp��D�p���{:���̅�Yښ�D�,b/V��1s�_�w� ��C�6�C:�`���0Y���j�7l7��CF����]\b!�ۙ�T�,��*Ԯ/��:G@[UL$���|f��{?�l��v�����9�W�!�$cO������-5���c� ����d�U�X��:��w���:3��x�d������g�"Eٷ [��[Q�\2���YF�Zl�3����r�+�1����aD���o����}���*8���:}���Ѓ��H���K=�1f��F�r��rC>�Y2}�/����B��v�nw^�.\�7�?��?�Fr�7� ���j�S_��Oa��td��x��sK��SbO��=�s��R�A����2r�A���EU!��r�ȕ��b�܋]����?g���9E��^�a^�~�̙Pf�1	�)�Ϲ�j�F_�$}���� 
�P�a4l�f��������!c�`�u'C��a��2e�{�l�ȭ�z�Qk�}�^��k����v�y�+�M�;�A�� Gͳe���T%��³�C��E'RT��]l�T�kĭ��U@�hܘ&*ސ�+2z�3[�J/���:F�S�&cg�g�|���!�����C�J>�����f���,��(������B�f�kc��p�JgEA�ˍ6LRaV[x��p��-��?^�vw�&������Yw��]��>�?�vz�C������-T���E3q���<E�0�nv��5E���r�!��!)<��/U��Yy�ٮ�b�^p�|17��e#sYʹႵ>^V|74�}��V��x��i�4�b��o�j��Z���pyY�v�(��[���F���m�,�=o�-���w<e�|`�]C��_�/������ϼ����z�g�x|i���˚����o�дKw`ɉ�2��R'	�A��[\<�i���d�L�g.<I��PCW����,������bm�Y
_�`��dm@i��U,<�l����x�b���<�kŞιa��l��@�)��,��g��(�Th�@�N��#�Gh�q��#��?������o��u���o(�y����=D~�S��c�o������[;�X��J5��4�uL���rL<B��Nr��a KI!=3�j-����#i���r���Q��1���aF�m4ik��������Y�𥆹��Y`�^���F�e��[7E�:� g8QPb[�Xt�n�ER��8�Z!��\�Ȧ8!f���;߱�Zr{���l6���W�������?c����v�f�#dJ�f2o���*4�%��ǳ�Y�-�[�0#�I��^���EV1�p5�7�9f2��d|_�����ܐRTT�=K���1^�v�ㄾ6�Z����u1^�"�9e�1�N$w�LS��j>�������Wl��K����w�͌�u���9r�;���ͼ>����lZ��TR{�r���l��\��WZ��3��_���)3i![q��]\�|�ҙ�r��Ls�$�dv*1|�,��!����Q�%��@Ҙ�i��]��f-����n(RbL6[7)�A��sn�ISU��Z�X5)��$D�.��C���?�w,��-��ު��=x����3��e\���v�#�?�_x[�A�S�dÊ��EJ�Y����� dP����)4f�3EP��M�C�a��OXM�
�=��,.�Q̀�5[v����d���D��/KG�D�g��x����T��.�W�;�X��^N:A��\��ڏ�6���=�%D^5�LK/�.��;�o�#�;��u�,�pQ<�/����CO�T�ک���}e{J��H�\6�����fQ:��Ő�R6���g��X-7��~-���F�O��rZ�xsb.&���(9���[k����6�uF���2Ђ��`��w^�w��<?''�8�M[b��&�ı�c'����@��@X�@Hh-���^�K�U����fFD���f&A=�p�F�]U�~�����yP�3?�P���>��C[\�^o>~�u<���¾o��¥}�/浬\t�[����a̤` Iq(`��3����w_[����=2��K�~�r���n���r��0��O���%�5�,�bH��R%�D�m1����6�v}®L� ���b\������0ppxh/��@�o�3�����g���ۃj#�G�.��7a1­���6S����g��nX�82�������i��$�u7����<�\���¿<+�`�,�{��ۺii�����ji6̨rA�ac�cxx�i���aa�s�:"��0(��Aa��M�K��I.`YHL:�����|��G�Pe������`o�`0�Ơ�O��I���J�u��i;+���3��#��M`��7��u�g&��0X�W�u��x+6u��.]�.1����M=k@����я6_Q��d�[+_�%��M��j0��V��@�����Ig�|�@���M8�����e|\xp�m!����i q�r�;��f+'�N�"��3s:�|8��tb
�l����|�Y�<�������3PX��D��$�ԯ�$2�����o܋��_zx�7�̎��B����O�Gv��j1t���O�5<��N�H�o<�va�w���D��x<�0fN�&�k�j!��9�o��� �X�Q>U��b^8�e.	�`�(ZVfp׵�x��[�F�)l=���Aa���)u���b!c`�q�
_�zh&8�{d�e ��ڂ��`������W��2��ĜK6����3�W�������&�|�O��>��r��p"p��$��n)��g`C��w�j����5�4l�l@�G����q��S,'\�'՘�ϊ�&��\���U�9��-�>V��g&�ͼ��\1�p��ό�J��gSQd  �	:�V][UM�c�qG<r!A�QNd3�o�ӭ�=1���Ɵ�ge!2>�9��拄������RUs��;���I�� ��V��	h�1-�0����L82��0����[YMl�!�~;6�?0���n[������S(svdc+�.��l�(��[ +��&���7X ��� n��x�x|�0\̂N,,`! UA�Au	
Zt^p�^LϽ������}c��WO����o��oz�Z���N��mN��	(��ae��N�XN�)Uh��1�"��Q+�ĝזӇq����y�7�vNM!P`�f��U½�����`��Ίږ߿�~*�����&���Bީa�����1H���Rk�M��y���ؼKx�:�:�T݉j"�J"é��ד3.Y3����QHl8@i�B���]�О�s��oc��� -9`�����5�1�Tja� mm+�C���d-ڰ<�ɪ��7�n�3k
���ÁT����ȧs����9����@(��:>�TB\�|<�'�N%�؜Q�mش*�9 ����vO
dX-@�c�]�T�dj����h�k.�m�Ͻ�¹�z�l2���5��S�}o�wAϑ=�e���N�
02��*r�*r00z	�Ɋ6�^����X�ѡ���0�N�ί@`*��_�qc�5V���dsN^�AT����Z�B�PXTܴZ�@�UˁG��G�G�YĲk6��$JY��,��2��f���(�x���	��lV���r�!�Cɲ��/!2��⭺/�Ǜ�����}���:~8��t�mǷ>6��۾-O����y�:����bI�p"�)	]�0�����c@d�7H��\�u�csj�Κ	�G+�	6��Ǻ��Z?���48��o���M6���#����`���x�һ�-�%���s?�,�@Nc �e5Y�p0@,QS+�T`��J�4_Ye�(SXU��9��D����'/��ƿ�\���Q��g����X�s`�J)��
�ad��[��[���o`�xH�^ C���m��4��i�X)Z�`HpF�����&��ج�r.��l�SL1��g<X뛏���Xӗ�j ��A�	�#س�
Ivj0��S�PÒY=v��$�XN�%6`)l�Xm��f��
Ua��4eq��≀��C�=������QVTw��W\�����V�
X�e!�����h���o�uW�j�fw�H��*A�h�i�Nϐ$8�1iͤ��#�[�D�@��Y= �&�@�%"MV���M�0���h�l�N�Xդҙ*0�Si���#[���X#,J<V�5T�q
f�n�A�Լ��X��=��h{���k����ҳ���	`��S90�dA�wp���a} A#Ҕ�����HXĕ�`�s����N���G�;.��sum(���qٵ�?)������� %����(U�][  j����-{C�!`@���6̣�E�)x��цQ0���q����M�Yg=H�q�3/ *sx���Ԇ�	{؈�a5��WO���8�`E�ʝ%َ���k
��[ ӈ��A�#�i�F���Evx�I��:��,�L��<7%��EC.7�d����v�R��ҧӈ�ܸ�]�����)H�$���4*I���'Sg?1i������s!�u��&��ܷ��r�G�Ҹ9�J�|N�f)W��h�s���:>d(i��LJܘE�6C&����4��)� 	�0� f\0�]�Xx(���ր�n���_|�@���M�H�����c�
7q����T3.����%�l;�6��¾Z��V��_~��y�0��[ �p  M!Mc�:L�,�T���[8eGQ.D�N�)�� �N)���`�OInA5���IN|55{��	�/�}&������ atnv����z��\<�4�T��ZA� �XX���BJZ��
]� Q���Y�9�����h�0J@�*�#���d<.OUUF�
a]C�Z�X�1�
V�a�(�ZU�"�<h�ER!+jKl;0*    IDAT�H7[���Z���Y@�x����2��M�d^+�~�]���j�{�|�����4(����l��A_��@rI �ff1��h�d�A,���L�G��A�,�H�DDj*�I$*ɠ2�E��e�cκ֙�7�.�l��Ɛ ѹ�W:?��?�}��֊m!���z\f�4��͖6�_@D:(���w�� $�ª/S�N�
��-�H'�x���3�"RUq�*�.@Je��a��9L颟�L���&5���I�B�9T:M@�]ᦾ�]#�!/8�X�xPw���)K`:��l�b�K~X�S�X� �'����ft}���4���C%�.�,LPa�O�,�
��e<`Ņ�(�v��DX[��4�� G I��PyI"Q�N�
�AU��3�q�Zg/zdj���I|. �C��۶>wQ����̗Z�`Dr��U$�9� �i�+�*V{3�R�p\�*��W�Ly>vDZ�5�6u�?Ԗw�dt�}����������J��"�xȋ��ƨR�a�-��{(p&���9���� ✆�nπ�2�0�V��H�������f[vh@I��������t�������Sb�n���Q�ОO9=����np��1~_�h�I���F5n"-WZ�t�x�=� �3A��f��`����I�
bd�aV�E�3�'�1��o�,�Ⳳ�7�����W�\.����R����&� �a���N,��"M�ѲjҨ.��֚�v�l�Wpܯ"3vN�qM1�-�Sw��?s���>�t���)H�.�Ui��0Ƴ����K�
E@u[S@���Gfq �c���OV���*�_�����5��"��cyEܽ$WpM �M�%E��E^PN���!�?��
~��rn_D����U���љz��e��-���V�.2�1��tJG2c ���#�AԐ��8g���H ��j8A���D'??~�e�/�e�g�oCQ��w���ߘr��5���(���w�@��D�Hu��
�*EA�$#]��� `���@�T����L�Epܴݓn�F��g�S�y�J�/�ŘQ�N��ꅆ$��Zm�sI
	-M���!?��z? rP`J�5
��Z?��o��X~��Rh�������qX��T�W)��5��$dвn���زA�}�pui�s����G��	�/���W}�no��y3}D~3����Jw���b�u��Ms#��R �,#�P�4�yA5�`]Vq��58�a�S�p���@�+�A����8{���k�9�����#�k��k���oI���f�|[:L#`DQ*��n���=�]-W*��`Q�X�� �"� *�9��nw'��}z��RK������R㩧��託�tyĒ�'�R�Q�,���������-�,zIBs:i�5t��$���� �$ȠQkh�9S��n����Py�q����U�RÀA2h�*dYAd^3��=�˿��E:]�P/�n�x��ĥ�:�L��ǥ��@���'�K}��ة��=��Y]`�!cqS�߅�"��i<*��UI�UH*k��/5����?�q�ww��@���Y���G~���Q���CDA�C��֑�� )5���^�ÿ��8�U+k�]�	n�M_�u�ҿ�L���|�u���}nT�ܪ�U�W%a�*W[	M9h#�(��r��5/E�N8�$Y�	���H�vy �d���#+/��Q�J�Uj^TuT�	"g0l�q��O��<�Ё����I�`���;C����^~,Y��5_����Q�]��k�.JB.�:2r8�O4CK��Su�Z�,�t*�nUqǶ&��_{Ɋ��n��Q��T`ߞ�N�۾�-D�phe�Ԋ(쥐�����F8�8�Z�&�I3�.��\��L�9?���Y��z����� �PsՄ<+c�u���M��*�HC���U�	�ǐ)�]�=_��BѰ"$�J�H���J1L�tl�d)���.**�g�	m���P�����ֿ~8��}�">{�S����Ē�J&(�N��`I �� �񠲄PYfPQu���:�t�|�W��Oޙ��KxF@~�m�w���Z�П%�(��*i<���&���шf\H��q�	���D�:j�֜��:^�H�rq/A�7�D�N����>u�z�����(QA�d�$IE%$ �:K�*��ҩ�ɐI�� 5]&=:㧵q����"�Xz��0v7�9oͼ򤧻w�4���?���k}��r�bH1�PW7�)��	�!������Q�:�i�ċ���ÿ́���p�����C3�����Υ��A��|�����e�
��<�N�UM�([�`���p�;���x�-��vce87�|-B{7���v��t1{�H���U�I-#�S��>�ŃkKc��j
�*���J�C����X��ˮ�>���ia��ؽ����{���S��)!�&4
y`.��3��SW`��#�U��5Qn/:�ǩ�ٓ���i�=Gt�y�Os�?{������]p������^R�]��� �E]_��6��ОA}uU47���O�g�pފ��rh� �Dn�����,:��{��7ˋ�(�#�$�A͝"�(�fQlI
����֋
��Hu<�~��.����M?������ܞ�/��B��i��gtD�u�bA�O�!�J�H@*I�5'*+���W/X���S�<��8��?O������>$+�c>��,$���㠑��@�z��L:�Ha��My*�+��m����/��y��g�T�ϻO��6u��7Wz���G妴 I�#7k ��avu)08�����@���4w�%������١��i���?�?y��W��uU���(�V�7���aR0>E�� dO�@;¨Fz$��<1a�e�|ޠ���`�u�"��ܷ	]p|�{��W��ץ����v���������A��wћ��n�G�ġG��ɽO���֕'���&E<*
�d�\��p�=EՁ���TK�l{�m�%kƏo�{.�ʚ`X�������K�����D1��栱�FMёLzQIs���)�Zg=<���qs�P��(���h��+�}���>��r
���(9`�6�(AEպ�̓$¯�Ϟ��i�h��|s�n��z���!���ӎ�z�^�ﺶ���� ��f��e		ȁ����b��YϾ���θ�� q��6ױ-�����duN��������� xYTPE@��z�ʄ2�+���E�>к�7RTin�� $��~�z�wG�f8�*r�:��`h���7@�P0�?g�˿�/�a$�Nv��׫|���G�T}���/UE.RB�lm�zEUa��P!ݭ��殙���7�����}ŉW~:k���i��~��t�au���jHD4>2JF����W|�y_��g�T�r�|nÌ��_Z�VK�}D��ej#,�s����
I�3�����K׍_~���w�F��+�����"��K�^N��(�Z! cl�2��d�p�c�=�/��wéz�1S���_����+�B��}d5�w���U� T�iMr�w��}�c��͡��>l]��Y�/�U�;�#�7/;��և�Z���C.TAn�$�� 3�D�v�g\v���n��9t5�3�s׳-�y��̡]?��B{�-�/����V�:�D:�J�|!1a޺�_�o�g��s?	�����n|@.���(z֤��8�\�Tx&�59s���p�tg.OQ�6��������°Gw����Hj�Z�5�����^�ؼ��=G|ƀ�����_��n[h���g���ܣ�Z]Fyh�>���� ��w�s�|���e��n�gd�����{w��R���a�%E���N)�����������v#�}����������069�������=�����<��M��ԚN����Q<�~>��?���ֹ)�m�v=۲w�{˸��5N�>�!D\PzY�:щO&�]��Ԣ�u����	�Y��6/w�����.�NA	�4�FE��G:�_���l<�j�@":��?�:v��t1����HZ��n�R�vN�|����v��c�Y��k�O<;��������^�R�$��������?Z���o#@�?�Kïz+�o�����oU�Zr~�W�d��)�/�7}ɟ����/=G+`d^�:����ν�#�q�f���%��el���v,�Α�^�sa�Ώ��r]9����T�Ck�8y�d��c�B3�`ĩq�}����FqG�����?�V�[!�	A1GS�0�K/�Ћ ��G/,��� M��-YV�����ُ��9v>l�h=�������_���Ε&2�)	�AnO�'~���ŀ��olH�8~���U��� �Y0��\��i���������|�9\��ǝ��[V��դZ��H��}�~�h]�:}yC�tC�ӳcI�Ư�Hb:<� H���O4�^��VXs���( D�л�.�!u
�����\�����=�i�	'{?\V��#b:4�
�P!)��d4�@���׻y ѣ�Wԫ�u�u� ��y����-����au�ٷ4@�]�}W֪�����"�b��ا��تp���9x��Gs#���.\W� j�B��N���	x�H�ѝ9��Z-�7c2tBK�$��B<�\o߬ps3��ˍl�ۣ�o�V���$1IS4h9,�������=�	C&����Xgwߡ�<�?�}2�@*�*R�x,q[,�6���s� ��gF���S�r�+�O��D]ё�j%���L(�77b>������r �Me5YRe�v��J&n�DR�*��3���D1{#Ǘ�P=T�dI�\.߿G"�U�H[C�C����W����pd�F�,�
C�o�R�[���9�X�5�/}I �$�n*�˫i�uYVx���l<�'n�j����CW���`@�4;�6q�c}����= �����̕�0ۦi:�v���>��F]��K�~����pdH��2�cK:��5J�9�7g,��`����M|�[��4���Z��	<GV����ZV�Tp��!I*M�[c�[����c� ��5��?ٝ�*W�V��j�
��M4�w$���;���Ñ�OAIRT�v��N�omiI�n$g~�o��>?X�ZO�f�RZM�F:�+�Z��	<E���准�C�{z,��G	d`@Ȳ��$�-�N�	`@��~���|?BE���d�
� )���ժ��}:L�`Dq����J��(��$P~�eY�H�x,yk$�����C��Wy�����4���\���y%��R��b!�'{^S�+�"dLĀ�T�$�w��ĭ�p 10.g��漼⩀����8�����F�?Q@����\�#	bL{�$�D�p���& F� ��L��raCip*�2_�x|O�b����x�C� _�>NBE�"�m�D�p8�h���	����3�W�r~Mѭ@\*����x&��Q@��9|U�Zy���T
��$���D���1�H�.g�rS�+ޏ��K<W����g���82�$ D�^WI��}<��-i:�æj��2~q�
��d*7q\�~��V`L�<_w�<�Ģ-��B�GΩ���J�q� �� @$�V<��~:�>'��8[5:O����ĕ
4C�J�2�� �|A�`�D�ɿi��63����S�bZ���WZ���@��p���$b����̡e|����(�2��7���D[��� ����t"Z5�GFW��z�[o ���Z<Y�H��x�㼿$X����r\�G�����v�&I��L%���������B'#�}5
����`�D�/��0�VP�q\��q?���~�(�uHy��ܱ��*��
N�$II0�FB�;���M>�` ��W��
oY�4���׉hzD��lo��R�R\oh�i!d�$��#�Н�Ȅa�k���}!/���~��~d@��ШV���.ϯ��������o0tB�e�$/E��RMN� H�ݙ��W\m ��D����:��;��J�'۹��O�>R׊,�ɼ��'�F[j�U�]�2z{k_)r����X������XK���ݓ�\Z�]�BQ����MD#�4i�c�2�0\==�n,����x0�ÑdL�=٣K�\����i��x$
�h*ޏ&�pvg:o���k�>��,�����D(>�>��wt1ϗ�ȘG�,�u�v�6�����(���a��]�PxX'��'P�*5�����pbU�����ş�$�ؘ�6-�X! ��w��r9��N�`! ,�x:	�J7�s;�<{����j��`F��HD�b������T;+|��t:�ER��G�d��d�^B״i�@b�N��d,vw<�l�P��8�{�J��N'�vX-�"����R#ȩ<$�Br!��T<vOc�b8�z�����1�$(�Bn���`�wOj�lO�s1��`! ��`��,ૂ\wƸ�Tέ�!���t��=�ߝ
N1N%ۛ�\R�� �$I=�<2�������4�c�p���#��F`!4M�jZE@�ܘN$�a�aG=Ǯ-W���n؇�n��� ʥ��O���$51F@�/k����T�?�k� � ��x.��1����v.�8n���6 D� 7�≻����A�at.׵��e�4u�X
� ����C�����c���P�Lo��R�+�WUe�i!�0ȍ�d�	�FV���0*�=�����4uH=����#�l�Ē_1Z�DQID5q6�я0���;���e�ٟ	�����x>
ߑHL�l䳇d!�œKK��z �%�Dl!ZS�#��E?�9 <ޖ� �F�C���(��h�\��Y}}}�KJ�������-�q�l�FF�KK��z ��$$�1���5�Y�<��m�̓��*� ��x!��l����`s��e��^��)6 H�i���<� �,����Bv{/�"����T�G&�ue�TxLQ�)�!"��|,mZ�s���|ę ��^�F1 �: ʅ�Y�@և��hKE�ag#�y�c���R)�����-�x<�F�L�kY��\Q�p*%Q�H�y�-��C���m�#NIqy|/&b񕍒��b!�L�{E��[D6����7ـ(��V����*I��u�
��H�'k^�}wCD�\x�ߩE�"��[�����0>��P]���`h��"�ue�+����!(�٘N��l4�Ƴ7_z�{@��eL��H4�l��w�5i�cX'�J���Ȱ�Ъ��~1�2
�T��j�B��1ޚjbL��)t6 ���� �P�ý)�L�&64�bH>Do�kY�D�� ��ĸ��M16����K�El!FٓK��"��1 L9 ���Tc��t6{bi��}LU���b(�c$-�Ň(��e�*� ��1F`�� z�'�}�*�4���#c �-�,.�dI�NX�\�zc:oFc
�Й��>��Ҍ@�_l	��h�I�����3��M}zck2�L]�! r��+s��GUM�n����FT&�uy�T|B��Y�C41F(tY� �|1G�t�B@�rS X���\���͝��/����˩�"�J�݌2�@��m��}DSe��*)vc�;R��;�\��"W1[E	D�O��jm*Ȍ	" �|��l��aU�0 dY��N���@pD��
�A�Ĺv؉H��T4~g*�D@�V_���R1�cE��Z�-��p�<҉)*W:qI��?1
�������M�ʱ�;��l�5%�o�,�S��5�-���G��E�r���*�B �����O�ok�Ojj]�&@c*����R��HX��Z��tz���T��{)W,��څ$	�JA#�O'oM�:�j�c�\1sC��w�$������@4��Q�n(�*W�]�ʏb�����v2��5�j�`�㼿�a�\1s= B����y��� ����P�kY��-�ݒJM�q�
�^  �IDAT���,��ʥ��Ȑ%IdY�K�H�Ѷ��m�D�Dbʎ�D�u���G���]-+�ˇ���1B��t2yK<��~sۘ�z��[-ɢv
,�~%�#�T�m煉����� ����QƄe!�+��U2;�DQ`Y�+�@tekkc��Cs*q����y��x?�J/��A�(��y9;��k���Yf؀p��W����v��R���a;����&�S �y�C�� ����3W��샢$@ё �p�_�0�,�..�Kjun�!T���0O~7�h�N�4��q�_ Q,�.)��y�<��Y�"��w�Xle::r�)���]\�7����`!,@|��%�:���!���y�C�� P�(�W���C<�ͥi��eY @����1�\������Oju��~A����_��w�M��8�/gV;3��Z��<W�����PK��F��� D�j�[8�B|K��:�n#�T��ߡQ^ ��º~@(��2�7"����B�\@�A��._�P���� ���X�ɤ������z���@�˙K���:�/Ϸ,��0���(��}��"��E%��D�Z�#� � ��d,��d2�� b�F.�|O�+ �(�z����<_��˸��b�;ӱ	��<�;��+n��;���7K}/�j��D���;M@d����[@�,%˲���w�R�*:~. ��s��y��H�V��$I
[�vƒ�[[���Ne������/�X컨�����/�4˘�pn	�b��R�*:	�R��|!�`��-#��4E'�#��ߖ��;�ag���;�u](d.,��U����\���,ü���iKL|��� 
�ޙ�r��j��� ��)5� �I�cw'Sv�4r��{_p�K����b���wCS-�biZ���tz��F>��c[>W�#��    IEND�B`�PK   F�X
� E  8b  /   images/f891a845-194d-4c25-9fb6-ae7593a7f9e4.png��X�0+**�SE�����EOlA�[���&]=5��P�f��	Ho,�"UCG���;3����<߷�w��̯�ٙ�~X��e���P	�ta~Ւ����\����B�_����{�I�{�っtA� �7��!���e�����i�cΧ����g���Os<%��lѧ��@�@8����#���Ҿ���<����O*S��C�;�sG_�iK��P����F�ʇg�]���_u�O\#8�ϼ=��r�~H)���\.vu��g�1奋7�YVz�������㪯,�RO��~78�K�ݭ��#3�3	���.��@׺�W�����ر�	��DH���+�[E�D��G�h.0�T�Tn�"b%�� 0x���ޢ��J?��Ԛ�$%]���'F, �ߡ 	�qIR���"�=+	�r)���V�L�[�xuPД%������O�*��ф��`U��W*1�@8�[���1135ā4�~lX�m��-m홻p�M��>A�0��Jc�c�z�����2M��ayp�8�_���<ɓu����F�KOOW9��D��?>�?c�)�� ��aD�w�73%��$GB��D0�6}:Ƕ��z����k?�"bp�'ש ����ؐu�
a�c���֘P�7�*�����=TԞ���9�?ߗLtz5�	���k�	(��q��
��۲�1ث<��Ȉ��bs���Ww��V��*m�0��F��f]{�����[���=�W���{�p�% �.y*�R�O����?l�B�:^�X�Uā�8o�y�+W4�<����*��Z�4� �Zv��8�A��(���dg�_2���t�<��oF�?�$��hW���A�rrQҐ��0��{U����k�/ֶ��iP@�aҧ�:W`s���N��ڛì��@`�چ���#�r���$�����j��p����(��A�Z|e˙أ
j�aO�A��zW���j�Pkk��J)�N�M�����2�I�d�=�gQ-k|��J���0<ߐ>��s+�����HA����!���sF2��?�4;^������!2�&��B[��V��u�I���	_���O�tW}{��9���5(X����'F�.���hU��Z����t�Ip�IMJ@���~��|a �
)d��Ǜ�<��B�5�t�)(2�-�""1�ݞ���4mh"��ꑊ�ᇱ��6��'N�H����܎B��>>9C������T�C�@�0�/VGp�˲�i�g�o�dpp�֭[��V�ڪ�5=����{�7of$@;pxj�V���D�O㴭�n�����Smq����k!�WIID111������_�Ž	Sn��j���%5�w��"�MΙ�z�t3	@�������"஖Im'jkM�J��\z��G���llW��ī~��^����xy��ӏ�u�䌌�9��/��#r׆�[����߲fEBcf�`	2�kH�7�����&'�K��ޔ���:�[$��,���)�����\:z�W,���=�l��U�2s���խea�1)�#Ȉ���-�x=(��)	�z��7��|0�2�Ja����kB����� A���<���iO{{�������E�	��ę'�/�\��eM��Ww����{w���qJnUU]�Y?��j���eMҫW�'䌘e�w�p��\̑����z�}n<`�F}J���Jj�Jqj-����e�Ә�.�y�͙�� �GDܬzjP�Ť5���� ����{��XW洣��B�u\�Ӛ=_�^�qC��H���@f���ܹhm�[�Aq�]MkC}���s���)�R��ɒ9��z6`���筭��n�=��?1"� u�xq��>m����i�g�G'+��=�:���L�'�Yy�}h����B��ke��;��ݺ*�4�`��45�˵&콧c��|:� �e+���Ы>v�@P��Nn�;�Yu�8P���Q��c��V���&�9^�ß2�}�~�*��@����q� ��AT�Vh/U�ɣ�:���iB����g�U�ML0Wbc!u�}5�.���п�Y�x��'��At����'�;B!�I͌�ɭ���ڞps{ݩ�A��z��ٳ��������m���LE[K��J{2���
�k7���`:�~������zL��}�&�l[^3U��=feպ��H��e4�8�[%�C�����W�yq�<�ߵm��<	ܦჃ慞ڤ�c��$��Y�~�~(ܕ�������g}n��s�*l L}7��ãG�:ݹ�Rh���r
���s�T^yS:��D�	�Cp������NQ��ϹS�X_wbsz���[�$g<J��ڝ�	m���:�77w�AG����&/Qi��� �M�7��G
��rFm%��|MR�k��yq�EoS�z��t�[��ݯ��i"��Aht�]�o_C��ѣg���Y\R�?�����ص{_�y�Lb�IHcfr0����"̞��_�ʬWs���RܵAл�<>.r�$�t���m�������U9�ܷ��z��^���i:�!3��3�~�cq�����NQ����7��{w�;��zHW�T?jjjz��h�3bbu����&��{��N�����S�%���1�P�/����h��V~�[����Rs�ܹs�����=\c��;a~a�y��y �]D�ҕ���=~�ԟ���
 ���7�"�V��'9wz8�g���{
� ��(��8���ܦt'����	�uɶi��(z����G��F��s��6W�scֵʂ����b�>�R���knY3P�ໝ�-Y�ɵ 9��/x>��Γh�Nk�|�N��v���?����KW�|n��u�z��&���K\��q$ǤU
��*�E�-��@�86���>���0̂�R��R�3��S}�m�c�E��?b�{��0��Do�;~�+{�� ��_�|��I�W�ԭRG�1Y}*�֑��ё�<��ѷ�7dv`unJ���-r�U孲EE�-!!!��z�xzu�!HD�P�O��:���B��q�n���$<���5�<��1-M�����t���ͼћ�.�T�+�|k/��͖8z��Gו������ƚٷ�te�9�7t���\�h�zLA�I�����/�
�x��u/^�H��\ӷE�3�y�T����	"���Z��������M+%4Duuu���E�$n1�UtL�����7A�..�Pn+��0ݭ��"�W3�2K��Ύ�97���:����MI����i�&��2��2Ը1,���44X���Š>�	nܧy�&����w�Z[�����z���a����_+�o`���>4���O�LB�>�#󧢪kjڼ�'�����o2�����[f��Y�7͹ᑑ���KFG=n�X-GL	=~�������D"W�ϛ�v�,R|��0SQr�`(�%�lnh��N:�j)m�Oϥy�{=�V3619��:��9�	|��"�P퉠7���\[A���2i�Kf�B����:��PBqHG���Jz?(���\�n�֘�;�][4��$�N���`��(�ӂ���pp��	�����=7��&h_�	�id!�	����Ğ�Z��2
��D�24�\h6Gq����tx҉�K��`b��z�v�A ����&�Fg��#�f]x���39:����LoR���3OA�7��� {�6Ry��4�.���F�����PwB(煂�|=�G9���gDz6,�=6��v�j&��QhS�����+|�J���P;��@�dN��GU��̤X.��x�}��H�;���x{|��R���^�	sQz�D�x�x������Z�t�����k�����
��:����D"A��2WKI2Υ�\�+Ґ�X%pp��ñ��?8=���B�C����D��3��,k�|�Y�֤O��(�at1+o�ɢQ�>�Y�2d��H��[��I��H"��y9�����#���}E,Cň���/Yŧ�\m���v�c��zw�!����Z���2@L�k��AL�|��@k�V8 ���9F�A�I�C>�Tmqޛ�j�2�����v�!'D�UIy��U̠y 1,��� $��@�<N��H[]�2���eyƆT�x>Oh?�٫����<S%?~��i�NPt�Bf�W\���6R1.�ǽ�'�U
��aϜN\g���� �ĸk#��#�!��Q��gC׈�nH#P�]�f���A�b��CO~��Y8�D�Ho��(�J~T�μ3����z�B%�ET����� ��u��7$�J��GYp����8ĳ�
���e���	I��<L�����i
������Oc���p�({jB���AJ�nٲ%��F����߀pX/��3�(Y��ŗW䂩��������<E`Ùp�q��AJ�ϥ<�~)���=�_��d��"��=��`�=<6���{9	pgZ�<���MNx����t�Gȷ���,�hU0|� �Mּ��6fE��@��|���9Aqy/r�M�����^� ��r��W��Ǩ&� !�T�d���Y�򟳠[A$� �Bx�\��Ho(���7~��ُX""���4ģ��h�*���p����^<����y��D`��Rp{�:�}�v/diC�.?��I�A�4~l�R��u�7[�;��o����K�ۆh��G�,�%�cA�7\[M`^�a�aM"�BԯQG�x}i��!�k~��|'�ćM�Y
r�⥸��1�@�?�t�RhKN{$J�������m
�M�+C%f�{w���ǭ�������0)<B����櫬T��Ъ�|z��y��^�C�p��]��L<�v��Ǝ�A�� 
Tpd>�����A��w�&����q(��[��VJ�Zh(f"������;H�UA��� ���#�f��]����;�6N�\��#q�o�Ft%��٨��t�R�#[��t��Ċ�ED6SPxEF��7���y��گ���,� =OhĭV��O0�.��Fʄ�
�	�_g�j$��!��w����J��C���-���'zG�c�/𒒶⏮�D��D����x�_�Wbs
�(Z�k�]/�Aß��y�?N�ܫ B��GOή�W�&���QX?Bf�99}3�����y�
���f�T�f��b �+�1�T�yS$r�E.7g�3B�DP����$5�r����@�����~�O����A(r4mGOj��H�`{o.]�����"RP���b����Yd2�/�Y�Jh�^�_0~���B��������� 
��|%�C��M�4��C�'�:���37>V����@���з2�N���8����<ovl����.?�|�37��^6�s�R)xwA�t1FP�$ά���[����:��l�<���iWH�u��˯0z/����2�� e���D��������>��������6U1�8�Qȇ`!�� ����91��[4
/(;�a��Ъr���D�l�oP��j<.2p����N���( ��d�I9��H?z���s\�d�,�JsI�7#���`�*�/k��QhzP}�� �ol��Y	��ޓ�J ͷ����[�r����"�Y��z_� ����]��<xy���԰ ˃{�%�ʼ>4�3�����P�J��aR��g�b N! �֞��̬��;�=�	\.�
�YFx|��.4�Gj�/2�29�r�t֏�D�Y��4I��ID;��vVJ(��&#�B� }��'gf"of[I��vHNAa�S�N��F9��ѐ ���i�3�*sf�~�p�Ib���N�*'6�X���e����3{,�*��IQ�b���g]�{ ���o>���f��e�pq��������qoEQ�*�D�hmmt�hn3��(B��*Ǌ=&�aF�ɭ]����D���>���A�����la"����=��mA��=rf�ķ݄��s�hI��[����g�]%��(�3[`a���>!�a�$s֫�^��d��`�%��x֭F"����H��a��2�g���M��X_�-��������Y���L��)�^H��;-/s��Y�/�6��<v��g0��Zb��h4Y�������_o�oo��lf"��̇��^J��~�XCۉ��[r���N���#��Po��j\s����l�?H���i�晟"�?�|�߄��_��a�Ԋ~�v}��Fq�:i��������l�(�9��Nj1�䩈.W<�ES�c"""fڔ}۔�4������ʛ�Z�ʉ)S��b�ڳ�f@k���n�i6���bR+�����驰�!�6[u&TKSi���ֹTO�F��	�mc�Z�0¥�-����3=�>)�l-%4'�G-=ط���.�RjS�_5>�%���$-w����h�ʋ^�ۥ(λ�iP圼���g?I7�ldޗ�>��w�U�;��lܴ��F�v'+����������S>lNr���C�DD�D�U�`N��&��I9�M�T9�}E�����p�Co�`DVc_���ܓ۫q_�gvMfdd􋭼��G�9ԩA T���l�$�����f������맲�7��?���㣼�{5��Y�C�/�.X���}�1�1rP�5H ��_�7M��	���mɬl��[�~5��UKLL�q���=%�Eܩ	�5p��g�*L6@���??Z���-n���3;<��(z�[�Lp{�躝��^���'���Bje���3����L)1�� ٺ�Z'bc�sl~����vr�Y�󬡥����"{�r�ϖ��������L����Ó��y>���V��,+(t���Q8�:��y�=��� �x���(lr�m9\IYMTx��W�>��4��ر�t֞�z�5^9M챱1��n:����N���I�G��R,#�~Ǻ����BjQ������|]�Z~��k�"e��~2���K����6q,fU��H��|���>3^[u�Jk#����K�:�X�-RaK�"��a2�&�E�uީ�f�ܧ���ӯ]�ǝ�]ȍ��"�/��O�J�z�{;Ȫ���\��ku/�����3k
���Q�X�`����:�Y��Ľ���w���z���3�>*뭨��qā�U%L��4����NC�39 T̺l�ɢ�Н��իU�٪��WpF�ʯ�g��M�
+ا����t�� n��M�B�/��=D|а�PA��j�=�>�ʸ03=U.#~R�O��9��2�ӑNY�r��9NRa6�+������Q9O�U�]��%�{{,����#N%_���#��n8#�������1}Þ�)jwϩL8x��A��'�x��m��&��/�����~o3s������~nL�Î�j� �)jm�Wb���\�g��DI�0'�G.���/����đYB{�)��6�z��g����v2��]��7��<<g��ϝ��bM3T�\�	�b(\Lہ9�t��І� �W���!�<u�P�CJL��Y�9b#ӫG���kn�T;P�$��If٥��7�ߌ�mF�t~)�q�;��O�+w_��rPvHͱ��( �ۼ�R^�2Af�}����,�!m	����K���� �(e(�i�����^��	�暸҃������b5pL�6�˩��E����6yX��_w���(*�ӧq�`�傖W���CV�@%^��D\��%��{��-j7}[$�%�;1��HS�pNBx��]:Ug��*�!���ߜ7�ʬT�zXU4L�W��1[���yl�rB�xW�]��U
�	/_Z�}�"����O��x��tW˰@@�<U�+s������{��b�ϙ"<>h�k�	�p�=��/&첲�S�N�lTؖtɋ��e}�a�׵�q���~rlK�X)N�&׋��4�:/��~��aђ�⻡GH�r&[�:�k<4x�8O�5t�`�Mz\���n��f�뫂rZr_�rޭ3yZ�4`��[���A���Ic���5D{Dn���=���E�h�P�C�V͉\�����\���U��]�u�Mc3�?Q�+ʫ�(��lMn�)�n��BPct�)J���y����m�M�8�v�	zc����ҽ�(q`�Q��)��M�ї�ļ��a�����ooo�<f}��G�?bT�ڹDk���t��~J��	G��:�AO-�;�!�jD�x�'�yF˭iHțW��/
�[�<�̋}�M�u��xw�'�fj��������i�+q���� ���~���o_!�nM/�i�V�:)�&0Su=|�U�o�W�-[��؏�iW�b*{oI��K�H\��YuZ�ɨ�� �dC�^<C��'�>T�q�^?��E�MH��}7��Օ)/z(�4�e�ɑ�]�tr�1Z !@ȷ��n��k�Ė/�9�H�ܳ���.�
U�$�"$�֥tʱr8/UbƔ��gk���!�Hz'��`�}E���;)%�2�%W)ǧߪy�]���G��ð;Z�{Zʰ���1�-P�W����Pi�����4\k�-g��X[��4�9Qn��;��]�e�o�a[u�[�uV�A�G�k�F�O�k�в6�c@9���l�ԭj��Y�ޔW0��>n����q4�1:.*�'G;�e��#>@^���y]�	�VLRK4�I3R�M�W�T��4��Y�O�P���� nN���ˎ��1�M1b��I'G�n�RV��d�n�6©�e�2q�:��A�}�Oe�9����T�DO��U��
��֫�(#�\��]�`�z������J�s����va��Ï=퉍Iii���p�t�\�օ4�`��`_�[��1��{g6�M�+_*|�����)@,�'_��as�K�X��}�!���r���d֐��L��ܙg�&28�Qĭ�d�R��*	DC@��Zwp!�,E��3�M��W��k�0p.{�����6p&�,\��qW�#�h�,�{V���ުfӂ��n�z{��D�
�{�l-t8'/0�~�,kHns�/ρ���
o �ӻ�>q�o�rC��t�K��/A�p`�\�/�5��o�{�?�!������bJt��1u���ђY��3�닸�"o��o �����������$M��D]+����Ns!���b_��L��Kjy��2��f�?aE��km9�"A,�]<��Z�u�J�	�/9�ڀ#�R�o�����bQ��g��"n�`Շ�����FZ��;TO�"m=G�9����2�Ժe�50���?��/4��D����i���Ο$�\	�t�JI�I�jd�A��F�狱�Wj��x���.�pBr�*�!�y]ҽ�i:���X!�a0n����Ǥ��H[)��k���E���3װ ���y����m����s�f���C�)��	�6x�,� ���1&��Y���)Y���&>��{e��f����*��-ñ�E�(�Xd��걌�-h��L�6j�\ �KnFD��.�`H�����e ��U|�a����1�f�ʊ�jf�AL�y���䊥��o�ЯR�����Y�7�[O�4��ª'܊kB`U�����x�Q��PǏ�!Z�"��_�S���;`|�g����f�$h�iJO-��}�n0�CWΟC8�D�*'��/\~�~3_PȍG�MT����C�.�� ]=~���/*�M\�:>�S ����	L�nB����9_��s��B���m�5���g���H�y\Ψ�Gi0GSpnK��*hy�` O��T� u���=_ߟbB$�rB �)/b�J�16��?-�`���L'�a%�MX}�
;}�L�Y�T��Gi::�����)��p�|�	��N1b�����1�/'1���zi���+@�M{f���Q����M���m��毤�(���֗M�{�'�*�f;����{��'l��@~b�{$�ѽ���jsJA���*133s\��Z�ȱس�J��t����U��
�@q��D���3�cp�f�DN��� a��=� �Sz�_���9�s
d�g]�0�@j����_zBq��͛3E� ���1zy��6������H�)�r�Z�GH���������Ƥ�6K5{�:�+�:��w g�Z��le�td>AQ��ڣ����6���3�y���O��[��/$��l��Ξ|V����9v�y<|+X<�'ߦ����z,�4�ܽE]:�G��sW��\��w7k��n>�v�3gq�yӽe�3{��1�%ŕ�t�Қ�q{z��|���ȯ�}G��z��faa1��X	��5۟C/nq�l싉�*�:�XNf�l�M~R��ē�0�A����>_���JsRkG-?�ײ�u��A�QD߫$#=��D�A��{�k)����CU�@�v�w��O@׋Y}?�t���y�qh��[�aa��~Z�: ���b����,+�=���}��1 }��%���E���g-�#E�<�� <�{�Ի�F*˾򩉉Isj�B|w�`���8�i�:��_3q�*Ǻ8D�`�k���<O�t��D���՜�OV�H%S�����L�}a־c��������q���?5��y�`�U�����:���T�Djg����]#�_1�irr�\�9��پ0+�Ni�˛�m �\�%���t�a���H��{�&;����M��q���xJu���.S�.�ɱ��� 1�3�~���MA�6�� �1�j��"g��¨�Ck����Z����j>��|�^Ė��lB3}O��s�E䶽���J�� I��a�r2�N��\wY٧$ö<:�jޱ��Zq))C�7���߼y���5ڧR�ޟmGjm3W�������˵����z��Y�l(�3��kR��p��>���՝�"TNN@��f���Y�����]q� at�t��kA�$���KV�L���[�2�=�N�t����z��菅<� �W�bc���T>�>˽_+�>��Q[�,�I�"���>������l�����|}���������L+�x���*��i ��v���) $�m�3�Q�|)�ϊ�}IP��Yz|���M�i��W��� _R�"{D9�Y�@'�-��>v��U~T1P�~� ȎR��-2�< ޫ����й�2>��5zq�4n_����OC��~+ZR�3���~��-��k�Z�J���ő���&��:���"�8�V���Цσz����j�/%�]W �ys���@IK�]G��2_1�џm���%ǋ����K�KP�n����K�����k����w��_�cǾ�fx�i�GH̹����k	���>�hM/-�N���%u�n���#�jl�^�i�y���Gt&[*++�x�t�HZ}�V��,�ٰx���[��(ҝu&?��d+zܲ�U�2������-	*f��5�]z��}
�+�[/K��Ƚ\y��FkK�I�������������D�*ͬ��3"���#H���sf_>�6���y���.\P%YYw� �|9_8�@�׫ͫ��cH�6Nv�I���{��7G����rP]H�R*{ݸ���'d���L���ۺpu�?�|�"�} ��A�n-�pS�A������}���U%��kc�a�){l3ú�c|�K�H9�Ŵ���a����Of
^@f��ӌ�h�D�d�o������3�cD��p��Q|FBFF,�EԻ3���LW��O�[�G$z��d�ⰣD�]�V��|��}m�]eYϫ:�����n�n��@kʠs�u���,�_��4�{�ӹY���|�"������t��['�E[$��������l�����s�j$�O^AatiO��6�ǜ��`��1�^3��k�1�\{C���珫�i��x	��O�&K���7�1��=N$�k� 5����\���[ϔ��'Fz��I��*���s�H&�>�Y����w�q�t<��77��߀3�14y9��-�\%�t:|��wΜ�a@���g�]u綤�OI���������N��� ���x�;o�ٱ�$�P����Z�锑��9V	�;c�ϝ.���P6��:/�U����Q�1�]Z��Wk�D{���D�w6�u,Ĉ2�A	`ȏ��8u�VZ�ynq���c��u�SN$(�
*Al��1+�����rܭ}�n>a5Hl]����S��ʽE�?�XOٹZZ���F��3�έK苍���m0V+M?D+�J�I����7o&�J1�)ҕ"�	\DP�}�,��u|{��G��Q^�$�ɫ��g�3t�~���1�	$�����'�#�61
g�0|����4P�+p7��Q99����.~�:=�T�TH��Θ�h��7@�.�Qm�/�����Y�E:>� �pǩM��J⦂|�]\ mV3��M$چ�Ѻ��7��,�R�ط�9B���ęԪ���A��s���D���V�[�C@��dx�t,�T�Ax
����T�rsS_�*gƹ��m�)n_�{�J��z�A榦�T�쌚������X� �Ⱦ��W�#��	�Bi/z���>����{||ϵ�>�5ݟYB��o'U��~#J� JN W��<E�%�~�d������*+�/Rw�kc����֧&y�\�D¾����/?�sf+蓧"��	��Yb��u�.���:�@�
�g��k.���S ���(��dV�tf7�!6����	�ԏ����	Ў��\a�>]�3;�*���ε�ӣ@�I ��<�����e6c�*����?� ���Cs�]b��I�����>]����AIN�̏�{$��=];�{Ԓ��.�L�˩!:��]�XWf|^n|7�1S>�q����p7p�?�������Ę���T��C4�Ϸ�	���O�Ν6�8���@��#����(��1kמڤ�댛T�A �/{d����8`��xP��x.B߽_���#�:8�c�3J��|&���szoW�S���T[ַ�Ո�����Fkr�`���@I���7�s)�����T;�ɘF������dD[6��.KZ��)�V����St���c���NQsB�a{���RͫA���x�:����|5���ͤ@�Z��ק�#��^/u��$�#����=�����5�So*�Ϛ��r�h++�ss�M^�	5����lzE��vڠ4h�$(�a�����[��/5o����h���r�Gg�X�E��4� I��w.��z�pY�V9�ɽ�'�������L{��7/���f���B����j�מ��>i��36�_V��A��V����x(=E��^�b	�~z���N9�G<�4����9�A��(I����/X?���]��>s���ي���?�}+z|!a��,1�1uGn�}����7��:��'�p��g�0F;kUm�p/���~��-���1F���Z�\� d�� ���d9_\�*A����6w������wV���=�p���^W��Y��T�+w��:oO�󱘽+��y� ��<l���^*�k;.�ӕ��^S�b���(��h���߿�e@{�8^�7�fߦ'���P����W_F��J\F������k�����	�u��M�؃��$
q$
y�I>��� N~ϯ������<!��B�>��maY���C鴁Q��G�g�?���TE��� �Bb�T��qC�μ�㔻M�6��j�O�q|b����y�ˠ�h�$��b���_��ӽ�����3����H\�k�-��D�}҇�T	��)��R*E@�������U�1��&2��p�#�^[�	�/��t:}.��Lꭧ��}G.V��+�yN�1S�&�Z�XX>��~�5D��ɟ���d�v²G,���hׁ�:���85�ி�:Ytl�m知'/m�x�������m��}���J�����O\xog��r��);v�4N�q�4f�+��'j���'�p���'&Z������~��m���&���ڕ�h����ObVd0~�ߥzl織_\���ľ�[m��N���n받茒.��a���G�YV��;w�o������	w��� ����ʣ�V�pc��j|����z{����[o���Sp���ח���8�휥�
��w�Ejn��$�����b'�w��ZpY �)��{��p+�<������7���K|TL)1�X��Qk���3���*��g��;����Z��O��'�` ��{��������WB
���������������	�O�F��;�����eH�w��÷D��c$�p���C�:[��������p!�٥%	'�" kK�{x��4b��OB������SE2>��غ������9�ǏwD������6����� [\&����}�D�P%A����O�V9�GG���ّ\W�C�iNQe�#&��
N{yM�N���ʏE��s�Y��j2���O�� 
�ь���&������w��Y"	!q��☞��;�6�.�m�ᔠY�|-I��o�Y6������5D�:�p�|��<�M�nSY��O���n~�'7���q����8�:)�,��6i��qT
�J�'r���"��:o�?�ѧ�b=��i�F� �w������ aW"\Zߔ��u�w��~�g����d�	-��w/��~Jr���0)�|�*��7���_6ߠo!l��p�EBxMV��M�7��v��ƌbMH L�ғ�� 
��ҿ�H��b�&����x��CR��5�E�
�lX��?��Vb�.N�$� Q�7:j��X�G1�RN���)������t�G$�/��b�~��{3�ג�Ua4��4ݥ����q�<������`w�]�22�Ȣ �)������?~�@�� gz��?i���@��A���Of(�����:鸂� }�_:=���#�t���� Й$t���Y�2���AN-o��9�Fn���}!s]��,ڽ[X���x�
ȌM���̸���<w�<�;t<f3ns��s��ſ0tR����9�F��޸���� Y�}{EI��K1)�F�d+Dp��T}}L	�2�3��G(�W,��������﯆w�U���$��L\L ���8��b�Y���7��P�7���x��I�oae!��p_�]M�g1C�70r%���9[���L�6H����a�k�#aT��g	e�z��8�Vx%Z��O�@
�K Yt"�<"�J .���P(5-��-Ĥ0��Q�%%�[�.O�.ƏC�r�|at�\�ĭ(�֊r�8�V��,Ӌ�|�uJ�$��)ɡO��T �*� ;2���蠼�g��Op��#v������7>���K�R�@R5@��R�94A>M���׵�oZ��,��H��?�@��S�K�������cA ��.L�a�,¾��I�}~�]ܹS�Q�m����5E}�ʖ�*�T��9?C±۶ҨtA�%�0G@�>�eEB5E�fRÏ`��^���;�O�Ƶ_���ˠ���eV���e�2�[HeG�C�G�U�cN�sq������q8���ʁ�$�h�T��Xȭǵn|Į�x	$���p�O3��r���o~�������,��T���r���oF�MҬg����K�!О�N"��:�d�%.Z����������̡�����A�/���ɡ��%H�/R��54Vϳ�h�,�~��&�vW��ͽF����R�yΤj��<P��3�:��w�Cg�E.�h�%}t��<�zzz:ʬ{
��$җ�_��ÿ��&���l-#=dRݸ\n�I�5E�JR�eM� P�Ŝ������1_ĿY�#��6��v�{��ݲZ#�E�h��3xX�����%r��:�1��?6:Ψ����N��kzuo�����?Km�kjM:.m�|�!]��O���
̕0dG�F�9��V���t��+�:�8��,�O�Dr���Fܖ���t��ms�*/�lG¦:<�6�;N�>@���A�+�~�ԵА)8�8�fB����<�+R��|b�X,�d9����>6��]���~-�t:��?���)|F�M�������1�C���pΦ��/���&���m�L�����gu��rRS]ա"����tN�0<Ҭ{?���S����BE�p���aY����3h`����ƥ�j�؊`��<W�M=��U��;fv���#���p�#?Omj��˸7����G�ϝ`�NDlK�t�O�l$=�d��/�euMm	���ly���##���>,0 L��	K�ފ�(�?�}Ƞs|�`�!��jA*J4�3�;Ε�>dK��+�W��c�����/�zlQ�λ>�~��K�"�̎̚tG�GO7�����kz�O���֛��]H�|�m�ۯ�����+\�~�b@?�*�n~���"uz����
�AB�W=~7!���-|��-���(���%%W&��&��b-����ݰ4�1����XLI�2���ln4���A�Z��^9'��8���ڟ=��_��Q��8�!�Z�W�t@:�f��1�7\������&�iΐ�{���Ux$�]i��{NRژZ������$�b���y���G�f�$,��"����܌�߃�[f��:ǹj�`���c�ā�HKbH����	�)����������`1���&��b�NdU���&�i>D��p2�m4�P�d9���2
�]�����/srr�R�p^�u����"q�#M�*!L�iVc������Z�M-6B�����"�9��%��G��B�+��f�x�����u����)|2����f���-o���a;9�@YTT�D�9��"Ә2��:i�����	���6k&�/=��O:{yM��ݒ�.�_Y�c^�o��h�N�Y���������F�~d����u��Ǐ�H g��y�D�\Ո2|�Jvo\*�5	��(�UA���S�(�ڱ��uk�*�m͘L6�!===A����R�C_HKO'; �D�,�#b\ �v�n��^�C4f̎O���(v�	�!���m�Ǽ��JY�+j�S�ߦ�����ȁ)�0���Sm6��J��Ԥ$'wѫ���$ma�O�kl��n�4�煪���¼�p/���=k�~U ����U�@#5.n�p��[��9Ʋ�Թm@sy��m�9���uuuc� �M��A�l]C��!�^
��XZ��^9Ҵ�RD������0F�8�Тlo\	��s�Sg����~$�ٿ�JJ����F��i�To_��HGA�d�W�b	فfݗ��GR9�3Ӡ������ӰVl�U��˛��+�~F��sL5�$4<8��"��r���S.�^�}\�e�~g*;���B�e��G��էYL����C�k��	�o��!3�g��Ќ�U����@��6���#d��p�0q�d���}:�v�N�VA�UĘ�RS�FM��I�2�?�۴�o%�Ԧz���{�u����� PK   ���Xg�	�;  �;  /   images/fb3f2d9c-813f-448c-93d4-6d887e4d49e7.png�;"ĉPNG

   IHDR   f   �   ,M�{   	pHYs  �  ��+  ;�IDATx��}	���U޹����{�tO�>�F���%y`�8���U�@0UvA�	��(*�J��P)�
��TŐ ���M��$[��K�/=3���������ޜs��_���5�=Ӳ4}GO����������ׅ��9����9��A����v� tSݕ���!F�o(�h�8��(U��VO�z���G>����ru[�Vl�Z�|�pB�:�zK~.7���|b�op�\�n��}�n_5�M��t���XT'�֗��������j/���XZ��UY��͞D��(i��f+�C_ű@��@����Yw�\�b�W� ����R����ᯝ��v��Y���/��h��f��RR�8����S��pOuf�=aeiOZ+#W,���f^�0�Ab� B#=%��(Q��W-h�g
dT�F5��:���|�����g���=�=8:�ߵg~�Ï��u?p���ꟙ>����n[����������hR�� �s�>NpA(p]	AP@<"�"#.Ci���F� ���#E*��T� k��m�gv�܁P���K3��ї������>�_N��8�z��0�ܡ�ą�����Ͽf��;[so���N�Q'��\���x.��@R ��	H0���.�I`bI���F� ���H�$I �|�-*�+"�v���j'^<pl�����v����ϼ��=�z��a.<����yꮋ�N�b�����܈֋EB�# �{�a���7�HH$��N(� �-q�@�X������0<6F�A̓��<?Cj��T�Lu��N�w.//l�T�h.������/�y��C����f���JR�SO|z������O��jTz�ro.jB/rF	��D$�4�����[�$k�%8���$,�x(��H� ��s��'�C$�_�������{x6R��>�4��Ps���م�۪s�w���/�����͚�׍0��Q���z����G���pT/����/8	t��9�C��cT�(�H��W���<�	 ��gp��!��Lx>��N6��u�	�bO�ALP���!q鈞�L�jI��6}z������G���߻k⾏�q|���u!���_�{<p��'?]8�`W\&n����$�����
��p\&�t�Dс'�a$&��qʉ[�tq�`U���!�bb(y4�m��D�k�,�H�U/@ei�R^�q�]��/>�ѓx��r�6�0g��Sç���{f��h}���u���M!�\���H��ǟ27�\�P��M�F�0K��0Bj;�4��	�ӌ	�q�
�X���)Ii�;x|����ŠB�Pm��&��=R�o����6��.��|�?x��?��5Cm�J��o���o�&���/���]��
��"�'�E�k�=��y@���.1�		 鐎�ߤU�Ff��W,�H�1����?����A�&�;șD8:׀	� 	~�uKw����*���B���������L�Z�զf����<���>|�g�E�8yk�
�@��"Ί����	e>N�`�Wx�Kڢ���L�A=㢾p"0gi�C6� ҈2�-��4s���H�����xd�xL\d)�7�72Rk��ʝ�'~t�U�]8������O��|n�j�צ����>����:q�#�:Ӑ�B)�� ����<g�x��O �IK���PZ��	&V����Oe�@zE�"��Q��sF��$�n�M���t.�_�r`��B@Dt�y����ʃq=X�|�?�+����_����5'L��W��~�[?q?ܚ>w�0e @k��LP�
�r(�"�QXޓ��P��$yB3�L&�FbL0�w�ETtLj9����0 �o�#��G�ȣk���b���hC����M��F�����(N�M�xs�t�S��_���}���kN�������O��X<sp�kAŒ�J���c�����Z2I���~`'�Vp`ŕg�> C�(wc���c�9�!�F�8bπ�~4|��d's��#�[��'~�����=��)^����5S�9=� ���8�+��)���������!4lp\S�L~�<x�[_��x��=EՄDX|p��49)�+�s���l�8l�V�fŧ(��j#�����Bi��
,r3��F�2���M�^d�n�&���1��5X�I�(���;E�NK��	Ҵ{wOij��O��?�4�xa�sw�s�П�}�[_�׍ٙu���I���hl�����]�+��1�65�.mջ5atgW_N1怰�E�Z����hKxm�Y��]4�j�����ip����b4�q�c�V�,|�q�d��?�7�y��~wz#�wM�x���O}��'μ�ֽ@�k�'Y��M�k���!C^im��0 �§!����He�B �!4#��O�
aRm�tr-�:߸u����NVGj5��|-6w��x| U�?76¥����'����?����kB���̜~�C�2�ÃrH�Ns9Y_��9l�3K��.FPU[3��3��E�S[0�`�ȧY��eV}���`��_����5�s�1����lW	퀏��l�G!t�n)iWn��]������>�؋yd]!�N���>���S_���Թ��NQ���i� Z(^��)������
{���	dq���F��9:+��"�[�CL+�` o++&3���,��C�W��5t��H H�ѽ��ҁ�$~K4y��K;^ }v=�xU	C�����;������5�FA	o�gW��<��3�q�Hᬈ0����Hɂb��hW�9�^[�ɒH�>t<r�  ֠�tN����y)���k���t��p���C��w�UZ�wϞz��s��ou߇���Z����\�;�S����R҂B�V}b���D���e&Ա
׈Z�B�$��g�@G�n�CR�O�>�}�p;#���U�"���҂a"��} ��zTjU{�w�w�(\c��aL1�t�赖ʻ���x��a}��S�ᇓ���U#�~�9o�����ɷ��ZŘj�xÞ�K� l3��� �dq�\�r(X�/I9+��g��xU7�����|< @z�m���!f�F?D�$Xm�4�е!
y��p���0Ǧib��ɔ�Ayd�\t������ M��EA��ZKOyߩ{O��%/�.�Y���g�tN��:��9W.�)�	dI^�ƙH�6h�a+ �#AYߕ`ģ��g�n'���:h���'s�k��B�B�O�Nd����H���Р�Z�:,���?e V�ޭ�������$�~�-�`������׏=6#y$�t�4'G/?�@����FQ�!�B(r�;֊w������,iD�(Km\+2S��6ɂ��&>�:�'�[���]����1b��@F�[dŜ��3�˃	c�t�=P�R̝R	cWQt�@M�Ǧ�k���z��{���Sx�ܦF�;�{�;�|kX��n|���A`���p�t2��������b�I���[�aXl�za�G#�1$�h��d�Fksvʈ�6��DΦk|a��+��K�	,j3{�a�$���� |&�w+H���z|�giq��Z����&Luzr�2s��|n���d�B8�F����n�Ҋf+=�fe��ϋ9�����+���Eb�6P�����l��1��8a�3|k��q��v��ݖ0�ڼi@�
̖�2;^���$\rx���~�n�\8���_�뽍+����O�k�*�S7�r]\u�cn>A��\�<�8�VDQtkI~xZ������F�@ibC>+i��X�%D8R�81B�X%��R��N�Xɱ���Ҹ�H�z��j��N���O�̸:�,���ZW����"x!��(Up�&��k�Pr������s��O6�0p��]]�}�U]�I�0��Vw"L<]9d�$k=s���HS�g��L(�X�4$��Ajh#�b$y�(=�4�4�y9o �c�֥z"�(Fs8���x9z	��~S�ӑ8t��7ܱ�9�9����16x\\m� ���(�D��"�єS��k��#x�Ħfn|���44�}�
EN�*M�x�}�U�ae<�:K v00bBJO I6
��d�]Pi+�[l���L��!� }]�q�q5 <'!IXS���0����@���G������;F`�' �/�w��o��hEduҠ`��W�)	��F$3G��g��AqQX�����8u����a����Q�a�����j��n�����H��IGPBE��b��� �u��EE��ǢFWX~�8���0�W�.Ñ3e�]L`��� �?�y
�;5o�?��ta[	/��<�T�W.�g'��N��5i��,(8X��=7��-�]�G��m0y�W@
=s���g�L���Ak���1���r���Dg�B���{��؟���m�NO�����oە��EXߖ���I���q��J��"�21������tC�zA�l��!s�f������46�ϝ[���H\��"�A\�1r�2��9�rszs���7�g�ੳ.��]x|w���P)+8=P����B�+�������p��HM0��{3hRZC�eǀN�����ͪ�<�'�fH`c�����s���z��c�&ޒ�ti	���u�� ���=�N�Z
��	�`�����jp�,���}#���ؽ���s���9x�����&��j����#
��ug �z)�ƅ��1|{��K ��kp��E�d�m�e`�/F��eE�)�1ݱQm^D2bU��8�o'i>jׇgwh}���E�!I#_)��N[�|@V1q�b�9Cz,�س+&���S15�>�Q	���vQ&��!��@i;�p�̓p����ӛ��.���AWC����O��B�yA"0x��}�k�mU��b��N���&�+�� �(Fͬ8C���MPL^b�|�.R�ۥ�Ј�Z��m�%��C�S��M�Ə�o�ӆ�h��v�ܣ����mORN�e%i��J�o%LK��R���A���2�QQmݾ����Qq�$0�,@;N'x�����瑘%߃����E$���nn,�Ѕ7��oė�\����Go3]�\	�4C�W����Y���rvaj��6q��o�8_BzL����7���kJ���8���n�Gq��wv��WA3�c�ghM3�N��cdƈ틂jí#y؇H��8SS�U����&*E���(��g{����n�Q|߅� �j��2"���)`9��@�L@;Xy&X�4� 3xU�a Ftw<�2�%�%�K�x.��$׬���8
�5ƺ	��c��7&�d��S�7o�1&?{�W����Н�G6� �CD�@.�p|%��/jB�^o��ܲ&����\(��|%\��w�ax0�y	��"���+���AE`��Q��//W���l'���G�ۏ��vb0J�>e���/�q���8UJ�E&3����ğ�4NW%]�U�c��漯�c&w�����t�����9Y���X8iNgB�Ih���)6a"*�ʵ�2��p%�KC!!�B�:������Z���=��P���n�ʥ F�Z��(�=X.��p��4�D1��u��h�����d�^2Ѻ���Ў�+���g�D ?��!mk0�z���-;T`i��2���Y�~�^�iX 6Uho�T�����j�+�S���m� 6%�
1$$*y"�˖�b��B#��Ÿƪ	<3>G�C�-l�x�� �C����=d}��� !�;�O����y(@�p���"�$˼��8�V[�rJ��69P30��
ZLj�4)Qʆ
tVnh\M�%����
�F�T�����aùf�q˦Z啊��`�f��J�0O��/��f"�R�g*K׺�����q{�Ԓ�Ó8<т���Q����w�}}�K��8��-|�Dsb>�C�M�����;�m�X
�{�y�x�v�����W�����j{l�
&�ICd��Q��&�ȃ^a��MDR"F�Wd�p����h&4̉[�處!;&����HĈ�U�b�E9�hm����G���3����A��u�(�{pv�ס�넪Q��D���"*�gg���+�0�D)�Sޱ#�P{ z��W2�T�����;���m����Wd��a6C8�o�l�l؃ӧs��
ʞ6�ʪ��-�lo2Si"9����y�&���PdIt�˽]	V�����#�:ha͡ayd|	N ��o�$zp��~ؽg��\D�6��-�~s9/��RO���ED���G��^��Po��4�xOl�.�$\��y�hK�}9�4��4G�w`�.j�{.;&A�A,��H��5ƺ	�b��\V);"�Ũ����V��o��CpI,9J�J�!���LJ��h��b�96	e4"��PiF06S��G*�F�ޑ���~h$)�|bNM�Exs�a^�tAs*D��6EF���م�@�Ђ̒�M� M����BX�%&JN^O��U�����H�M|K3��>v���k���M�4/S�u|��V8}9%��[&�l	�2Y+ʪc�C0*K9�I1��ɔ��(��x�t^8o�~꣱���$��!��Н���C����
.��JH���<�M!2��H���zp���4�G�*�wV��rR�c�dz$s�giO��X=;&�C@d5��h�u#�s^3cf݄	�i��2~Y�"̦I):1{���6�5#�F�*j:�P�n ���6���ߦLH%PI5����B�h�Dh߸0SWPn��F���G5����d0��5��J�A���	wd�;��\��SM��*.�"Gm�*����8mf�0���L���d��S/�np	�}����Ū�^[��1�3KL�>+x�/YL6��5�	�o*z�Y��-�{`���F`_�)E �����H�"H/���7��=CЅ�+h����;D"�� ����D��j�Pp�u.��)����1��˄+�R�\�����Q�cML�q�[��鏂�0�NLiMD|&�#a|����T��W��}0Ο:^qe���Kx/	Wz����"��\Wo�e��L֢�2���s�SQ����)n��<��ua�V��xTm�c��"1���O}|5���J�zPx���=�K)mU�؏��7Z�Z��S8�5�/��-ׄqpR��&wr���\e��Ҧ���������N��I��W�+u-��k�3�.#{�����A�-�K��s8��9�Eq�Bj؛��k��H�!�1%x1N�buK%�f�BQԄT�����S�@�	8b������� �/�����v3j��� ��'HF�yN��& �G���Wp�N�Ao1@.t�B�I�"gc���u5?���=:1!� �|'�wy~=W��
��6P�z�p9N��߁�$)�/@��\[+itd�eޓ	'�tA��v��9��g/ ����8'0��(������5`���Rw����F�	��786�-˳p��4���<��?��]�(�lK����cu�#�t�+M�:U�*���H
�a�T,�W�|ENG)A�L餎_X��i��kK�Bow�	
���[:�K�6%�l��8�d����Ҭj��T�=Ca�B�����~
%R��EY u	����K��z(Þ��&N��xN	SdhZk4��l�ek�Z�&�(�')�ӗ(A��jsW�������2D�%	6#�:l��Y���-��60y�0����3DT���+K3B<r��2��i��ɴ�k��UJm�%��Ѹ�ہ�y��J��i<\���(;.�9P)���<���e7:n�X�Q�rޱ6e�8�8%�V��C.�c�Fɤ�]b�3��1�4��	�!������PrѦB3-E������d�Q8A��ϱ�V�Ԕ!�C1Y����A��|a`�3m�0]nT�y��t�g�vm�C��Z̯-�׫�2i��(pj)��h�j\VZP���&1�b���sh�����XLĦ�X�@�u�x�&ݥ�f�!,�R�gnUHQ��K)��Z��ws� �[����n�HȦ��/'�,T���\6��K!
�g�"�5�q�����ȡ���+�	�!�POɳ��7�K�hwܔh�z#�.��	��Dc�@sQ����8o�᎗���񡢲s������Z�C���p���}X���5��)�D��i� %�K˾�Z�������V��B�^g��?0sz"pi�2�''2W��h�3���}C#�����͆��z�z���31��#v�zBZ�VmC�W�"��,�Nr���	��2:�?I��:?ST����|m�b9q�����e���Q�+&�S5Xc"1��a�I4G4����4�0���Rќ�0'���(�X��u����2�E	�.{�CWܤa㙘������݆�{o�Q�̺t4h{xd�:S�#�w��(�v��T�5fYp]��,FȸS�~�׎�x��$�ë��";n��S�6KCX׻�p��V�@G]�� ���v�d��N"8#�y�ia 7K�Pi�7�K2IV< �QfZI��[H��f\�����\qߙ���g��v��L�\څ�HƈC�h$1#���"�_�L|������L�c��n�p�d8�Fn�C�¸K��&�#�i
gBUY�����$��,صJ�R���J.c�͡l~2UP��'S��B�Jї"�0ٰ��u8xnD���D�
�j��#����Ή?Y�4��:��O�5{N5+�\O�$Z��c�q
���#�.�D�ULB�"� ���S`��AeŅ.T��s��uIG��u�Y
.�ǽf�
ߣ�g�|B�=�t#��h�?Sn�;���!�Kƣ�����9lP��%�PX$&��Ƕ#u�v]8�ޝ7��=��K0h\�2�8R��>ۘ�����a{Fq'W��f�����f�=�skrK�)[A�H&�&� ;�r�Ä�~�ƀ�I޶���w8,�����.��H�
ٹ�`7�0�G��t��X�dE�\b�<w"��o�6�Et�x_
�� ����gGw�[S��B����Js`�ӳ��1�z����S�e��S��P�ְ�M��n��eb�r�H^g�d��bʘ���2�*l�����V�؉Ҷ�)?$W�(�L�[ƖYR�&�$5.Mu��l��11L��D��Ϧ𗂁������p{�	C���������r�h��j1��Q��l���Qsi:c�dRe��q�l���fu�`�j�#T\���p�]�
׺�{�1`2Z��s��-l�l#B3����R@֧��¤u'�g�J��=zn`�>�?ㅛQ
���(�Ln�w��F���I�Ѹj5�;w�./�v~�G�Q<P���#LJSǹ'l��˞�:����%l����lj`��DK��r��n�*��[��I
ÝY��.҃��8�WcJ�;_�BCm3*��m��q'B�p@�4y��f!H)�.�m��̞�w_�W�0⮟k���_>]�:}2m%����9.\5�v�4Y�M1�?׆�؞�U+��f�����F�i;ѩu��)tB�����V%�12�+aT��R�� �8Y����ur�W�~a��0m��I� v��Ş�=û�z�-{�TF���ڀ�޲4q��/�5���bJd`��K��$��g$EMA	�f�>+V����J�m���'��bz�ƃ�z%n})��� X���'XQ�q��f&#��^ �NZǈ���)Q[��S�t�ێ��v����qu{�l��)���E�����N2�<�L�f-tNf.M��%�*[#��:�P���ڢ�9N�7G�Eg���(+�SG*��Ji�{�1Ft��W��6�$n��J�{��]#����8��v�W�0{!�A����4[��r�!i�D2��U��%i���u�������؛)v�n��7V�\:����LWA��1�1�I����je��v������Δ=��|w���]{��C������%��]"U�S)N'"O_T��W�	���޸x�J2����.�Y�
@G��ÿ�`�W�l��	3��V�Y�:q�°�-�R�'��q��y$���N���_)��W��J����\���8��约���}�Ċ&e$[GIk��M�$]<����t��/bU�m�.%�X���y���_�x1��H�T���G���H4	�ㆱ�#8#D��s�]�oh���J���cЪ��괟�ʹ"�<�}�¾J��Z�t*�mYXX�z\Z~�m�s)��%�0���IG����W
0- \�Uڱ`e�`�d�R�-%�p���
�d��S����Ƽڸj��;���#O�
����"��Eh�� N��]�HN��/��L/k�i��ǭ^���
f:�Z�	\�fT��k]*�lQ�}/��8��D���{6Fd3��e��crf��ϵ�K;:���f���W���~���n)�����.ȹ��y4�y�#���mC�q\�WW���Z��}�Z� K)�����f@IَM��ҭpY�OfֱlrHV�M[�lG��)�O�{fdH.s��m%/J� 窧d	%�^]�x�{�/W�0'�zl�≗���Nҝ��B�+�F\�B��<�>��'��(�=6��N�.�2���iaVq�iN��n!�Cu'��f�^�%R�l�r:�h�$SТ���ۜO�g2p�#�u�s3"�Z�8�R؁R�<��YF�.�"r��2UP�5Z������ė�f^7_����g���iu�IcG�\�I�n¸�7�r����7e�P<ĕFz�ss���%��՘��R,��P����3��^�Ĕ�1f������rR2^��ٓ��5/��T�
)v�,����7��	�$I�dE%�oFe՜� YZ�b:cࣺqT�Q�@�4�>����b`R�c/��=KS>�ʷ���yW��(���c�b��X�
�:�J�P̟����3'���e��mڳ8G���2S���C`�IX��u^7Nl�W�{#JY�0�A"V�$E�# �U�0��h�ʛ�wR��F�L��}�l�5�e��K�
�7n�֧ν}a��g�
�-\u��5O�>{������}�v�Z��)�!�Hnq|��/@�W_�f���#1YK�"�5]�^FCN�|���b�.G i˒(��_ӫ��-E$�A(Nb�"�īLI��~�Z8J�[s&��.@�&��#�H�;H�q
�K��rh)3tN��D{9�L'���&[[�h��(�IK��n"�"A���U�k��ݛN���o���O�W{� �{
] AQp;�ز�/dsJ�u)��ʡs&�_������m�&�z�Imz��Y��o�/��٬�َ�{�4�s .PMQ�@�-�BY����)��P!8��9�
eӓ�W{NMT��Nr:Rݦ�>x7թ�@��Q���]����trȸ��nm˩���8TЫ�iZ89$T+o Z��_�p��+_:%���5��'̙3�.�>�a]_��ӛBO�C}B�81�JN�}Y�j+Uˡ<��/�����il��v�xf��;���L?S^�U�s���iXߩ���z��	�.�Qż�m�E�ET��������[+2<�&	��y���&�Q�1�,I�6���J�l�����ӲP<��{J3�Cݨ룮��xkua�G����tG����z��M>A�:���ř��oWG���|b��S���o
a�O|���?<�������N0���娛Rh�)�:�B\va���K��C]����o=5���_�G��啕ZC?����x���B8?��,_�7�w�v�S�4�v�x�
D�W:��T�(�4�l�g=a��JS41e�g�O�$D��2�n��9%�-�9o�~q�w�22�@󦏛���r��cG�GNT'�W��~$V��n���J�M�P��]�Ęj��4w`���w.�xh�״e�Ӝ_�͟}/4�G���Xм�n���Eꀻ��c���74�����o}�{O���xKu�euپ���.�?�byj��U���./��j���4�;�{�'Um��U�'M�huR��;Q��B�-���F)2o:�Rl�q�1�Ou��\�5\q���"g_���}�&�}����C�~z\�+��d<_�{����]�
I��G3��
)�[Y�14;v�����	�����?{r4^��y���.B���R��|mu����-�;����O�z�C'���5���p�Q1���¯��,�r���Z�b)����L���(,�(*$�i�c�� 8ti�V{�,��E�y�7Ώ�Üj���G�8O�}������{���yU�.��nW�?(@T�B�TD)�@�D Ԋ�N����K�:O�:��0z��?|���ve��ϫ��:t;�C4#� ���J�d�x���Y�[o=)ZQ.��kp�5}��G�n�8��="�&�Jx=�*��t!=?�7y��G7��ٸ���Q���w�����#��L����^���^�W���>�ڨ�����w�-�/��W�#Ӛ	S]^��*�=i�]j�c2[B*tE����ж3�n����C�vͶ�=�ȣ��mb#�D�֏�y��o��Lm��fkf(��"�2sO�oe��f��By��Rk)���X3aڵ�Cٹ�OR���[(��F�߅햆(������#������V6m����8��O������� �����b)�bw��-=�r��8�EK�_���L!C�b%��$B�3�S�����\A��N����w���(x����>Ь=����υ�F�s.��<Ӝ{-)M������5FŮB���'���>�-��9:�*�JZ������9�͞�Y�7��z�G�g��w�8�8�O�{�q�O���J�NL�Pǁ5�5&��ǎ�φJ�[�v��'b��B�6#�A���7|�g�=�p���{:s���T�8����Mꭢ��ܚc3k&LO4� 7�
���Fm�U�(����{˳Co��u�"�hC�{�<��'��*���$ʏR�4�%�@ \H/MM͵�1�����n��IT��e�*h���Sݷ������x���7�|�6�������.��uM�J2,���n�C�����?�W���¥�D�Ku��r�
�C{<�����P��q佃����~'�|O.w}��#
����`A�k�T޽}�b}~�����ĺ]D�X���GO��z׿ن8x0:���9�L/O-ܐ��f�$���y��k�b~]����bX��j�2���d�;p}#s};o�z~��M������7:�<�slj��ۣ\M��F�b�t�K]vW�r�uf׮�ZcO������ɤ��i���3�����[_#W�?ʛr�G+�m�_n���e��N
I,�ܒ?�oR�������Xw<�k�����^i����V���t��\ǣw/�+�]^��4NPp����m�WTۿz��0C�����o���C~����'[��&v}��׿t�˧F��������/�5�ݲ&�?�������_���NnٕR���w/\�y�n�8�/�,����3<8�w^QӅ�c�5��B.v��n�EΧ��[C�@'^���Lм̥�H��rx�`��0���uS��V�I���59y9�k�	üH!($B{�����>�M�R����\@1t�l+�D�k{y#�I(!�\�K!}���κ	�yM��w��}FA�J��·�ؔ�k
�ecc۔����1(F�j������ lme��Zk�V=su���[��5�a�HP�q�����l۳+�W�E*̎ДNI��=a����0�$��#��qbWP�u>D,m�,�t[�+�q�
S�P�f� ��eTRB"�S���y�Q�[	Qk	����G Pp��VA�AǪ~�������xl�0�n����ୖ���!Y�.�Rp�y��!%�3�yt�(�>��͵�� :��!pɩ^���~�ȶH��Zy����K�`Re}���!����[l��ɾw�"����o�!.#��.�A���AAC p�[cd���x��s�`l�c�O��L���!�兗:A6/ӹ�D��8iAo�a;�m"a��kP�����J�P�E�4'�&P��\�AvU�!"�)�-�h��ϵ=4�M&��p��c!M4oё��ށIC��C$�t��~�m�c���T�|�)�M:���0B�RI���$�^-�)e��ѲP���a��pM�?_�-J�u�vDeZKG2 �U��chx:�0@]P�z=����7[�e6T�jGxܠ��A�U:��	�m�xa69Q�a���$�&����Ҷ�4���� �yjزB%��F����t\-��*��C��a�T.��aV�Rg���a8d��tc=1y'k�*L�t��u� 	l����5�ɔ����g8�n���y��u�q��8�l���V�'L >�8D�CO�RśO�qЙ=F�-�٠�g��Z�R�}ph����	�eŬ+=�����>oչ�1H�H؝!8��֙o�1c��B=׆�uO���+���W��@�*���Kڃn��4m��mbD�ho��K�i4���ұ1î~�m���c���^��YG�on&�%	~Bl��.������2�ƨl{=�^E�f�*���y�J��-\�MD6#�����1�>=
��f*p�jj�׾'��{@��(d=�[�e0NLG:���&��Dk�Άc��n�B�d _��lh/:6�c�l;$���"�J�5#ۊ�&%ʦs�9։�ж�[�*=�Ӂ:�8fvS	��\��[ye��UY����U���J]ʆ��Eڸ��uDv7B)e��J�,��+3�jb��`cVk"����f��-;�dǂ	 �O���"K�u�����:�Ni�M"F
f��`h�\�1_m�a�������iTE�`�!J���r6�Mr�LL��v��`��&^�mi���9д[�<�K	Ds����?�)�i�e    IEND�B`�PK   %�X��%� V� /   images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngD�eL\��qw������;�ݵ��݋K��www��Nq�b�nv��Μd29�I���L2��r�H�H�
�Қ�{�^��<��9�]���r�53�g�
�ھ&����$�O[g�����]1			c	S����##��/��!Cj�pNȈ//��#PJ@B�qr�Lp��-~AJ��h��g��ֲ?���+��5���9:d9{��#��.�>j��&`�cbϩvac��]��o>+B�Վ���	C�0�����E0U	��1.*3��u/z�a ���ߪZC��{��c�/�C��/���U����,�x�.4V� �|��a��Hbd�|'G ^��*���w�~~5܏q^�7ޙ��uF���{z��Ls-�7��g�����n�5����M@�����ǥ�b|��N$+�MO�����7�ਓ�Cd�-ϐk&�{������D����AUBC)����7�&D5"��GeG�˖��O��W\�����e������1}���>L�v8G��([�D���(������#O�BZ�C0@��Cd�I�z&�je��q�/>��ە�[1�,��(��dxc���y�*b5{��8�:���)0�zGUj3N���yb��A6}�ϭ��&�Q��XveH����ʈ{��`h�(���c˸����e����Vg�wm�j9�E�����=�o0f��	-� ����~T�"���XӴM8&/��~���X�O��T꽴B��>�����<D�ՇS��K �������M��!x>����2�qb�2�;CD�=F���ڀ��įTr�����*F1�Z���͒f�?q:��kk!E���j#�>�x�Vmջ�f�%e:<PK����5�NsⲂ�Ж�t2�2߂8����D/��+�3��r?yE�� ��B6y�Ő{:߈������ ���X;��D]��\��,B�r�|н+�g�_��$z�'�*D�O]��9���a����83~�C� �j�j�;5���r�a��Ë��E��O�H,�2N��BF�x�B�0_!��_فU��7�����'0P<ɘ��1�J�&�>��A�X0_�9Fb��Z{H��c������a�����D`�i1�\����(������#+f�*L[��f�-��K;Ǘ�)���ys�	F�L��f�.�Hs���������f#"��fc�G���E����Avt_���;(�f�G�j�I7�*�E�՜��M>݀q�f��\8G�h�P2�(�Jr��nB�]ƐL3��Fuj�]�&b������P�t���+��R��Hu�?Q�UT̀6P�7���H�%�n�*�����9a|�%��
�h�WCI�#�5g��&�;R�a�$��*�؀FSSs����l֨�����TRR�]��������S���� d7�BVa�8�/�Q��ࢆ�!n �7rЙ��&��\V:i�E'g��:NΕ9�L��+w�0�j��@]9��|����Ka���A���+�&�P��S�h�3��*c]���ꊯ0�PR�Isר� �w(^u��ׂ�=���G�K*4I�\H�B3�o^r��)䦋	/	�}�/��7P�@�r3$�h�����g�TX��,L�׭.���rf��7@"'qa���-�B*y+�E��Of�Ks{�US9�xzG@2�Κ(<}���b���)��Fv*�^ w�eHyV�7
��)���h������_�cI�L���'8�g��8`k`��O�X��/kA�͌��fT1�o[}z������*�kE�/Z�����W���@�W1t9�5�s>m?~e'�U��n6�C�����I)��xN��1R,��Գp�����7�u᧰�{��y�������e� 'RC��)��F��]�sᄰ�����؜�؂i�Bb��FFѼӛ��厎�2�`T.g(\FR�#?UR�2"0�V,%��^���P�ZňNQ�0�ҿ�5��x�&�Z�1�1�_�N�X޿Q��5��E���f��ce�#�Ki!�~aW�tZ"���"��3���>ڡ�3��{�K�&WϨ��Ց*)�\=�?�;����:�=�� �[����v�
[� ����gfe�N���+q
	G�`�����n��]6�]�hCh�d{k���8Kp&?��m��*P���1�01e����xH��h�]ۤQ�	��x1mjoz�����)����:���W�J0�Z�^��h�ؑ��"�|� ���2xY��n�l>h?���!�d�=���B+l�i=��N�C�&��o��,����38W�-((���/��y�x�FP=�e")1J�~�/��>i�P�9�s9���z|.ypL�@=��܀1���( ���>ӏ*A�5�5�ogrQX/���>ܰl]#�aّ��<���̼DOG/6u���^�濜����̿���u8{�����\�o# 1-Am�',o��Ao�|��ifUX3���t�
󏼔�lL����\5�'dk̫�o���	�H[��btM���u"(���������W����QoF����>�D��GC�MJN��F�ki��+y��k��>@ڇ��~8|�gNʶ�r$�E[Y|d�2�P�2b2��b_��ԓr^8a�M��vchn���8ܼ"�á�_��{p�_\�\mwǻ���uqG�vƦ5j�=u����Wh��/UBL��ocE��N�������H��x�$>��tgñ��*طZ�_g��DA�4���}��t���gG2a|R��?����UB�eb�_�SB�f*�{��]-P�JÈ��e���y�|#]b���j��1F�b�,r��;Y.+ �#Yh����kH���{_:���F���.�"�Ɨ�иfӱ���o���QǑ>�w��bZ}�Kk�T�J2�l-��Y�����Uի�L��w]���s		��}+��ӓ�>��>zv��L9��Ug��V�*B���d	�+�ڂ�� �E��f~A�?�Z��"I���_�[0��GFk.����X��&��R��Ieƭ7�{��lI�F�ǜ�3LM�X�;�)�>���{�V�9ԓC��w�s��,��ڸ�]z�5TiaR�9�*�%�b� y�-��1r3�?�A�!$�jC!�����"�
�����m�ϋ���	��x˫~�5@��W>�P�꤅�Ռ�*�d�eW0Y@����`t��T���/=������|��u)���\��
cl���/�_�C)��y^~I)�:�\��>�f=q!@��O-
��*�/��PZ-�ݢ?T_j`�`�<�u���)�x����r±n��x��t}��{�c8]�9�2 ��c.S�S5 �ĨS�x��,��Q�΄��?���e~g|�<{�9��$4��/!��~�����������,��4��W�vh�hf4�Wb�8EO�1��<�������c�G���CHM%Vgrl�BQ��P��^}��WP�����Ы����`P+��~�r�ŐR
N���2�`]���@��B#O�Ex�*c�vv��#��a����=��/Nu�N|N�}�~^ �ԫ�qp�|�V�,<ĕC"��Y�|Æcv=\!,
�w�e�	n�����-�5B��8����5������C��*�!����ZZ����,����H3!�9X%�w��f<~���U��Ʀ��0h:����y��ף�s�"\2U�]��{zP?��#I*s��L<�̾T.�r�=܅8g3��E�����>�k�x=\v>�B�;S�3����q̵>M�]����X�>>>�#�9��1x��#�m<�!*i�j�/.�D�����B@�%	AM}V����1	vl읾X�E�
^^I3�<t��wN���JgR�1����Kb��0�^�ܠ��(=R�=���M@��wt�r��ʅ�Q;yd#(T&%��/������b�׈si��1495r�����I�_t���)M)O).U�,���k�A�� <�և��^��� ����C��#�L�[��f�+Ð�<��'c�7bڸ�&�^=99�����E���H=O͵�>���e\Q{u��l&f��Zwc0�an�&b�P��U�X.|F�"��'Qb	u�^Ԉ^�'<q������������J�?��ʗ�	�Ȁ��OlP�z��2��_��Iۀv˒��2"\��g��.�	K<KS�_�hG���wn9���y�������B�²�9����-��N��dR֘Mw���JR�`K)����K 1������}���9H�G=3�MzsT�U6S�_�h){�>��l��͋j��{�\Cv+vVA^�+n7���H� �#�t�h�������ŕ�2q�$�P2�h~~�\xZ�����p	��t	�(q��%�&��d�߻�iW�.x���^�<�V��2ֿ�8�`[���mc�3��e�e��o���⹾�#�v��"Nrjj���b��`� �� �q�2�+��F��1NNrk�L^��;v�@l��o�0��~Y�����96�2�B��������ﮬ��/$80r����-P���N0��\�큪���^�bM�T�P�﮻�yv^I���r��%-�}jj����.��`�Gx�@n�aM�зg8'�5����(L���࠸����?<[���
A�GCd���W�?�p7��X��T�`D�~�D5�#*3�������](Ϯ֑c�A6��]Sc�����W�������(Bÿ-ѧ��m55ˠ �<V�\2�^��+�����ڴ� �hZ�%�0�1����o�$=āҾ�yA��>c����K��9��۟q"�:�NZ����< B	�4n���Bػ�^��z?�Voj?K{CnoyU;���}�LJV��卒m�5Ӟ��	�-������J�z�G�,!-�����l�W�(~h��JO̭<�19�S���.Ȯb�6���Ijy��'�
�0�^N�"�䜖�إ)�IL4��`� q�D��[g���1��,���Q��	*�E2����������9�2�V���g�`��nn�c�R9q�ɦL���P��c�R���;RQ3mˆ�.��D��"gKd�F�>}�+��	}q������zf�]���@���GDR�̟}����Nf�,��vl|E�MS��U(��3���}���
�G�����f_�"�ʔ�h��>LM�����#�fNF�Hp_Yu"���<��2��`eU
�`c�&���584�Q<�\��N���heov(jR�L�B��@]�'�<SW#��7,�������n3��sJ5h
G�be6�����O��]�XJM�5j�	�hh��jeU�֫;��*@�9�ޕ@�I�e%̩E���i-U�N��XZ��򔯑��v��S􍄆Нi"Ź�0[q�VԅJ\���:�ߤ��*�PNV+�� �4�K38�!fJ��iI'�$I���D5
x�x��������;��@�ǌJ�N g6�f0UӮ��<�!��O��j)�[M
8yN/�ҋv���Jlm���_�9�� ���lg��A��������#�O�&?�I#Sl�� �.�_/�!l����|�LӴ��6�ֶ�e����^I5/./c=�~qr��(�o/֑�'��ɢ� ����?��h�㬈d�GTǝ�,�������M� ��['=���}p]H<H��'~L�{����U�_M|\����y�����>������L$�Y�����\������6��|���ꦒVi��� Geu���^�����jvmfjwV	���@�s��.y,HbE��[��K5���T�J��c�!�{=�=�G �c������@7��>g`�]�J;f��X��X5u{��Jd��jo�����VJ�!����)����]����G��b����Şq��yx��Ơ<k?�j�e��+���g?�\i>���e�X�m�O��y7��0�"��cFɨ��v^󰦜�r��a.Z�'bUYjSfP���.&�̢̲��r�`�O�Y��d�eY��V)�q�	S��}��Tkf�����wE��k�_�u��Da��=�v���Z��P�k�w��ޣ��nf�^��ز1*�dM��#ʃ�,X����WO�.�O��
�%�'d���kq}��Ԯ�,���kV�\��v��iN�
fE�ld�\0�gY��,JJC�t�U�����P�y�~�m3!�>!�N�j̬d��jH!*J��C$Y�Y�~ւ����=�,(ɡ;j8�z3�T���F�� �����ìKO�-Mb��L����w�+�-��L:�9E<2"賨��"�[���!v��@��,0�;D��d	(�3�qF���k%�7��8Lg���R0�HE���������a&�}66�a� �f��sq%tEϮ~�;�H��$�1��*��%�����i�k[P�� �:�ˢ��	�p�̟�<�]���ћ��F�R�#�,�!4��Ѕg#nکgB�Ǆ�1��6�k��JU��g��+P���6U��`#�& !�,'L���M(�H?�&y�o� �_��S�,�t�#�kJ9Ws�2a2J���ڵ�eE�igC=+`t̃�|���l��P����2��$c�9B������D��� ���j8EʽU�7��G� d�E�Ţ<�5��7��&Sb�^���y��9�V����˽��������Vx�'x�|\�߫h�����0�����෰L���*�?�~s}�}=�哽�|��E|E5�u,s�����-},��������kr�;�vT�h��(!=S-�>0��#�gll�沽�g֨$4B���9p���+�$<�n#��&@b�Cր�7��}nl�i���ML??[�`��5�{>��>�%�P�ƯԬ7/ ��ó��y8�,`�J!�'����lj\�c�����p�z���Kc�ˊ�LU� �S��}�l����9q7Y����I��i~'@�B*it�j�N`jÑ�;�}�7$Pѽۆ7I:���a6�e�g`C���Aqإw�!H���ƺ52~G.L;?�*
�m�v�
�1*�{}������HK¨���D$E��Ϸ�HB��̩IIH��%D��v ��.�iό�1#�9ڍ�)�h�r|�	��6��0��+��|#�o����"��}o�=��j��@Rs�T[Nm!�R(d�Ij3s���7�6أ�ekbB�'�d���pLJ��d���ϳ7���q 2?$��rx�+�f_b�ߔ��)���0c�w�Q�6s8�tOsj�Ec���Li�<9w�yf%���k"�C�[$����-)�rr���|����:��r> �{x�O��L����8�)�=�z4������l���݉�AOҢ��]eM�&ޏm|| �|���r�hj�r�?)0�NOn��G�
2���W�$���G�%Z����>cO�f�{t�.P�­�+����p4Ϙ=�� �ue����Ҍ������|�ɂn0mlO�}
�X�dx�%��9�,� �_ð��f��\R���lKl���dǑ��+n��L��x]�3�A�Jxr����@��BN����@B|wM^D�-����ѥk	JU���ؐ��<�ѳ�&��y�kp*��M�i���tt��T���M.����������i!` N
�tj��NP?ص�{��?/0��0�8�o�]��W˼��������'f":��/Q~u,��u�|"�s��8{��Pm�I2�w,��?��L/�p�����n$((b�]�޿��gLx����~�3y�ܠ?��A'�	'�7;�q9a�C쎉���kaÈW�9���-���z9A9���;�l��_aa�����t�� #p*0QS��*X���Fc� w��CJ&)
]���f�
���W9T���7G�K��7���G�/L�>?lU�|�<Y�[�a/eC�U2Y���D[�+�&t�O�r�/^�:�)��o����_9g��̆b���b�����������l�b�2 |�'����
��F�J�� �=��%3,*�������$��Y|�oҮ�n��[�D }��\��h��yC��և�IF�����{?�**Ȥک�M�o�"^�k8.3Ӗ~���`T��O�u;zGێ���?�0%����a�t��:�̜sp:��O�$��	���j��
��栌�T��3Œ�>�~���W~���n� 0����Z��Q)���ݣ-�rY�ɵfR���=����|��/��~r��<�S1��V`����r�����R@H�����vls<OB��Q�f*:JZ|m_��zo~��I5W�A��1kXm�M��W0m��M��Ps jB1Ϛ����O�Հ]J��_��uuS��)�Q�l)_4���ccj+%"nm��з���D72u�R����tol�RPBty8+�k����ā6�V0H][1�!����M��[�&��OD?o,Ǔ��	���cV���U�t�3㝼��Ҫ豙I'��U�^����6-;�S:�ݴ�n���g�ͽGN�,�C���(��>oUƲ�����eU�/�~8���<l�םVNl8�P�r��v�J�AY9C��NZ�m+�=0u�!�ɕ�zp��!*����mXh�*W{YB�م�k�#�;}�q����t�T�2ad���������'���Aݣ�Ĉ_[��S�y��+����ý�7���I���{Re8�s/�����,kq1�{�GO����pa�Rfq�����K}�^��4�Hu���r�qb	�o��#�c2&�_ç9����.�18���鈌��ʔ�X��0ڳ�u~8���i�5Ҽ�k�It�3¢�M�qJ]R�L�9��P饣������qE�Է��ӫ�q%!{]3[23�FB�F
�;<��	J�@��E�c�)�(�d߀b=�^�"e���QfX��j&���!S��ݾ:�\��|?Q���^�3�UhzIA+��3�1�9t���ϞǛ���p?��o�D�;�:�_	�.��記0���:���aeej���g���&F)���#��A[
J{m�	��]���I�e��b�45%=�|�	�<�?e>>�-	�V>>V%�L�
������9��A��~B�Ɛ�Ϣ]����3X@³�g�M���`#�*|�/[��c��pG��6�ϑQ^��������?h67�	[4M稢M/N��qgϮ$K�h���=�η���\��\���	�v�#|xݚcm�w�P��b�Ȫȃ�zS�3�NW��1�|����b����}�*�u�;����d��3��H�|�SD�j$&ng^t�5V=&Z�����0���1B��*'�S9)��AmF]�k�W0C�x�,�Bb�a	�e��U���F}~4ZFtQ�K�Q�Q���i'��"�T>o�3�m+k�=,UJ[f/Hz���W
��-M�����fA��K�Hiȱ"�i��`�>�qr��X;��Yː9W.�u�mA��7ޜ�%[��ዟ��қ<�/c��?�G�,���^T��&C��g���e��:�ݾu#�����ꅫ<Ui��,��'
�������
�%~��^�qM��v���cj�9lJ��,'t���d�N���U# >΋�p�p]Vk�Т�#;M?�b�OH4:�BM�X�T�\��S�ŞZ�;�51|D�_�L{B�\�tQ�K��������ڱ�K�1��Դ«�[*���e�f�����B_�����&L|�7���@���7`������FiD���~,Sd�L��@
J;�?U�q(w�V�G���q�-c[qlL!�jJ�17�3������019L(�^h@AXq<�%���$8O9�����>��1>����PE�1���	"���>��3��B�r���0*�ə�T3��a��(O
AƆ���Ba)l%�Z�Y���lp![�Y^T���:+Ꙙ��r�l"ٛ��Ԟ�,�uH�,�q��{+�����i�Kd�qBDU��.�k��- �"~�y�5����Sۇ��,]��(�����~H�l�}�M ����fB *6�#1)I�]�n��[��?�{kS�z;,���w����F�����5�ǹ2��\�XE�Z����j^��F�N�6^�d�����"L�r� S~���-F�kj�[��M� !�Ďr���߷�F�9�Q�+��-�hq�Q�u�8^#�zE������Vʜ�}@�cB���Lr���p8��a�(VIhV�#7�z���q���E�ۃ{��,���P���Q�T����K��e�A+��4��y�����B{�,l�S�7�����?ڰJ=��M�C^��f��ԙH���w�z��n�5TҾ���z!1?2N��?4ax�$�ə7`V���҇]��ȍ�8��"57(�%�CT�����L3yka��%�7p/�/JA�X?�}=$���H[y���9ƴbU�ۡ�§�RE,�y/~<���㔜j�����1�
��f%�C��*v�
[�$�j��>N]WGc�{�*���Z��c˕c
�3�K��j͒��=�l���M����x��f=2F�0�$w[<S��$��E�T�(t��X������f�"��a*��x������X���tK$n|�=��@<�.������l���q�|�W�;�)Js��:#ԅ��c��'�|���'&֎ am�-���@N�6s�IN��2�r\�i�T�A�lӜ�~�>U�A��)�����c61S��,��(��h�u�d駂�MY<A��\�9�R�
7s���F��x��M,���2.��Ur��x�.�5���w-3���8�ܿ�E�+$��e��q�c��F���2W�@�۷e��s��/Yq'�x�wq-�1��ҵĖ�����(e�|�έK��{uH��l�|(sQ�������k�΀
ve��=r[c[��A�5��#[]c',ׄ����qg����T)�3�f�t`Ѥ�ɝ����Bب#��zcٚ��дޕ�K"����Xɚ��@'���.��G�����0{DzI�����Q��TF����;��.���H2'~F��Ӷ�O���Ϛ��Hx����b�oOc�/��W����ӄ�fv/���ڨ8�\�X=/3�
ϵ<���&� ތ�:o����:�o6(H��=�(\�e�&��\GEb�Wݬ�ܯEg�+���?�����QP�����@��!��P��M��c��g��e����Q��y�*�
�S2�ր%)tT��ǔ+��J�����+2��4��م�q]X�0Z�ݿ�'�}�	��~��	*�`�x�4��W�o��~��+~�:Je���] ��i�:��*߃�Wܽ��L���1h��:osO�`����ʴ�T��;Qx��(�.d�W������6�P:��eWСν`ҏ�(L���#�8v �ˀ��`���{&�+���Z������ ������׏ذ��аu�R��U}���JD+7+w�@k�U#n�x�A��xL�;F�V�g!a��0��XWۻ۫�� �;}�|�	N��s<\����8�7�@UqP�_��H�]�g%���;^�)�3�����_����=���ٝ��Fh�3���|���2J�{Z��H^��0��^�o���H���S0��L�8����Љ(��ɲ��	���+��m5E!R�(�\�dp��'����t�)�4��H��v����G^{�x�㿭N�'1�i�����E��D��B�X�(�G�s�e��t�ԣ�*Mg$pL���N��۳JC��͛���ᤸ)�L�R	Q)��2��p+�<4{-�S�j�Ɐ2FN���^g��;���b$6�NO'�G�`E���Gth���ac6w�1\�\��5��ZY�S��y���r�o���G��*Ŵ�e��%�9 �W�:x�����vq������m:pwQ�=.�L;5��,��q�&%�?L��W�w<EL���'�$z���
��ԷS���O�S�nC)�:�Q�#mR�P���L�5z��Sn(u���o����5���>���<O���R���L;m�rt!~�c��Ś͏�4�7���S�;F���1f	M^��uw������(K-�������.���,Ew�YWY(�Ǣ�d�	oЃ�
��\%��z{�=^T괃{� �DƬn̪���n�?�ڀ7��c��{��"�p��J���O1Wf 1R8F
�m��9����Wp��\R�uJ����ӣ[�P�soh踠P
2�38ԗ�����(	���{5M�eK�O4�̟ņ���O�Cq�YԴ��SS!O�U)>6��l���O��rϝiR�-2$�*�p串0��a�za��{�wN�q���j�2��<���L�&�}z�`��>�}z>o�N��m?V���8��}?���`a�H�ɸo�|nxEN�������O)ge9)h����Ǽ��)�����͌ZR��g�o���K�k�P;�̸�$Ƅ�U��τ��8P�l�f�;�S�RV���]7��Tl���XZ8 �,}b�|��|��7�~�w����+�n��]���ˍ��W��=�U��Ǩ?$@\a��.��4��`K�Cl#�7a>��mn�<���r�j��A��ck@�������0OR���Y{A�xS3a4֮:,^�?i�3���.S�T��~��S����Z!��mB}lM��F҃���l��$8Pn���2�rQ�)�J:�ȯ�t�K�q�>g��)�)�(�|=7�Y��XExI��s�	C���J:B���a�>1N�P��d���}Q��s�(�i���Xˌ�4#���T�? c=�|��stǬ���}ڏ㮵Ӷ�o��Wɇ��I{�<��X'޽`Tׂ8Xӏ.�~��J]�����e�S��0�ۅZ�����E��w�k���&��m�&g� 6gr �zQ�y�\�L�3�Y� $iMo�,iP���
�������e�DgӨ=IX�8%�5T⢂�gП{�Pr4��T4bd�P-�}�Z_Z!�j��"���s��B���^�>=[�����hY�{f�̈�ĝ��W,�G`�������j�z�� ��=�'�����PR�������Z���S�8㫵;al����%�zJ,O�3v|w���du�M�M		-վF+��|��Av޴
���]��V*)��>n����l�Έ�/z'z_���z��.l��_j�wIp|9�|��B�F/���p�{�[���h�Ϊ�J|�/�� �����[B�Ed(���D��ߝQB��p�]��&�'̲Ѭ��*��C~Ǆzf���4ヱ�&̒z |��G�9�Oj?�^;��e%^�}o�[EE6ޅ��.������4r��h#��f��t~�n�}�|��;�"vq�w&�������ǜ�N�3�V��>�����F�L��<�n�|r.�7
��9^�8�S��^����ґ�O� �4�sO*PZ�2qA�lY~�߉�\���F�j�B�����D�ѷ�H.ʤ2�!��ųI�]/�9J'd�$�Gz�;�K�W$�KIj�ņ]ȝ���/��hH�P��x IF)�~���6~�6B)q�G�<��j����'%a��
͒���^��<�3��9%�]����S����%`�z*��Ӹ|9E�����Bk��YNJr��nu�7����|%~5�<	Nxâ\C� \em�rw&�g\'��$���-_<c�ωuA$���;�KƲ|��n�Jh�5����
��# T�i�#����>��l��/'K"�� �) (+R	5{ -l�#�[���}f�퉊^ <0>^/�[76s1p�=�j�9	)�-7��M*����+���?��-��%6�~E����o�F�}`��H�_�����~��N ���>�'6���itNI�KB6���3�<k>ʖ��/�1��R-ͯ�-���^L�ӎ���v��4����5;x���'FV�t�ySR��!e�"�5%����U�M�r�3��$�g��3Z�p񄿮('4[+����y�%ڞ������fv��_傭X���Ҹ9�Ӛ�����jE��a������8x���B|����n�O�Q���E� m�r��sc25���a� �d�	��@e@�
��D`R֖3�{�F�Q��@��3T��E�r]р2.���$���BX����9�еM��!�/4ƫ��I��#�IG�X�x-��H�0f��_J�K9���L�Fv�	e���#%v�ǹ%�������Sw�r_\z���g�EU"�EJA?�|Nx�s��qq��!m�������ϴ����=W������y�BR��ZG����196+���L�{kR��_��/！ίpW������o��ޏkI8aN$����i�f�#�Cت���𵄣3?�0h�%��Jq����5
]��0@Ɩc��(��}��%"E�o���&ι�D)�m���M��1q�[�A�Sl,��lݡ竵 \�:��p����C;�7�0�3;���F�o\���~I�����q��6�,����$��ٙ����흷���Z��~[gI�=�*fJ��� �"�J ��5a�rU�M>�ϗ�#����Ŕ��`~����og�~j-fg����)Yz��JϢ�2�=%���{�k��$�W:�4�f)V̫k�
1�Z��%ª��,xs�H�o#�qZc�G*#�z�~���*Bf�TZ�:��5����5I6�U�/�|
H�me�9і�G@��N�gџ�|+�7�}�&���C���<Ӿ3��*�yd2���lD8R,=6��Q+EM������q��=��a�b�MƊ��06@.C�o!��t�����N_v���Vs�#Vťw2	z' "�tꥏ}��%]}F� ������#��ڨW �*���
}%h&�JP���s��0I�Vtж��nKDjG�lc���x0麟��:4obd4|�L�;O��QG��*%S'o����Ǜ��e�+R~ ؏�8�=�|��6��5����ڝ��߬J�Q��R�� ['����p����G���E��a놢����Ze����l�~U,�f�3�P�|��3�F&�  ��9<��Oj��W�e?#��Ty�<�	�]���%�y^��pgc�U-LO2,M*�h����\{s���\G�]�����qٖi�����X����{S�"&�^�i�PNsIޛ� ��x^�@��k���[e�g9��I6��N��Wo��3N���_ⶢ��K��`U�$��TV�� �v[8^w�_8���u��F�rَ��~���6e��;,���nv��?��bFF�o���s����!��}��e������D|W�ӥ�m���d�Ad�d�p�L/:P�	I�_���vs>)���j�.�!��OX������,����g�ca|��ct��ac��%�|�K�&G�Wr>ߟ�+���`�8�H����j<�D0�ť��rq�7�O����v��4���(����u���9���ﲁ�~��kA�s�b@)�qE]:`�5��܎,�gDZ}�5����.Ѩm>;��,�G79�Qr6(O�fR��/Rp�_���r
�PC&�r��^P:F&*l��XF6����+�L,8F�G�>�"
SO�gw���7�[��
eFy�<�l^����>�3j(w�Y�x&���X�%���N�r�!!��6�"y̝���zt ���6{u�V���@�)�Y����;�z�b+�w��ͱj1O�ߘ��[�Κ�)5=~%��OJ7c��sE�l�>�j#���\Y��"�F�^K8�z3~S
~fnr�c��V��in��%B����m��{�M��cگ��֫��ߧ��}h��J�VO�!��ۗ��� ��Eְݵ�f9z��V�w7����"v��8V�������Tר�6�ϙ�%3<�>���Z]�O����B�h�_��\єm�.���|��<G��`�2��ő'q�,�d6z������FVo��UXc2���dۣe���IN�LK�V�ʹ�6إ����KU�xA�6J�m�CY&�|x��"������R�4�>4\��ԥ1�]�GVhhAo�Ԙ� �Af�T�6��c<����tU3����g�7��SQ��oF�&����PԵ��l��4���F2^G���g��K�Er�/z�a�u!q�M�"<��z)q}4�ť�Z+��37
qf	}��a��\��c��n��谨^��	�;�fu8��h�b�x�Rc�~��I�I��#�L�VX�g��m�p@����K4�MC��Eb���:�,@ӿ6�u� ���`Z�):������"�H݋���H^ 9q��Q�	&��`�5�bcc�{o�p}~���53�ݫv^�FA�o>���W����y�o)��r ��ǐ�|-�Ģn}�UZ���{xse�Z$'x��x��Zm���Z��	�i�ݳ)�p�����2�;e0V�F��.�d����.
f��㣉e+:Fj,e��eoIҳ�t�������=ɝNNt�N1U'S��9��>p��3<z���?����|�ҭ���}��?����p;�3�q{��"�����ȫ�p�晆F���A��շ���;Xi��w;8:ڋ��D��h_k{)�
��S�17$�1�3b.��r�0~K��J��<��|w�x���k��s��{�Ê�k����d���Jϖ��p�o$�P0�@��M�N��u�i�����%��e�P���JfW q���',�)6��V_�Yƿ��o�fg
��s�:A���*+� i�ű�]q\�JCͦeS�F�&�.��~�+��U�0�§l��%����	s�K�Aڐ�,:�� R$Cʜ��d�a�/�H!�6ġ2?3�R�E�[�?�N� O�^��?�����ߘ_d�1&Ƅe+)7@��ZM��P|w4Jc�͓#l���������_}�oߥO���}|������&��h�^�an��k7�ƭ;����Q�����ӏ����.^�����}���QES��HD}Cʽ�s<\��|��c6�1�L���/}��V�������x�⩈�H-��;2���M�#IQII�(���Y_��DM/��ɝ۷�0=/sh{G@��OޗyN�����7�ǾU�R�#�l��Mq"�9J�q.ݾ�\������4;����������O�;�P}�� ��L�lVAmJѱ��M�UQ�.b��1
)�W��Pc��p��%J�.��mafV@�^!CDF�E�et�뒖����"o{	��rIE��AP])���I�?�@��"�T��8��z���E�.�Y+��f%,SbG+6ݠ#^�D"�k�QmT11?-%v�����Y��&���q�3.�T���6�HS�/��3�	(k���HM��JEk�Y.H &+qcq��X�X����[�Q��|g�����Z��;�0�'��8j�#�?0hy!��x��]|ia��&�O���'x��!�J�f�)�d<�V��Y��;s�R�m��s���[R �'}���Яܑ�eٌ���ʓ7PxE~���� kTi巽�/[}�mnIYgbJ_�Ru����zUz�����V�O?�ç�0�8����x������|��w�x{���&���U��ʗ$=+��Ə |��Vg��������b�����/��`wGr����9j�^U
٨�s�5��7*�WD!)��b2�ڹ;��᱈�nݺ���x���BG���~�����%HF�c.u�b^������Ө�dcoWG|��¥]m.Eg�r7��{U�u�-A�)�D�
�Y�J�%�X#;��]���y�Xlt�[���>�v�1�w����n>�.�x�F�/�gLu-�g.H.�z��@���Ѫ��(T�X�3#��#Q��z،�]�8�B{����� ��Phl�z��M1�e#3�u�(���0��)��^�|�o�ۢe�f�1&��#���kbCQ�*W�B��R�s�
��a�`W@x��������krk�;����P��&*F�~��ﾆ�_�^�vY�����)���q����^��o��V&��9"��I��i9�8($�l{=}���S$A��K����+7o���ma,=����=��e��jbnv�SowDXEG�����4�,õ�=�v���'�$�s���"n^����i)k����ǟ}��}�ؙi��"�T�������"r�(������X������Ա���Wp��u���%b��'���h��4��� ;�ڝ�2�E+ eo�Bp1����iE���ʨ�a��s�ٝ�ݷb�0+=��73>)LA��c	¼�إ7s�E�wLU�X���2.�sG���*�d�9����/Q�")Z��Nҹ�V�./�u�:a�XJ*4r�9Yj%&�'�bn8ϥ.��ĴKa�{���X����,��W�yݯK����J��R�K��2��BO����Y���Q:���+����_�[�m�FA�{��ş<{�_��ޡ�>�KH�R�@h�Qb1�EX�����k��ʊ䋲�1�~~k��j���Q�F��EU�҃�eY���s�w����d�����l�|؅�r#�(a�y�(�/	̉��/��zc����_v���|�5����1,,-�Jz���(�
�5���q��S���Gx��48x�7p��=T�g��Ώ��G[/��;B?*�y������կ!sudai��@c"� |s�&�77������S��D&s�|p�Q�����"���0�i�]�:A��0�v����%gn߹��[74��>��O?�/>�f>�)˖���	��Q\nsǎWe�i�+����M�%">O�^�Ad1�(KC#⡂�*���� ���Q)�O#�F"t2H�1G�41��߸��}�_�\��t4ċ'�� �Za�N��"Q7ǎ`,��p��iI�P)�o��G�p�\)]��z���I��NGup���Y_�n�zP5M��$N�gFãL��)��(da>�����ƥMcbs�..��7���w^����w%��3<|���?�v~'���0GUk�1=>�v�^�.���xnǌH�E>�N��rw�,í[w�ͯ~�����o\���w�}���p0�ݗ�T�V~�/㛯��W�]���?}����\��wn��xCꚛT~e$z,wR��v������&>{�[g=T'�1=�,����n,ߔ���/�����|�����Ot����;�o���5TÊ�27yi�����:���c<�B��OO����5̎�HZa}}M�����H{B������,�Z W��]'�D��C)���x��)�x������������>~����?�Ѡ'�R�����ƨ��+K�R��*���>�'aJ��]E�Ϲ�K�7�'���Z|��wt��YO���F����t�ũ.�0�h��DU�.�K����.M"�n!�.��e�t�*�Q.�_>�B�#_�u���G���a��YJ�ؖ�cnn퉎�_F�q��TE@�u+��c��v�m��T���wc�%�R�{�s:\��>2�,��*��Ca8N�4�JDc�Ǉ���r���^�� ��ߙ��������?�y��&��ȉyʪ���&�6��=���������Ǉx��'8����̔�?�dG'YP�V�fi�A�/��i�ab���v��C6�Nz��
��b�@�>7�	���J[��h4[�+�n����_�\Uc������
)�8=>������_}k�{���#|����/}I@�Uq�;·�]�_{�ճbÀ�	A�Q*"�!u��Ғl�Ψ6�RV�'��	��u�y�c8�X�?�	=�\rzA�f�T�2��� 3�qܽuoܻ�z�"*c{'��@[��e��۷�`��u�[�{x��g�����vѥ��%dk��격�l���w���h��r��[��"�&���*�"���Ar����t���I���9�*ǖbh߉�F9t?�m��\�����rkY������;[�/o��cY�_���s~�s�ꜧ{�gv�R䊂iB�HÐ2$Ң(C@����+ئeS /ŰK���ι����bW�^��8����K�6�U��zu߽���s>'���&��.#zflP$�"��!�6�"�L��u��j�O�Kt&��h:��K�es�Z+�.-	+%I��<��ӧ�Q�͝��M �	���� R�r���E���¹�8s��{��O��l����U��'?Lgk����2��'�	Q2%���_n�Z���2�ss ;���<��s�"|���;s^���{;���WX;�A�Z�S�}!�WO�U�D9�ƣ�����������8���qD�d�r%�A��U9U$D���B�����&�w���t� �;��edd���'�����󧂌9-1�fx`gO����,N�$y�7V�ƽ������m��nbsw��2C�`};��X�i��c�^L�(dt=��BFA��Ē}[�&Q�����k���:59#�H,���[���-��P�dh�	�_��]3!M���m�7�AL]S��ߍ<ኚ�N�t�ku�M#���ʲ�+�aC
�QS�!Q�ϓ��0���lh���#���֎X�6~�JM���][;�7�OS�L���Ҩo�1+���zk�C!s�C���ֶ�w��E���y���8qb�DDA|������җ[$M:��:��Dc�Fԇ�'f��\w����+�0}�e�䒪�侪��W����&�jvwD���Ӊ���y�����Ww�_��k����j7]e��:���khu�s�.7E4���1=8�S���K��I���"�v��79wht��#
�%ȋώ�'a|,�v\�XkT�n��iw����3��o��EN9:5	�_ ,8�A��6X��_���I�t�B:�b��R���w;W�_�#��t��C实XX��'��"��m.�u.�2�[����������fL�*�4�ov�wֻ��<�	_X���R�wo�ŋg
�p�!&B�B��P�d���c(�f���A�`�$pSn5q�����8J�9Ұ��q`;}�;����+�V�bp�A��ӱ;Er�G����Bh�d���R�,x�2�0=���_K�df�y2Y�ƎٰO�3L� '�b��KZe�)]ˮ=:�`$!��\~��E1��������T�����"Ѱ��:�CG2�~켻�%1>:�X$����+j45]7jU�\��͇�����6窀;fD_P��B���qŊA�%a4j	��F���LV����!��N�<��'`��ID"9A���l��ǟ�X��F��� F��Ba��7٣$%c2���[�*��70`d/�Q�юɉi\9}W.��BO����s��m#K�%��M���Ϝ�;'Oc����#᧋pp���A�s�,�F�eցvC�8C�o8�9��͹�G�>NiҶ�h�#�皍���Óh����Wx����Y�#� �Ο8���Y��^��%���'$�$$V�ɖH�\�\�rUu��à�J�8���=,��� ã��#*М�ɂ����M�)�))Y!y�Huۇ��e������/���.���s]W p��r���D�{���ޚ�y��Lk¢D3$i�š�/i]B���? �\6+�U!�G&�F�J�AB�\��0Ƀ�Y_��u����;_Ci�q�=�"��ςd~h��A譜m��ș�e�,k�[3Cuh�T<ɴ�y#�]u�~�L��u�s��ldx}�=��'��8�/��p�AᗫW�����&q������R ̀�r���h�o�C㕴�i2���C��V����V˫+X��p cã2�3�3~����^��w������g~�Qs� �X�(~n��yh9�M5O�����$�F�џ��R�a��sl���C��͉�9N
"n��P��:8����ߓD"���E�[���%x��ۤY��M���M�i����&঱��`H���ju�k����1���o�!���b��ۇ@$��?�cs�H���/>C0���y���#�0��w����ldS(��"�IX&!$���a�}����9�E�^|x�
./,`,�@�p�����z��ƣ	��c~|3��z�����lEӮR����l���#<{�
�٬����D;�C�|p�_`��l{GP=�G��0���`�+���0e�*ʘ+82
I��Ml�Y��40+B�&=�����{�IL��oeKdf�h�l�	��.��q�ǯ��!�=��l�����g�H�>�����`�l;�rP7^��Q�4d�879���1M"�Bmժ���i
#�6궝�ϰ��N;��6*|J�.�~���L������Ôdv��_����~�I^������^�����66���F077���i�xѓA�}?2��_oয়�DIJ|Nȩ`H
�\ȝF<y?'���8b ���-�l���{ldO��Ջ��5�I���74)��M�4~����qe�$��QH�����{x[{k89?��ΟW&Q�.�������C�6�ҕ2�D�B!4�Ad�Մ����I�k�מ��ۚT�~���&��"񇥇���n�,����(I��a��}�u��&����T."�:���m&{�k0�s�͸��P�(b$�xz�
���B^v�l��>���C(���f;��Bٸ�p���O=�ܦ���F�b�\^(`�V�n�T���9��"������i��w�8���KX^^F�莟{Ә^�����[Y��&q�E�"kYzZ��l1����B�,�q>Z�o�WƮي'�&ӷ!h�N3	�D�>�&�k}pp��i�B�:��O�8���7�#�����sq�I�Vʨm	]%:����	8�HH�P���$�	��O�e5��dz���QN��:V�^ck�)b���ȟ��ƌ?��-�����ɻ�k�t#���{��'�%у�Z��y!xஶP�ˠ����8..�cvr�p �\�˯���9r�i��O�bz|B�vn�"��#u0��}�'���с�UC�^�$,Iu�F�e�	$}�A�٩�W3�mf��	��n�����XY]��������S�0����x��)H��o ��U{��t���?��X��g����9�gw�Ƴ�+X�$�",���6Yd ��b��&�^h��� �6�.>�t	�0�L"{��;wo�ٳ������1>0��pjz�������I��b��d�q����=<_]�Q�����}�ҟ*d�ŭ�����J��2��-i��lm,��h�lHÿM���ے�y�s�w��z݀�����z�r̴*I���룍�Q���#�C3iX���wg����ʼֹ�a���0��+��}eVW�����E���SSS�����+��!����4�Ƈuؒ_�]p��Ӫ��'>�o�ږ��N�����|A�Ʊyk5�b߯,�as{G��p�_'���: �.�;�4_�l������=C�*���!��"S�`}k_}���"����h��%�;1:������)�`! "Rn5`�zU��u�{]�����sp�8��Γ���w2i���r}�(>8wg�1C8����{7q���X{�����˗U���gS�<��ӻ���歋Z���l�<6'Z� Z6��8��$z��D-����'q��-��F�E����L��!%���{D�D���ޤ��T>��l�`�pDB�É5����{��Hd
S�؆�f���֚�W,`,��.�h��$w�$��s?;9��xRF���
}���Ѵ�P*DCl�X�Y���U�U��d�U���%ɈiWl�H d�4��y��Ǧ�>_73�9���'?�	n޼�X"�P$"�!:��$�,3����h2H���lk��oMÆt��,����4,5��G	�$_��=��V�nH��U��eul��8>J����X_ٌ�ę3�;�C"U�������U���l~]���J�g$B�5Wc[���g�j�ᇃj_4���=�	@�� �o>���kZG�Y�����=�o�\'���f���/~g9w��͚7G�Ntv��n�զ��M�d
���͟�œs87=�T��c��"�ص��9���̌���LV0;���A�%��MD�:Ъs\��S���6hdnP�V$'Bj�4��v�t�B���1���x��	�8F�Ş��j(�JXz��K	�P�q�"����:�(�g#�rav��B_߿��/�a�pu&��\�G�a��$�D��JeGeh�w��2��A\;y�9�ف>�l���;x��)\~�:װ/$����w0;2�����&%"D�~8|.��up�}�{�    IDAT(ʘ���k�ULLN�l�����1n?��[�+1�جi��̆�Fv1	
|�5�������єOPÇȰ���a��Ci˄���%1�tBS��H#LZq{��2�M��L����m����b$����~��������q��+'�m��&���Q�:���Y8&FF�)�V+��(�e3���D���}6zf�d�I�[��6��\_��bm}�;j����Յ������I ��(Ei��Ζ^�4D��{51u��n���"[�akg_|���,�n�X�V_@��;|f]�*��x�{x$�]�ْ�_*�G�����8�����_WN���.n=}��4��y��l�z�1|��%\���XO/Y��q�ܸ�6��qrfJ����B���<���6e<.�ЩZ��խ-l��b/W@��؈��N�>���q��,�,���GX|��}�$��&�QJ���E�ɏ�j�Fn��P ��"WW��qx���2���u-��������F���+��h!�W������u�=Ṣ尡Ԭ�P�
�f�8�cJ�(�@�P��ξ��'��Hz�v��6:l�>��Ľ59���DdDRe�8:��ޮ\�(��j�
�T*��C��v�
K&����#|��������3��(�F:�%I��_K,s3�����-�٘b߆����W��V�v���X��7֘&J(�����Y�0�~�3��*	���k�C}r8;J��!I��gV@�S�U;��NN��:��^������g��ܔ̍מ�M�\���-�$�+���������
V77�p�0:2������w��s.���(������;�����7ocG T��Fz��Pi��B#S@�P�ɉq|p��?��|�/��au�%��>JI�l�	Ny��p� �r��Z���D���H�#���h��M��:��n7�s�o0r	����	C�:����r�;�XZYų�/�G��A,���p��5u���O���a�3p�K�'����N�{�ȕr����ѯ��e�첣D�:3�U���ՀqHP1����lq��<��Ϟ��� R{[�{��>{"ؐ���7�]��3�G��Jl.�'H&���<���n{âps��&��14:�p$����<����a�\@�ӐIm
��ܖ���ʌ{sɦS:�nG�0�j�	_Qr��I:E�=�-�=mHF�.�F�I�v��0%YѦY�����F�;�FKE���$~��{2�	���g�H��$"�I�x?���A��LI��ɂ�!�ߏ��AL�%�pr/K�C3Mt�<R������X����s ��0N������HA�x�xB�C�3I^����{�jU����t����`o���y �b��2v�v�駟jj�K8=��7��gWr�c���#�bp`;[x���RAQ��BV����Q\?w������	y������%�ڐHW��.^���Y����u�n��
�k/prv�/��﹓T]���4LIht�Q�T�cWc�x��v��v�%19=��/bzv.�/V����GXz�LM��P��$���196#��p�/��O��u��\�� �"�v��~!"s����B6����Yl4c`�S,�X0�=8In��yҔC$<�M�q7u�k�B<>��Ԡ&���d���/-8W!|_�7�i��u��,2$���Y�K��Ѓ 
h�LBٳϱwt�ׯg��B��X,iB2><��x_P��'?�_}�b�p47�]3���DM����Q�f��G���5���o,)�9�=Z�5%[EX�im�ߵ�0�iC�f�y(E)eȔ���eQl�������~I%�T�~�ѝ����P��!G�����sC��J�"�bq�	^�|!�U���"�e��jM�	ዄ��olmaswG����؏G���/��s�����G�Ϟ?�'/�F�w�?��X Z0m�F���(!���kWqfa�\Nę�WK8::���R�G�u=K53g$���[�$���� �b���岌�q4��4��c�pfWLU9;�bg�f�6�+2��S�������\��&���M����M�x�.�������s��$�M������^�r��˶z�ʶ�v柒hd�o2���fː�0d[Y�v�!��U�����S���s�����ܻ�i�ߛ�� a�J'��0?>%�jfQo��i:�5�P���:���R��R�NΟ���(��R�n=���O�a��U^+�Q��b�!��6��5=8ڷ���,dS�[���V�,��?�C2;P�l�?o��v�F���%k2�ŀ���`,��!f&����D)և�cS���?�X$
w����Ed�S(V�Fl^���b�����%��u�X�����F���-nw�h7ʰs�ީˍL��lN�~�ƥ�[mJ%2�*�$f9�>ll����k������%���4]�ϟ��sg�JF$�dF����0�"��4����d�����O�Sk�Fc�&�9sJ����Ɔ�}o��GK+˸}��`�|��\���kbl�.���>����Ζ��$f�k�\v%����х+�0;��d�v�������`kw'f���3��w�]Ly�q�����q�S|�g�˸�dK[ȔF{p��i\��N�>-r%u�O�<�J��9����L���v�܋�I��S�t��6p\(��M��b����*�Ʀ�R�X[��������z�1D�>%Gѿ��?�=j�L�����u�<{�3�k����c ֣�.'a6{t�Q��$5�d8g����T����Tc�{��)Mx�a��<�e�C=k�Pv�Kś�!��C}CH��j�y_��/p��MaN�(� CC�OR���{{�U^���5Q,Cl�U~�`}����l��_U�ߞ�%%2�_�Φ�4�&�_&���Y���p1�O��'���O�ŷP�%��rjV�ŢS�9�s�����ava^H��۷��|Qk*!ᰮ5�
>�ܭ��H�?��
H�N	(���������Ͻ��_�n�/�����o4��,HJi���0�@��U�p��2��~������
�^.-by�!t�?���1|67
ق.2!5��z35�<n���'��&\�v�U˩�y�F j�� �ł�>��F��R��r�%;�T:�6�Ǒ8�C���L��X^]!��AxL
.�[�ھD��877��7�l%����s<�X����Ƞy�������e������I{�B�f�9�/���-��Í۷���C#0�p��[����	�ZTR�CG'�ب��DPnV��z+�;8�eQ��EV;s�;��������-ls��9�$�Jt{�n�.4���/�/����[�HN�v�|���7�td����<_��X�,o���ьx�K�a32������U;��F�}�09��~�=�&zhv������!2�,r�V�@�і�s�oP��I
��k6>6���D"Y�v[�kEc�kմv����@�Nc����Q������˕�7��-m��?�'�����ށ�#|B]����-@�Z�6>0���1�\�"����v�j�o���/������wo�������!�Fs%
������/�D��@�^G�P�nkhh����+V�N�?��s<_]Vf����~����b8W�ݻ�q��g079��'ψ��~�!~ 3�:��<������e<^z���jp�}"^�zUr)�)��/���x���"� ���0���a$�I��)��#�<W)�ZU�������+�tOr �O���Șo�jU���{��\�:=FOx&�X���|�7���N��k,�ϟ� ��A<;1������f���D ��{��'�l3i�$ucq�s2<8���ii�I����v��d�H6/wڌ��Y$b�ߏf<sj��͗����ۚ�XP�AŌ"e<^/k����5��_��T3X�[F�%Q����͎����{b�����l}=��K,q:����kptt�t6���u���z��Y���Þy�햌6����(�%� ��H$O�(���!l�7qm�5 ���������!�+y���~�C�E�$N����P��߿����G�G�n,��J.�[���/�"�8�f~�#�>����@_ ��x"La(�@&s��Ϟb��K�xvs�k�:r��n�T�BA�4|��z����r��$�C����QP�����0�/N�v7j�2ԡ�/-ߺ��+�]؝�g�4H L!�Ӈx$�K7�j���1��)q{�z�C=I������9D\>���7_ai{��c�m]T�v4��*"�H2AMRc;�M:��3m�+�7��kW��$<�ߧ"������Lĥ�k;TxǓ�ҟ���y��Ʃ��J��"�}0}��mH6q��Ua®��Cܸ{�<���j5�K]n��ňr��ED�R��`��q��p�Q�����wr�1��9�')����T+
MWѴ�>�)9VV4�K)�"��$[PZTi�}ft�|�L�{G���p�>�� ]����6�嚈V�N�VՃ�&����FF��ᠳQ��lE�8(��nWQ�=&_���嶡�"��*�8<~ll�J��i8�#���(�Սu�ri�)�	�&��̟w��3��*�n�"�FkF��R^r���/�w��6}���J�N.�Pq���C�r�K��/WW���&�������v�2.���߇T!����%��z���`8*�h�^�>=1��c�����je��bztT?=8���`x���� �G��٨�:x���ŕel�����H�Եk�p��E��o�ʺ�E8_������<��&�z	D���e�)�'"�
B?.�4	S�OM�Q&#k��g�bfrJ|��i=x��mBg���W$�WK��i��D�
���bT�X_�a>/�jafN�������
���G��e3r��^�֢����zi��F_O�ٴ)	Z6f�Y)8�Pq�%�J��*Y�$��P����/dB��b	�!UPo����)c�M��i3؆g��"jL��N���oEZ�ۅ�"|��!�$.��e�dV�`3e��<[Ԉ��*��oM�d~����%
�4&}ZhR2��a��&�+i�M)[���ZU�ao:&�8�#�
�*���+^��di�����.�����ɑ��<�?�������?\�����wVs��>hԂ��y��;b��^�"��@0��Ӄ��^���	������G�AH��D��q*�|� Ȁ</r�N�_#K��5,�h��B�a��N(͌Φ�>C��B��.ػ��j����:#.���e�`����y}��$z����P�Ţ"|��y������4���!L��|�ݾ���]��(2���5�dS�jNu**�y��c�(S3�.�����û��`$��7��!���"Ls���a�Ē8<���z�än�Q����,����:v��||�LN�#��`?��� ��ZI���ܝU	]Ɋ���dx�&Z3���.>�7���a$��{��Ƈ��?o��(43���X�t������Z#��)�~���j=� z�𽹓�k�g�Y��R�zIh��ڶ&t�����va�O;���!�%�#���<N���֑F�eX����@���_zw���wn���+&�;wp|Rnd+���T�!9D8���gu�q��%132��!��mM����BN���Ѿ�:$g�SGr�����DB�n�L6�o�0��,�/����E_��N���2}~�&�6V���l\6_$O^�]�I"
���ʟ<{��O�a�� cC�<����1$i+��XIb��I���6�����t�%�R���8��=�<N�8%�eusU:�G���=<w�,�G5;��È���Cއ�L�븘A�ZUZ���M짏�&q��E��=!|�Z*h5�� ��#Rb]^xY���њ�l]i��ż&�ͣ}s��j���<�&�U������sMY�^���=��t*�f�&��Y,,����FzdT�a&s��g�/�noc-S���d�H�-�r�χ�ׇF��b�(8<O��c�5��V�4r�����2eYK�,ãڒ'};�ϷIjշ��*�oO�1�*�Մl�߆��asʳ@pt./v4w�2	Qf���MDѤ�P���v�iD�f��i�A���#^F��!��P��z8!�C~��kM��Z�����WR2��k�zݲÁ�h3c�"��ϛ���������/����F5 BZ�+�"d��}��� �_�?��9 �N�ѽ�x����u@�͒�_S����A����1�RBH��6����J�4���{�<Fi��$v�>tG!w�Z�Z�jS�,u�1v��BpҎ�{z���1nt�r�Ih�T�E��|dbJ���7�\��?���2�HUJ�;-yG)W��C��nC;L���-Fk"�m�ۇ�����K����=>7���{�%��C��Ņ�S�!{/j�^(Y
@0�G�)-̎m7�����`��+4;N������?�����G�#�yx7Ʉ����>�?�ǩƄ����"QV�}�?���ɜ7!�4$�����݀��+v"&O������:kN�
<��c8�ڰS%�U�Bf��Ű$��O���D���l��O�c2E.T�9lnn`ms���ꠏ���K�{bG�*ƲQ�I�#C裵�����#H�$nd��t���Λ�o��p'�j�Q�6��t͚ҥ2�������� �}�jA��Ӆ�^6���zg&5����b89:���!�N����D�Mds9��~���-1g3�c��xo���B�d���N��BN�`w8G8�@"
_8�h"��d?�N��i���~�[G�ȓ��v���~���IYV�Gb��0f�������踈Y�Q<*_hR6��(&Z�<��*<Y~���{�����$1�7���q�G�++�߻wG׊�߅�Y��z�IEGf%�C
|�m��V[�dJ��޻$����*�g�N�MM�"�mȡ�$��X��	*��@.�����)}�a6-��y�i�[���C ��mKĂ�^����%٩҅�rBJ_tޑ?�A�c��,�bE���ǵ�0Y�<W���������mvD�I$�o(+����8��7��;Ϻ�I>��H���?[8��מ�N5��lM�yGlM��d����ǀ�͆̈́�y]eHM:�:3������m�χP$�t*��,�m�6�V�1o�	���!�V&(��X��A�?��9��'O5lp�~���1��<� ���S�f����X����=�ǏoU��?���?z�<;�����R�h�hb"�����IH� lscvp�p~n��
��ܺ�;�n�L�?94��gW�&{��5PoT��Ã�7�bn���ؼ��v>�V��3!R�y�-�N�z�AJ�BL�͗H$�`JJ0.Ȑ�Y`.�$/�7�VN��!�bzxc�/��,���}�3(4��,3��i>M�2ʙ��_�<b�*��{D�����xC��� �g��K&��n|�"L���y�V�����1�?*������Y㱳~��7�<«�רԻG�x��u�N� ���p���`3�C�e�m>�.��}�B��N�g�P�M�i�A(�+�n�G�)��oMhe��P��a�A��Ņ��܍����%��yO�}%�$H�}�K�eآ&�p}jc��v'��^�����g�8�F6_����P ,΁�h՚�u}4A	e��K!���|p�lm�ݔ��)��q`�O;�9�3��v�X�
aa�{�і�\�\�Z�9L$��E����F� !0:W�G� �J]V��6g�,�m�ۘ+݅H�r�K��>ؓN�Z,I'�{L��<d;]�P�E�{��]<���x�h�X5���.��>��|��SGx����Ҕ��4ߎ�׏���0:�~A�]��K�/�ʧ�1��w�P".���=�&�MN�V/L;��dK8��d��8��Fџ액NN�˯����C=�JI��p��$J�`L�J�(Ґ^?=߹.a�J{L�)R]�$L���N�]��9�PY��X�w    IDATe
�ˮ�+�D$
'�T���S�Tnl�^�T>�Uw���BVN��a~n (@׿�dGg�x��9�,>U3�g��ף��Z����ƁȊr�U�:�Jq�i��95��~a1aa�Z�k6�|�����W��9ck��oC<�T��*��8M[�Ħg;ˍ`,sj4s�TK�dA��$lV6y�LH��/[{�ad�s�.�\�X�˿�v��:�|Ǚ,�3]�-��9�}m$`��pre����F��+D<�X��qa1�$��Ŝ�R���g���,L/jE<Bp����݈���SM�J�͐��s��i�w�\��|S�~�۵W���������[-�m��Y���6��Lm���0�^Gb=��k873��d�l
����[7�ɥ��ux=�Vjڏ�qI'a���c�\��EǢ`���`'��V��q��fsz̬Hڳ�M�+��d>�n0��A?��z�t����FW��|$�����%�L��/����3)�ɝx���\���ǅ��pH����@�TA�����n$�e��PwH�Oǁ�'������S3�	zQ.�����D�	�H� �ϝ.�U�+�֦��s��7"�u��,����}d�U�f޻�Μ:���^T�e�����/�z�B���v5d�6y�9�	�X��d`�]���e2m���uho�C�74;GP�����4&֒��&Ꭾ	2*�V4�v��@�&P�#�`:փ�S'0� �t���)��ы'���\���T(j����!D�^E9_�^3�rc(�@2B�D$���lʫvR7ܨ
�Q��I6S�If�����P,W���\��Ad��s�N7��(�i�>�h��)������X;�:���LLa�!��n�����|���}�JIP1�D��Pw�!�]��g>Z�0��B�\B�������%�?�}Úy����.��2�*�ӂ���I|��u���J@	���Wx��6������c��xA�q�ȵ���>Q����6vw��I	��?u�N�Rq%q)�e�aoO�>��7�֎��"���ф�0�I��T��Kb�渎�M�P%7�s�SE�Ĭ�'Y�m������C�d9J�_��o0ɤ%��QJĴ�G�qI��fu���nY�Z-�?}gO���̂(n޽��o��Q>k�k�vI�t��0u�JW##������LS�}�3�{}�O<O*�l)�E�E�5��X�*ƙٛ��NXh�`d���0�6�L��T�kHy�}%Y��S�M=���aak�U��[;e� [�^����<�-��۟k��2@30��H�&&���L���l��߇hB����h/٬��s�FM�`A�����k*.H��s���'-b�d+V�|���ѾZ�R���c]�.?�G&~836�?~����C��"|��;������;��[.����CW�6�u�ޢ��HQ�����Q9֓D�Z���.��7�h�7���|������M眢�Uu��{+�o:H��Z�N�<d\r�2v�
wr����ś��D�n�D�X0,GBq:�Db���4��)��)á�:���nv�ÒӕK����/?�����j�x��z<����5�����ر�	Ӂ�%N�v橺���_�.�͡/�G9��N���(V+�$��ŉ�)�Ebހ�	��ʭ�ih�$L����k,2���(�
\n?>��Ν;���A��e�}|�ݹ�M��v����:�	���F����7�d<n�DMX�q�{q��
��e��4����O�I�>����u�V�P��3�j��f��,��dJ�,� �ͮv��'gD���9L��;�ȧS��_n� S)
�b�r�RG�f����͉�S���,�Q�7��2���0hA]71����Y��XX����(r*�J�:�����x����N�#��"����M� I4�y��EL�K���4&��亡CIDCƑΥ���c�p|��!¸:���V�(�#W=t�b�@�~>�	��`���3�|�
X:{���l`��I��ך�����)}(F��
^�z��+�d��K�c���pX��M"Bʀ5���:�QY6�$7ɺ�V��)�ӂţ��2�Y�X�5���_���f��A��'g1�7�kC���t;���m%��GOa�ze�P�U�/_��+�/��1f������v�l��L�x0�����`93JqhlT|50U-G�ITtq��y\8{ss�ܾs_޾�c|p�ⲩi���\�q*��S-,��΋�d q�ǐ��㺡]k�[vl�0�&�4%�x�����+�H��>����|��I`!!���lk0����)O;k�8���Gk�k�n���'�tɲ
.?�ϟVV�C�q&�ķ����l�m���V�ъtd���h��DX�G��YR��A67&���F�afq�5�>�ү3�Fk63��e�[,��\�L�^7��Qv��afd�?Ώ���`����w*¿�����^<����Rq.�� -�ݍF�-�W�������&��1�����&w�6�6k��?7{s��7>�܋��")X&C׃�4�խ�4�1庲�Z�c�{�3�~�E��6_0("�f��Y����t��ɋ:d��|�L��_����>�S<�XA�\B�;��XDi4�G6���x��
�G#����R��������~�+'N�/@!��g_}�[woiZ
z���%㜓���#��&7�	��8p��{|����39�J����裏ELB�^T���=l��ȵڡ�����qN���PTr�r��L�]�<E�^��E�xD�""�Y�#舐������v�FJY�41���!���f��|P�~v��azZ�����PW�f0��G��B�� �+�9�C�rtQ�]~9W�m%��*M3�94K%�I�k����m6���-���>\MJ4��Å�
��ˍV݆��kMEr��q�inS��/Cbp�^���`�-#�P>��L�b��$���c�o ~�!̗��a�e��,�������0��F�Eu��3��Ǝ�lF]��NE�-��`7�B�Y��=�i3�`��y>��r�^-ac+;�88N	a�5�'W?�j�Ұv���W�X]_ū�5I�Bv7����"���-�kj8H�a��4��6ﴔ�M�ǁ�a��.`jh����Ą2����cܼ{K�n�dG_�|M+N� ��>�.�K����|��Y�5�uDc=�����{�pU�g��z����O�N��N���+W�U/WQ-��(����V�^.��ƪ<����!���K�t�"�g�Q����R����z�[�
��1:9S�B��55R�$�rFo���,��l���Pn05��kp&&��"��Qa�M[+�x(��#
i��t���UEWiA��3`V~}+܁EXE���ZE���ZRC����M�o�`��͝�_G�=[��E����a�p�"��a���H٦/���A��"��D�:�ﳽ�Z�.K]�V&드 N���e�b�7���&ǅ���X�;�;L�,�e��0=8��������w��NE����_�ꓽ���.�N��**9%$���p����۰!�������	���5Az���4&3��T˿����C�_��{���MKH�Lh�oՍ9�p+�Q������o*�ӄC<^�������`W��Z�1#VōՄ])_`n�!�0� ����m���<{��t�m�^��IL��`btD;�j���lI:e�a���bm�3����ۿ�Kx��	�C�e�d���Ay�W�:v�I��:fd^��)aw�1!��˻���XB�c�/�'}�KW.�-&SʘfT���&�$�uZ�:3��N]�f�r2���]�w�����i��D�7!M*={	�ӭ��J���T�aa�zyĚ1�
I�d�Hq2<c	��U����AN���Cb�Ë�P�&�1��C��B��˯���>D���k����c�J%6l$2�)��
y4+e�p��%*Y��g^��%�9A�K[��H�ǖ�jN4���U#�����
L����� ڛD05���\�pG�\BYx��E�855+�O��K�ｉ 8l�U�X\z��8�t��By|z6Ԕ�e40�G��C�HĦ�Sa����������q|��{*�4�aC����r�
���g��<���1����v��$�{k�.�B4��KUI�����h$��*udD�lZv;�ՊtԴ�É�i���}&˝���ܾ�#�7�
��N��KWpn��
S(��
�|�k���.>��s�G�j��~|��G����ܹ\F�)?�����Z�eO/Ν:�3'O)�JhI����a��M��q��?y�LnYl�������2��ܼ<��?z���
}`��Uj�B�U��|mCҧ_���4Hh3&`��l�9����څ� S��p)�2�����O,�$�Y)b�|y��H��a��\j�=ɲ[P����5�J^h��&^Yd0�g{��ec�w뾵��U�4	�jMB���1y=���EC�R��5�0�y&�ĈB4v�W�|ތ���]�{�Bx�q�5�ҁj#����gW �����Y����Z` ���_F'~��h4��Ѡ|��{�������m�Ŏ��ڎfӰsw]Jb<_����.���8=9W���dy���҅��h�@�Y�˔ŏR��H��~���iɚ��b%,��];�t�}�:3ʝj4:7e1̓�r�Q 4�lxCқ�؃�#�J�5&г���X7��:�����?���{�6�8,�Q�^7Qv/j>�|N��X��?vy�"���EM�	�D�*}�)��sS0(%!��K�����a�|MCk ퟩ�#$���b+��A��|��P����\d;������8(�P��<J[Gp4�FX��0��Q�Ԓ���  �X�Vw�P����O�5����4 "�UH<�t�l`�0pU��c��Ώ�3�%�c�J["�R�i�я���T�H�|'q}��⽈�](��jm[rc3�ßMC�Bc|C��b��
=��T�Y�\v�aȤf����v�|n��i��F����>��:�tt$i���
�$�!�"�ܑ��M"��q�ݔ4�³�pz�i990������5��2�GGm$ݭ��@*���;r�fZx�X(��ĹPDE��� �f���ua��=�C���%ˡjucU��ԁ�����P,�c G�pe����]��m#ߪ(��Nf>���k,<��&#��\Q���H��{U�v�$����yL����p���`i�9��u��7u��N�����NϞ�=�:>���jT�Kv���%ܸsW�*0X,9	S��޵w�[�g�"�}�ӿ�ͧҪ<nɌ�7fx� �f[H�������6��VT�	��U='�.]����%U�A�����s��a�ATK� s2�	Ul4I65�s$��Ź��-w��/�{��IH���H ,8����%����Ȃ��x̵#������v��#����XE���3R�E�Z���#�v���lM�V���1���p��;��h6�f)S�Ôܩ8鲉��c�o8�ڠ8(�ɽL�2�+��|���LT""��|��aq��)�%4���*s���w6������z`hP��,ĩ�c����(׻�c�?:���������;ۿ�:��j�f�;TF��G�뀫�F����Sg�хK�8=!���S��rV���F[!�,�
q�/�
ܑ4�&����إ���b p"Q!6S8X�Œ3�3��Go�A`W�}a!������WU�s)��3"rm�Y�)��Cwpt���!S�i�\���q�,-f�٢$��m��b@����jf�%i�L��6�9�$|ea^E�\���/���|-b��X�0���u���K�&�xvd��u����vSY�+-�z�����ŋ�10<���~z��xtG܏:�:eX��$J<|mH�6�_��_KP''B\�ܻ��F]�C�,�<p�X�0���U�n\=���p�%��d6�?��k��_5X�>��\�Ȋ�5��1N���<&"I$�^�JE��-�5���`O����[�jؘ�C��;���1rGG����H{1�����E���aA���;J�IA31��a���a$��M��K:�L��IȺ7���>ɱx�0�!J��k�u�m��o��L)��K�G��l���>lPy��ǚ~���R����d2"+ٺ��&z1�;�O��@�?�a��
�Sک�>'s����Ѥ��4m!\����M�|v5�$.Ҥ�h��M3�d���q>W4�B^�" �ɯ����t5�3�3Ss�E�A��vv��=}��ɃM�S8�,�G&՜�����ޤ
&�S�<Ք�_<�����^���r1�Q����s�@/�#�^�,қ��f1|������%�}�H�q�#<SX��\���s:;��x�;�i�R_�4�T�'�KX��u�H�H@b�<Y�x�$T�2��|]\V(��Y7��}AT�5A4�%%�"�,��b%!}[�y�򹳊0��6S���`r8��(
b!��IR��"l�����k�'n��ZßM�-��3�����bN��J;b̽�x?"R��x��5�	5�n�Q���dR�H��x�2zac���q��.�u�s��ZC2?��h".N8&<q�Qȕ��􇃉�?|wd�[k��0�~�I�'�����[�|#w�n�Ӓ3TU:1c����~�D:N��p
�=��'O;]��V�>!�z��5�+P�VC�)���E�4Ӡ����C�alH��^4ª���Bl	��}o��J"����euy�E%[!{TZ���I����C���E�׋��1���
U���<X\_������J��kgG�)�{(2u9��X\�t��GV���pin�QƮ���W?ŗ7��*IXAB�}�����t&ep�>̈́j���n�erX�����]�����ǿ�ӧ΢o�{�����U��K�]v�����d!e��:`�S�3L�a�*�"�l0n<���;(v�.�Sz]�X�Z.��`:oq�ַ�0��$A��<GSJj(	!���7��֛m��-��q\[�T�I�UK�K`?�B�UW:���LCm��c��ݝj���Fl`�����
�R�J��&7vϼ�x�1Ӕ.qDX��jZ�Os"M(���Ԝ����G��ӭ�W�D� ��<x�hL)��zY;,�i�%�l�b}�.Pi9o��P;��e5q��CT��U��˘����ب]t��tJ����T�����`��s�����u�=��3ҁ�7�#�涺���[X�]G���z	�6�-Ʉܡ�n�����C!eLy����*ַ�`102��!��OM�`~t!;�J�8:>ĽG�p����i����?�~��pB�U�YA.��K� ��/����?�'@3�t��P�����<���Y�n}�
�>l��)����+X��Wc�=2ܚhKJ�BN�7���7�d�j��W�j/|jnA���Ǹu�.^������i�^��k�����#�����|ٍ�-Y�
����-�6��:Di�"�~��N5W�=��6�N�;bL��$�{�g%�o��b��$Zu��i2��-����A?�A����-k�2c\��.���F(���%��v�a�	S���HY$U�vt,�cG!�.8�ߢ��~Š�th`@M����.qL�$��V_ڽk�wkh�3ĉ�X���� s����r(U���w#��ui��N�_���|�to���gS�st���?m�Ȥ��%U"�o��8���	|x�<�=u
�j	�r�J^)Itw"���"lZJ�Fv'�$a�h��W%R��&���Mk˺�Ī־����n��@�!��t��%]���1�-��V�����PO�)�Suj��&#�D���Y9���9l�-Қp�W_���
��4��� u�M�I�G)! o���FWy�����f��Q-೯�/���|���8]�alY�(�JSx��Y�]+�/�4�r�"�rkÓ��G�����	o�ᳯ�"�[ʣ�.���[���CKRd�F�,��w�)��pic��<��yݜ$gթۣe%��1��Xl�h�9Y�4�l�_���Jx�p:�.��]x�%"ְ7��͟�
�*o    IDATL�_�'�f�jU2�6���`��$c�a��E�R#W@�({��b!�)���+���#�L	3t�����t�+�;i9I>#[��T�!���HD?�$&tgl5� �5��t����&E�"feCE�ו��ˍe�ln�(��M%s�iSɤ$��e��UQ�}YF8cҊ��&�*�I �ۏx(��� >~�}�d����ʨP�S��	�#�	��c:�֗�����\�O���x�i�5���K%d�%���q��3X�Tɸ��.�"#6��J`a|
'ǧp��9<���W���=5N^{_E�7��r�cL`ux�������cx#A�1�n���㓏>VLa.����
>��΀׏��5LOL���8���3�^��|���y�fÝ��q��#5*�rA����%���I��ݻ�bͤ5�.�&*��Z���0�@�O]A_���"��\�/y6Rnǟ��l^��ݨ�p���r�d@��Ģ��������Lm�i����pb�&׷W'��^���J��CW6���]��o���?��|+�ؘ����=_��������5X� q��c��谆�x"&��b�w�Np�ͦ�h���^C����gQ���F"2Ҹ�^�70��&#�.��2�ޱ�ٳݑ����!�����"���~#s�;~|�I���ዝ���9�^����E���eC�ޅ�넳֖����i|r�.,��V-���+��m*�ّ6��J��Z��cq���I��)�R�اƔ��;�F��ZS�6�ʕ\��0F�E��{�H�$Q�W(Q���UB>���,�ˬ��l!�(8p�~�����PmTD��!��q�h�v��|�j����vUx���g��]M'�o���I���;�MeUe�,�}w��ތ0 �K͒�\,�%�����}�.A�+�(B/z�YJ A� ��i�m��.o�\Vf���s~y{��^�0lDǠ��dݼ��}���i�W�w>�'��FgS=2�8�ݾ���/akkCl��C��in��%�Ѯ��$�G3Y�<�����Y�@4K���}#�=<�"��ނ��Y�u\�wk�$�t��^Q�p�^%�2%`.��/����fu�l`dʝ\<���)�#?��0��q$JX_G�*�\�02Ȃk�\ZS �,*V�����5t:#�3���Q��F����5AIɸ'罐,g�y�ǆ�M��$�<��_F2��B*��;�;"��@�`�w@>�DL���-���Zu8q��R$g�X��C�6P���:�y�4m�r���5� ��fe����bU^/vb	wv�uM���c�4��}���y�E#B#<Լ��
���6Ԉ�P�� tOc�}�뽴���%�l��.:kB���Y8)Qډ*'�Q}��+��F����&�6f�N�ɳ'X�XB}sBM-���ҽ����ڊ�Y �U~xh�C�i��ױ������S���`���{�w�V��"g������[k�8�� �ޏj��a��1����@_�����,�<}��/_���b)��s���O?����w�фɿ�rY��T"F�1&���ǘ���z�t�A��r� ~���h6����3���n����Ҍx�Y�?�65<�/�)p~��)˫�tG�k�k+~��7���no��O��<2�<d�Ƥ&	��#�����IU��j��L�Gb'�?Wc�c�Ĭ�������LϦК�p��cl�I\i*x���P��f�i`�wV����oѬ�$�Y������'��\Y	K���,-x�H��#@Cc�d���W&��;�2��Z��ZW������O���j��2��
	��.S2��"�#.1�nq;�4�W��o��s==߾N��U���b&>�,��DYĻ��_��HC[��_<|Gv�������x���槐/�e�(�V������� v�q��T@%/��&2���0��J�!��=����.C�1M�5�Z�BWO'����&�5sy�-1�N?�\����v�y�qh���+�]�'\D(X�d*��3S�g�H�XO�0��JlKE�@;~,��s��괹PH����}�!��Ewk3��$�޺��/)�	'JiF:{�V]�I��d�V2R%c�FI���*��$��A�k������������$|��m|y�:V�	�]� |�]7w���Я��T�������V�$��u�(��� u�pE꠆�PN�K[F��g��gқZPw�$��d���,Iif`S$��r�j����݇p�w�M�
�s) ���"rB3J�hd��p���T@�1�y��w��3s���)�S̢`sʤ!PU�F�R;>��B��$#���^�K�����9ְ!��mmi��يBlx��S��,R\����������m�[*�'��0^��ֺѾ�H&I	4�	�ֈ���"�c��C�
����6V_�j��ih��Ϋ`m���5�	m�c�g�=0�û�ʿ�Ex��ܾw�?Bm�mݝ��R�G�Sj��!{�6��LN�3��zxۛ��nDWk;B�������յ��-�����!���v]�v4��#ˠ�͠>X��()����􃞞�����N
�ĎX��!>�$L�d;�7o&��_��B������Fs�Z�u�0�Ю��ZF����	��?����s� ���c��A��'t����_he��Bcs��:��`�Y����|rf���%�r(��t�g���!��ʬl�Z���/N�SS3�wq��������
q��$�O�
���NZՂ���Z���ϭ�xX_˚�9	[֘�ױ>��ޑg�cQ��X;ʦ1��0Wz6�ET" �F��af����w��	v���ʋ�ë*�lny�)�02E>mEi|�".�e��$�o$�V����Q��{T�P�Xq��Bl����zo�g�D��������m���l������뿾�rm�/�"k�X�3("c�}u�t��ܰ�:=��7���á�!�q�x� �����M'ڄ	�pRp��R�P�ޔ��������	��/�;Im�m�$��P�u8Q��b�7�dJIv�݃��!��5c���8�r���h�����N.�9a�-��aڧ�����.�jMDp��=��c$�y���X�cɸ&q�l(��^ټ����N�c9��j�{~������%dp��������B}�hW/�j�h�W�X�2wMO2�(��Rī���oh��S8|�7i���:n޻�"���Q�^�E�Xj"�0��irJ�ǳ�K�P���V�06'j>[�G��ݾ�]�3&2D�A�'�r�t���������g[ŞE�X�~���|"�������>��wA@�zO�;f��4��Z�{���/�I)Pڸ��nC.�B>�BA�C�4x�l�mm���ַw�=Ї��N�ܷQ�K�biqQ��'���A��C�82�����5�1�0I��嵍'v0?�|a�4H��?������*�t�ٷG�^�mM�Kd�W'�*��I���-]�5�	����'�JX\X�y��Iaav��B�At�7��O�O�
��-\�qEZ����Z,rgvptT{���AyG�ݿ��7�bbn
�Z��w���f4u���fd����.M?k������9�C��^0P��@C�}��.|#����9�r����I�_KMH��ɍ8jk��hC�e��<{����DCk3�ڟSj������y�&�hb?��/�@���*^�����Cq��L�((Q����޺!k��yJ�_�����,�/�kmn66�Du\��Q%��YliC( �q��$	����z�Ɗ�f�$�Ɩ�3�w����炎��㝕l�FI�Йd2m���
�1��M�u�깤Y�e\Qi�Ɋ4��}_��3YN����� �߳ɔi�;�,�C�^�0U%JR�Pz_�0����!|���+���v`cc3s�X^^��м&;"[[���|��I�����`�_D��<��5
m T���Lź�&��A�*�RI.]���Y�U~@}cÕ���?�N���oRO���͊���������0Y;���H�"����9��n ����E��#GppxȦ�z|O����k�>��eH�h�i��<�+"e�@t��i�}*/��ܬ"��Q\��Ig�+�d"�n���;4��F��g�(z���<�b�RV_W�`u@�;��	�&�y
lgRX�Dp��S톺 ~�{���&���._��o^j:ɹl2�H1�d[W&<��t��E��
�b"O���ۻ��9߸sUE�7�5�ܗ�VQO�:����y9gqJ#��e�zWcq$��H;w5�Fp��1��Fxk7��¥;71� CV�s��0_�Յk�$�IC��b��I6!t�����e�W���,u���eqbQh��A�L�lZF�**L�!�~�2�0�8N�>����$�I$��tf�Q�;tGw�Q��ӗ海�_\@6_�ٳg1�;���F��{����9m��f�)����{��k\�{�H��C�5*�bN��TRi`/_����I�tu���C����Z�}��%1�z�=��_Q/ʟwl쉮'���aM�<�_����#y��KI�Ǳ��2�XZ��L����=�5�R�}�bȍ����T���-bmy�^�3ہ���~���jAl��ܐk����$/d�ٻN�Ɓ��j�޼�k7����Ե4�+A2[cKzG��>�$0a�a<܂�Ɲ�ρ&�(�0���OӤ��F,��Ҭ�0�#F�-�Σ��#�}�e�z��B�|*�<�)z�f�[Ե4cms��r�c�x���m��,�������0hˉ��eO_:��QW�D����MAx���ǃO�^��U��ӭ(���V�<3��LoiiBs�IIW|؈J%@�?��Jx=_;�}q`�&�7ߑ�7�J6�a��DKX�9�Q
)F*�˗��ڵkF#� ���'��J^�/�k2�"�ZE��U�M�66�V~gl8�n6��76�F�oκw��{9�jB*���]F�P�RI�<��Ta�GC���?��
����������4����s��]N�2��gC#�[;��֮a��$��,�o"Il"
��dTzH�Y�����Ư��Æٕe̬,bm{MM͗;:���;-�E�?|���re���׏f�L�h ܗP��/���E�9���?�����Q8���Wc�w�&ތ�Qɮ8T۬,͎�v]���-��ÈF��@�;}N{X>��}���>����d�0/�Nn�a�f"��a�o@T��eu�G����VW��� �A}CP����);�L�l���]C<�7S�*������wT�c�|��_`l�)ޮ, ﴡ�q#+b�u7f�B{M#0EEEXl_�v¿��G`��h� �����ʗ����*�-�Z�,�9]��$�9#D�z'��R$�7+��L���Y��	�;{{��b#��kwoૻ7��#��p��&a��<pޱ�y#��D��YYv�4��Ή���Մ�"?�0�y�r'Z�T��I^dYw57����L[�m,��be}M�?�6���M���c�˽~�Qc��39�����Gpj�4������꛷nau}U�O>������0�9%+�tO�@���b�_� �����FD��C�ȡ�z/���q��<:���y��=�3g��ȡChmn�K�$d>܃����ž�0f�,��k�n�Hq
c�������ך��C>�g�8��kx��^�v*.��������שqY�XG�,��,������TL���x���¿����wqm��a���,-�9⾔������߽��"xp��}Ϧ^���]�=X�l�d�|��|(�ɚ]�<h	�S�KXPNM+�jO�{�e�J��3
Y�]j��=A{�Y�-���[wY��,�1Mv���E4��bm{[E�D������3�����W�����O��ӻ���#����ӧh;�թ�Hl�m�\��8�M({�Bo���w<��/�f���WV���k�)���	o�g���&�F%��
Ɍ��	��!�ǲ7tQ*�f�C�VrXT.]���W��\�i�d:���9U��i@�,p���YŖ��w��~a5���sXE�TS���l��a�[E��iYlhc>���+s�����n,�F��F�p������3�����Uli�4;;�fju�!�fsJ�"B
5���C�����˗0�8�!���FA���U1f�����J�p(:m����m���~���oη��)J|������Ĭ���^�$�"L֦�y�Z��[��z�OE��8::
g>�������}�̾�^�����[���^�	I�b����ے.�݇�~�����z��5u�|C�$�q��ʦŪd���)�ɠ��I�e����p��)M�4`����B��rϢ��2���tYN�>B����!t���}�5u��#��?��O�0D��Y�ܱ���tv�n���h�b�fFoځ:��s����[Q.fT�/_�Z�!z��>�������o�о��8������ە5,mn#O���ԉ3�p���c�yS���U��XW�-8Zt
�S�>�?@�Xsh�Zf�_��~..*1?F�F���w{�&	6Y�w�b��R�B~�٬�3��1(�Nd[��҈�u�@��f�"t�Ke'����v����8�:��0��5ݻ���5�Q#�u���@��4��oU�31�zp6M��ܥ{w�卫��S2j8��0>8~�K΍[70��gg��=|��GO�a�V\�l6If��j,��Ng��"�.߽�l�(��ĉ����<}�B�luC�w�)a�F�6�f��ܧ��7;��ɤ~v>#,z�E�!���1<73���Z��Ceg��7;����!B�$}t���9*����7p��5��y���.�4�u0�ʇBI��V��� O�S��*��0��nG��^;���^x�.��Q�ќ��d������sT����
�.9ȕ2B(_>y�B�0�Am]�G�D�jo�ƹs�p��1�UT�'^����sl��ERTw��~�A��h�A�@&�֮1�u��6�;u�#��N����{hH����e���7!?���]`���l)����ѡ����&�I�/,(7ziuE׎�3md�>��0tSS˻"�B��W_�ʕ+j���-��U(�/���W���d2{�"gY�0W1�C��^�
���hm�������L����U�0�����X�9l����ȳ�?�-�t���h@�D���Z��F:gHb��i�&��#���=�KkH�˗/+&�r+"d"��7��*���*P���6����`��LH��󶣽��]���L���MQ�E�O_�����,����kg飒�qZ��lQi��9}8�?��O����! ��ċ�>���ya���=������]"//aB-ܵ�c����/e7�_�{����E�䏕��dV��7��� �̿��;u�؇��&����	kj�o۱muQ�(����]lk+��5)���I��g"�ƕ_���1L.��q*�r�r�"��a�I:�y����儇$�x�7~x��>����J��q�2.]����%�׸���7`\�<>Y��h�M8�����1����Vװ���H,��
'����s&�!UL�����1�i�h�|*�$�)Ɉ��^X�XA�"+�4,/4��&����I�D(hlA���M�<��Ł]{��S��(_u'��|8��o'�|�\�b$P�P�|�{�F�߯�-hzi��ܑ�p訂B^?��۷���3u�]"޵�Z1<0(a:jo+��`r��p*�Ć��7�����؊%���wX��˩����������##J�RCGS��!��#\m�����#���10�����'N
����i#I
�;*εȦA4� �M	_{&���ʊ:vA����
�
@novY��a���n�6>�H�*v��+��\��[#E8{���ŉ����S�߇c�|��i
�W�Đ���2��4��p:�a�or<���QSP��N��}]=r��c��4�d3i�Y���L�P����z�~z2�Rtg/_����"���	:�    IDATܸV�6�������=u'�FCm-�-LL��/��\��a�0�M��FƼƴ�d��fӈ� D@��*��[�f*��a��Z�C���R��}eu��&R�t����tV^��HT4clX����ʤ'���������c�/�o|ml��9���>�`2�Y�	E߼ySn|"R���6��pMƿg��ݚ���ʓ,�NH�&�o�U|�~�/�m����mlg��c�%"�Ju`^�
�<��@��庆��Z��Q�ْ�ΜDgw<^��.�6����ׇdW[)Q,�l����hm�R���;�n� Ygk�����PUS+�sW��{Ss�[Z�������֞��7l.�o��7�	���O�=/�xzc�c�M'�^����m��[2��J�x�0�3>,���'�0��!��}da�و���G$/v)�H�ry��Oeae�ʯ~�+1 �f9z��U�0�0/��$'h�@7�6��B:�����#���C8���/��X	���d��l�\u���uj�ƽ&��?���G[}��|}�<z�XK��m��.U�J�@�(�KM�ׂli���pUف\��sGa���l
Wo|���\��FX;�Pu5N�=���.4Q�O���,�M��r*f�'����6"q��=uF��辽�Ғ@�O�o��"L�'�0eg2�O��t�F^ci���f�-�Ĥ��׉�DN��]�5�)��Cسk�",�v���;����ثqL,�c#�c�O#��tŇ�t�v�w0���#�x�8z��0�d�n���5�k��f&�n��O�jkk3|U���`�afs�x8��3�"ۭ�oi?t��1\<A�fv���ܽ�ɉ7h��oatx�=��L\�k�"�Ѫ��a�߹U�K%0���{o_˻���ǙӧQ��J=1���}��pfmg��!���D*e`~:�2�����bi��p�Ю�b�ǆB0[��C���C�lʲ���y!�"R�a��h�I�2���>,��
�z�4#�@J�8ue%'��hnihe�C#��!�C��,���9m҆�f0mM͒��m�b��[�KE%��PNt�0�9�׉,H�J+���jyu+kX\Y����4斸��m�C���P�I���~��߫{mt�wb�޽��)��\ES�]�;���&m.�,����%llG�{q��q���`����&��$x��%�8dg��!��ؓ���UC�g������1E�M�@�Ը�$�^]M��4U��1���5d(c~cbEm�w��m���?�ZEٜ[�a�����tK2�#�\-�8���p��C������CYMV� ���7�M�^l�H04�m��&npx �u��n9ʏ�
izS�|�Ue3�u�������ud}�TM���
ei�YCFGGU���&�ʯ����9T˴������������OQ������'�s�qr}��wJE$Jyd���εÖc�!��M� �tt��#�e_�L/��	*d������V����G7G���@�l#c��KcC�ҼQ9	��z���s؈D���Юau@��yA���WI�N3��67�����Jxe�o�j�`A%bymi��/�I���Y�0&21@��>��4�"��杫����`T�ܚ�yM�f�H��ts�	ji[x�p.%�غ\8������A>����_a3������āÊ3�km��0o`�V.~/� ^NO���x>9���(�Ξ8�ChמQ�w���{��f%��b�������T�������Y�|mv�S�鋼@�!���勨a�����Ÿ3Ԃ�#�51��`��;���h&�7�s
��\^D4�R�eWt�W��ع��3��gƅ������g�p��5���aF8�,�]�Â��{;��E(Ԡ�0�H�0"t� �G/�c~cSz�h<���~�s�=�ɞ���7�x�x
���I���!�d�I���6j��#�@�	L�󳘋lb)��f:!���|_�/|�l\� #�v�ك��$
)�Dkx����g��/�XZ!��,���{�*+?:�����,�mL-2�|N��D�λ\�4�����^D��PW�Y6������A˙�2���g���W � �̜.�ux�~*�a�Vl���✰��>��<���k��_�����qqJgr2�߈�ى���W���E������EOG�����I���?��҂�ǎ:"�����<K2P��Y2"�q�T!��]��a�>t��m>�SoU<�5~�>{}�-2�ȧ��U?mQ������U�`��F��0av�v��u5uj���}[S����B<��U}_����(�40.�aB��=ճ^�|5�����ZM��C��D����������5 �\h�J���e��7y�1�4�6E5�D��s',0y4J���]�34�\�"��� �f(�%96��ť����^6�6�{��%�$��r�*��*'Ps]�L^�:̂�#�5�-�-m��������Q�o�������vc�wX��(�o��|��C����l�� FۻT���= Ǭ�gO���-,�� W������FOG��O^d^`�&��I��#{���������)L߻of�W������HtK�#@^���&5bB�#C�8z�jj"l-�̩@+�I3���'1ԼHx��
�`=���Rsح���#���#�LT��=�=N$JE��-��W�q��GX4������D5�)�c���]���ϱ���*��M�8�� ��z��ܦC��'!hn�([i*���<z���Laay�9q椙���ٍt>�n���;�_D���$bѦ����aȨ��$��	��Cb	��(f( �IX^�����X�m��[��ZW�\,���j�]C衵#�|N$��tR��)��a$��(� q��@�!�<��
L`�j��ǹ��q��1t�7`r�aNq��!Xx��(����Ѧ���)�#	Bl�b��EH<��"O{T�1�7��{HOK-9���[7���C,//���Jpd]u����#�GC�ΐ@�ەڥ�.�ى&���Mx��6��%�ƃ�{�[T2��c� �W�w�>x<~,����o�WK�V�H��H�:(��,�r�%Џ�aB�"Y!ꐌ�#2U�j/B�T�]���J�����p���O����p�{�2r�=���sC9��n
���s���2�������V,���L�N�S�	�ρ�`��P���m+W��U\v� ������;q�mE���SL����V>s�z;;�����~�˿�=&FFr/M�~>G���ic����{�`�Λ9ů�0���x6+)��ٯ��՛Wx;=�k@H�丵�����TȐ�l��HP3q�^���=b&s�e��N�ѡtdsV,}�]��Jƴ�욄)W$��������wE�E��6��"��l�}H�(�Ŧ���(�[0�!���m�D�v�֚�}��OM�"6a4�\޻��9X���"��	�2a.�y�P����EzP��u�6�`v��Bz�x��$ƨ�b*bi�E�U̡�R�7]��9]���

v���x�g�ݍ�P��]�m��ӎ����6�����͟~^�󩍕�zW���CG"���9��2BN/v�wⓣ'��TN�1���&ṙ)�s��^��5���W�� 	
�Wf���?�׫l̛�o`��b�(�*5Y�PU[�n�Kv?���x
�,E�)��N�����CsKH��m�D������Ң&�x>GU5���Ξ��������	��;�N�q���~t��&�g�,E���.FX�p�)�D�9	�%Թ����8sp?v�t�V���_�����zv[�$+����$�?$+���:�n	���^X_���"&f���)M���ELٻw�]����L��g�.��,�0��k-xɚ�Ⱦ���������Ʉ�(5aes��A������kT�}X�[c��������
�Pʉ�@8takM�Ӌ�X߉"C?�bI��E�6q|����m5��p�>8z��A�}9�[7�ʯ���.���]����{!@r�����$���v*&�#c�$��m���Á]�p��Y1��"�v�1�nz5�Uf�t���Z!�A�OG�<�
��/�];]�:��+�:| v?�8v��k�~$cQ<���d�T���z�u�V�]�(H^�t,h:]M�dcr4K�`LB��0�iK�X%[�k�V�aH%���:�2��l��W�Y
�I5�L�k$l˃Բ-�ME aA�c�:`X��&X�)�1Qr,">�GX�z�]���ڂ�S�q~�8��]��s�(����q��S���Vi�L�2�_\���
�k���S>{�z������7���/~���U]G�R�^q�a�͟Ŗ/�'[P���d3�A��d����CM�t�����3�n0b�?����5�'�UQ�-�7�8"܋
���hg�������4���Z&C�*�u^�S�v�Tlk�����7A#,�*z0E�@�f�7�͎�:��]�
yew�f/O�zSFޗ3�4M�I����w;��I�$�ɚ(w��0�%�IaN���4
a��p�}��G`�B��\�0��J226��̭"L�d��Ы��<#c+�n�٥�՜SP���9�K.hD��l>��5��i���O�����"��o���g��1���q�\�N9oRw�\�Þ/Ù����n����;�N��}�1�t�9ݻ�����2�z�����S�`˃�7z��Z�������a�<|�Ϟ�mgh��� 6�#Z��ͩ��UFJ�Ig��'u�yM-�=xh?z{���_ZX�Mh�"���EAM�	�x�I�!ɔ�[)������w�?xx�����"� w��Ln�@��o��é�JvѠd��Fw~��EM»��h6�"����X".ؑ;��`=��*�^M��x�r��UV��$��Lbyc��M��v�9~Ο3<�I�ڽ�`~1� b�^j�+9�d�Z0'wN�z@��\y`y8���i�u�8q����B���+/�|2���y�]3�����n�5�i��*�O+�tRrja��֕��Aw�|A��T��	���T�?<v���}�wn������H&�����	��=����+��H<����v��S9E���䤢��&�����v����]Ѝ[����C�}�Z�z�<h,������$x���r�v�0������3kh�/X��WMIG��-<�}_I-�*?N�?k���@��B���["����9/%q�3݆�&��]tb��vE߭ưM�ɬ�FؕL�=�yr��d�?��t�5w�p�쏮c�9;�*P<�,8R����1[�No�,R��E!�	9�S�*���i�XS%���,��b-���2�Ns&w�^t�d-�lŉ(�����Сk��4��r#�����
ghkiF"���So���_b���TF�+2������ڜ���ĕ[���!�>`�M&��=��.����jf�=��w1�l�cld-d��+W0��2�{�ŗ��7!J{PQ��RR�_&/i��e7��#d*{�|^g&�K�>��]���eɀ�"l�o�H���=洊�?��3��)�j���\.�N)a}���DkMgvas^�BBr��ʲ�.F"i|�}UպO
�R��̚��:P^���@Uu�dsl@3i���������0I���!*��1$2DJ��sJfT)�\��2�6/:�������;���"�W7r����"��;�������(��|�];a��6��;�E�ًB"���Oq����L��E8�؎��Fݐ\��-�}.�B�e"�pǘ���<~@r�"�GF૮Ѣ|ym�^X��=Ŷw���#Q�7�So�f������my����CA�י�99�PS�ڂ"��@����ى��?I%�I��û�y�6��y��Ӵ�E�D�U���C���� ����R!�������s�l<`�v�T2�)NwV��/M�:�Fh�@�E٫�sX���N�_8w^�p*�1�ʽ�x���d1�۫"N��Œ��R�lX�9!��Q�t�,�l���gَ}�C��7�j���M�hl�������)bVwW'Bu5�ȋ$��~>|������-�z�FA
of��������\����|��I���`v��޽-ol�GL�i5c�P�l�Ŵ�d׫��lS~�j\�$�Q�So���]��:�T�i�@�3٬�n]�[ڛ7�!��;�!���Ԡ��qfh�0�)T��Vj�g�M&��zޖf�kj$�9�� �}�lF���CLL�B���A�67*��!�ds����Y�i�b#�儔HI3KdB뙴$��}^xU2��5[a2��愬)��MŦ��DP,W yÂ��ŝ���<��	��!["�lvφ�c�étF�]	B�TR�KJ�b�&UX��Vc��Q1̹��A�I���k��7���̤Y�vPb��"�aJ�l�TFp9B��s�،}����3�D�jij��z�5~���a9�$ȝ�?�(d��:�����GJ��Ћ;<~1�H*��/��~�3�����2�+7�+�:_�km��#jX��ӳT`����n5��^����eFx�S��'��"gJ6Y���-��2ai�	�!B������4El&U�	&PQ�`����L����Ǭ�m�����[6�|���_ϸ2I���S�e`銓��
rc�d�=ͯA䍱�K+�������d\(w�%�O�1V�)$]&^DT������St�8F�5�{�㱸�|��#�9���üb6]F�a��BR|U �ߙ-�����pW��n��?	���OϽ\Y�˩��3	I�����C���]'\�"j�N�56�'����ǣ{�{wocq~V��e�`5v�J¢��ފݻw�#����@'���?�s/_��]I�/
'a^Tv5\�3R�E��<������zd�]W_+X"��ޤ��I6x$5����zt!����5}��o��D(�O��G��Q�̓��q��<�x��ێ��������l&�o¤]�f�k�N8VD��Q>{� F�:��&4	�կ5u��$�g�C8N�!&��@(�N,���KJ��Lf�ϟ:�I�6o�|J��wnbbeEE���+¼y�;уZ�ue�u�!͇�d�b��*��L^.L��ط_L���l����Ǖ\��]��}���Ӄ��l���#D6ԙ��܉�c����}�+�m�Ƣ(8\�0��@���Ȏ>q
���X��Q�~�lL�04<8����Vf�4���<j 9�ӷ���e\�{ӫa�ӈ�p���}���E�C�|�2�ܻ#^���!?z�v�Q�rz�'a.�<c�^%E,��fV��z�-f«�3���
���ᩳyk�؉bl�)<~�'���k��Cu���V�a2���=_V�+����̞e�TJ��	WךL�Ps�D��5&d'=x� �B��_Sl%ҒS�BH�v����-D77�O&u�Ry c�e#��
�u_fsy�3�����3�a+{l���/�jq��a&{�9�{qykE���L�ij77���.=�D�h�� ��-�$MF3h�El;�C����Ο��3g��X�x4�Wo_��?�bxI�2	֡�)$}�v����.�lǃ�P(���l�"��������a?&���JNe|�X$�Ӭ��Y��r��>�$�]N��s2%������6Cs��&��%i	[��}@Mkc�Vrʜ~��������a�-�˰���h��x?���H���+��w�s�o��ZP�;*�JV��7{�Jm�Y�77����4^�l�p�Ďfַ���a�Y,	��~׸�e��P=5Ȑ1�a�h�t����v!��w��0df��fP�}t��!^Iq�����$]�����?�����;�/����?��^;��YD����9	�p�����F|��\8|�dϟ<ă{w�^�S�� �;Yd��	�Ji7<00����v�\V�'-N��5ී�zhH��UWIwL(�Ł�Ir��'�'��n��o$:k�5���sBBө$�v�{{����~\X\���jiş�����n�&�ѓǸz�:��G�e�0�K�a�KJ3�T¤bM�%Ih�D�e�>�p��;;�����k_��_K*����0����ѮQzW�u¨��    IDAT$�0H!���S7����E�7^\<y�Ξ����(�s����y�<4�Y8]-��i�gcE�o%T���(u���t���pܛ5x8�� ����d4��%R[Qd&��7:e�r��>H/a ��`;���ך�T�ZZ����x�������9]ȱc/�D <u� ><u��i\���{7q��5=0�������?"����4٧
��Ц�{�go�����ѽ�����"�|}��޿+^��}{qx�>����F�`�_�N�s�h�L
�TJ��s�K�\]�Ld.��u�(׷���T
o&���gx1�K�M2�hj@SW;��Q{�/�����Xd[��0k¶�����֊��VIo�������V�`F|G��U��6@��(Õ,���N��C�k�1y�D?�H,���E���H�,�:.x��K���x��9pMM�: g�sx��%r�2�^�X�K�a!$Z��XDKc�B8³�}9���(рr�S~Ylڋ������h� �bb�������ʢ��E�-h#B�ޮ��&�3�HmĐ�Č����?����N,�gϜס�t�%�޺���x6]I��RԺ���e�#}z2-r�f�9�}���>��),$��
j��H�}f�4�H���I�M��$P�tF�ZX5�2	�BW��Y��B�~�>F�Ε��!��	�Rl-=0���[���ኑ��8%�P��O+X�c�^�Y�lxiV��2��aB��D}�~8��Y0+`��I�Ne�$Fv�e{)�2�+Zf*{�w�bNh��5'fʣؼ2Տ�8%����˃]]�����o���W���K�9�8�r@!��x`���*���(;��Ј�9��E��ŋ'����==D�	WUaqi����H)omm���d���it��d׼�����5�������;�N��H@��ɥi�7K"�@uM��@+P�J����Y���s���$�ˍ��z%Z�1�����ֆ?�W�=݂��=0E���]vdx3x�(p���XE�0�e��"�i�/�W��|��'�c���DT����5��bg_H�p�e�?:�[$���u���y�����a�7n��L�\Ю�ܙS2*aD�Ͽ���"�4x�ގ2'�]��Z{6*�Ɇ��(R�	��.�m��8}�:j���`{uMc�"��*�j���10Їֶ&�3)D�;��)ѿٯɍ8w@��r�
��)���+�2����p���55`ei7n_ǥ�W�1��0�Q��5 E�H0?\�S.k|hY�ޒ����q���Q�6:����D�$�pxW�_�N��zǎݻDګ&���Pf��hv��l
�b����x�8����:�p��I�L|�[^)�Տ޾B�1��֐���>�MbHr�~�ˈ�@�h�j��x�[Z���ݍ����%�[�����9��ő�CT,򊾔�SJ�*��wN��t`W�<r���16*D�����[��3[��e�l�T�s%�4qz=�� N<,8�d��o�x�9\�>�kHr��ē:��]W[���ҟ���xp㶚^��`�~ʡ({���EA�\y�Ķ�v�~��ϰ��h��ː+RGOBm�פ|���l-� ��͂�_>@,r6�����Q9i��<{5���ob���D�4�|nleVK�Eͪ��LV1�t6��ˁD{nJ��$��"y����c�!��J�Y�YE�9�4�7j}�B��"\��,��j�̴k$F�^�2ڰ��ռZE�fDYK�l�Sd>����B�F�h	
eyR���H��j�@m@�?�E���	[p4/��>���pT��VW�!Ǿ��٘(����B�s��˝:v^G!EJ�*�Jl�:"�!�1D��	9G̿����`uu�\�M_vw���g��߾Y�_|���//�x*�~:��.�c:b_�����W�p=>�p���ݍ�E��QBD��VL+h�@��߉E�H E��,�l�ɸ�C6����2��hf`�wt�P�v\�ë� ��whO�ݯ����4�1 IP�iBF����������M6wcO�+�hl|E���I8S!f��b��q�y�(尣��by>\8qg����A�	ܺuWn\�o�t2-���`�6��c��4���o��YXT�- �N"�����8s�ܯ����[��������u�����ܤ
4H��(��.pZ%ZIJ����$\������H{'F;{0�ցB4��u�����*)!iim�����G�UScP�o4Ss����9�~���d�I���4n=}�gӓ��&<��./��هs'N����+K��]���������'80�W�Ry��/8=&H�{0���ڒQ˃�/0����:m��Hp4�Y��M���/�ե��^��G�{dXE���Ȧ���E>��
��3�1I�\�Y�E�Jj��o#�͡��߿��kC��|-n����K\��Ȣ�������ܑ�S�w �)�i{c�<�rPb�4}pɱ���0>Mc�i�b�`�NEX��l�X"w�HX��鐮|�[jù�;e���3��p)�G��憊0����>���]�7�^�������ʇ�Ls���>���g�T��T���|��;�4qz��?�B�a�Gl�TŦ��ӈ67������~��?��������&4������≔y�˫��m ���M#O���P.�l�����}_��	�����%��ڂ��^x^CӥS���1"Q$2匧�b-5��1w¥\��FS���	u!!��;坔X�|?ؤXE�d�А�3ް���_5b.�Zf��
xPz�9O5�W^��Ѵ�Ϻ_*llM���Ng���y��ׁ�4�{�m+P0}�-�&گr������q��g��ou�P!Bʔsq]�b��o��ѫ���m<W�|�VL����ϐ��k�&���9�<�.L
��@WO�|ݩ_�x9�`m�/�;z�����_��'��|��N>[^��ɍ�w�f'�Ҙt;Kv�sExv��e�@�����s8u�(�����s�Xʼ(��X��&��DM���M����<[S�m���$����	��D��Q��u��&muq+ka}.��#�!k����]˥��f�`�i�0j@��:�\Q�?S sﮮn����+��yܻSټO^���"-i�et�"�R���$Ex�Y���l+YDΝ<���w�\����k�v�
���C�7����t�Q�iT��D4k�������"2X2����N��A2�Qƭ7���+�ZY�������_�a���A��́�+j\	��!dT"wN��-��-��m��ӇV��
HD"2E���"��G&w����^��]ax��
���wL,���"�����>~��/_`�&���)�q��\8u
�!�����ۊ�#<G���=ؤ�<r�k"���i�u��e\�K�����a|fZ�q._��Ƒ=������v���|��)6����ߋPC�r���T�QΑ��5֒"��$���Ƈ��g�����a�^ۨ"�Y�$����&�Ø�Z���El�2H��HR�������Gqs��5D�7�����pC#��Bb�S�G���$zy)�~��O[I�(C8�I��3&���&dh�H�b�V.''4�ˣ�,��$;ҳ�����<��:���K�1��EF�R���UN7���ؾ��58�d�������눗r�
5���M�%y��.b���c����$R���U,Nϡ�ʣ��_+*�O�8�ǎH��f���4~��/0���	�������kK&�t0T>���D$�B<g��:5zz��ɛUӣ���G����! O^<���w%w����vz}�(�@�hU��G�UI0?'3�'Z��L�(�>3�E�����<����9�L�ϕ�^xߑx�g�8�DZ���4�����"lHa��F�mp]	}���:�Wh{�kU�+5 Yk��?g<��ͦ�Q���ڊP$���|��w�A��X�u���k�H�#'��vtYtre�{�e�d,�,���V�Wx���0͊өk�3��2�g8�ҷ]�"�j26.p���Ő�����@�?��v�٧�m|�E���c��?~����N��4����c�L�F� W�W� _�.��'����#���x�Ϟ<VYdhR���7hmC<�*�3�5� �QrY����®�ף9Ԡ�-�Laiф@���ͭ�X2�h���bjwm���b�$�/� lzCt(QII,��
�
���T���,��?�$l�4aZ��P�.$琣���2��pÝ*�gs����8{����	��_����������ޡ�����䋗�R�Ix����� ��	�!���_^�'���GU�i2��w��M|}�2f�����1��Y��h#H�''d�����0���\^Ը��	����C-m��؝���XZXD4������E׍�Ԕ�q�ǉtieI>��TB�:�0���9gM��T��>{"3�|���hCU-N:,N�ˋ����&a������k뀷���U�e+��I�$v-�0X��y��U���S+�x;?']kk�YS�����e��8� �,ڧ�w���.Oݱ����v�8����4B��n>�a�cy��௯G�m�b"���Zu����,p]^[���2��I���X�$���x���6�3E�b��0����"��w�����]��9��1��+*в��$�9u(���U�7v��TX�b�����,O�|�|�`e!�o�Mr��T6�NYa����˙)̭�be;�C�p���C�݁]�8�� ���a�~�6V�[@���.��kM����%5c�6'�R��anr�X
�U5A+�Z�q��a�>ym--�1s�'_�+[:؛�;D
��ƹ��{)c\o�TH�;��kkj��K<WZϿO?����'z�<{�k�n�I/Y�)���e�ݰ͹[�����ޝ
Fv�$�BX(�UX������钉���������m���F��IP*�n�be0�3S��p�o��)éSA����W_�:YN��	�aZ�Yk���`�J��g��Z�'���誙�}�7����0�����[L�Z]5CA�M�U`�պVD]��՚z����!�i7*ZT�k3�Ͱ�]��<Wˀ�>�&2��l6�U#/������c���WÈlms"���P���G�l~�E������+���������I��@�xz�"����ޢC�,?l�W���9�=~T��ZxY��AH���g��<�����Z���Nq�ABC.��5ux;�U~�ѓ�fw �JH�`+�n����y,��1�?{���a�dS�?ӛ�E� oB�*^������������ |~�B���?Q"��g���)�P!'{6$��4�?d��bc@�R�ݔ]� �9v珝���{`+eq��u\��?�N����ݧ����w�2�7Y]}����RQ�����$L]�����ԙ�8r��`�[�o)���f_�i2
��nN�=ѭlzfF6�4e��:X��˫Ԣ������A�����5�B��f�9=0^WZ��3mn���Kk+rBc<d:�ԡ�i�gx���������x�j\��LAE���g�é����+L����|���,��������87<�8���y���+��l͝��][JI5�,����;��p��ܿ�ETW�1�ׇ�{�H���F.��^��6��~*��/_h¶W�li��&���0�c;h
��Ӌ�9B��Ǜ�����B|�[�v��
���#O+�`{eM�!`�hy�t��cxh@0t=a;5�f/G�)1W+�O�R�I��\��ؤB�l%��L@�"n+�oC��]�Ȝn�i�@�a6�g�S��4(�]]���[%�-�����C֯M֭��G�Z��*����k���%�*�S=zw�BϮ!�l��)�"D�qyIG�H1�`CG]�\ks����+�ܩ3hj�G�֡3��/~�D>���:{{���N���ѝ�H8����fd�uWK�,<_=}���w�ݏ>�G~�"���c\�}/&_��fCϳEV���8*�e%�q�d���X�"QWDM��E;���p��H��Q�,�-"�Շˣ��l,K�Y`�P�Cu��BHdRȽ��Ҙ�XEXT%t��O�7�r�����+�W�AŠ�EX���>I�V�0��	�����~�1�M)w��ц3�b�&�02?��"��$s���@���8|���@/i����KgRx��&''uO�֯���ԕo�zQæ�k~�@�/%�T�-5%U�\gzA�@xo�.-�������w��lt4����饡�jy�(��ܫ�V�7�Q?�9M-͸x�4�;{��,5��$���,\����fZ�9�FW�P � ��'���N�X��[fxٌ�>�Yc"�tf?҄@��re��ԍ�r�r��g1��>�|�7~��������D� ����ܾ����)��]��ȶ8i�)�L��2y��|�m��\�=~��ޭ��ֵ����W�C�����BC�-�'&Q���ݭ���Z~Չt��Z�5���ؑ؝7֡�Gp��	���gܼs��^����,
����{�ؕ�Wb����9�Yd1gv�n�;��W��a0l��<h��_��o���7�X,�4��G���f��3+�㩓��ֿ7�#��.��������[�
�����X��;:U�g��p�M[��=ɋ�����]��&`W:���6�'�q:���(H��.=yّ����uDKg�v�k��[\P���Ɔآ��vw!�ڂ���x93��3��U(�7E���]��&&�ceiO_<ŗ���Ozw7w���]��<����҇��i��0|��<�;;�ux���EM/����Ə>��P@��_��w�>���"�	=��g1���ө�Og$$6ylΨ%�ZYF������x9;�l���d#~�G�����W�&����kL�/���(�� 
�2N�22�(g�jB����֌��l�cW0`&)�ek�"L��u���F��E�M�Z��Kl\������2EV<�'Y�lb���2�`�H�2�W��+��7/el���+Y�|ܐÍCg��B6u���)����q�K+������]C�p�8arm),׌���Y���k�đ�����,��)ܾr���'�2dc�������+����Ds38\� JN Ms�bA+	jp����\dD��%d��������mܺyS���1�<}���9I2�@KS�TcqCZc���1-FvѤ��'C�m=.�M^י���3� �!�M]ɗq����T
�hܘ��|*���U����i�(*I8]r���[b���k%��n>�4L�2�Qئ ��T������[[j<X���"�D��'Zm�3�$ˉ�Œ����:a�U-��PNʴ	=7j�1|\YlZ����r�&�4O������//��(�/���	s�bɄQ.r5@B�K1��)����c,ml���8�}����Կ�OΝ;����������ѿV�Ȕ�D��YwR,�ܑt46�0����:��T�B���t��^Hn&t{ក�{��*���m�#k�%�K���Z��q��$���NM�k½�)�M��>vU���{�9;C�"�J�gj=��qӿs��-�1���o�>��ׯt�V�C��e�&I��<��=�*�1��KYC����uܸx燇E����]|��/%�hmk�~z���I��Ʀ�C�u@[���Q��'�H��+�q��+�/�֭[�t�"�������+,n����9�&2Yz;NLb��f�L&��20�T�X��}���D��#��7W�G/�=�Ծek���y�pY�@6���7w�hǲ��cX���gf1��ۇ���Hv����^��`lnN�v�qw���!��;׮!�aqiϞ=�����T(֡y�oX�p/��3�;������9,/,cue�B	��m8�f���l��?��4�������������\]A,҄fh�g�(~��nfj
飔i=nL..biw��fDP�yu�0��?��O���"��7/���#�Z��92rd�8�^d�4�Ul!�Y�A���i"oki��5�6�/�    IDATƼBdcG��eާ,X\eЬ��3v��%�W�K�a�^��FI�3+M�:�h�X�.�׃�J���>�drs���=.r
�}��g����/���x�Wp��WIaGF�ʘ (@׿����G��{3t�
znJ"��O(��1Sfj�Cg�9�J���s�������m����,�xIMR���;����ג�P�Sw�ԄhcR\Ƃf���8#�-f�g�P��p}8��S����׮\�ّ�bOON���ӧx���I����Tc{i�Nu�J>G-*M:8��=c�Z����Ζ<�9rG�b�B9������r�����g���f����`¬j��.s�hj��֔� Kl3���� �� ���k�]��)�\b�����/{*VP�`���;�OH&c�c���?�Ή#DH�g�qEHF�zl8�&j�k��q�m���O~"R$������rq�S�h�	ܐ�"������ǐ{�ۣ�P�o� b��6͆=ӫ�o.�:�;9�k+x��o0��w�5��߿y�~��7���-��o���I�7 w9n��A����H�������>��w�Zu2��á�Txjؤ1#�D����At�C�|��7��b��]ݏ�՛ǡ���]";�
;h��I{դw� ��މh��UQ��Af7kUgސ�X鷻st���,,-�F)+�<	��~U7��0NP{�e��c��}�n^�"B�_y����'���d˄���u5�'i��%�}�LB>����P��ffG����+�s�6.������op1���z����:e�z�i���*��~&-���o.v�-��j�BW�^�I�ӈW�����ԇ�B1����9u�|�Y��b�$��7$%E`xF�T�!������A��r��F<x�K��^^��Y1W���AoS>�qw�]7ExaO�<��_�"��;��#8���J���5�<ډ�w������:��Puz�7<��ǇÓ���Y�G����JLZ]_�w�ػ7ؠ�q!��.`C�N�X�E�����%T�.L//cyu����(��o=�5fg'~�'?U���ӗ/p��}<{g8�t.�/�a������������N���G�i!Ad�VʺΉ�0zj�azixTL�v*�U�3�Q�edh��|5����v�5��$�
�7�ߒ��+W����"���t���]X�l'E����ɽ��]=�:2���gP+�87�Ͼ�{;"�9B~1��D��@�ʓZM�59%��]s �tk@� g�� �3��8��c"p�51򹣞]^�(�r��8<���a5Q���F�L�>[��0�$)K���w��M�"+�O���G����S�Ex���w�G�|�������}8'F:�)`fc�p(����uMlI�DN��r������x,� 2�iw��_ �&჏)Jt���ơ��;M�>��X��1���-Q��
��Y��I�Jh2��ba)Tj��rQ����B�"�3���~�l)��,�$@�
�jYX���?��8;:��&}����ff�ͥ�8lNTT9�U��B"Ԓ��� �sp(.
L�~l�Y��Y˯ҼV2�miԍ�-L.����"e�������ůc'���y5��?L�,��	C��/�(X����HE���Zs��H;:�_?@�%*�*%Dw	�Pv-Vj�,�a\��w�Q;� R�I	Pԕ�o��'w�"�Ԍ)/j٫��>�jAʢ�[N=|�Yl��$�m���c�`��<��r�rSSl���=vE��X|�F&c�;`�c��ګ�]*��+Kx;F	̊
%�7�+�p��yM6�ܻ��~��U�#5�X���}��F2N�P\��J��� ���l�`�d5��ś���܇]9#y���߈y�"|X.��v O�K�������~6�,Sp���ђl���&���$�Ɲ��O���	y2+��7��R򴾾�"�)���Y���¼� �d���h�삷.��=��a�4e�e�B]�:��2˯�@] ���9<~����R!����_f�a_g7�Z[��ݲ�0����5lm�bmmC�3�����k����A�l�~�?�;��������ԛWҜ��������*�蒤D;���GO������%�o�'�d�ut�'��7U�=�`�/|����W�$�Ǩ�|p��x���EH(��GwW��X�Ȱ�*?ɉ$��S����
w�4�Q�N8�|���C����eCfVCN��&��\��rA7$F�J�P��\�k����M(���يh�*<H��^�� 1���\��)���ζ���k�4H	 	��s
�֘�0�E�!� %^|��KS��Z�F�љ�@51��H�i�r�}}&_@U���R���&��X���4ծ D6r0���!5(U�{I6�4b��n�>|�g/�J�S_�@oO~��Ǹxn�r�"�WRz������^��7�w�������G�7��X�X�y�s�L�r��|<����?���c8b�(�����
Z��4Y���&a�i}������z�
���Fey�����xlx�Hs�g&r�����|lonij�'p�|�E�S.Qe���������������)T��3s�	M�|+Q�"%�qgN�kw�,n��D@=yl�u䘴��S�h��.5�\��"�*�#4�Y�����y���9���_�����/�]z���?�/�L8�TWn���&���e�)�2	xd�ν!�"�������):��8��H�}&�W}4�������/�J��bF;Aj�����|L��՛�EX �L�x"�6���;.+�]�v�4����2���^O&E���M�+E�]n-��]�(ז����sr/Lw�|��<��+UL�L���g���c���֩��폔������_����bgG�a/��x�X���rA��\�?قI(��<I6Ų�y�^>?�k�.���K(�ڿ��.^-���p7����+�t�pIY�����.�2|${�èK$�[� ��Ó-�}���$��=�20�S����R$��Q
kۛbV���D{gfHD��Vǻ��&�^�Ѐ`��L
o�~|�=�^�:5M�j������7o!��annZ~�_{�<]�<�d��h
��W*)��tJ��rف��Il��{` �PP��=z,g�����[���P(����K�{���q�lobxp?��S�w��ZSGǂ�Mx6�Oލ��1�(���ܼLIz�:�?�M�|�:����o�ᠴ��	�^��*���7ݻ\���7��#_�q��h����ZA�퓯5�=�C� 
����7�Q�}�B���uŰ�H��m&a�9�A;^S2r�C��$&R�HJB��T���ɩi,�.+G;g6
�.�9�O._�پS�<2� ���l�h�Sq�4+a�Q�b�D�t�0;8��t}PRƵ5�<�8��S�+�ij�pH���!]-(%��H=y�����vB�E^N�,�z��K�J%�x��}��&�	�����k0�8�_�$�T*-���z>Z��w��K�c�f�vb\����x�*..���hT��z�����3���?��\�h��7���f&�&op��lC�6b�^����!x/o��K��]��d&٠~�C纃2*����$ςȉ�!;D8�ز��YId���G���|�v� �ݩ�~�������[�Z�����ذ�y���X4	U�n�3i�̽0��T�Ј�����T��N� �ld~u2i��O�s,��j�ȗ��88���������������K�����^�.�O������p���wӕ��{�-*=�F���5Z��a;?�V�!o�0w��l����2�:3N�071a����S\�s��2^Bvʁ��}��G��ܵ���nE�}�A��B�e^��k}���F����d;������وq����xW�ɚ])'>���E<y��>�N���G�n���[�t�<��#=��'���-���<x]&B���o�B�/c�.���y��̡��A"��*���x��}}/fg��QxPP�'��ok�]�L�S&�	)ҘD4Q'x�!o��:��r�|��,�q��0Nw������`@QbL����������zA�5�D�P='��wS)��2����!��
eM@���m�������ɍ�����ܻO����&���D��xvԄ��jH6$�H�E �n�1ь����1bu8)��Iaum]7%ؿ�[?F���6����=y���$�b���ę�a�ҁS����k���A�����ށ/E �q1��O�!�+f�'?�M�������_����_������ '�aE���b��:��Ԉ��Q����DLV������Y.+�룦��B�XTҋ��5K�
~��Ѱ�:jz�e�(�kg����AO���H�G�?fs�k�\�f����+,���)�9��*pa�4n�^���A$}Ax5's���{��V�V�n�?6��6���!,����ӱy>�|2���)�ϰ����*�F�)i7�(��u.󗔮D$��ɟa\{���S�_>�W_�����1�Ώ�E{S��s�K.YD_N�SJP�O$E��%b�l��`f~�++:�t�L"w���ɺ:$�q�h���>���Klo�2�-A��b3Y��c�����C��=�b��-�v4HO~�umM���[�,Ҝ^�|�xs���.Ml������c��dz�ϓ�$�̒��,�j�Ô#��d�?��KW����M� t����I��Mf>#߷��F�[��ʅ�ۿ�;������=��:�*c@�v((�u��li�:�S���2�:�f������[��f���G/������3ã�8w�������.2�#��+��	/v��~ͮ�:C������Q�~�7��B�,��(��c,�D�	�˩��Y��/.��dEs�L�w��GF�B�ө�"L��.Sb���4Ic*�V���:P�P`�2���s��t��%+�U�T~�����a��j�M������C��E	�xSܠ���+�|��=�g�+!O/�B��\���.��%��L�+�p��`"�HơĊN,<%	9(�4����{��<|�F&����U%�UCu�$�:fN�*�ᎆkI�AJ$��:��C�,L�J��Σ��`sz[��F&�7�'�y����K�snhH2M�V�d�Bx��>_����R�X<�E�ZF��;�E5�p���\��O��D2���2�=���}���#Ч��k�%�5�C�����2֗�T��O�@�]^E����4�OR�H�s�~�?Q` ���_~�Ǐ`nj��z4�r�I�b:�JL3*��><>F]}��v�N�����*䱸���s�XMuȇ{����V��4�Ѱ��X�Y�|��h�o@?m^��0�
%6P%M\����	j�]d�ל�	'�Q5��y�o��bmw[;a'5�t"��)�C�k�=>˘�a^��4�b���G,�T%��9�E��7���B�''T�e�Hß4	Gnv���鳸6z�@P�/��E�--�0-;���J)��>�\ˌՐ��#�C���<g*����*����2�}��ـ9-Jjh��I8Er����0/τrM;o�*X.R�VRQ�.��/_���_���FC"���j�j%_����u	�CE�Ɋ�O&B���j�����r�Ҍ��V���)}�уﰻ�o���;=&�Jf1��1֛J���>��R�,�g�5�|`���_��!���`�[��s�/�K��?��qiK!O~���9qV><Й���n�dI2�����&1��F�I�.Y��X�v�&���Sm<NIS���&밗��������|~!f[͂�Rx���'��ެ�pw�PCE"���=]�/�_��`�����O��������7�����{�#�/`��Y6t����槑#����9:�P��=��'?�j���E��C�P69�nȰf�t��TS�F��Ho�
���4v��s��N��r����A̴�b�l���w��d~�ߖ�%�f]p�_��,��[z8���%����!�t"rr���B�|�.��� ���!����W���7X#����+�p��%�xa���N��%3�%�.�T�I�{�(;68
'��4lS�����$%��~��Q���gO�v�Qq��!����B;f��9�[�ڐ�X �xD��(��9]��^�S�Y�"Ru�>1��=ݤ�U�K�����ކ��aߘ�K?ev�iN����������}�dOdTA6#}����!ݕh��^�oܸ��hD�ݗ�^೻�&��uu�������A�k���WJJ����ց��vh��݃�ww���!�5�u����}�V~�K9s��Uߐ����o5֑F�B�N�J)O	0�������U֓�o侯�����*�4b��5�1�jWGy^�^/��:�i>�Ќ��$�D٬V���M�\�jc�A�<#�h�AS�&�D�d]\;;� 0�{��d%;����|�|��ъa������6N&#�5��{=5��}�k��C:!�]�
Q����&����E�da�i
%���נ|��;�+�{!�$p���9�4Ҝ���s��E�PC���r ���8��keT<�gT��U�������F�����18Ѳ�}��Ξh')BU:��Y�e���ЬF�X,K�����n~v|/��`�$�`sg[�1���7� q�ǂu������[�똛��F�`�P�_4S�b���b��K��f��|�`cO�z-�,h��Ōc�����+���,ȿldP2#����5^rg��b��cw���َ�e*m&�"ɱt¢�C ���9��9�R�����?�M���I4f$���8��B8(�0��,3>o7 �O�8����σb�$n �'N���<N/����������1	�՛��y7�'뻻gΌ����i��8վz��}���m3NR�6DͰ }N��J��`����N������S/�P1I:�]4���mb�����z�C����P�([sog_$$y,�õ<���b&�ޜ$0�NP�U�ν�%	JD�LF=;d^$bZ;$^�f���Ȭ��м��فI.2�ښ[$�~����յ5M:���F�O춮]���-�=���`�O�����K�iX�Msai8����f*M��������e���bbzJA�Ufor���b�_$O4K<.��6egڲ�>~ޙ��K?J��[}"��8�hЁ������Nt�4��q S.c�����3'���û�	,omamy�U��p��C7W��\EOc;>�v?�����^�|!v�����0ї��^���"D��;�"<�{K`�����W��o�#���.����������~�c�$��������o�ݣXYY�!��>R�R��]�!b��v�^��̞�}���m�l��|��bzq1N����M�2�#{9��w�L�PE����N�+JKI�[:hQڗ/�%:�k�\ N{JS*�#-%)�a!�mr���ڡl��}̤.�4)Qf#��H�`H(�H ��'�w��<��n&,�+c�D��JM�NN�t�FS�Ijkh���:N�r���ߋH2�Xs�ѐ�T��UP*���h�^#��ȗPe�{6�ƈ2 �	�1T��}�7�f(�P}��P���oK�rުCʏ*}��6��O��ZQ1��o�'ĂaE�� ��K�/$󷬘��ѱL8I�eO-+}�noIA��G$
~�Y(�hѢ��ś��R��C�X�����|f�U�Ȧ��mm�
!SѨ���E���`!l4>�-Y�I$3ot؍�M�V��^��8A5r�Y���6�u-�˒8�e�����g&�X[ش�6�J�.H���7�����Q��H��ω���H,�X2!�#o�/�H$�D,��#�9�]|�<k��{������ZM;���ɗwƧ��dko���������.U<�_�l	E�Pc����N��8	�\���gF���}cC�O
i3�����*V*?��u�L�D��^ڷYF�>��������/��`���4�T�C.��ô���oB��`���b����Ύ�C�D��߳ ����
$�ǋ/����Ds�{T��    IDAT���$�ˉ�T�L������Fn}co�����w8Jg�'0z�΍�V0<*%��Zic��OȈ����[bxj�m�Lh^��`�$�]p �66�@:�V��I��C�������P2��k�'�z21��&o0`s�� �{�8�����	Z�T��1]��0��$����.�\@�R���1v�5	3�����������'v��cr�)��V���N|z�~x��b쮯�������ϴ[��A������A��FC����Pʞ�Za����"&����ǰ�>���.	I�Ώ��D�����/~��ϟaai^�u_O/ΝFc<� 6J�hB������ߓm�F�DE��vḔ����Db���L�R���/�$.«��}�zN������Ü�����\M��9�2ycѩ�kY�w�<|���0"�{���oe�*Mˊ�NԎ��"�qи܅C�h��9e���������(�Ed���#�����
V�װ����Ў�䞘ϓͅ��$O��46�����:��ܿ���."F�ea���'Y�N�?J��32-e�R�H���C�W�.�Dk��2}���LmK'�)�T�i��EO��M�f�7��/ٷ�d�*���0�U�2!�\��H��q@Ř����AM5r��d�{r"�7�#j�����HN���z��/��g>^����JQ��a�Cـ�r�JŖ�Ѳt����MN��8ĜQՠn����
�]tMR��nd�Q3|��Ҷ�Թ@�����6�3�>��;\p "�i������q����J�,M��:Vf��iu�� t��n�	�c�43������s�5���/�� eb&�;2�0mH���s�������_��>��鹥?���=30t�Ϟ�`g/�"޼y�������4��P��
x�!YM����P�`������PW�����+�'[*�����A8�ĺ���"LX"��zs��ꄑ\��')������qZ��I�F�ds�2���.�^���W�j]}��*A*%�H�/��B��<��I���О�\�";򊚉e� Cx�?��嫸s��/(ğ����O�g<���d���<\9�0N�$/����K�|�90��l'}���%=�\�"c��N��`���Z�X�ign;�9�UK�$�󂿋�Rk���L'�y��-����v��OF�嚊`S]������hko���L�tJ��,<��]Z��o1�0��׫Ʉ,zu�̡�9�Yߊ��_Ǐ��Bk<���-�}�?��ϰ���t6��a��Op1M1��poD���b�	�!�Ig�x��_f�lNE�l� ~��m4�b8����{_���[���~3����[O[�^��\1�s�frQ):9B@���` �jYьl:��VDN�]ʓ9]�H�f1��ZS���PzS�dQ+�;ɢ�Pu�<�H�$�9oE\ ���'��E��;QbB��0.�����mHtG{�@H{lMƉ��&Ѥ����"��{��H�ڭY�ME&����2h��3��B��捫��p�GM��ن�h��B�!��8AE���M\��T�\U�f�0���>�;�p�q��fe,<�;�UUv��� \_gt܉�8��p��i�_%�����Q��h-bO|<DV�}Coh�)C򷦞�n�9�r�&��d.~���."6���JES��Ȃӽ�eY�	�f�Ntr=��'�Ֆɥ�\4��f�s{g��v҂������X�/���E����H��s��~���}�b2��Ĝ��(98Y��z?)M�UEHc�u��H�:��PH:�Ӷ��������<y�k�Ow���ɍ�=	�������ƣF�IU�k��w!�����I�����ٸI�b|k���ۺ������{��U~��v�q��[S��vsggd`hD����^ŷ�������biy^�v��O�����`T�Wt���hE;]�8%��"ȗx�U������}$�v��ڪ���u����A$M�X;����*v��t��a�I���сn6��O;:B�;�d� �DN+b=���
��E3���:2�ޓ�|n1�d�kU@��y�$�L�Lk?�u{7��*�$����IG84|W�^Eoo�Il*�����INR�Q6-a?���!�{?OjB��#� 3����,�v^������)j�g1�����W��EJ�JƊ�a^�j��B�����^ռQ���xwv����Ε�;!aj�>^�pI��L�b��F�И <5��I�&qx\H��X^]�ӗ�057��!B�$� �\(��c�����p{}��=�{�
?��ϰ��&8��j����o甔>Ih�VD!���R:�;C�@�0܁ �vw���,o�ݹ��?���=|�͗�����޾���'���@"���l��j���t C�wN�/��D��'qD#~���Z�zx�KE��q��,r&#1L"�� p��(��4�f�O�:�&���&�"��޹,�ۣv_Zb�K�2_3��PA��d�]�-_�`Zy�ވ���H��'tNv���A�{�J�eA.B�Ti��uc����#q$Hأ�܆���i3[��o��H�־n����)G%�a��f����W9����N6wQI��@rI��@�y��e3�t���͍��#�z�~Er��8*����d�ZX��R����=Q��&��&�*v���(NVt����hOˈ��sk�,�
�<�Xȍ����d�rz��[��b�/6������ЈL*m��3q�4FD��\/��Y�W���;�bf�mˊ��w�Zw}�#��Q-�a+���f�ƖgZ�W�K��W�����W~�4�Z�mkR���6a���;>���B�ͭ$����S=7i�ɻ���Jy�$3���u���5�I{���	�����$�H�A�N՚�IyO������*����D_�w�������_�{�"�W�޻�va����?�;0�ё�8��-S��������d�@t��]f\����ӣ��2���=��k0�h��Je���=8��e(B�>��XX^��N���d67�����r^��ڎ)�z��d/Hhv|⍼��!�/+�o�.e����w6aq��+f�`ѢN�<��듍"���Κ��01	X~����6D�1cX,�|���Wx��!2�._��"L�:ulS�x��9������z-܍:D�8]7����=�X<y�����$SXD���!�V6]��r��L9�m=Ȁ�$���cJxp�<��ʖ��?�U���DV3B}��++x��ӧ���b�o���ql��I�q��%�S#���ku�(��i�s����4ӇύL.���-�|�+��888T�J_�L�2������z\9�ܺ���vlo���'�{��.'��,ǃ��.iػ<,�8*y9N*�(��� �֊*c�|A
EɎ���ik�+W�����}�w�o��h����� B�^�ɹ^%ZQ�
��$�_, �#L9Q8���o^<�	���ZTH`�5���6��2FIFh|V���{��Ϣ������T��m�_x��[@/B�u��&u>WNQ)F]z}�Ɉ4�!r�I�T��x�������0�$�Uae�����E\	FL$��{h�K���ȉI�����/0:ͯ�h%Q`����i�Y���2-H�5��)�k8aE��+����xx��A
��m�sey�K*zZk� �N@�Z��hlo�~�S0w´���MT�����+(+,���S�,�c�Y��KdNqS̽m&F��y}��@6��(��3�T��!P�V�sD��O��{Xޫ�������S��UD�N��T�/d��'k�\аA�$vӤ�{c�϶��-oҹB���������K�f�%����Aq��l��mb��v�&�lO�f�����s��"��Y�0��3����!�#Y�R�ޜ�����w� �\�?~�>��t�M�:��|�S�Ǩ0Q)_Թ�)��7�����/Ow����:����.�-������hW?Ν�HW�����gF��4#:���C�č�71pj�\�L��0�ۃ�d�XTP�:�bIF�ǺQiI�ԅ../`v~k��s�?�>р��p�ŋ� �́�/(�M�i���������*[�Ei3&{G����� )!jjk1i>��J��!���irrRP5/��9���r��4������}i����@���.��?FkK��"���\9�k׮���QR�t�G�{��,�ܯ�@.��[*�;6��5	�O�E/d3���R�W�����I�Ɲ��<���c˦��4b'���KR��=���H	[�9�s���zF'.��*K�tm�*�o��cG}�ЙӒ<���R�Ģz�Q�!�q)c���������nʉ�
�\�.� O���h~p�
>�s�-M�������w�����]��gH6e���r?JȾB�a���!Ӥ���8!�p�����������@��B�x��/cva{���}v�����qFꑠV(�0���<�S�H�f��h���1^�L!G���k&�U���d����)�@��ɒ�դ�%]��T,�4J���2M4}���b��*#� �AI��4"�%�}����Gv���s9�t�k����8Y��K)N����� 1?sN�ԀsR�#:=^���$�)WTX%�c��r W��|��ˊ�dQΔ
���,��Z	�4t�!�� �xE�/�$�eCJ�OB����S8^߆'_F��Jޠ(rݣ	��Og��ނ��445jM�B����L�dF3�xp���e�2YpO�8��n�i�Y1�RM��Y�ݮ�Y;�0a%�o,�D�XXK3~PyOr7.n�=��)�||}6�艜h�[S��؆�M���ey�K��(f�t�;����4���ő�L�\:3�g@�"�5��ưw����Qq�'k[JR����Q�<�l~�D!�w8$�(��:�Ɨ�k&�[-�(�+"�,�)J�4����C$�U��[�A5#8ia�ح"L�=O�ni~��7~y�����������ͅ�S�������gό�lO?��^�|���caqFTq��I ����퇣iR;;t�-�H�c�g�tw|b���N�Z�prЧ"L����4V�����#;ƈ?���Ɔ�t�LɠKU�ִE�#�_~�<�L��.�>�$x�t&�����S�$i��?���eO����>�:uJp�4w�t�j�0��vvΉ$�d�*A����M|��^�}��j��E|��GhkiU<����=y�I���+hiiB���vujzB1u�B�\��EM�,��<@SCښ�������,�����A��lj�k�z5� �;���"j�\�܉�a:w}u��s%��"0�I�zbL�9ʱF�G�O��aic��ں;����^Y'=���ĮJN!�]䌯,����f��)Qc�/�}�v�Ƶ���t47 ���٩1|��]LMM`�###�~�&FN��Z��4�⠗:ꪢ�8����X���]|Riٜv6���i��!���1�N����
2������vt5����gN2:���0��W�V�^&-w���,nl`ugN
< �J��})[a�=���aw}/���J.1^��J.'��B �f
㵡ݤ�%/]�K��kN1��4�75!M��BH�����0��3y ���bEBɋ�ߜ���J�Ƃ1)cb�K%@���@ �hL�?�1M�0n\������F�RT����,���{HMc�"�)�pt}gm͚�K���E�jZ���*�q�7�˫[�*�Q�P֤,/wB���ɓBN�]�zE��a�	��ϩ[��@�;��R�;��3�W�&ZU4S�m[�B/��=	��m�RY�$�$ه���E���ʇ����Φ7?����'JM���E�r���4˄�m�^��%�"���X,�\iq����ks^v�:���q+4���忳�`��x~Y���mhZ\����4mM�Ĺ.㺲d�EI�#;�+�P �(I�!�-lΉ����9Fb���e�JN��ݨ�nUN�
Z�r��7�x�����Xd�P���\ׂ˃�����m����:��{t���٩?]�ٻ�yꔊ��SC��L&�n�{PNçNK�wy����L�=�����DSC��(�[�{��?�^,N[�����R��҂
����V7��t�_d&>C�i��ɛ?�����o|�/�r�v�:��$G'i47�"���u�Ԏ]�zE����.�s#geIȩ���ʊ �H4����F��1�䬍��z�F;Cބ9�}����Y�߾~��zx7o]Gkk3�v����k<|t_Vn��4�]����Ύ����S��\�X�uwu��E�
'���=]���{�.Xp�1�wir��L�~��J/�x<*��ql����ur��/j�m�=��ۇ�|ZI7�={���y�9�s�Ϣ��];U�}�Y$����H! L�#'x�(�8o iv���>��/bll\{vBњ9V�h���+������nmF1s���)|��g{�ZA.\��[wpzhX7�C< #� 
�2�!cyT)a����V�v$�b��?��ۈ�V{'�|���y9�I"��hFiҒ�!�	�� ��\jO]�>>����I��<�d��(L��-���>E{�Q�A�oRG�c�mNݹ"�Gvt�$nF���<�}4c�H�a�(�Z<�i�Rߨi5�i��k��R��.'$)R�����`�a�6l�vwT����s��i���Ʀ�cQ�77#���^��[0P=B���H',�
`mGҭ��ul����>��Ϊc�mͨ�h5�v��a�)t��"�-!D9_����%��Y
�G�jѩ��:�%����c�Y8������I��<p6>$a�J4
0�}r�Ss�Bl�����r�"\�A����n�ڃ����,C�lN�&޷$։�a���GV4eK���Yp�Z��֟��.���O�k��X�j�X�h{��n��Ւo�&��?^�,��b�x�qn֋6����������j ��0�9�>[�d���д�K�i?o��4݄�e)��e��}D ���{AE��0�~7�=�u4"ܘ�I5o�0�U�Y�����k8����F�,ǹ�p{}×�m]�k)���ޥ7����w�p4e5�*��������w2�Pr:��8���G�OJBD��x$����C���.r����=�bq4�����͐8�E3NMarl�����"q��t��=j����M�!H䃮�v�?~�P����]8�?$�����S8�~��w�81vf�����M��@�f��Ό��\I̊�T|	���?��q�)n{S�}��\�&�RWG'v�����E������G�T������cܿ�5�ǩ�(��C��8�޸��/�:8�Y���}]�x=�Z�����Q��1L�%���gR�դPkʋ�7*'�S}�r4���VV�lv�.�O��E-���>4ExzjgϏ*6���;�Mj�I/�?a)�[�3�[0:%"E�sr�b���
:���2&'�������a1�����틗��۷��Ձ�I
��*c�pr�A?�^��"L��lN?�0^0B���.'v�y���`���ۻ�Eb�m��a\F���R�S��n��$����|�ɖ,��HQ{M����#��v{]H
X�ٔ3�u�m[="�L��R�L�Xu� ,�r�ˊIkL.r��*I�d5���;�(�g�"o�9}x(*Q ��i_J4��5�|,��V9KL��kcaJ�M���̞��P�csu���ƶaI�)��!�ԠX���&��t&"I�>�%�[�&��x�EӠ�����,V����F='����&Է��8ړ� S���Q�=���&<,�$8�&e�W[��	xpx-�m�����M�7��XԸ�"Fw?���Ei�U���V�䈐�)NڗѲX���)n�,�=d3�9Mʷ�L�B�,0[֔�4f���຀�9%Nl�������)6�t�c�dg��3��f&nQi�|��u����u����c�f�t�i�E\��Y�-/i�O�.�|�����&{Jf����Œ 	�!:d��������7��f}�bA�j0hiK���4śשF��P$f��B�E��	E`    IDAT��z�Ӎ��%������&�ev����f����/8�GS�*&��6���=z}����W��_�����޻�jz��Vv������+��c����C�L��H�8���։��3�j���I��(� -@ҿ��i�S�����!rJ]S#�O!ZW'8�y���Sx��-֗�t��5��%&}��\*�����Q�����A��������[᳣�h�w��sZ_����2���084$r�h�Pç12tZ-�����s᎕PV&s"��7jli�{�RHx��A:���QZͅ�p��Miei/���k<�}��p�������L����x����XF�tGjllE4V���^�wu�3�d���t��J��f5�~���4���!��v�P�%&w�=]��Q�{I����m=�\ 4���͕+W�=���5�g38Ȝ`veE����6n޼)�<����2�wЉ�r�"�OrP��WV�PΕx-d���tN�c�ǘ�����$�66���ԓ�p��e|��G��@�� �����ݻX��Uf1 O���E>�~Jr�j�耟��N`���,]�*%gr�m���e� q���9L�L�ū�x���Ѱ
f"QC��?����}��S�R��I�(�a�#�|G���'3�4�u	$�!��S�Ā�
�a��3d��C	yr�`�G&�|*-�4%54���I{e�r�lV�d-u��X=��ܨ�_K+��Xk�H�N�����=<|KE���X3��E�ϋ�)�y�d�7�4��T��^~�,�r�Q%Y�ij�`�m,�B�E���f1ɨ��-1Q�)���f$Y�i�i�Ś�TIj")*���+]@~�'˛`A���j���?w�d%90<��x�Z$-Ky��V��=�_����,���Hy3
Z�e�N�~���D9�h9jY���U��>�R/bF�a/[���az���*��M>�	�9�\r��_��_��0��ڃZ�!k55�lh[�dO�r2s��l�zn��S�!��M��:l"�c��EA���KKI��X��r�ˆt�"̿�jQ�y|	��)cqK"��p���B���C��@}_'�}m�6D��u�"̮H,p	�)�t�}�9�{��.(�.��%�_��v�������.�����������~����[�|�SoQ��$�h�o�P�0:�;��Ҧ}�DՄ�j� r*bܗ�����E�I/��_����v�F誳�����i�ќ�$������D.}bE�uI~�������+�ya�9{���*&;��Z�%Wb���T�澗���ޞ��\��3g�h��̄������I�0IF�`mgOE��F88<������o`�o G�x��%={��S=�y���ڱ�0�ׯ����o�Q�&��Ճ��A4�4�!��P�S&���W:���t�LL����tQQfG�M����8���S�Z'���|>�s�#�v}c�8�8'G���e�/����5���iϻ�Ej���+h��0�JE6���4�n�p��hFS��_�T����7�h�K��VVְ�L��*��v��q��%|r�&�:ڐ?:���8��w�3bԓ���7��A��X ��prx���!tvw!�!�r`�����>vK���CwK'�t��G�^1������3LNO���$\��S��d�P����n�N������&���=�{�D��K��~�G+�x0�D8�x ����M�-D�J&[��/�&�?j��Z*)��
���&goG�����T�5��c�$G[Q���i��IJHmdY�	�ӈ��m&g����a  ;?��R'GZ�:����(��soG�qK{�vĜ4x8�!Ɏ�i��$���BW,�|(y��V/lmbfm�;pFC��4 �� x?S)��0�1,&
Q62��"�Zބ;WB�hz�"��0�b�]:w���!����+C[$���">^��*���[
S�x�Y�.����=���ԣ�U^󖇾�V���ӆ���ELa���\(�g:c��1�؁&aH��,Δ~�@��Bݹ��}�~��q��b���<5������Ţj+$� sW�=6'�v����of��wr*��P<y����W�Җ#I�|��ߖ@);�<���9��T���i��csXd��a7��q��`K=�mI8�Ȼ�(��ɠ�3��I��6;����"L� S�x�9h�'��$���\��~�N���ğ���j��YܗZExz�L&:[�0�s
�}��jL4���h�OtI������a
�޾�-�a\�zݽ=""���bsu�h�7vL��-��`�\�JAa�4��P�b,�_�f6�ٳ�p��9�݃C��j�(4�E��/��g�������;w�4�a������E�+p�9V&MH��?�w�"Q�nqwL[��#畒42xG��x��<|���~\�y�������������?W&%%�$kjlFo� z��u���_��ي~Ɲ--��V�<#��޼$b<�9�K8�?����v��F� sr"�����D�
���&f&d*B���ʲn�Ʀf�|���t0
������b�xPܸuK�$��<��D+j�]&�C{O�����h$a�e5��B�����$�D�������wcX���A{��yܹr����X^���$f���/�$�q��p{��5,�G���DK[������z���`�v�p"
���CE��а���r���x;�
�K�Cn�����B�[��Ox}����8ȥ���[$�E����Ǉ0X�AD��$�\��T������*)�,yz�uX2�TDJ�� ��,��"\��]�͂~��O���׃��6�g�4���Ʌ����4%�/i�F���\^j3� ��HPb��$"���9��9�7��`X&�*���O*?��:>_��f3¯���#�y�A������d?����
^�� ���*�� GЇT1��ם�G���	��Ȃ�I�rY�0q����ו�Md��/'B2�y�R�H�X�qܣ��i�B�4�4�
�
 ��*��NSV����@������h�]�(�f����|~�,₣?9�u���'�ł�_��ω�E��y�D*N���!϶�|��R��<!�!�N\D�8�(1`�\�b��>ɶ�鵠mU�x�:�=l�'|�l��Ž�=m�\!۞υ�W8���I]f/V#`� fd\$�)���4 2ɟ�ǲ]ɢg���
~��"�&� r�����Ei�U����p����B��BK,z�+^��)���˯&��luw4��"��š��K�3x��!&߾Rf>���l�BC�a�X|��$���vaso+�;x>����r,���(g�l���m�-/aiv�Ô�ԭ�l��"	���	�MM�g�P!�����)/@�.]AgW�)��ct䚞�D(CcS����g039�s��	�li�c'pd�l3�������ޑ|�$�`,��8��vgt)�p�>�u[�	=H9a�p���On���+����۷H��$��ȽK<V����ho��ޚ�!�=__��/_����7lGo��N����$�r�0==+�p{k���6���l_�>^��&�W�^����"i���FE���蒼�TA�ZV��<tnݹ�+�.K�q@�)-3��w�{d��R�HC�����UCt1{#�qDNU�[_Y���*�6�dzn` �=]��֗����o���+E�q���ݭϑ����u���h�^���h^���:��n�=nl�2���slJ6�tG/.�9��b;X�X���8&��tpW�ܮ@�9]u�*�_�n�㼞V���\�0��"��j�w���&���)3��*�f�01ϖY���0�er���q�)�6�|�I�ah���DB���v�w�����H�p�{,�o���8^��D�l�r�;I�>5AƓ����~��-�&�
����3f	n��^ēI����g�g�Ƹ�&�(Q����>���9f{G�%�\�B�
X����Ζ�z�d\�'l�)���V�|&ސ��,�H��=���
�'"���C��L�ܝ�7p���*|VX�>���=SH���t�q���U�C>��:���*xOª*-L{UKw/(�֝N�y��?�A���5�lwmj��qﴜ��Z3��"Rytk�H��1r@��eA&���ME�E��4����e3��b�=QL�%���ޛ��G��ʚ>}~�>�"�dmsӰ�-5��of���>������gaN�D")��ޚDTj�y�XZ`��V��D��~����-�cJ���>'iZ�)�I	_���j��,���r~
��"JQrn�!�"�!G�����j�������WĈ�{
!/�>�ےl�����ǫ��*����J;����+�'��tm��}>������y�{�c��k'�"|��4%�e��u錈��	�?[��*¯������C�֝���F4�,�Lc��;LOLc���]>Y�-�2��EBF/�}���}>}H,v�����c�͋��B{�jEE�;,^0�nWr���ԇ��E`ymU���G)��0����l�锜�X����'L�Y�}���n��`_?����;|��>�{q���ho�����^����gG����444�.ـ��f��Q�?H�����S�]�������ҔN؟d�����Exwka�/�.,/.!���p��(��u���L�9	��������� �g�Q6�T��������yD�as�}0o&�,�,�r�"ϔ/MB�|1�tG	��#�Q�ɀ�yEř�L�.?�?�Q������mAO[3j��V��Sc��ڕ��WؘQ�{|�����u�����|p2@� ������fu+^�^��cOyʡj��+ofᅧ�U�z1#{fe׌��w|m_]��RKԁM��9g���|߃��$�(6������y�����P�����I���٤O�R����Ţq�tf����;�}P�U��¬��x���)UIy�-y*?��>�q�ͅ�.j}w����¬*Mkr��1�T�Kj��+I�ԕ���GͿڒ�d �Q�!&$%Q|	1��LQn6<��+%7f0�#պ�IG�P��̱cf�����Y9�-���rfN�''�lfNK�ht����&�Lp:,5I$�L���=y4�)��h~s�uT0H�4�V��I�����)�5b��-�k��g��2l�\|#�we�eT�E�^�hvg][��R1��J�ݶ߅M�6fB�A��1������9e�a�a6�F��$|���u�u#_���g~ڇ���+ޙB�*W��H�j�{Z��w��C�I��o��қ�v�.>�R@�BJI���k��m��iIU$�FX�ts#8��o�]	�0O�;�J��#ސ�9��7�ȉ�d��1q��b��C��L�ތ{��rnl��M&S�י�y}$Rn.��o�\�h��x�)�L�,��܀�9e�ߋ��L���Iq�t;�]�f�0�ɡ��bn� ����dU��+���!@�m�_����ão�X��^���#a��n�w;�s&'�yjN�B����Hļ��t�#�������/?�v������u�{pPׯ]ӹ��5=�B�n�G������Sg���mO8,)����Jfȋ��nn���d���J���L�\*����=kk��7/
�b~��Ψ+�J��"���4�dHb�c��ۯ�qYi��d����F��A_ʍH�cxi��ʊ�g�zM�g�����ukgυ���O�=���V��T.���s��[o����u�����{?uRo���&Ɖ�[ѷw��G��Pk>{�F���BJB�]6o��I���W.[�EA~��;L>���ޞ౉�:����={aC�y5��{��o���#�n�0���1�{��)������n,p"���49;���A�:w�$��t�t��5x,"�Ż�Dt"���fKl�Rls:4	�2�_x,�0�@sL�ݙ�����?���VV׃$�����EK�o4;0�=��.��+8����[oj����
���z����7��9�Oͼ��涚�e�q]=}�S�$��W�je��=&B&zB*�ʇ�R��]5���}�`@��n� L�V;�z�R9 ��h%o�Q�n8y�V>���Ο8�s�z��̠���w6����g�����f���T�����:�P�h�L�% ʞ����U��Q$�)	����}��	���:���
2F
<�����u|���뛛Z�\�V�l��xL�\V
qWF�TB͚�*{�k5�Y+i��0瀢��uBG@Z���-���dS�	�	�N�"��$t��y�}�Ξ8��L��4ﳢ��WY���	�}0�5�uC�ryu)�\�F��杽}�����N��Т��?��u�A�x�ϮTpk6-���R� ����6�*�{
����l:�"�/�R,r�?yd]�/��O�]:�,nz��0�I���`�ơ�!|��~�@� ��֜�W������@��������Y��%KPu�@��)�|�����a�%ց�^� $)��}�S�:oh6��{�����4[��NBje▩��`]��"�;�Y_�}|�[^��� �>�/��h���_������0	������W$JxoBf�z�5;f=�|��>�DO�S,����"@?��4��#[8��0�:���O,�r����-�l+���?��wj�����7_~����J�/�|������D���d�{|v��q�07��{��\���tT���}�L����B�-�"Y�t�]łS�p¢�{����Q��(ڷ�l|�HE`��y-��U_�K7��������U�O>�Lc���	���hskUw�|�_~��,-p��NI�s�������N�0��y��i��PW.�O������:~�68W���w����MrA����絻��SgOy�!���+--/k�Z$Dm��Z�� ��2e����5��ę��N�j��RX�J#�vt�m.]����� ~��{�fArHY���G��4P.�
������V�4F��8!�Xx���t9$x�pez
���i��i�	�j��aw�ӣ�~�M3�hz~F�^�,h�BS�[�����>�LLʥlPQiմ�����e<�qH��嚶���j�����M�g����6�@*C�%��$�@ZV.WT� )�ҩ�o��-&U�4�Ng������JH��6���fϿ��MKw��]�y�IE�� ��p�ZǊ�(�hĆ8�C�;�t6erEx��1u���liuwWS�nn��%m�l��%"u���q���^�k��L��q�!�lZ�Bg]�|�nӅ�ʞ�`w��U˞��-0�ᕗ3�s�6���h��ճ�ލ�t�w�.�+�ы}E��sav�m3�9��Z�{)mm���/Ι���<�^�{�;��uja��C����ޒ?b�q3~	�������A|���tZ��>P_O�'B����-ܔ�O�����,������Sk�m@#鄛O���7i6h�{��X����k���;l�)�1'ja ��Ղ��C�N��a�K���!{�P�.@�{W�N���#:���=�ł���\S�� �v����V� 9g(�L�9�����5���/4����LDʧ,���A��I�8o9g�F���Wq��9,����r��?10���,Ĭ����o���73+�W�.¯��d��ɗO����1;a�|8�����w��-��{�{H,��"��!/����Qm�[�D������Ą!���W��n߾e}!�&đ-�N�@붵�J�XHG���_�4���f2���z=ة��1�P�)d8`9��Cχ�
���B����pzt��q�=���"7���Z������>x�-���M�t������ǎ2<::n��ѱ#A���>��C�,/��m&�egΎ�N�fV��Þ�Ϝ<eO����2�[�0�xK�;vn2R��2�V*&y�=�f�t�v�ӯ^��ύ=��=O8��`��?|D����ʾHu�)쎶Cʀ�G&R&tϬ](*c|���r�    IDAT2�v�y/@,� �"�
V�!��_���C�@��ޮ��_~���U��9d�2�N4�	8��Z6ץc�Nh��1E�)'(�+5�/��/Wй��z���n.k���N>׷�51r:���s�g� Ԁ6��1� g6�v�F>�7��  �t"�m�C��MFv�P�����Zq`<z�0�'��zS��y�������^U`չ��yEK����s:�_͖ʭ�Ӝ����
9̚u��֐�b�p WV�`��0�x��@����U� ��Jɤ*�J�[��M���{��i�fyc��,Z�H*�|k���LC���/2C�&�!1�F��nԵT�1�L�:E�C��Z��.�nj��+��c�f��:P� �t+�7�_��o�Й��� ��.���n�3Y�4�;���Ƚ�L���f���QЦ�ʥ]�nnx�\��P������4�@�L��	�n�~�={�/'�RsqE�<3�2���x^�l�3�׋�)��@��,���t�ۻ�d'ܕuscr �0����N�)E:�P_W�FF�}ZY^����?��u2��&N�Iޥv,S�Ʊ�Lx�3^(>��(�|p5�%f|r��#F�c��ɇ׍i��49�WV�}]���ĭ���>�㜱�h��\�yC��^-����[_j����DX���n\�[-w`���W�����I8W&SZ!�g�{�{������3�(�͝�.�{��߼ZZq�v���AS�s�t��o�ͭ/�����U2W:���:��vVμ' �Yҫ�yͭ�*�ݣ2iF-��.b3���܌>��}u�k�>��Qw�3s�
D=�T+{
GT)��I!a�'0�F�Kn�:�}���\��@β�6�r�e�s84��P�Siǰ���v+ѕv�8�f4�@/HM((ཱུMқ�����@޳���`�O?�Lc'-Q::vD��|��~���I�IDS� ��ӊ�c����q�"�,ө�'t��qO��~s�$����!�
,W�}>��g1��K�c!����W��2I�/=��ԫ�9O(K�~��ι���=j�04:Oj,�|>�aGNp�xCw�4�.�ن���,�B���a)�5+k5$�E�Ц�@c��4�-	� <cyQw���g�/��F�m<��N���)����[�����S?y»���5���6�5�7��g.���ok�حrs_�=��|�;��s!O�}rtB��V0��\�Z��E�f����������Y�6} X��E0UT�%KX�P�a��l�c���7��4�hl�OG��4:��Fmؽ��,hiv^k+�����B�a���.E)L�D�F��)�LCe��X8��K�FF��L�=7���|�39K�q�d��(ՕS���ؿ��7q�p((�)�-�4�\;l+�Ʉ���R�=�:�$�\F����ǖw���4\#���(Zj�<��ꆖ_L+\�aR��VD�FX7.\����a�p����f���:b4�ɔr�`o��l��˴W������� I'&&���֗����fi�|&l806��8��0CQ78gн�c~���f��ٗ_�;��0��M$,;Z�b�쳗/��C
v��CM�ΘD	zǤ�����=���%E�)aH�Já��$�����B<P��H��F�47���h4���Ͼ�A]"����(Fcb��t&(��.��"�:��v�`$��Ҹ2F�`�CFc
��� ݯ��������c��t������Q7)�7<7��w>�����Z)��wni����H[�l0p4E��N������m�E��� �B$a�����pbp��o_o�ON���[�r����jq�rW_�]���M�v]K�szp��[��e_(j)��c'�&����"�4 �V��=~�R�dJ��\���?йsgm�����O?��~�����b��1�ϫ��Z�QQ�������w�>~ҍ:6~�M�_���σC�8o*\?�G;{��]��L�Ň��v}G��3��=0�z����G�e���U��\�9������Kk+z��~������ѱa�n�蛻_��_�º\v��rC��*�f�7+-��G�F�-�/�?V��O�S��/�����+w��9;p�!�� ����2���L3 �
��P<���}~�Yߵ���Ke�,/;F��b`xXgO����$�`M���v' ��0���	,
*)��pL�AM��_����T��64��G��T<b[A�W���T�Z��"�Ӡ�KA1���]4�fXO���P�6�17�d��n���w._���yGC����*���=}���>$i`Y�u�	鄶'�ֿB����t,=@.ܯ�{w���#R+H����<:~�!��.���[
�+
ժ�\�HT��.?�Ѿ�ND��L2+s�\[7�]L�:i3�A"nb�QwpE��K�83(�r��!����ףQȓ٠A�U	Sh�����Q.�"<xtT��C���R��Ǝ�VW��KLX����;F2V��0;ڐtO�(慬�=EO�[��wE��F%`�c|adS{�Zx>e�!�h�*�0M�q�7.\�o����g�S@��������^���T������/P7�l������DhqzZ+�s���Z�n��>���M)İ(H@Ս>�g����$�.�_߾�$6t�>S!�K��ď��Pw�f��Z��@Buc����夝ǐ|�D�'�f�G���xn3	��i�Ȩ�<d����=�
�$+�����ps�b�Iӂ��[o�冔�t�իW^=J�(����g
�^�t28�0�$���=A�|�, �r�(n����s��d8o8�v��922������v�Q+y'��n��
Lt�!�S�5E�Y�I��mCT!u��T����ha��3	��۟^����^\�T��wWtpP��̔�|��j�J�5�5�ѱ�q��h{�D��x�hP�q��E�ƭ+%��/��/tbb\����o߹�{h{�`υ3�(���:�3EY{�����t�6��K�����������~���#Q��?뼙��Y��Z�{U�S�@���H"��5:0�j��'�
�9dӅB:��$��6:��~�;�=��7���#��\��o��/���A��U*5CVhJ+��JX���ݫT:��hH�į��ޟ|�\��ZZY�t�G����R|�0�1�o5mx�ɍJ1O@�ù(���0!�W/����?q�M?(�h����|a��|P؟|}:m��t4�l,���kS ` K�Ч���;t��т�gf� �*�vN ��jے���ϞjqiY���FG�[5+��٘�7x�@���@&R���wT�.���q�{����f��{���[_���\�h���i��kuw��%e���{�dʓ,�9�Y�_+OK����A�d뻃C�Z�	2�Y_Q�YV�ZU��PO"���]=wFC=����AC�3Z��5<
�S]:k�{_���jM���ql�TY��bq�q}�V!�1�`��I�@_�z���MaNS�����KUO��V���w��	�����]t@z�&���7z�G;5
�-F��/�o�ؕ�� ���|e���Y��]}��ȿ:EZP���7�hv�4k���c*��m��,�p��UZ��3�s���MP*0�q��@fv�H#��ɉq��2z�⹦�>�;z⤛�|h���j����PA:����546�d���W��ͷ��oy�D��=�H�d���;y���8�������B&����\���W��&0�m�@��/��@3����N�O�=��|���ڕ+N���75�B�S/����:��P�	y������~Y/^<��;ap��&M�w���J�z�)#��lh
?�p�XPO�ǲ�/��b�Y�@��=h�	���67\�9GG�G\�3��ڏ���4���m�鉰-kA�@?8_�02�{��~��J.�T>��l6������o��O�������O��/S�K�u�u���y��BMM>�>������V���ѩ	�1�1"���ۖ&�ե������\��w��|���J�ǎjd`H{;�&���\S�N�"N'�D+VWع�U�onn2����F|�Z��C��i���1l�l9P��n��8t�A��70dx3],(�M���W��7 �3'4R��;m������-/���g���ub��{���j��������b��ۭՕ5��<��cZe܈8Ds�9j�򅜻�C�	t��<�ߑ��g��d �Jӓ\����h��M�
ˬ�6,�|����Z��>Ϟ=k��}P_Ө 4���D�.Q(8;�T{�v�œ�G"<k(�L
��kGJ3@!�=	��T��)�N�\H��f��&E�.�`@]�EDLV�J��Y��ĕ!Sx���z@>g1��}��7�[�S�����������~�i,�0��^sOB4a��y���"���
bX����)��-۲5@m�f�F"�e�;�^w~nV�uEu�J%��5���0zTg�G̈́N'qM�jvzJ˳3����29�RI7��XB;�������,t+��+�J����m;���NG���Lv\�T6m�T�?������JZA�ҕW�+�D��l_��ł!n��/-�y�U=�ƀU��DL�B�C5��d�V6�DwAIHZ���jf6�خ�������K��t�tU�Z� A2���Ķ��W�J�RM������\��ǹ�?��?W��[��_qQ���X[�d��8�9|�˛[�x�Ό�k��G��f�����S�d�2~��0M?����J>wےG��щ�8yR��^=z��)lw�����=8J4 p":,硱Qb��Td�:z�F��+��krf��Z��D�DR�0Lb��2�b�W�"��J��ȄΝ:�b��ɓ��ȥ�I8��NOz���-��x����KW���W�8������ܢW��CZ^Y4�ȳ���a��������}�4{�8�O��Y��/����g~��݆��_z�� �n<w|.x���s���?��@p)¿xG/6����"S-"U#d\C��ј'��"̔�c�z>��O<�����G}�՟���۟���'?5�|Bp4lP�*E��ݯ-S����j����1�w��8!#ӑ�^� 9n�?|��3�Σ'`�֜�����g��@���bR �o�_LX�t�� .F���#J��N\�P�($�< ����`�#:KrD#�v�˚�J1br�Wi����m��|4�l!�ѩ�K��6.웸�a�S�[h=9��a7�>�G}d������2J�]ݻW��/�_3O'N��ܬ��ww����=�Y9��U��Φ��z>_י�Iv��'��v�	l�`��4���ú������>¤��HԨ:k���`.�P���0nz�W4zd���p��IH�=X�����AX�X�7r1�c�U�0��ް�?�JK���o���	�֘��V�� #ܣJUC������i�[A�@.���p%h��� �f��K�l��ҕ��FwC����bU���l��="Л�m_�ti~��wM�b?��}�$�6�h�W]�)������h�X�0��P�h{sM�k+��n+�fMx���tJ'`w�+�EZM�R���e�6w����O&����,8�N���JE�D[��khX�B���x���ǰ��#�>VSq#W�h�ˮR���j]���RŢ���O�M����jc/�6��x�_��i��0̻����U��V8��/�]T��e'8���B���xi��N ٭�݀�[iXB�0=㰅�"����╆Ch޼vUo^y݇/��>�PSK�ޟ^{�M�ym�&�χ�9g�5de(�}�:c�Х��i={���4X&���"A�7�5"#[6�����Ǖ��֣��t��}���vD�|�g�`�10��Y���0:\�,<��Y?��S'�Y���;��ޱ1
E�f�6��b�k,��l�ΌOxG���ӧ�{��w�4K0���q,��"8�� ��N��勯9:tceն�����1P��	�����=8����9�0c�j���MG��� ]�#��$�Iu[�tJg/����q� < �����y��7�������{��)��kG���7��Z�Y橨Mb(­p�;/j�+&b�a�?�I�Ts���0f��Yg
���������?{�ދg?���"|��Ew�/&�����Nn��{��:꜆���+�A�\�jrսG��rnA�%�0�29��'?�ٓ'��]� ��xD��:c�꽳�t�����t�̴�~_m�w����65?7�����(�,����m��$5td�nLRa�2��t���V����B":4�pf-�՚ai|��I��7��,=�{��޽~S?��}?��Ү���V����7�3$�4~�@x�}�(�a�M��h�C:�Zϡ'�'�cO��Z4���,Ԯ���0��&c�E�]3qqѐ���]9%��A�I����$g�5Fb�/�8��:�1�i�I�I*M��u�Rv�1#�>��f�b
e�0]�]34j{B2^���/HH��(u���Z��I��s;dM�5�U�z���CC��{FD�A(�˱��L���4����������s&
'�e����C!��{f��,.�L������Jő��݊vO�y�E�mo۾@�r�� �B>D3��H��X��D���P\#ٴٿ�J�Ȕ���̔�����z`�g2>H1�	�c݄�\��ΞV������1��m4����im--�'�D\�X�~N�x�(H(���qUk-픫Z�+yF�Ո�L�Z�߱�E�~r���ܰ���'9t|����Ąv�+/���V����T\5��T��\hf��m�nkm#�P.���R�Y���NÄ~r E��ɓ���z��5'O���Ň����'_;��gO*_,hku]�dq�]]\P}wO�O��XO�F�=�OjciIs�AXM&ig�C�w
�����517��ޖ{���ѣn�(�S�_X�N�
Î��h��u��[C�G]��d�f���D���O�SA~4��מ"܎��	$>��vX�Hʓc��i�f?z8��h�Pn6����iV&k�
(�@������'�D����Ea� x5GF��̡�ý���ԉ�Zr�S�!��10�A*@g,���}�C�eryg_){�75�J�[�����O~�S쩡�ܿ���u��j��<,��0N�<�LÒ���+�	7ˤfE�����cП��~,����Yt��ǭO޾������_� �$|����$��<����-��]D�=���'t|l�&��8���\.�����sb�Ly?��! W/���#C�c�H��~��"�(8��Չ Cg2Uy��k@�bQ�T}��LNiueŖ��6>P�����	�ᘬ�߼a�7n�q3])�/�5�0g{�$4�o �"�Ih%�th7>pK�t���!�	y��楫�˟��>�RyG��>�����4����m�]�����c�}���cZo2��f��_ڱ
2�fgB�:�+�����!K4��Qh����tT�W<���I�a�)�ceB�,n���x�;\�%��L�D9D\�H��C��'1� ��_w���V#�'S��ŕ�� ���*�D��x���GzttpD�LỨ6^�	1����p�H��!�Q�L
m'���`���F��m˯�U��g��}���ddavF[˫��ܴ�t��ם}%B����S���Zo�Ϗ���8�51� qh7��/)Skh$����ɘ�q
K{�[z9��{s�h��nC�A�c*�BZ����Ɩ�ї��{xX=����+ssZ���>�XD�����9�/Ř\�jG�H)�ɫ\kk}w_s�kj���$��ޮV�ƚ�kjC&1�HG}��\y(�UP����АR}E���c���Q,�Q,���ț�Z��-y� `[;���xͯ--����v�2�ׅ\&o���g��7o�ʅ׼�@W����Z�&�i����#C�p�5[������t���CC^?w^���䴿�n�0Sr46B����'M?��l+f    IDAT�:� �	�qi���}>�J34o[�L�l3�?�< �U+V%�|�. E���8rtL�N�u,�a�ta85&a��@��M�,\��jݙ��?��g�)�L����zxﾑ5,w+�&�i�����	s:��Y��ft��Ο=�� ,@ӿ���b.)�|����(I�|_�@�+�G����`�0���y?�{`��x��{&��u)�=�s�q��--�3�7����O�7:��PS��wKS{A�$��j+<:g8M���ݶ=�a&a�z�fK}���C��?�o��̟���E8_(����t��%%#=zxO��!E���mr�/�SO�G'Ə��7,����bR����d�v��o�ʵ�z��t���Jň�r��O�b�%S����6j&���s��VJ���鼝���\˯��*�2ᰊ�L�	2ɚ�^V*���#�����ßW!ݝ~��OjfmU�ق]���
����5m� F~)�Z= @Db�
�m��o�����G�s̓��������8����Q�����4�M�&Q�T�ʏ�LN���Rؙv���(A<���BM3!L��N(�c=�pg�Ŏ���	�μ��yL�%�F��!
<L,]�3��{HW.t��2		�7M� ���20��a��ZM�m\:�����C6�o�[j�L.�؝�������5������Ⱦt��f T,�gj
�4�8/򨠭b�j~uV/w�$�4��G��/�4����9�&iʀ����@ɠ H�؃��Mn��k� �*i �[�p�!^�}�PW*����=����Sw<�L<�f�jr�����]�˽���V;�(���Z����֞6Ke%����*���i�]]Q����\N�=E� mˤݨ2Ѳ�!�;�+�DT�Ξ��T�Q����,��& �<1n ���&�d�i4l9R#U��㾂
cG��S~xH�ޢR�E�!i���LИ`�u���^���>��zr��;{�ޠq<�pT֥�g�+�a�_�[=�|n2SW�n�wӶ���^��4�:�ݣ������'4�7��tF[K���㨗]�!e�����V#0��Ou[�ۖw���8&8�664��dLo��{x~�ݽ���5;�5ba�5���Ő:�9R�F����׫��9=x�PO�&Ռ��s��l��K��u�B��9͕�t��K�;ȞO?�� � �'�e`�?����E�Ƞ*�����uI�������4<�AZRZ�ˆ��3X�g�U�3Ӿ�![�d�i�'�7��o\�J�����ŵ�V7ֽWF?�D�dBGG�����9��p[���+��]��AC�D�E��0~�V_���� CP�x���J�Mx'o�՛�~1���O���E����������k�|A׮������N�鳇�}�/�ww�g����z7�"$�Z�@_Q=��hz��f!il�(��jys�E�ĩ�z�ݷu��9=}�Xw��ѷ���.t;'�����'�p-gJ���0���:H?A��n��X�ts��w�=���F�$����0#�٩�#7�m�t��C}���6C-0��?�f15�{kqE��˦���aBR"����^��;�o�'�`ȅ�:����TK+��f�}��06
�c.n��V@��<�6����=g"�HR@�A�8}�8Q2��S�5��4R	�Y�t`��r> lx�βS�76ִ���Z�b�"�j�zlsm��k���XT��>}$���:0�m>7����=uI�	�� ��@s��?$��&�����@G��u��Qvt&a&�ΐz(q��ަ]����� Ӊ*���R�%L�"@輾���)�n$<5lhn�V�W�����ֶZ��z�q]+U��t�7���LT�;K����3P(8�Z͚%C��R���j��׉��a��A[���6����1�A�
���=LۻZ����Ύ�p�I��u��UcoW�����z4�WTw.m;Y$%�u���"�{�9��W֋�ymV�~6�Z�����bj[�n�y/������OQ�����U��c��W��w�Q���!�i C�HV!�)j�}�n{j[ZXԃo�hciū V�Z1�ۺx��S���YkW�w�R�>������}z��w���K�\���e	U�6\p=�B�P�+�mY�� ��:�0˗���\H�[��Z�F�|8��jE5������޽{Z�[tW�����f������(W����An��������B:d���Meu��]���'a�Y�ܗ�����	N���9�-$����m[Qbt��iO��ӯ\�==�,�i�������B#d�z	����ߐ�G�,P7��>���3.-zEg�~�1�$��Р�g��>C���~�����{�S�'wV�A�p�IS�M�eP#�C�!������e"�m%���t������৯���_���ƷϞ�����kx_�|M�x�Iӯ^����mֱ��a8�wdxT'������v7�T��4zd@�B��%���/49;�H&�ͽ�ַw��;7�����B:���?|�����-�ƺ?BÝ�ޕL��'LMm
#�(
ց�Hd񾰯XЉ�����hbd��0h/��@rbǐ�e,��&����������sݞ��|��]8���@;����VU^߰-�<@��X�M Gyk�E�G|���N+��zzy9�\���ޙA���G*ż��^.��d:��ń��D��	K8���q�r@-i`��L��L��3Iy�.7bF/0�H�Ę1�m8N2��1�7�����<��9����NE2k��ίL����=]�!�P�׀�5�7�*�'��-�x8x�h(ju�=�60�ggw���c`b��N8�y:����,&�8�)��iH�"���:٣b�f��H$��������t
��Е�LM;_x�ù�^�+~-�����r����q�bW
�a�tǿ�C�Ol8��U�W^H$5V�ֱ�nP�����uF�ݴ�B_��2�D8��NC�S��fG�Yq��J���RJDv���Ry_=鄎�i��K�LRI�1�گ���(��R���v���K���/iO�@�J� �;��0�MpY_N�w�=TH+;<��谆ϞR~�O��~E�)K���~�#q�"+�M*�2@�}���z������Kj�*
�=a�Z���ɓ�~��n�������w���=���.��n���.�=}����0AX��5�!�4Ec�����F�Ϯ�D�s�6�����A���dj���1_
6��"$����w���²6V7�s��
$bf������O&u��)��x��e<HB����ZѠ s)VfX��m���t��(���W-A����W_�]����R)s'Pl�H16�N{��3=��Y^X�Nr䦰��j��y��4)W<鮮,��}�^X#OCR��f��Lkgg�(��ҒM����@w�iOL��	�2R�~�����qU�!���z����v=�	c�d�p��3,q��^G��دyw�QG*V� ��\��b�����{������z9;���k�����+&j,�����[���O���LiM���i]<s��J�`1X]�G� �|N/gf4���h6�խ-��y}�����;7�}��W���7�u箶I� �f�pe;g������)��a�z�i���4Uw.�������.��
*��}W� =�ܣ�E�oW�n���+=�}����z\�P9�4)�S0�PD�VH;K�Z����~U�(QL��@�SN��,�������S��1z��x�O*�3R,ң蠁sv�����.�-��I	�SO{�;�0��1_���f1i˻m�r��U� ����g�+���Ç�ꛯbP��Q"���@6�X9�����OCч,��	�Ə6���LR(��ց�ÇV��������B����r@9q��?�ǎ�sz��L+h2�A��혶�{�t�I�i=���E��3B>�X0�q!M,B7�z�g���2�[�����{e�J� ��Z�G`�v�a���)@�n�����k�=��ha�eu���M$4��h8������V��_+G�Âm0�L�}�'_�����7��� ���>�<���NT���%t�H��z��&��FD��i�DxP^\{u�h�Z���f��u�Q:P�	'��<e��Qs:(�Hp2�43	Ez
�S��:y��NY�IE4 ��'KA�� ��Y����T�Ӡ���\^����\ZQ�TV�gl���N���˺��u0�����a�Ǎ�-����K����M>n��u��憹��CZs|"����J�j��C" {N����c=�=������4F3ഐ�\�,	�Wl!eu���B1c+<8دg/����ֽ����ߙR�<�X3�\"Ƀ!�A���������L����O-);�qJU4�\"a����^?{�{E�v���%��3�~?��)�N�Ja�	���z��p�� [�?t�x?�e ��W/Mf���oha}��C�C��x��������?���M*�~}�͔�<	S���0�bב(y'����Ύ�hM,jAa���~w������7�����|49�/_�-^J�3���M�u�RѨf_M��_�ޝ[���*��"S�v���Ə�����ʲػ�k5�X��D+�P�Э��u'��
�����^�����oo�y������T��F�v.�C-۝!!�7�C+ܢ���%Jf�N׋;ԏ����L�0Ѡf��L!ì>�#�4�=Qjw&���Z8�h�U�Nݧ|�9�\��J� ��icnіw��Z�����w,7߸�����:ylB�v�Lfm;[53tn"y�X$�R��*��z��$�0�.LX=�ФS���J�����<_�`꫹����5�#zd���i��S����=y�<��V�{=XݵF��?��CO�	N�^��h�aV<�<l&އvUΩ���I'�D������9���q{m[���Ɓ�T.��epV*�L���y�J���igk�D
%�0��JC��֡s�E��T'S�{'���<�C�ƶj;;j�1	��2F���3�4�� yo�b����	r���B�F��j8�'`��a�A��;Jd�ޫa`���ܬ��KZ]Yv��ԋ���KD�)���r]nL0�h���*�j��K�}] 2����JU&ڰ�ܯ����Ե�W���6�U��>���+��M\�ԙ�QO��o��2J��wbL���48q�p,�	��p���9�L�}��z�Ȅ��<��bi���FZ����b:���A���.&L��˿s�'d��#��2R�4fav��I�֎�:6��WhԘ��?T	mȣ�IP��A�g��'1�z��>��aex�Hã�p�Cr"��"$&%[�[�}�y��
�
����|��~�{UPt��#��u�TBHzr]��~���yW��.��<y�-�W�T`�y��f,g�)_C�@K2ԯ]��;��*s���3zo�q�#�?'Vl^y.�����S4��uD�D�;�jfn��3��4�\_>~x$�]_���9��d�ӿ�K=6n����Ջ�m��������	�UNy��X����Tm�<Pt��8��|�wǻ���%���~���S��jv��"�����A�z�T����o�r>-�]4z��
Yt_�6"������?ob�}Nٞ>g�n���|��n\WoO��˯�Ч_|���y����:�9 �����}����UW�����57&n��g'N�ıq���P_w�{�V�����F��X�ӕ9ݛ��\e[��k�`q��fH�xFGr�$�"�uD޵;��f�C���Z�~5;��W�E����u�؄2� *�V�(ly� v��N�
ņƣi�x�bK���.4�@����8�!�i(�����ΊL����äG1���DMn-�2���e�,�;��ɓG.�x�����F�� ���&�����	w�a`$�gZ�
&+�H^���q8�k�=����7eP1�̎�(���@8y��N�>�޾>�:������t*�C6gW#�1���_���b�fm_��0���4�6C!�+���x��h�l�ݛk���E��w��
�(l5���a�w�Hu���#��^iw��L��V*A�^���i��u O�G�E��$�گ�����-��*�}�Twv|�>�����|/5�;H��=�9�����>�%%��t��[�}E���7ʪѰ���+�ʨ�k����~U���Z�<�^S��O������@��D���HF��Τ�/(=<��cc*�����'Oͼ�U�d���|P��EѡV3@Q�9�V��`�%���{��D9��o�q#(�K���/���Y����(t��Yɰ{)F_;	՚�T�bH��5Ӂ�t�<߭C:�������R�{��Y�xe�s�(�F���ȽJQ#Y�Fx�Z�Ԍt����׍��5<<hB�/~��>�����Ҁ��xD��d�Z��!����h�L��5��M���'T
}���������ٜ�3@�=�V��5	|���3C$�(�!�	�����Tr~:g M��㍆e�7I�����3�7����W�6#�������0;Z��L�������}Mn�h�YvX�����AgܘxhȺ6T��Tu��"�u¨#��;W�|d������?�ӳ�q�z4=��^�-^��v�7�޵��
59��E��O>��O M���5��9:Jk4�Nqŵ���ì_>���ʆ�K%�{=	�u�u�vw�����Ol�M$TTIPJq��$���7e?ā�_�������E�!nM��P�� ѹS'�4#3�q!�i����̔��N��ƒ�J[Z�Y�)��j��WG{�4�3�#]=�g�#˒1�jچ=[�q���e=y�B�}F��1���[.��d�0�̫���޴�9���~��	��1�@�%�AX1Ӓn���dɻR��t�}J�h�^�] F'+P�I+���֮��L��a�p��i�\W�\��¢&_��˹iw��C��@@�H,�1`�t���z�̞�u8�P�$�t���혀�;;ndV�����冫	iG�̨X((������������m�G����҈�$�1(�%�r`�A�N#r�Tfj�}f(��ZY�h�Zj��ԫZZ]��⢶W�=7wJ���~`�!RØ���k;f�Ih�ݒ�'A�j�IKw^&o6��O��$z�R�H����n�GX���0�ȧ�&���� V�z1���͠a������zyOU�����j�X��.{��L@*��%��gsj��ڨԴ�S��ڦf�6�^���;�T� ����a�0ۈ�Ů7�T����H��o�蠺)ty� �}'�f���a�Q�AA(¤��,�
�Y�O��Q���:�/�v0�h�Jӿ�l���˗=yQh~�ѯu��CM��;W� ͱ�R���M���Z��<��)�K�>�	b�y��!v����1�C*��I�"dw3�� |<Mw
�Ѭ��k344��o��k���*E���Z���wn(�Y?�懞��X`���)��E���[vic����#ݾ}[�K�P�'�ɚh��{��l������|n/tL7xݜg\Ok�C2�N�o2�WmA�qH2eE�?�g�h�l�f* 4+˫�[Zpd�e�ɔ_���ȧf^igO�d`�<~�'�/�?���U���GS��Ji�#�d���0�u�I؞"�h(�i S��Xo�?�n�d�ON��ww?��`��ϧ��.'�Y�u��^?wI��^�L��{�����x�ؖ�y���8ݪ}9>����IB)��_��Ɩ&g���������{z��Օ��S�>����\Q._��ɤ
���c��և-�����gz�౶�6��ID���hܾ�����������OjttȨ 4S�WOug��V���+��Z!=�3�'5�=�	�M*�+�����I�l�N�����ԫ}��_i�o@�_����ƕ�F����'�ի)��v��rȲ���&g��qӅ�34;�9v-(v!w�LT�ݬ��Tx�N���    IDATA� �LL�@9@��,o�&�����0vdD�x�2����E=�L���'�h.�h��ɪ�w�T��
�:<�3�.�/�ot�uFr�q�ZMX��z�pu(�
E�G�ĉj5���9�s�6;��|�S'O�l!��5PWi���������\���\r�?;.��'a���8�G��!0�I����L���ʂ� ��*�׽�B�e5��: y��09ˑ�m���2� p3���.kv���	|ł}\/���jjonk0�ёB^]��b^��r$jL��{>L�7����Қ���L�d�Z������e�j��Ǯ�;=܁�1� B�EY���������-͐�[%���"�d=�Y�`t=�R+��A!�F�}*�Q�ȰR�J!�;��	W��S�-�l�t�;gy�&]h­�G�����nᘆrE��J����Vf�nA�{M�!�S���� Q3��s�Œ�K�%Q�L�v��
j�x��b���x���l�Yi`�O�0X���L���4�k�
�¸��<�4�@�O4��+����u�Q�I:24��ǟ�^����+X5ID�\;Hj��}�.u��6/�z�τ�/_X��5�{����9�h�Z-�/ہ ME��f�05鰰� �r�}8Pat���`R��ݰw�� 	��3ל���߷'|��L���E&:��+�׏~�#;}����Gv�Zm�8�S�1�:��Z��9�
��:����8�i^���;Gs����ޏ_�ɋ����'��|jn�J<�N�MݸxU�dJS�^���;��G�R�3gu��5�)�ʁ+��%K�!�� �.����K���u��s�I���[�ľ�+����g&�����ku�ƛ6����J�@Q��
i�T�_~����w�:e���iػ�.�����u�����˺x�Lp=	����n���G�7�B�LT��M-�l�J���˺|���a,�}p�)��T\�$]�h���`ls��([.�����k={�ĻI��}O"�9��� �&5q���9��5��_���]��I ����C��[��Δ����/���A�N���'Փ*�M����>��w����ړ�[8I{�C�Ý�!,�`��v�@���6���I���M8�� ����c�IQ��z[���f[�qN�� �->�ǵ�*���O9�4_��5 ��Ҵ0�atv��)����"��R=ᡵ�������VVTZ�R8�\��p�}=�E��I� k�HX�t�$���VÂ��<�i�r��1��:9>�n<T�jkzF�f�:ᾮ�r��
=E߷���	��������l<Q����ˉF����7ٲ���ڒ��}����]t5���V4��VL��o�ii{O3�����j��}��X��\�Ƥ#!��:ܓ�	C����
c��UL=��ң���	�F >k9�M5ZĢ��������#*���4�)�Pcs[��n�.\��]���ₙ�t+[�k�À{���g}r�5l�1v�8���~�?& i�؁�>�|Ûl���ш;;=�W)�ܷ@��OA�=�&��$}ܣ�P��J�^���g�o��6�}�Q�Y��C�%$+�`|��xKo�D�>|�X��C�/��7�/���f�l�TV�\�󋉇�;��^����z1���?��N��ix�Qot��|ft|P�]H�6Nxa7�u���v��?��N�9�Z<�/_<ҋ���	GC�ƯP78/��qX�魀��{���hZ������|�?��?������W�~o��ϧ���J}��Ε���턿���9]�xQ�νf��V������(\!g�r��si�{.�o���+ᙅE��轷oz/A���+=z�@�ZC�Ν����!�F�;�h, $�{W�^���}��~��o��bc�X��-��T^'��ҋ'�������{Woݼ���.w�w+Z�Z׷/��〉���+�Z��S+���3�����K1e%e�H
�\o2�t�gisw_������}dx��ӗ/'�����^���{�dJ=�^����#�
�}�إ�gN��wnؗ�� :J<]�ǀ�����{���SW�S��#p{'�I �%:~�I����g������ǎY~`�)� ���|�>���;�0�� \���0�N^�aW�ק��>u8ɘ��Dv�L:5����h�iQ �q0�w��e��LF���5�m����\�t�.I�鹫ƒ�R�f��'<	S��b��?3>�.��i?���yJݐ$�7�k�_���
3z;�SkwiM��M�vJj��-޷AL�,�F�jӰY�̀pЎ�0��Al(�m��/��?�b������*Ѩix�W=}����@�	O94g�r��!���Z�tY���F���v��u��z���1ėL'���/tI}��O9RrqmK����]��������ӨPt$ p	�1�V��W���9���~%���W���P:eG,6�ޓBLt�� �7������^�+�B�栤1�,��i4S4$��k{qI;k��(��E������d*?�'������r��f.��)�p���EG[8��@|_@͎��yL�M|�	4��~������$G�~ќ��
�������{�H��Wb'���0�MUVeyo����tO���H-��(�A _J�A+,Az$ Wt���j��\ΐ��3=�1=m�My�U齋�p�ovK��~&Ѭ���̈��������%y0^��.������(�]�k:�^�6�٬pMG�o��^}��p�ӟ��{��H��s�;a�ؤ�>�W�k̓h�+�UB���d�5�=��W�y}�{�;����^H�eAՄ�y�m���m�Wh&'s:���6�|O��9ɟ=52"b�O������y<���N�l��!�~�׌�Au������G;a�'��G#�����7��G��"��o�����?_�ظl��n�XX���۟���Ϥ�d�(!i$��U-���ں|FE8���G<��E�����6V7�9�a||/��^�q��(��V�t��
GO���)Nvd&�v�zL;B��.��w�y���/���hf���:��?&���&k�V��ܙӸ|�<Ξ9yh��j6�`������6����p��F��BjpGG'098��?,�'ag"t���!�@�ü�>�p��m�����`d8��ح�M����`{wKf,D&�&u-�l�n ��EL'�;�΄�T|H��{zh�.#��2�0�Mt3S.�jie�#�C�'a���=~�����n�5���a�qA�$XdkU��l���<����l]A��R���D,8��7�[��bC-��剰��âc��M\�ދ[�qv�MT\�jKA��h�'Ο>� %Rp����߇א׏ё�>}R׏��m�C�6���h�O����{;�\�B�E�Z�N6c��(�fP�Ϫ�(U���al�pny��e1��ڼ$����t�ǘ�sJb�¥Ku ��,|v��p5j�Ej8��!S���DhP��Bvc�}���Q�UX�d4�)�� 	st(��Q�����~2�d*O�/5ʆ�C�dź������W��p7\���-�ִ��<pz�����D|t��4��i��X��A��j����t����O6��5Ԥ3��2�vKEX�[�K�I�5%%�]']'F�QLD�P��P��Eh����UK��:���pL���iڊMa���TJb�����Z�Y	Țr6�E��7��3Aݣ��Y�8��Y���\�ƹ&��g�o�~��'�X��<�X��/�j~����矢LRf�D:��1ם��r1�A�E����_�׿�5�?$^��ч��fS��&G�]�������43z�۹��q��Ӕ��0�g���m��Ȑ�"��	g\�h��v�@��;2��T�C�d�D��:����N�Ѐ���$[�ǎ��s���
��ob���3K��&}l�Ӥ5�U�9@���0@�z��ɪy��T 87���?{����ῼ���G���~�IG�_��W�>��˅�y|~����3r�p�4��v�*��!�5'a���Ćh?��+ais�T�-�9����
^�q�hD��O����nZ��Gt�p'Ș$�FMS����P�ȩ�;w��ϑ��Y�˫����`�fO�Ϙ9'0:<���05>n\�@�IM��Y�Jak��̿s�*��4��ܧ�#�ƥ�wrT����E1N���4`ҝQ�O�I:�����Aqo���2zhi=�NbtxLPha����5l�n�Afd4��7�3IF�
	��$I8�nFЊ�������k5�o�T:����olf�?y���d�#y��k�Hs8��Yl��hJ_Z�8�}�8�!�}���О�J��[2ٌ�=�4_/ah^C�s�j�ޒA ,N,���&Y��R$a����c��������A~dG�a���5��0	5���������&�p�!K��J,Y%�ƽ�P
�Qt�^dj�d��e���h��- �*:�����gqpQ:�l�Y��K�#��nC42���X�,�����bhp/���萚�g�������&N�L!EW�dL�t�&�ޔ��ag�n����6��8�]�5e�����y���pC_q�C_��7:��_:g�o�`~c�fe��n�N�jU�o�>�lN���GH�������$��0z?�7.մ�6p��v�u���.��IƢ���-y��L~vW�N�hǉp��ao��Ca� 1������x�Q�N.�I~o�T,&1�f�"~�I�j3HY��V;`�M��E��g[��w�3'��(���3�|T�٨Z������ه��-W7���պ >$n�Ax<7��>��ܻ-�n"Ud���aW�aaf������/⅛ωiMb�tY�y�y�m�s�\5pt��F��!�b�3�1�#�|��\�n�
m�f2�4��4$658z�mݗ���c�����F�/���G&�͆�:f�O�'rF�Ro�����5<�la���hCr98	�(m%k�:��w;��U��0�_�t��U��ht�w��W~��/����̣�������A7�<��/>������Χ�u�IL?F|!�N�"K�V(ckyE���&?°�p�Z��X�ޕ�o%�_x�h��A�K�̗�v\���ݒ������v-�*���m�mm`goO�?�0� �j4�F�&胃HD�J%1<��~�v��C���N%��F	K�]l׋�t�8�f�Gf�ݬGN*~x��PׁAo �Ǳ�1L��h��3	giiE{�p,��`Nw�jw�Qvy���<"�s��E�P��C���g����%S	�9s
��&N�4�32�F�F���<V\���3���8q�����X-��x�	��x�W�Ūi*�!i��d����[>�^�-J&�&V���2��-`S�{b��_![������)��iR���+E ��(� ��F��RI~��ϞW��?/�|A{�j�����#;~Tf�,�DH8��--acuM�����2�:�p1�+w�l<(O��#:�F�V�n!��BVp�n[�
:�2��"��:� �X�(�zC6�L�!�CxR>Җ>�]��� "
�zѴ!���1s�w�6�ٝ��uL��qlrc�	L	�⾙�����P,�tNOO!����Da#�X�%ܺ�����:Dc�TE�u��p��f����d��0f��F��Y'�ͦ���A;�J�H	Rd8�h:	G((�������)��b��Ă���N��ݢ��ՔL�S���-(�qqo	��J�����+��x�l����g���S�+\�ɻ�9Ò#�����	f�3o�˚0�+�����H�&���a!���ɜ���~�w��BAEV�'�&V��y�/�d뀠oz�����Ϫ�!�������~�[��H�T�T�W:Y�$UI��҉���щxL��*2�I�T`�t�E���N$��"*le7��C�Yύ��W2���7f5\':�K�"������Rn���b�8�J1nlN�$ ڃY�"��v�T�������lK�,�u�ib�u�I�#YT��j�SQ��|QEX)p>?<L�r a�g~2>����7���_z��;�~�����;7{n\���.\G<����y�9>����"�]��tj����~sac}US��'�'�K�e��܅��\����<%6۫/��P����EM���g�U��v1:/x���S�nnJ?\�4=v)�i�-r P�a�S1o	Ocɤ
!o�a�xL�/�>q�B�k�SG�[��Z�`�^�~���˃�q��,����gv!�q`���#�pjlG�#p�;�9�"]�U��Ѱ<���z����=���8�]م5K�]D�a�o��6%��z}D{�h4(x3��3�ޔn��Z-R�i9%� ��� �!6�lF��� ��Ϟ�ѓ9�{ʰ�I��Uo��c+�g��n�r:�*�b�q��fO	|չ[p���n4d�]I��%���o<4)�i��i�V�3nRMD�Q�;wF�H�`+�f��z1;}TL<���!>��ށ���CI=z'�ϊ)�B��,���ťÜf�H�·�$I�-��t�q�G��o�㰏��-�Ū��Q?(�����}%-3�ͮA:hɬC�-�T'ܑD�\xMN�]�i����q���C�9����L�����q8�����:v��1X�e<��;��`N�u�}ŘL$�_�����F�(h���krV��υJ؍�Ӂ|���Z�P!'D5�G��F��B��F�}�>è�<o�XX!!���z�>�ܱ��0�-d;��f�!*��e�^1�0��>��{����vZ�R����8�r��;qjt#q�29=+�vhK�c6O;{�Rn�p2��j��b��ň�;���`a���ܠLa��]�Q˱�P��p���/[н�bR*5-r*eAa�A)>(1��O��N��!_�Ŏ߃E��Q4*=���>�P�R�,�z3��~�+
Ԩ
�&�������B"���/�j,�6�Ja=J.;�&W�E��$1�)�����X�I�j� ��b5lp���
A�g"f�Z
�9���M92e�쵮�L��_W!fs�{��lp��:�70����JN.��u�1�E��涅o�����J9�Ea�Leh�p��]<���?z�o�����u���V_:E�e���x8w�~�	*�\=�qdd
��38�����9y���89{��#�R����/��r*���l���x��o���o"��`����Dr`>rd�k ��}d�������{��OLY������d^`�(^'��:��D��%D�Mq��qAx�D\>�$,[k�������-�j�9z���0N���IJ�u"�"����83y���8}���=~�ph �#i��S��������G���P�H�V1[B5[��E��i$cq�2��F��C"��'�� �9@�@��/����-�L,�FN�}N�Y�E�A3�3$�+/.����eɀ���ܠF&���,-�bnq^��'���%ԁ���$?Xkj��z`�S�&aY�Y��6Tg��r���t��[=ԫu�K5_63|������o���WW��{���`���!x�N���+����m�aae�hH�����Wp�'W���e�qtdS��$�Ɉ4Äϝ]��� 'ǐVG��������}:�Ѫ���A���J%4�A�FWa}��P꡸Jc��fQph�dҴ�+u��hA���d!�Щ�Q�gQ�g0>����(���cbd�HHicd���/�=��rdDV~�TNm![hw�Ћ��Bm/������|>�O�(�څn��6�-T�����I��������.��m&�ћ�#���8�o�^�:B&���k军�I�4QP�C��F�{W�ψ�����6�m6	2a��NѮqx0������&����"��s��)�,���'Y��bQ�Mڒ�Y^��t;Q�V�y���%��C���    IDAT8B���A���w��=0�|&hrA#"Y�����U���i8"�,΋���3Cs^�n�p��Bx��^O�c�T�/\�3���0�n�޳'p�E{t�dA��a�ّ H�Ib_��rC$2Ò(~N�v
�=���4�ύ��!
��7�˲õl{�$�%3 /@п>R�g�LY,"ۡ���/�U+	9"�Kr���ך�%"	��PZR�Z���&����nVe��p�P�Ѥ"�k�>�,�����V�Rf>�O`y*���?��o�K/�߽��S����������_�v�r�E�N,�-�������]��+�/b0�ă������R>���q�a�e
�<V.�[
�n2���ť�����/KC��a�OW��U��=z^M���sx�ͷp��Cao0���pt�M}Lmi�����ź˧"�.���>d��K/��^����ˉ�O?�A�*&�1�J'v	�I�jM�L	����;w�qqfg�u��_-���R	O>B0��kzt�f[�����\��wC1_D�PE�ƥ�1{�������瑩	��������DM��������m�Z(�xpy5#�&�ǁ������,�$�x]H�G�ռCޝ-Y���H��
�H�����JM?W�P�͇�?�:Av�F�k�eLRYQ�˽,a{³�bM� j`I�1L*��ٳ����jnܿ���9^�k$9�4J�Ν:+xm7���=�����������2Z�+����U��H[zdIf�6;[VD��`��Q$Ɔ��Pj5������M�5��	g�)͐��-1�ea��M8H&��g���M�4��l��e�-<l��8ba�E�F�\�+���D É�)̌�K^D�7�;�r�e����PC��E*b]:3�ZSA�"|���#�0Yh�JYK�R�n���V���L��wt��!�����`��e:ѢTm*62�Ix�5cO�C�Y����R�L���L�r��Ld�R��CE�W>��~US�Zy����<� G�
_��s�GqbzZ+�<pY�I����4��u%d1)I��Z.X|� Ԍ\���A��"����������3,b^����>G�o�}����R���TZ�!P�7�>�B�� 2��BzFI{�t^P1yL�3��ke�azdX��w?�����4=��L��L�|����#Q��t�0����)�*����,~
��a�[��j��]�i���oY|K�1o�Ԁ�ޚ�5��[v�*�4|�$N��IL���{���]�N�h
�*��FU��jE7DȢ�'=h�!�Z����D�z�	�p'\N�f�8�������������/��y��w�=����/��r~��#n�ח1��5J��X|!w �C�cx|������������X���
���k�Wl��|��M���;}!��K�XYZ�A�"<Es&��(���O~�;w`u}[wM�VC~���@�%Fe�t�?�9Ą�9{P��׿&��x,�"L��:���d�%t�������.�]ن<����(A��"��ҧ�fpbbR�Yute�p��=��>��'���sv����GOa}cU�q�P��(׵��$|db
�OnK�^fg�����ZV�R!��ka�ǭ^;�}(8�eHF�|� �'�E�#a����L�o�C��C:����&�s>�S�)�h�v��a�M�A��-��D��gXo4dr��8e*����DkL6$�.�he��tP��Uũ���Y��N��~y��
������O,��,����D�'�V�3���'gp��1\8uI!x|�|V�t��7�0'��HzV[p�$3��&���QO�#������a��p�) �1��J��dq��Ut�7l*��MF;�AYa�d�i�W��q�L��5j�	#��e�//�E�y���x'�M��Ԕ�XY��@(2�H >=���(^��p����E�{pz�3�nk���C�"����`=[�J��n~�#CLN�56�n<�.IN>�~N��QB����t�38�rb�AJ���h�(�r]�R�wʭr�r墊���t�4�s���q9�7�ˏ�Ӈt0
���~��$�x���;/�,�F<�O�>-2&�-~��;���^����o���؉��L&vǸ�qW�&���sx套��9��*WK
��C"� c�q��~���j�Nv���������L(���D��C�P���Rؘ)T��Ej(m�\:�5��9�`���m<�����a�rs��F�e�clM�&^+oyz|G��%W�~�	_,�"Y~ɏ^ς�vb!�u���lX�-�z6f�:\M)R�rϳ����V�K�4�K�F�4��CS2'pL�ynb���c������,���Wzm��n��4>"�Z��E�v�<�h�S�K�F�����nO��1�m4���������/�?�}���'�lm�f��"�����<��ZÓ�����wQ,�{$���vx�8��}	;�7�#{��Ns}uK%�����_j0�n>�kW���񻱼����y��c�*�nO�j�k�{�!��ck� NJX����3�t�Fc��E;I~�Q���aM�)��u��%��H�L�B�X������m�pY'@�-/��}��Ȧ��r۰���&�C��h<���}�ի�}��]��ff���wc7���8��AU<�:hT�9'��G$�C�]�ѣ�1�!�K6&�����c�,m�!Y�6��IÈnGהM�UN��g�+�WJ�R��g�ݐ�#.��Y�F�Ā�`x�W*r�bP8�Z,6��^�X	]�Q�MR�a|��Qɓ����I��n�`Bxh֚�+*:�CCx���x饗0}dϞ�?�)>��M�)�Q���ݰ_��$6N����S�C�c�;�51l���tE��i�3SQ�X$�H�O&Pj�5}�{�D7������TX�����wР޻XG�\E��z�6�,�l��h%&�sb��&0Js(�`R�c�aa�oM��.v����U�^�����0�L�a|tJ&X>16�$=���Gt����{_a$�QZ�H�j�~�n�d�E�nlby� �=�HX݁(|c��MO�5�B?U6p�,k_����|����#ᎇ:Q	2n�T�T�hMf�R�L��Ԍ9d&q�n�<���e'K�sJIb2�@6/�j���zC�9����Y\C~y]ֲ����x幛2S��̝''�@Ї��]������s�rz-�##z>ⱄ�ٚVJ���2�l�0=6�+.��}]�,��=z D���U����ڗr@`AeA���/M|F��5a�g2������2���ǥ�`��@Bzٽ�
��&�ѱ1�GF��?���U��6}N�q8H��U+�5�x�OJ�Xh�MDKPi�,ؗ�+�[�ėwX�/�6�砷��	����bO����&��ޞn�^�|�/�|]}s�Hma��$�������5�P�=�|n��xJkm��\��y��[ɕ$y$)�ׅ袲ȼv��Ǣ�����"����G�=����կ����ի��K/+�wso��ǻ��X��$��*�DN���m$��H�"<��)J���GjZ��N?�T���k�T�B>�-�����r&&'��r�1��6�߾�M�^RnP�nL�	k"q�l밤�
=L	��K"EȔ����rWC��iGf`�(�����c$u>����]3M��2�;}!w��B�%�jEjN����?@��!�=�׉��u<xp�KKJsi֛�a��(�J�6i����Ј��Jp��%�:u�C�ڟҬ#C��2s?�l(����DNTM��-9PjhP� bB�EvU�jU4Y�^l������)5s��
,N�wj�)Éx��&=nFF����wP�5e��?S!q��m�Re,}.E���պlk�~�up��,���Kbsr*|��>�{�=���4Ý�5��ȩ�zaI��A8��X*��㓈x|�ӊ�RQ-'y�K[H?_l"����W�*h4���)��ly��6��u�X4y NMO ���ˡƄ�|M�rNz�������6�|n�q+��F�b�r��i~�^?ߛ[.a,,��>ʅ'��F���022��x��3�9wѡ��x-a�|���%t�����M���h֙��~���LN��U�P�dޱ!��F�N�H2�ܣG���b��*�1��!��i)�t�FYL�e(Fk�HM��;uF�g���c�WM<�95���率'�0'�~���ȭn�wP¥�'��/^��-]+~�4� R�w��w��.���c?�����K������ur��p���e����<r�Ͼ���%9Z]^���b�i��-ޚ̬�_?�V6�,�������k/���'Oʰ���>��<F�Nn�R�#�%S�"=:&̃��X^_�>��5	�y� ��%T]=4<�"A��>�鍃�i`�Ŧ)��6�MV��SDd����灍��^eO��Y��u��l;䩘jl��Z����F��ߒ�h��Y`5H�{�������{>��m3r�`XD-}呓cdIU�Cȕ�7��Vn1�Y������+	�ٓ0�5k��$���"�����[O�������%hv��k�������G�k?�Á�#��i�8�6&%@��yc5mA�,����ev������;;s�hH��ӧs��SG�jq9;����g?���*e�ռhY^��P�bN6e��i����'3=^y����s��磏��񅂲{k����D�GQl��uPp�iy	K��ۃ�z2��B�/_���;	����pz*�G�O�K{�Y�O�bsc}�LV�4]�z�.�8ҩA�b	dPmV���� O(�Z*�Q�	F��6ִ/��$%������k�j���6x����,�^�>�"X\Y��DŢvx|"��U�"!u�$51=��/K��i��nZ�1CDPk��$�PJ�ǩ���iT�oK��!��w��#�I����񵗟W,e����'�}�[woI>DL��e�_�3��Cf)�ZE��BH��j㞶f�����H�!��fKR��nN���P��EX���{E��D\S�Z?�ޣ�n�B�R	B����\�6<b�tW$]ᤧ�	*nD$x s���+�|>�r�(ׯN�&�Db���G�G���K�p��)D�>d2�1��U�;=l/.���"�� �/�Z�䆦@�P�@�h�d��aG��K'�f���X�I����u�@���)h�Ag.�)6z��2�D��ڎ����\F0?O�:'f�98�y��&)҄��u�.�P��a��S��D�n<�
��꫸v�&���� q��^�ȅ�ݿV���ގ��3���ƍ�����'��k�j���^FE��j�B�������?���f��G�G���͎��2�,=}S���*���<��'ψ�E���d�(�9��9�%�%> �u|^����sR�Mv���2>'�cs�xݰO�At��_��AR$U2�Z_�;L�b̪�<��������Փ�َY�c�0�SQ�WV���>��w�L{4�pld��-8Z�zR���j��v��n���6�P�f_����6����$c�A�<5r|]]��(�ѦG�����B"$�z��#�����Oz�A|��|��=�����;��ɓ?�[Y��0�^�"bV"�>�������T�z�`��MR�K�� o�h�	�+����+S�ݭ�����
n\��ӌ�󸱱���%�E�85+	S�[�߽�x�{o�Rnʋ���6٣:S�B왽��vs�o��槉�`˄�K�)X�-�D��Ut�A�{���枆)!�9��X�EGk:��ɤH,��!ܾwc���E���~f~�s���(�$K�%��j-������Νq.w�d*.6&a��*���P�K=��m��n2|���h!gNd�W������H�����tP"��5��c`�����#'c^�s�[�o�"�����Qoij��A�'[�+(QQ�dPҨ>L� ڽ��N�bt+�����5�_�%ٛ��s�nݹ�[�o����:68(~ 'p��#k��~t�B�7��Vn���'�ImK�Lړ�7�!7Z<�/���m�Y��9�����!�~�G�k��D�kf��n�r�bܡ�ӕ���1Í�2N�#�ϖ�%	[�eb(���Q9����H9@�k�ׄ���Ňd:��N���s�=w
�XP�?�"��=��e��d�o���{O��ɣ����K��8�	�Cx�1��i��FR�f;١��r����k��[F"תյ/�N���-�ڨ�ܐF0{�+.��k��9�)�"LBV�֋^5U�0
�9�>^���&���bF��9�o��\9w^�==���O�8�@8 /����mq"�;�)�E�¥KJ�Qa�sM�X��ÙA$0��r�<��=��w�*��;~�,��*t[]��糉H��cqI\����Mѭ��ؽ��|P(�JU'2CC4fc|��������g�������Jș�S�4ӴC�N����=�ri�Ć�S;m#��*�e>³�M�U1�Ҧ�LSQ`�y 测���d�[�-[�dK�߹��Z?��2&��d!j�p������C�y�֤k������2��������)I,¹��٢V&2 �ҫdJ'.z�������D��?�����ߣ��G�+��ܹ3�x��=��|�;�kW���#� ��ǳg���PY����� M 1���=�-�'�/��w �+ �w ���7q��q�NL"�b{}]F�bNٰGgO�ۮ�'?z��wP�4�i����M`�u(���U}���k�S]^���I�3#�6a�$�)4Tzc[Q�{=�[e���UM�gǍq���M��k�p��YD�x����(h������ښ��z�o��������Q�ݞ��$Z�ԢLrJ�"[BI=�g�܅���}9�����Gg)���
�V�~�h�vKI���~(!6I�9w����
ʖ^2���4�����AF�U�lж��������Eo�zK^��r��L!Ȫ�u�m�O�����5��ۖ���e�b1L���[���^���c3�.����ǟ�|�&zO4�8mA�L�=����l���+��#rN�PC�^��N���'͵�v�6c� 1�%==���OބJp�B�"�6p���3���"zp�H�iv$Y"Y��ր�0�!h��a�;���o�dj�Ƅ��`@�d���E��p.#'�V��ωH,�T:��Gp��Q�M�*�����ԭ"�g�������]<|��B�z4��T���mӃp� ��L#�J!D�,	nb��2����Nm��|d�`�=�)e���kNt>��Z��&����+ݗ��9a�w�|� e�}r�J�CD���`��
�����c<>(��y��ϟG%���Ύ�3gO�`7�������V������`bjJ�F!��]$C�QڦRGr�r6zo��7�?��"�׃!�z��2>�a��R����=����^x�3�c3��۷���c�}���8���Z�v��#C"h� ��I���kk�v������������&�Y焸|Di
B,���w�-?�!l�PM��%[�e1�����ٿ��mdL�:B��������X��%��,�J��P�+=�����5��e�B��a1��wy/�M�דr�s8��������DN�M��?,钏!0���h$�����y�_��2�����.���j�\�x/����XDE,��ǽ����
�wvTN�Wm�Eng�U����d0���F���i';9<�!܁D�~�ll(Ԁ�N�x��G�]�$���M�-���|��.$9��~^EN"��a�M#�u:��&��Xt�e�T�����O�=M�2�~��F���̿Kj�ӭ)�ߋ�{�߉�.]��3�K���;?�7����sW�����������_��#���:J=�9Ш��nzY(f.^SB
"�R�k:l	�Ue`R��k	lv>o�AC>}&a�E��?L�+&���`@B:|UBٍ:�̎��	�q���8��A��BU&��#Y�-.}/    IDAT����O&�O{[�(zt��ĩ�@LR~F�G��0s����+86sã�ޥ��Ï?���O�C�.�#��F|hP������i����jE4�%8�M%1�(�!��݄G�����NLVy����BM8�� ��
�˹�����0ƇFD���{m�h���W�ڜ��#�.�Dq�W�tl`i�lx!G�V*4��X��P*��Dt��q a 9���a�ah4�x�C~���)��ۃ�O����R�er����4��iv���#�2������'=�t��3C����A��� [�ϼGx�s��Q	��l.''�B��@�F��	����A"<�D�DFY�}���B�P�t�ǽO�I�M�Ջ�𫯿��.���bw{[�Sl��q�x��p��}�2y�'i�K��PH�437�m�L{��`�����	��\�������c�Eoj>�$j��n���'@xS���G0�diui׮]Éc'��������w� D:�|�a䀔J$b?v�c*��P$���{?�YՌ��Љ��M�j�.��P,A��y��(r:s�[nO�:TLٚM��r��=9�8[��-�ѴL�PΟi�e&�@��4�o�y�M�q���/q����[d,����-�gl�����L`��0�v�RE{~������\��F/y�.�����/��������W��j��[#O?��ŝ�ߨ�{�|�"^�|�h}�~5k���@�Q5�F� �f�F-y���L�qH�7��@Ry���N\�.b�?��X_]�N���'f13{�v?���������^�\�	M� �{Ol_����� c,�,��;mOW~В����[>�PX�<�^�ߐ@�Bǝ����Y�-�4ӭ�9~/�W6���gq���������i�7��������%�ʡFQ]���mFm�S[{n�4��NS.��J#'����83���&i�O�'�\ل�����2���P��#�@�h<![��`���v���e��6�&��?~tF�u�^��斑��9�����Jt�^��mM��%����5�Ru�<�h����f���4^~�F�i$�t�
I�{��}|~��3��4J���Ht��
W!��X@�P�+����4Օ!HE$i-f��i�_�>�n-�[����q2��Z�l(s�D��3������9A���TP�9�^��ͫ`�!x�՚r�2D�D�h]H��ͥ��I8D��TR��GN��	��D�
_�}r����MM+�P��J�����W��JkM*��je���7�Df3@�id*L��'��0�dx��MԤׄ��D_�@��S݉�4������<�ˍ�V ���%���=���+L�=�j�7�*z��� &�&e�{�ӻ(�B�	�����W�(ݍ�0�������T���{o����jy����%0W���Icf�=�Aaj��R����_�=�S�"vq������ʺ��	�6��&�?��ikcS;��O�R&�����ÇD�l��?������* ����)���i�Ei����'�~��b�NC9荰�#c�pQ�F��"P�~��<����C�|</�B�I�&3���T)]ł��<�ڨ��lZI��kU�o~	��oň�g��"�����l�5-��>,�<�%���x��9��4#6iK{�>'�
�76ń6�i����lu{5ر��^rw:������{4>�o���WML�W��JE����������o3"����x��M�Hc���IbgE�=7�(�Fe������\ݮ���hOפ㸸�b �����rI�I�R�\���Y=>+x��?~��w�Q:���t���f
	�I&`�Fx�ӷ����p(�����~�,r�����{�u�ϸ�"���#����&�a�&�bOv!���C�҉s�p��%Meo���H�S82=�˗/"��`mc����xt��X���)�1&f"�sII*��йN��XU�������Ć�Ϯ�P(��#M�!1����\lǞ9�-�m:+�PdX]��6�NM<Hx���0�����L�y�$���0�HQ�Ζ��M��|��"�e3��Fk M;�IҐrEwbd�f�XA�9�ч��P�;;ړ�@G
�.xL1��!�u�hY�����ЪԐ�?"b�_ #��`�G'1�&w{O��Z��5!X.e<n�iY���t:e2B_mYR��o��.W�n0|�T�錶�-{��Ŧ�ð���HK`å�GB(�@$"=7�_l��0��>��[�X��fD�!$1��<pS�	�M��VK�ե�50�Q;?��>|b��uߐ�V��Ѭ3�DG�$)�'f��7R�`��\���x����f��6��2�XZ\��ֆ�qrTc���

Ӕ�`C�.u�� �����T��fs�l�|87{S�xr�	��w%��x�"~�[��sW�j��f2���;&�ڃ\o�߻�ŵ%�����l4��.���2M��ԑ�	L�09nG�&E���K��_���pʉ/�&��΁���O~!E�u����'ʦ`zbZ��hz�ӥ���g�� 2�r�

l<.Y���7|d'��b8�������ﭣ"81$�e�E�0��9��ueM�����Ğ&iς͉��_���f�k`���ʳ�.�bKsP����bn���}��gP��v�_&q�Lk��a�f�{����*΂�i>D¥<���զA�H�c�<����6d�kq}�lpz��'{�_�������������^5��_��+��=��z8��<[����N�y��%�v���x��`�<(�E(;��0��h\µL("�	3FX�/��K&(�a�4]X]Y���nN�SGg����g?Qns��"l�o�t�4X>�L��;h�;f/�縉P���n�FN��4+m�� �!�ɾ	�A2E>�V7'		���͟%�����{��5��z	�d���;2�?{��_���@��~��O0?�Tńא7�p�=lG 0�ǅ��&X�Z�h�$������.����x��q�%ذ�+���~�$��,eM�c�s*�p<�	8gSbv0$��u��Qv�NMk�����f$sb�U�G�5�W>�V�U�Y�eʬ�^��Y��'��i��U��iTj�3����p"�3�� ���m>Ԕ��sb-�˽��e\�N}�Z.��ujT�y�;=$#1��A�4m�@~��ϟ5����~��%�j��X�ݎ���#$�"�2��R*��T�]��[�I��p�\B�VL�c�p�-�-R� �0b'N�`i����{�k%�1�N����_N��z�~[Ey` &�V;�"h��=�5)|���4Dy���	�Q����ޛ�[�J���Ҟ��飘��Br|� ���l��\�.srJ����f3��$d��W��ww�4(Z�Kɡi��B�])�aؠ�Z�MLY{vzן8z��SXY�������׮����r����E��0,�\��v�6�->���:'Rj�y�)$;�A5�0FӘő�1�;yZ6���r'��g�����/�[���ӧ:�ǧ&q��M�LY���U�I�b�Y�rY�,��<��ZT���=9:%���(�͞���d�I�l����S�t�(��[ &ș�j��,l<ߘ.�)����~�&Pi%c�H~Q�M����V����0]���_�W�\HS�e�dG"��.���`+�\���ۺeZ�YgΗ_�a�������5�J�|1ڔ�6~�NZ�t3<���m�p�<���WO���?8~�dX~���T��^{�p�}���{�f�s��e|��s�ѕ��Ȗ��I2�?���v�E�J�N3�V[i�ܔͪ�N�
&��L1��<�6�WE��Eۑc3��9�=�{?����Ot ��E���,fv�����V��SJ���Ֆh��-S�j >���i�ϧ�$��;����K�|�h�da��eE���5q���E|x�n\���Sp}x��wv�q��5\8�X�>���R���؁��M��.5�A�<�F��su�KU�N��/�t�ѝ��'-����im_+�-"��LD��#!ԑd�dBM�7�An��h���,e
*_��<kdv�^�hb�v�KY��0eF2?/��M�-5�2��D=pO+uĭ�aDc"Ɖ�L.����ǀ7,N�!��;���a�M�� "�ZU��r6'�*�>ݧ�C�mٶ�hAd���Vޭ�Ma#g���0�Χ��n~�kT�5d��ni�m%�d���%��6�z]�sc������}+�M�OD�_O�Ә�9������؀pGL���Ť��d���Ɇ�׌ņ2�{�M��}��2�|��W*�t�Щsҗ%u��N����۔�dZUd�UTi��s/�a�M{�z����7T��Q6�&
>�
0ߟ�ljJ=��I�qRfW(���� ��)�����ਦ�����G�h׮_�o������﫡'7#2�������M=o6B�g��j�^���F"Q�o���plb�]���Db�g��B�s�V�@�{��<g�Ls���m���8v����D H�;�<�\�|���(�{kgG�8�RYlq~_��<@7���pdfF�p,�3#���d�,�l���^/ ��.�'�etfp��^�I��L�l8�]����BkPS�M�=,v$�ZE�.���ɢbg٩G�Hɛ�46Q�RkW���g��e�i��v��r�-ח׏�����ށ��H!U��r�������>f����p��Ɛ�S
G�������^�j������W*,,D?Y�����?��l��|�"^�v��U�hV�:0�'l0z���V4;H�exSБ���3RI@�>(�����	�� �҇` [k�_�G&�ő��8r|V���>��{���a�T��f����bTN�tx>��ԉ�%M��s�{�����!w�<h������jGI(�`n6,�2���VQ�7���@*�S�/��ː�~���ǫ/���gNj'�m7d0�/v�ܭkgm1�E��$���jE���Y���8S����o�~٤�&�#0M�d*�gvL�0p8���~��Șe�Mh��w;"�$<a������J����&�n�iŔ�~Ћ3b	Y�s
�V�7�8'r�Iʢ���u&�o9��0�h�2�����L%���e�IiJ"S!��C���|�	`1��)��Z�0�k���n82`)"�������^�=�,4N'�����s��"L� ~©Q�H��yOɺ�bs� �~�A tU����֨�[k��l�0栌������A�]2��sp��g�i-Of�G�2q5�bB{E,�
�ň�
#�������b��ҥ�	�=�/d��K4��`[�T,)v.�t�
���Yɣ@c!x�:���h�akmK���1`@��4��$L�ӸFԁ�����*"���w�jU8�I�����Q,Sg�G,���+��Ư|ׯ_Gv/+���,�l �����§����BlH�S/��~�&��I1��rd|/>C������{���5:�)������!ѓ1�l�I�"����
���͛*�$���x�tN*3�qP�KNU��������̴�|*2�ӳ'pi���b+���|�6��Z�`�UF������r8������"�q�нne�je�3�;�,H�#6g�Vߴ���H� ,v�ڷ�6�L�ӶI��R8�)[7�g��C�K�H�I�gz��:�t�J�����������π\!��s����!?�����c`���ŦQC���U���]G;����Gf��?�q���/��o~�"�����������³�j�X\8s/_���T
�jID��ՠiW��D�3�e�&A=o��)-��^6iv~��-ێ�O`bl;�ܾ��1{��;�����3|���%�glo ��ү��N!��)Ȧ=��|���W�� bѨ.(g��Vh6/�B���ü\v�hr��5됦�=�Z���~�����<a�);|(6�p��s��7~gf�!p�����P��Yz6��k�L�cb-9	�i��j�P(����,d�i�m�bl��[^�>����Q�N�/���[�����x3��9��=jux����)
ۇZ��l���J�n���九�0u�Y�$e&��$��V�^#��ϱ�".wO!c���<8=6��/��ˋ��m�����L,�~�ǅ�@L�/{ԩ7�8��C�S7p0�c��>N߄�d�iI4T��@42�BE�*T[A���Q������k�P�����r��f���&�Lx64W�u�ū`�=B����=(��l���=6�V*��0KN�;�N!�#�Nj�%���.' � Z����\��q�솇؎��L�twgK�;�k�H���1|Y��	�G�������uv��Li�eЮ7�jvԐ��sme�����$0Y�����~�����Q��!�dK�˨2��P��|�1z3�����eh�Fp��U��S��4���WX���1��W����\аt�V.!iꙩ��f�2��ׇ����c����nll�Ѭ	�'�f�}�̑dF�#>sZ�O�ّ�j<��[`<��~��m���"�W�F�rsh������X$�{��9l��#���3�^��RfO�D�T�]M�,.,�D����B[8԰9���8��xEd҄J��j"5)*�� �|�l�T�9�~�x�I�ڌ�f{�����8�pl��JR�Ό́��E�
��)?u�݋<��[R$�-jӹB��=��c~e���s9q<�a�o�ǜ���߼M�����Ix�tj��?���[۷��s����g�u�X���K�E�?8����>���W����4�cjt�x�5L�����f�k�=0/��I��k,�oa~~����>�d"�Ln��������BKOJ�4��1��=D��<Ŏ��,��s�,;�A���%X�9�<H� ��#�m�)Ά�y�	��c� �a�(��K�4!��l�h+ț�d3Z߱��l�I?�׾�M��~�N��@��g�RV)�]D��ecHhi��YŐR%�cdM�*��y��k�M�K[fKt8��!c�鉅���	�`����A�9��L�F�FG��	apNYސa���Y|6�=A�<L9�r�l��0w��7ޥ�֐(�2s���j����B�^I)�wa:��`p@S������xN��j��1bn ����$">c�μ�z����Ȇ1%�I ����`�N���{�8g�<*���"?��vG�~/�rۘP8:��{�C��>T��E�[��ښv~���
;`3����z���y�Ѹ��B�����zlH�����z�r�� !+��`�{��d1���E8cx0}(�c3$���N��SdT }�K%]WZ�*Ǚ�ݶ
�����D%?6]�N���a/��b㣚�y�6��2�'��p.�Q�m;�A��8Ő�J��f�r���n8�O�JGS�DD%�{;�C��F8�Ĺ+W���^åK���F�u"����_���ĳ�yd2��T8�Ӊ�hT����������b���(p��DK��׌���7��/�<�1��
B�D��N͎�ˇb	��9c�SAy���6�w�	�r�Q�A�@4�dl���� ��s�=��W�Hc�������m��n��m���(��)�	ߍ�6�ÖE%�+�	S#c8w�N=n�׽~i׉H��5�fiv�6"i�p9�	��*�.�m޷,�nQ�[k:$�����{{bd	��%)L��3���M�m����ʌߗN?�&�֢��b����]|�'?�����#|�H�{!b�v�&�(����m.4�tw������*�w����åg�M�P�;}�_��0���]�V������%9ɉ�4N�������4�n6�B�NSv�����g������=Y��=v~�{[x8��}�-l��"�#	6aY�TI�v��PY�����-�)y������u|�D�q"C��X]�����"�0�H:��Ԣ������w�q�g�]*�)�|D�Z    IDAT�����"�� ���*��ΝC<�C�R���<v2�����q�ZN U�[��	�RZ�GH�R-�˥�"��Q��)4,z��)A�S="�.0��F��+���$y͘�J#��W.�����\G�^��ؐ���G����3r]�0Y�4D��bf����A0�[[�(d��/@;�V $@ۿ�.��1@���'�}�ۿ���}AW"݅�H���r*c���VGS�������� )B�l���bKS��KWq��U$�)4�uxh�I�$���)e�?#&��'���!Vs�}h��Xg�ʒ�-��`aa+K�;��` f$"�DB1���k��=P��Y��Z���s���톟�����"g	��kS�8�
~��;2�V��C����	��9�#{��@#�?�sl����9�訊��ilHz� ��#G�T��$�Fu����7�����.�7�����}�=6'�ۂ%�q
�g��N&y;_��+6�^?Rl:�A9 I~�d^5S�rhQ����Kx��W��/��1�qbl��t�������`�'O�I���`����I��D>?�bA<e����iN�H��Zar��ȕY0(H����2�m�������P�Pc&��'+��!z�'��1:9s�������ԙ�O~�~��6�Pqt���a �C�1�E~�<?�`q"����k�0���|h���&1���I{���U4y�7o�}�##�3�Z��e�����X �XDB��Z�r��z��h��Ej�q�����ޖ߯�,p�K��n�Ír����-��;ocqk]*
N���?��Eפzy�j��<�Q���*�N�d�n��g'�O���I����ra���j���sx��ue�����G�������L(-����^���4���K��c�S`�i��2͘X�����Ul�HZp��e���t�)��w���k9u��@eWv���R��0�R��&>vXL��H�`'�cvj�jU�x�b�&�+;5veLᇢlW0)S<�i[:�h��!��8v��7'�@,"6��ֆ&an[n�x��+��y{���,;�����{S�uuWW�j7fgG�\��H?�E�W���%)	ZIDP i)��j֌�q�)����{���;��E�P�{(Twuefċ��{����k�	xqzr�O>���"�eu0����������7;W>�
v�մO{��>�ܮ�EB���-G*��$,�{1�Pk�=�b|tr$��lX�tw��}�v>���$��ch�������Ջ��.4\&	�S'W�q��e���z�!Y�D�r#�ZUH�-�lM&�K���p7���Q/V���C<���q5h4")��l���K�}�y݃
��z�ĠWzM0�"�B���&r��$�y��m��J�cYl��'c�җ�ń�
����t�=��i_L�S�h�3ٔ ���u���^�D��g�$!���v8�Z�Y}Vl^���y�b�?��<�;�:�70���lߧ���]�E���_�CNqbEӈ�bLa$��!M�eS���"%���E91�/S"�s��߅��A�z:��&I��pkGNj�vyO2J����O`��D����B*�J&g��LW��	CG�~�|�P#�&�fs��,�<ɛN&.\��o|��^���l&�]*u�L�����<�������#e�WVl�y�0.T�|��R!/��ӒA��]-a�PUs�r_���ѳ��t�g�yƝr�C��N��ռ,,�tub��f�,��m�Պ����^�u\�r�����O?|ۛ(:���hJJ��,])�9Y��܄�/*a������t�Db��}��.�
K+odJf�D��C�����"[�����"�Z\�(��L:�D�Wv����d��9�Z:�\ܲ�%�"(����&9�ю��A���1~��/�q��l��n�n��C�e�iC�iq�<#��Vq��F����&�華�I}�;��������V���d�����g��U���	���?T!��ux���!8��ˢ��"mp���bEW-�E�V�Y����XZ���i��c�:s�6?2�S�l��/~�c��o����&����\�a���@��aG�N����tx�x�ӕ�uS@l�*�4C�R�t��ִ�U�("4��en݀V��e��[�?�C��pif�{t��~�H)?�n�����w�곷�p�������Ճ�Ū�M��RU7;:c�	���pZJ��i7
o�{�sOD��x���-0�2��!� 9�p�(Ӡ�-�~uuY�?4�X���]6'd�f�y��/����������~�N��o�n�[�I��*�Q��w5������#�J�҂rK���W�\���)bEH+�t(�d����&�>���1��9P�T�?0�"|��5�
��<��W�b�l*:�����K��b�+X��u1�a�N��5A@V����Õ~���&`bf��I��]{���f���\!+��,�j��y�����:�eP¦�
b��L�P���C��	R�ԭV����T����a�=�G��j��KgT���x/�Y����3���Y50=5���HK7YSy�E�#6�G�+o򣃸���w��Ogdl�z�dJ���*�5�P/��������<nI�B��y���!��9��t�s��.L���7�����+z�D<��3�ךP����\�޼/��xس �Y����C�� �!Z6k��C��s�!�q�� ��zMӺ䃕�&7�L�Я��J���I�� "�v5�>؜-Q��)����>{���20�L1�O��o�.�wֵ"�3��E��M�����B�U�$�H���k�<}S���ǝ"q�J���f�҂i[nT�r��VmqAZ|�$!/I������NB�U�
���:�t�$8z�!���*�!�5 UJ%���w`��C#�x��[���X>�ŏ��{ۊ�%'�͔�<c�=.T9	�2���ӐS��v6:��q~l���嗒�x^a^ZP�q��:�"8:�c~�>��=�l�>��^��b
��DW�]��>�Si?#���UQ��p�H`��;G	���Mc���]Q�s	�~�.�wv�M�L�?�J>��nȶc'j%w��Vs�ɔC�Ƥqꪪ�(F�&ښѱ��=^��$@���	nuf&��J(�\�Ġ��B��r�b����~+�ϊ�E��3�K��&^�t�8��?�s�{pWō�51k4���0�[iT���|Aw"���@����i�e�RfJ�u���Ŏ�p�]����|�u���giZY]��ܜ)mmO]�<΢y|v�_,$���r�J�&�m����
x�_�5c����Ƈ��A�a���"4���A,��փY1EX�d��P��T��]c�]��~OW�����yQ�%�&g|���z��C�����ʹQ�h�8�����_Y�����xXj�.{P�L�E��h�GBٜ:�,L����Ԅ�`x�p����=+�}� �Y��m(�N&Ҵ=�
�pP�M$��c�ȃ�;�|:%])Mm!���>�P���T*�Y9�	�P#�T��*�&N�t`c澚��%�*@-~7�y�kl
t�*��`������ц�@/½�(ԫH�2��OO�H������UpX�����%ꃺ9Xy�Ke���Hʫ&I���ϭ=05�!�W��{{L�`�?6�������q��e�y�-<w�6���>��h2�ω����c��P�fDh�`�c�}xը
�.Ʀ���C�D�I�Ϝ����؂J*cM�f�#�ԨBZ֧j���s�fD�>ԝ5uDbx�=>�Ѩ�h�;���1B<��r����{����c~cU9��@@�,¼�[�M�br&�q{094�W���gdf���=�ݿ�)~iZ�� �1�yk��߱ȑ�7ꑰ/�{�(�7V�y��I�N���\��l�Vރ�Љk��C��?�+!���������&'���#��;?����Ւ,zyͨ aq'�� ��J�s�f�e B3��ь8=v�s�?��/}�E���M����������=��7�^��7�C7���c,,Ω3��e7��P� F��1�ݯ�7���H4�@�W�ff߹�����c%����p�����v��ţ�8:��Zh�<�ܔ?1s{Ɍ�B�fC'!����
�S��+[Mpb�Cl�Z�' �K50�7����"�Z��jł���&��o���m"�;d'	g����p/��"^�q� rg��ɏ�k�:�]�,+�]��y��O�qtr,� _��/��@{^_N�k+K�k�u�|��%ÊDP.s;F6���O;ѡ!��DºY9��on�@�����A�0��D"����nm�`��)��&���!V:��7�[3�]�������(#����c�#?�F]�eJ�(����ùZA�f�x[�E�R��T��ݽC$N���@�fG:[�g
���hu��IG9>6�3�|��	&��y���4]�)�ד-���m���d����I��'N����65�3���jt�^��q2%)kyiU��<\���3�Ta$Ȯ�nt186�+���M�-�<�RrWK�&#%��g7���aV��h��q��x�1ΰ�|Ap3�	���CMR����3!���&"��a��U�4��	��(��4�F*��@6?-�R��V6�8��!b�bYy�!NA���@���Ϗ�߇�ϧϗ��B���t��[��A(ځK�n��W����gdC�{�ި!�"����f3y?R
��Vj�>��L �>ֲ@lY��:���n96�\���)�$?�
�X�e�jɁS�t辒_qЯ�:�T��q��hgLI�
x(3$T�F�P4�]�GE����?���
����LƱ��~�f}E���?D.Ϝ��k�1=2�Z����M,>������0����Y�y���$o~�˨O�&���y��eoW��-�%��H^i�Ms`Ag������f?���*ZP���1B+-�d�T׭-Vn�)�C���s��ڰ�J��x+;��V�p����i��5�k���׭u���W�lښ!��Ϧ��������7:	/,,�?<���{O����t.|�������E�H&��d^E8�:����/փ��L�*^�]��;���1�WLߓ�8f�<��i����1::���S��q���0y���'89M0aC=�YZ���<���v)���p��\�r�j`k~��s0M�v���ֳ%�j�*�DAdI��"��v�MsS� ��$�LԄ��ݲ:�Gx��@Z�M�;�g�����zP�f���"~r�C�����7�.w���)��v�����%Ν7�`|dT,�{��ƃ{�4]�0s�u;첫䮜P�29	a��Bx8�H�@����+���K+kJt�u�<�;/9I6e~@����I����/��|�]<��!\ȗ����.��ٖjdB7���Aɯ�Ý}�X���y=|�!��Q�fP���7D�L>�|��@ ��W��C:_�I2�i��>�3�� ?��}���f��DZ,oN(DE舦ϝ��jKR�}v]��Z��RSדMR��'���i��)�U���K�����6�,.ca~^�H��&��ʲ`�}̩�	V�E�:����q?���0��z��?��ɩ��yB�D���n�}N
�<F�$�R+��Y�	R�n�ӂ���u�7�(,�z�%̆�ls���_�3\6��dy�I̟cw���*�,���$�%����i1��>����Y��:Y������d0A�TF"���֎v��X'.]���/��+׮�J?�2����ʎ����j��ҷv��$ʨ����ʮ%Q2��iݢhV�SX����*�o^;�S<E����h	3�U�e!K"iY�A_H;/_b~-��\"M�j�����Z���Y���Gx���t����c��V�JY� r�������iܸt	��hr��L�B�у{"c�%+߃&�f�X�6�y��[�;-�)��Vb��t�i���}֟�ĴB.x�����o�,?��݂�u?�lm�K���gA<5����R��{���I%ꥩ"�ˠ�X���̦e��W�ot4����7����)�4?p>���_ή/�W'�\�k�q��M�!R�4Vמ��?@��������^���b|x�<D�x}�rv��w"U�"�:�4�pq'T��Dq��%\�D$�"|������*]%����k�^\��/�|��������,�(ʠꕲ��i�L-���p�R#�X�!�������[q\b{� 0d��F�a!o2}k& �>�-%�>�A�D�j����� �فT��R�!W�ɩi���¥�ID�^�Sgx<��tR���$zb1�������VV�Tܹ{�M��K���B�����_���7q��+�t�b�6��-�s������[���cnvR8������GZ녥e��g?����Q��7���-o��)����ʘ�C4B[0�����熑���v���G��Q��^�+�e^E��yԭ���!�4�" 1��F�'�l�\�T%�^��w�l�I:���u�ʄXi`�)�.cA�l\�M�?l
Xp8	�,�PЁ�)E�V�`C�cRW�� r�j����`�	��'��סK%��x��A��K/alr1�^I������SF>�)�)X<�"��������مh[�D�Y.N,��JIbk�*P�$w:�[Zy��ץ���酻��)�b����YX�������	�uxt�
��7��	��G���ˆ|���L
gɴ&3}=�v�Zm�'l&`������X%�ׁ��k���,�^�0e��߸����ϔ�X��Q�G���k����ŗ_��J�>�J)��#E,�d,n�a�s���)	?O�j�m���_��eC����ҍ�VA�"�BҨ ��UD#��zU��4!V+"sr���-J��5�p�������ߍ6�4	b��*�?7������kH7*��,�Ӥ���W�͟G��t��Q<s��;0��)� 6<��g�׉��;�E�K����Z�g ��^|Q�X�B�������s���3@�|���'[S0է�+kuEf?af�ö�v�C��g �6��Fj�@�,�d*-S�#Z�d�4./j"N����p���� �8�N��H2W�^��m��,�D�(yl�{����������8�F'�?o6�~��/l���I:�y�^{�Y�'X������g��=����p�=Cw/�����=��pqW��\��t>-�탅�2���֎�W�K���B�����:>��Kn~o�=�Hl�r��U$���ؑf�����!!L��<d�6�h�ܹk<ȹ�6���(.+����C�����b���A��`e.���!ˁ*Ҁ���{��E�_`#�"|qfWƧ���O&���]�iڋ����R� �w���U$�LCj*olr�gT87�6D���}���\�|}�"N�Y���F��)���#���F	ހO_�?اf���Y���HS�E��@Hl�<�*u�?捝�礙|D�熇:��h6��t�k�
Q��2�I,�E����D��Wag�PF2�_+��]�8�C"�E��ό���pp�.������pQ�Ţ�f���1�pbldT�5�?��$�&=21����m�iH��V�������	IYgɄ�Ĥ��nW���#����/+��ׁ�.H��<��@P0�_חR�k��8�=�!�`H� �I&���s*̣TT�$��u�������ū(FNw�k��j�c&�i!7E�/�R�0������I�Wn'Jt$��%�8Bye�x##=;������%[�
|���BqK�BY^ D�ZE8�� ah�����A��#BY�&c���-5k.O 7�}w^{7o=�F�����F?m�ؑ�i X`�	`M�ʤ�� ®|ݚ�y_�Z��z")�FA�UD�شe�҆�Ns,�d��i�A��1� �RiАÐ:�^b�2��ȉ�ʮ�Ds��9E�lq\�./��
�V���G�t��d���(K����^b�U�����!ߋ#c�FO$�����_q    IDAT5-l���Ed&2��\˫����˦�$�Eg��s����l�lBY4�&�h12��牓���5"r���133#�!m`7ww���D�!��ޞ~=W,�DC��N�C:����������!V:�X,�G�r���0�3m���R�pm���&/|��|����Y�:�Qo6#N��3��|�N�-�������������8��~��ܸ�h  �!f�~�٧8��E1[Dg8�v�صŔ�JBL[[� �K]p��(5J
�fWtoa{�4�vS��^���.#$� ���5|~�k�Xu���N��54�e؋uT�cJ���������-�!�΍��<����.O܃(��N�EY1\|ht��l�4�R�J���H������0�Ȳ�!@��:w��6x;cp��a�y�6C�{��_�A��G!����{X]]�q|_�T���Ăm8�>��Ҋ�p/�E�"e��;95�T���M��
�`'��	���4�^�G�Ɋ��=YZTG<1=�����=�/.��>G"����e
H�®�2>�Fo_�&<B�
� ��i�6�hR��3�EZ�y�6v�,�������@���H=���:_M�Ţv��t���L
��9��/����
��^�`hj�9i�{��y��x?��Ʀ��<�������9r��j����_�MEX�2�O��D����)ߩ׵�$��ZN��lmnb}eUa�$D�o�x�y>�ڢr��rk�,[��}<p��5P��k�����x�8˦�*X]Ņ�	�7���w������4(�8:���U�Ǔi�gi0�R+}��{u�*%�
9�e���c"N�Dt:Pc
��h��`5����b�Ӝ���d�-�&>�&�h0�(�}�X���6rNBz��6�vp�8�J�ҥ���w~���*�e�QbD���V�A#H�jM�RVJNd&u����|o���n�R�
��R6f��W���iC;HT%a1Y�6e�:�h~�kkӤ�{QS8�Q='6ԩi���r��x���ټ�����el��qZ+�J6��n<�� �ܑ��M;�N�Μ[/czpQ�_���K�X��w��.cX��a�3�4��籷�+H��C�)uz�����iEI�ݻw���� �_l6� ��X�^�"w��5�������iT���5\Z]����ns,�,���]�U�"��,�1��U��=����ӕ<�=A��Q��3���o���~&�wx���=�P��s�g�$��D��?����w����|�E�����o����D�����x��MtG�����\�G}�����痦/�!���W�v.��mJ�*'��q�Lh��`�	���'܁.S$�I;�E������>�+X��c��������4�ӯ�.��������	�Y�l�(������eA7�F>W�������`i��=0���8I�|Y�ExdxP��V���s�d�ܨz\Ƞ�d��2�[2�k.���y�{B��2x��k��.��p�dB!	a�}���hﷇr������n>{.��Q�/~��t�CC�����O?�Cs��E�QeRY�V�/���W�cN�l$f.�`xtH�������2�g������u6s���{����ߍ��a�VIsH��rY$qp���`,u�<̂~��Cv�$9q
-��	��+��9����6�\�"�+����Y���͗��eK899E&���]�x(�!*���s�|���?�?���9P��I�H�J8�+Q���ZR
��v����"�֦����y ���p��L�L�[g����*��/��"�C�rh��r'�ɗA�&L�H$N�}�;;���Ws4�}qKR�&��[+��(~*��z0q�,M�kR4^�$D5��'g��֏��Ȉ��(0��Z��n��F{h4��|�VVf�%땺o"z��zp9�&D�J�j�+Z��H��b����n;�]HFoGlD���4Gh�5e)�\t���\G�(������=|�;ߓ���M���%Y���_�rS�Y�]#WA��6��$g4u)��~~-r�!�U�`-��9��>�����U}��+e3K�;�-$l"��г��U�\R��ۥ"̆�P-��׎���*��70�����	�+y�YfV�&D1�h���Y��D�׏������0:�AȖ�R:����alxD�z6h�bM%�����f��3����1��v�y>-����[ϩ	a�&4�F�����̿;35���5E2%b~��E죦��^sz�!T|X�����I��8��A���t��,�,ดE�V�^�j =.x&Ѳ�t�P�O7��n5-r.}�"N�_���?��F�/����~����?:L��Ь����2�����|��;H�&0�7������C�`�L!��g��p�ER"ugw_�=���ҕ:��(�]�!�xww����"��Ь�0�;���v�W1�ُ�U���ܣ���%����j�I?�����!I`�o�T�)W��y�׊0�bvĜ.Wɷ��;)���aBA?.]<������S�a�|���X��
v�i��(Y6���z�"����No�|
�~��U�}��/�^*c�{ �����d���ҫ���+�|������s|�ŗ8��;�ه�q~�.����g� �G����&��>�^��澁^5;{G��O~���]�h��Å��ۋ`$���
�wp �C������
���� |H73j�`�!���-���e���Y�f�JI;{|e?�D#�f�`�����HT�iJ���ȗ	�Q.U���Oѝ*#8�a�Li��i�֑�\	m�6\�xI��P'a���9���m�L�:&ֲ�3��Ǣ�=��ѐQIk�&Ӕ���ϸ 9��������Oh�X_���:�й�$l�����
 	��8�d��a�����X��]�����wj�y����4�or"W,�ׅ@0�����a��n���%WQ�w�t�V�OgQ�L�,'-=k�D�0(���s�2���Ҥ�.�j٘�	 ���s�uT���?,x���!�V�$��i��ۇ���{{�r����&lD�HB����Cln� ��`ll���o�o}�DR�U��_�2ￇ��x<7���M4�������^��H~���$-5y���B	��y�F�$M4=�yV��ӌ1H!����`o�z��AM�y96�~�'|�	�ͥkC(YNN�����U��1><�"���f�V�rz��Z%w%�/K\��ࢤ�RW���D\�	�ɛ�<c)����ds�s88:�/��BT�#�.�arB�|}������#����"$t�>|���M<��M5�{#o�07�#�I$����Q��z�h�͛75	�a]Y4^<�E�oB&Ldl3z��� ���'�ã#�$��'�y���WKs��
�$Ƕ���yi:�UO��:E�%�uY{Z��ɢN��C����O^���7^����?�����O�{Ȏ~���舴�qf}u	}�.��F�����F�TGaⲘ�GB����G�IF_=z���}�I����3����*��B��?���rv��Fz'�ӭC��`�>�Ņ9�����z18�#'��'Kr��Y}�YG�\C�1h4��䀻�O�����|��$ŰLd(.�}�Iѷ���K��Z_������=�{Qp;��Nb;}�,��/&G'q��%ܘ��NO�b����+�8����@���lAIA�l>o/^�D�Ī�p���;7-rw>����K����<��F�F�������Ç��Ĺi��廙��GGW���iRf�Kk��*����h׀���ޮ���
o:i�c [��w��Ed1k�#�ˋ��b&e+��	u�	֊�M'�L��eB!V�	�Xq�+9a�?�ry�O��f	g�d��`�-w_�"ҧi4�����������M�9a��}%Ř��
��4��%�N�,�ܥ��"I����ӛ�ʝ�JW1�l��%��*�,��e�@�-w�h� ������>/ҙ����.j��2�����������I�l���	��5l�X���Y$��G	�F�)�Y��?7P��`PM�`�����]��E�UF
sX-)�������bK�9:��S-�����niL�����5u+E�2��sI���N��OM���h��S>�,씼l� _,�677���C5�����˯��F�('1���PK|��G���O1��X*��z��A�#�|��\.��9�G��6}�U�iNC�K@c�x��uЏ�j;�@M�X8���.�6i��$�0��É��f^��T@eg$�5�������y=���x�*J����:�o,a1��x5�b��
a�r�h��Xӥ�PA3S �yj6\���T���+��,a{w�Rm�p��:�N���t#�I�p&+C��ǃ��NL�Mh@�B���ه����Ｄ�[�$�a/�m;��2b�ONNbu}MS/Wׯ_�u,���%<Y\Ԟ:�ˡ��:�5н�-?zF�r``;15���1��4�.�S�|��9��K�2��< �S�ߓ,6�;f���ZiN|&(�k�s�~9�3�������x�_�{�?�[[��d��ޛ�^A,F6�Ě&����;���8:�e!Ǯ�LJ���E�7�.(W(�4�ă�E<�9�A2xC��̳�u�:::ې)�`cw�C*�V�[�?�nw��K����1v7ֱ���;��W^R�e+F��S%J�:pt�B�~�N�:������P��]��K�΃��������ը�@��l,��}�;zp<�Q���Ӂ�ӎNv.;\� FFp��e\���Nwj�Qܿ������Z���.��
�

��m8��ӏ[Ͻ�חO'��q��9��>����5tww��g��a��x�l^����.�`y}��v�^*�2�Lp��%�b=����_�%�w���ڦM�CC�� �ݎho|�0|�6%߰VfW��F��X5�����]�Fb <p&`��U䪄���o�8>N�s�zWL���b����M��(��%�H�&QHM( ��!���O��gb��D�!��4��d�U�)�b�:��T���+8��f��'�S&���M�(O��]�Ѹ#�2��*�ZS,�_$ց��.J|ҩ�|�9qЖ�~�4�ozݚܡ������Ȁ'�@����Xm�*�6neu�ZXD)�C4�Gn��1�R�D,{�D5���P��P�=_��T3
&�I҄fW�g#��#B�MF��-�-�#~txc�����0�dkiY$�QO8����ĉ����k��>�F��zem��c��ҫx������;�s����T��P�O>��<@[�*�-�D+ч:\�AJX�{��ŸgC��;�iaLrb��Z�?z�D��N�y�d�i��������������Cp�vvt���4�U�X����Ң�(��t�E���&�m,a�t�F@]	d��Up�Nx�@�4���l�<�M'��ard�X���K��u�w"��4�F�PB�呔�Ŕ3�]=�ǅ�)��w��<�3�V��^�%Bv�٬��jjVB�t���ʲvݷn�¥+���"L����H�/���ɠD���5g����>�wwad|�c��"^O�����g��P���r�Ą�^7�~�U5;\���\����&v����t��?y��;�x���{���,���Y����7o�A{(�|!���E|��;�uFb��uk?L;4�8�	*�y9����K�^�ln
�>�Qw�$%x����B�V���2>��#�1@�Ql"P�!l�"w���aɣ#A|�508؇����m�wggc����n�(�,�<w�yd���Z��^+v���|��b͒yMȉo�v��,rү^����Q��'?�%�Ūχ����ύjȇ�ہb����\�p�&ϡ��5M�s����T"�f�"�/sr���>L����ū"*%�8=9D_O/z���W��\���6j�
&��1�?��'+�|��e����ܡ�d/�e�¹i\�x����i*��>x_y���pM���0�n\C�� �z�>�g�7MX��pI`k�٤�����AʝQ��E�;� ��d}r"�1
	&M�5V��U�	o���ë���qӲ5E�h�:��C"����\���-#w���~\Sg.�E��,f��}�9�k�=���a�YP4w�N�a&sJ��B;S;�ӱӊQE�V��
'Uv����{Mag��A�,�2�g���p��B��Z��B8C'���+��L����]��,|{���U)�Z��}5S���.���:�ى��>[Ѻ����BRLre,�4�������e�����\A�F�%t֘�����V���^PEZ��/�[փ�wN�-˧��\��&^˖������ө�T6L�	jwK)Z�"􀅎���7jM|���U�IEl��u��-O�F����p����ecN����,py]Y���dVz}���>P�I_bB��������\�I:�Y�>��{�`z! ����#��~����ڊX���>���� :zzQw8$�9N��Eb��=��F�D�Z=�Ã�'XI����5W |]���&j�J��p�ʘj�Í��_5~���ʢR�r�2ET�E4j��E���
ʉ��
������8�c2YYZ�Θ�K����6��KZ�M��ˆ���Pז�����kPz��Wp��E����K���c�	\ggjP3��x�J|�&I��C
3�����\�ب$�9|��.vsgH���q��r�v���Jj�tZ++a��'����TW����;��������~wnc����>��M���+��ɎNbok���'�:����kߦ�1�Kփҿ�i���e��y�X���p��!�+!_j��^��clr�j'������|�b���i�l�R���+�,ڣ!�t�?��~��)V�,b{w̚��s��K��x*���e��˚ x����^W1����ɳ3{hI7zڻ%�!!�7���z�q���PH�Ԍ��#[�!^+�YA�=�r�_��\?�g.#Bs�rk��x4��kˈ��|�1����3Wn�/֡��iK�w�b|p�|'�G*�{����T�N%_����I��h:Z7i�M��V�r:�ca��Me�X[_G�IB�C�E�����׃��Wq��-r�85��i�
5��rjp4�n��Y��V�������Q���Z�9�5�X�ym+�\H��^�;L���R��&V*��2Y�9��NS�>;L(��{�b6�)6�	���PF�m:l)�2��eȰ�Ӄ%g#y��? �D�B�D!�ю���ZrG�d'B��&�����*��DgZ+�Qe1���h��ށh{���������(���먖P�̖P���9��;���(�X��p��54���~��m�]�g�p��M"��7�ixS!��PZU�4�l��l�g���+��/��i����d6�{!�H�1V0���w�\k�࿲:4��Ԉu��Z����|@��ͦ�R���zm��;�9،�:;�̕M�{���+�bzzZ�&����n��ҫ�������gɉ�ߛ�AG{���|6+H��r�$Ս�����n�k:�>x������Δ��;�����ۜ�06����!W#��r�*FF���"���g��k��4�9��G�{�0}�d��:�	^/�Ο��W�[��x���'�{8�fQ�9Q ����s��}qmc˕��U�n��R�nL�`��O�����?~���2ur�t�L��	ȗ�����މ��1ܸxYߣ����Ɔ8+$]ݼ�ք�	9s��?8 �Q���w�,��n��)¯��._��旁-�|�
��S�c�X�pP�P�
:z���ۍ��q����w�ۏ�J
_,�a5q�c���\rz#�B��-Y��w�}�;P�L$���|ӎ����H{�������Ƌ�����������wx����[/+�d�����_�˖;���8j9qj`GM�"���`�&�<wt�Z���q2�T���u<�ҫ����>G�Q�$����w?yO��L��C��8M$�ߣA��I�=�0�x�6��vw���G��F�*�qx���Ɲ�    IDAT�qB�TGg'G��!3e�@Ns����oml>�Qa�:�.�`,� ��~���+��9���1ʮ��Ⱌ�f)�Zg�a �h�M_��.��B�Z���*�֖���TK�VL����ǹ�I�lN���!uql��#(��a{Gt~�xd�V/Tt�p2ag��Ր�5�[��yX0�.B��CJ}��v��hd9� 6@ɿq/�ۍK�����k*2�¼N#�b@�˩]�-AC�(���<��#��~�\����b�R�Ȍ�"��,4��And4�([��d�-�Ḋe!�����p~gy'*\�H�)�I�NW�	n�vv��}2<��G�4���HZ�bL���}�ji�	��P |Ń��0^IR�Sg�����5�-X]ߣP2��'�u�*��Qi�T��H	V'��׎];�u�RF�;s�S:]J[��z}�������-�����"��Z+��i���QJE���j�\Y��T���2�Xy�E�
��5kn�óS�J'-��4M��7�\+�$Y$>�>�uS�����&\���~��˥�-KUd@�#�.���RY~���"���gbb
}�ݒWr@"%�o Hƿ�8K�"����nT�c^,i:��&߀��,�,Ĝ��?�쳊�����_|�w~�s�N���yM8�	 l���/�e�o@��'~�8G��z�-�:���I[�����J�\�Bݦ���Y�^E�i������һN��������-a%���JU�h�<���̵�]��Sb6Q<?qF��H?�{���QhVt�R	�,��Hx��{�V���{��y\:w�&�dUk�׵�������sj|�2ط&a��ؠ����P@��%iA��o��n��}8�O?�D�$M�ϊ��dp�)�]E�r%br#��r������,֎qXʢ�u(���g#E�4�v�L's|p�k���S0ymv�磑����o�;k�x����ͭ-���Ó.�9	w2�Ex}o��/Q�f�m��������t!�E���a*�U7*�r��l���,��I��_�w��-LL��f�ci}?��?KȜ�L(����
��R�X��5�w��	ⷿ�-��>�<��G�J�́|����	��
z0B��C�,�1��J�����;ٖş�v)��eG����$�z:p����Ǐ�����_�E���2�Q���Vk�վ>y/^���P�j�+KX�^��;;vx�RAŀwL7a�ɉ��Y*&�˰���D�[���c$ɵT7!�d;�(��(��Iq�MP��b'k����C���*MITę
���Ego.^����u�pw�i��&��J�6��~Y��;�}����&���f��>߄TT�)��)�{>�-#�8�)衩I�]1m3�;��v��
��n,�k]Ab>w����>�BBW�L�h==�����dʩ�̼fʅ�d����D��I����ѼoZE�r	AH*�.���B�,ob�k$�J���$I���;���>��9Lb�6�����Y�rҥ�1#���!���E D���4�w4���92����"a�~�q˞�k�p���
*���駑+��l�bId-����
u�E-S
K��]�1��絑�(w�E��d:��al�Hnb�7�	'ϧP���&���6lTZ���x��� 
P�yS���B!̜?/r�řs�z*�4��s@4���KOp��#W�Osa��3��W�N�O�E*�j����ffp��U���}���"FRfÉ��ż�X8�m��ؐ��<c�Gi�¢x��-�Ǹ*��ޒg~"q&60�2����|6h�cpf
�ӓ��B����v���-�n�`�,.������p�00����&�ph
�Gp�gWF&1�b�x�P�l� �>I�\AÕ��i�[k��p�#Ԇ��nL���ʥ�z��ՠ<ian֤1g=��sA9�r�	�{͞�E��ͽ5	�\��|�U��}4��N=7Y�d��� �ˣbk��rh%��e�sSӘ���8�N/Nk3	�㠘F�mS�+"�<[�\�j���5H(��愻֤��󡎾��_����o������m,�w;��C7n���/�&8:�J`sm���'h��
Og�#\D�V%��Z?�T��d	��,8�88I�4����/��[o���f G	Kk���O�͝m��Ʊ�H�+��	9�lQ�F�nCoG���oct�O�>w�?���~�u������&�HH�D.f�R��J:�d"�wN����C�9���9tD�Tw�"f��,&]�h���	�G�l��wk/=�7�K�Ӹ}�2��b"�̮,`y��`N1o�4(�rU��`��r�|QBs���Nx��Ag�C)!n�8�&��'#�g���ܪZNI���3�HА�Q|�y:�}掄���̤�zN����f�>��O��ǩ��5� �A�7�>��ɒHj��a0J���M�<�rŜ:]�tz"�Xep�ɾeh�Ԭ��wƢ��do_����N��ds��P-�"JS
�t�b�e����r&$Y���<y(�SM�(6� ��YPfA%,�cljR��hg��V�����I?��L�78���ƏeV�i�߇E��B�lA�aʱ~]���M�s���p1M�4���;�pE�h���'b8�Z����'�GW��Uh)��i�'�|�jڿP#�^�ҍ,)�]��S����Ց�"����B��PE�-���*��t�$J����3�!0įFC��#�_NM6��j��"�Ѥ�w�L�7�^G����"��D{D�������a��L�tE+�u�YH�V96ɢ�;M�"���,Y�,������v��\�x�\��9GG�������nrlۛ[�jM����184��.�TԌ�""��ӕ�,���&"ݝ��r	�3S��'~x�#��|X;����*���4�(�k1q��
��&����;O��������+87<
�݅مGx8��rN;\��HRFR�����0D��hLŪ+ڎ�ϫ!&�`��,��H��>��Y�:�������%[�����k�z����[��ءm%]ٲē��=9B��ݶ�P N��T��012���Q̌O���!]+��Y,��T��^;*,�D�,�D�UlV
\����#�/��8�pi�����7���7^�����������ag/>B���[��#�:���2~��O�Q@_g&G&��J�e�R�"W|*�`'��EN2�<���0�����3���Zǋ/������c��$J�46�W��cvq;{�5��ZL����,�t���g��+����n>sM{گ�����u��y�ad�5lƏ��˜[	*,P�&JL0a7Dc�~��4mǵ�Wqvr���M�ڂp{]���B�P?�����������D6O{��n ��=7\�=C8?<��f.	�g�[]���&��g�%�Hr	o(B��y؊e��Uml"�{��iJ�B�yN�*wu�*�N�f"%�Ž�1v�Mr��QNb�@ZlNx� �<g��x������\MML��+��QWJS���[�'_x��CÛ\+>l��%ƀ��5�l)��2oYו��Cs�bQ$f���eu΄�85�x��X$�1:��>�(��(�F�T@�#��"ma��S/J��$C�-�N�S+I��;�S+]��X��xЪ�`���-Å��qt����@HB��!��}'��;�.�������U�{���y�g�ɔ�
<�l$���SM��sE�qjcB��g�H��x࡙�� ��F�
���&1�+��n�N:PJ�9�� �8�%!���Rמ����BANNz��[�x>;DZ(�i84��mK_dI�Z��;����ӠO��	ggBv�
�7�x`��E`�:?#�T\#�d����M�l��K���n|�\�O͆�Y
�|V�H��q8�[x�����|�wq�I�#�1}�i���g,&��ɉ	�~�7��͟�a��8=����J �͉�39>���ɀ��w�>G����Y�ؔ��YN�lθ�~��=���uc`r�Ã�B��PgL�8���-����q�⁊M�T5{ˠ��t��ز%��t��W���g/^�y{��=<~� �B$-ݥ�n��	錚V"[\�q�䢯��!����o��W$��l�����V��")�;D�TZZՠP|x���/>�T#�+ S* �0�8TpC^ =׉ �d;�ы��A�/�T���f�r���Be�I�����'%{i8����<��oBEO0_��,�gc������ML��򋏾������GcW�\��WE=��2X_[�O�CM�Թ��F{0"M/w�,�YU�y�2���T>`����N�&��+��[��f�M������>������������%B��
��+X���n;��z�V�S���*<$\>�e8H��8uf���I�ౠ����9v���rDb{WN�C<���1ɮlo���5F�\%��h�$`)ӎ�p�L�ǋ��(Bm���%<�\�v∫4= ��\~/*��/NA�� �G����S%�p''X�la3��7�=	h����rY��6�Lv�,��� �\S�Kbw&ͰfQ��r�t�{|~M �R~p��Ɵ����)�P�J=!j@�i���#MH2>�W���h���#[ȉt$G*�	�H�)���A�p	N��sZ/򰒑'Z���gy�'3rZ�5�����PnM´�k#

*�tE�0a6��XGZ�?�@���D����Dɑ�ý0{�\��B��Ⱥ��Q���J�r&!�md4>`�>:�N�GX�C�_���i�hs�I��w�$9�e8��.S؝f����or�CCp}ڹsb��)�a�C(��H�c	���IG�4!r�2IY4�!�	�9��M�-�2��Q���C���B����E�B�6�l:ihB?6Xd�Ҫ�f���9*���`��
�s�dFh��M�혮{�T�Ťx�g5	���ё�:T��v�_YYR����
����B�����h�N�X�$�`�xY@6���o�տ�A>55"�'�8�wv�����q�T����!�Ã=M���^{�u�=�wv�������ٛ��T��i'"@�6�rN�
r�Mg���m<XZP����(9(Н��2M>m:qա�o��`Á�h�z�e�r�9�'��>���Kd�C����^7.v��ZҐ�\b�����crNhq,kVr(c�o�C��!D�*勄^����阤?�K���RQ֨�o�P�E���I�i71����v�[/ML+4"]+��'sXN�㰐F��@ى�E�����]�B^�"̐_Ӯ"uz?�����"�����l���;{GcL�>s	�]]�W
�X_�/~��ꆆ�{156��?��%�?m�X��v��f2��}q���ul%?ˀ��Wo}�MLLr/����*~����h~�'�#2z�TBBN����vU��V���	�����M6Wӗ޵���e7��h����!�E�ҋ�7b�R�ѡ��	8�ҁſ˩^׺�ch'J�/�=n��Ş@v~M+� ����9ܚ����v�؈�b/q,h�Dݨt�)���v���I���N����P.@wjyA]�Ĩ�kTjbt�iy��C1{���ͼ�y��k��(T+���!'��/�������/sZ0�cS��a�\��(�����Ø:@Z�yi�����")�)U�-d%+��bϲ 2��]4���3s9�sY}��jn��E�GR�ۭC�v�,����(p�/�$"'���;i&����t��!~���c1�ӗ�:*U万*��F~��C��������>���2v�*�#����H�%C�S�af@=5�ĩ�0''Bvd�sZ׳D�D���6;JyDʷ���j[٬��Xh��ً�����i��1B�8~��`%)e��
S�h�X�c�p:�D5�MV4�j����Ô���ԗ�S�eB�[&"�RQ�*�.l�x=�w�Uh�*�������2��+�N�A�/��X_/�?�l���$�f�泷p��5D\>��o�����K^__�.uk�:I��$,iAr�=���;0�g�W��e���$9���տVc�b�I���@�_G6ql�)ա_2�N������{���W��-qr���y���s9u�D�R���\6N�W�/![N�w��Q���˛k���]��G��I�j�Ip�1ֵ"�j�9}�\��C1|�Λ���o `w����w?x�TB
�Ǆ���X�{�rC�F+c��I�ju�R�	�Ŭ@�8��0��Z��&�4����?7�P7ɠ>��PG��.8C~��h�l7�o~?rc���މ��1�h��2�,�M�R�<%�i��&�n�"x�򬠹I�8!F4�#'������ݿ�������X�����w�'��t���Q��w��1�������#*�8!�k�ȡ�ʎ�N8��$�q��Y�R���������Y��X�x����_bucgI
�=�����N�7w�,N̄�����EL��v�n���"w�ԅ�A����ÜP!�_���JG�����`H��R^��Jp��x;1�Y;}x����p*�(���OE�?szr
�F�e���iC�VA�Y64aZ��GpWG�P7�ݭ@u����M�PLg���	[�k����Q-���RL�!��\/I�K9�ث|�Ƞ��88��)��k��ØA0l>?�Y�H�\2	5�e����=&���Kh0�����N��1�|���(��L��B��B�t�x��͞���a&�*��� ?7_^{��i�Ű�!��$x��mM�,l����L�}�����"LD�60���(�f�M�&~�,J���ǌb6V��.�ptx(���^SRO[G�}��z� ��Ct��k8��W��9�a��ke]�2��/T(_?CM���՛z}<`Zd[��_��ܴ����=v�"���p�xd%��mB��P�ņ�Rd&kY��Dg�Ts9بæ4�E�%�
�U�n��_r4gSf��!�t�ǩ6d�_�|�)��H0ҦF��"�gL����ִ�Øv���ˁT�LɁ�ņ��7���~xۂ8cRR��@[D��[Ͽ�g._��\W��eC��o�W��y~�3��� HЀ�Y,�U�]]�mu�Z�R�W3���؇����y����y��5��V�j���Ѷ�-�N#u�7,=	�$@x���l���^w^F�PB�.��y�9�s3��}���y<�/4���H:�"���V �I	c�����q�؆{��������Y{3O��,����"�*���T�P �ty�/~�Kvj����RE�~��-}Of/��X�*�VB�.�&�!��׾f���%�G���{�΅d`_ /��Z��Ԝ����^9���zے��M���_����b�`���g?���'���f�rQ##�rug�KDw���nb�YW%k$&c���!R�S���:)�I87����;g��߯4j�?>.�> l}C�����������l�@g�̄&�GeD�r������=�l[��f�0�������������@�c��P+W�������o�����]z�������,�M�8q�^y�6�۫ L;��~�e@G�l��qK�ڌ�&`(��\\́�A�pmٮ�߳՝����,Wl�k_��ұ��	7l����������~^6|�;����IB�^��[��d���
���K7��||�,�O��7�xH���D��o�@��BQ�p�Z,Hf�/�j~�E1�E'u�����P��
��X�2��y��ٴ4�	C��ѸE��h-�N�U�?�sI�1Wp���ħ�Q���F1��D!6KAw>+Y��%N%
�A"s,���M�)x�n�������B�$b�/��f�õ�.�f�R1�w���atg�W��i�[&�w�#�Y岲n� 6��5$,[�6I�Pr�J٬�����gN���8:���: �P�� !�i]�)GC����k��YϘ�!yE��8AJ�D-��	�T̃9�_x�E��I���	�@�&]�x�1���S�������4�go�tR��{
����r���gIB PD��&�w	�əˮ�} ��CZ;�cT    IDAT=:iǟ~ʆ�S�=i4��oTX�xf�u���`�`�i��mQ%�VEnb@v��=�03`�DI����	�$x��V-�x��9>-�~�YEp��C%V��yNz�ՒHiV���鴒j�!����A�i����\�]B���Ϝ�N�)�����h�������]{�������4?�*���m�JEs���!̈́��_y���
�������)����v/jmR��^eёAȂ�1���O����e8P�T�ڍv��%����`�N&53�Ym�mko[�er�}������⑘ݺ��x����g���f	k�BVA_ɱ㿋Ϗ�;��Zv|�}��_����Y�@�y{o[hd�}?@���p��<����|�e��=�� �� �DϳF�*P���v��������[	����a�FF�4�����U����~�PR�0�n���S/����\z`˹]k�#Rs���Di�s�w�k�Z� 0��$�C�O������o��ԁYz��׮�����V�	¯=���X���l%bT�F��ء�R$��=��H��ا�5�\su�n���Z&gۙ�e�u{��/�׿�u;<9a�P�V�tpb~����ޮ>��j�u�;�-���R�a�SE��Yg,�����0\B ��] �����LX�]\1d�|���L���Z�����?$��F�W* 'ڙ�0q�v���u����q<���,&!�i�km�rQc4��p�p��6���Cu�Y���84� ԙ����ʖ�����T�jǻT+��kO�]p�n��o[[�7}P�j[m8��jqB	�6qH3?u�5#cXg��8t���d^[}�6�K`���NR�O�H��qhUr���9'�pM�|�UU��&0#�P}�ݷ썿��ݾ=�k�K����q����۲�S�3�Դj�h	|T�8 Q}sRWk�e�I�[��g�U�|������=[�p-i�qLh����8��O%8�wo�V�}���
4��[VAh!�(�5��W��˭3��Mݨ;7�!�I��>m�Ϝ�xO���H����1n �(����� ��6�9�܄�V([%W�8\o� �@|BSc(�/�N�y�x�&�L�E�d�f�1���)��������+U[͚T�|�B|�-i:8� ��ez��*nT��I�>������G�J&	���׷��V�n*�>���ҽ�N>ٝ�0T�h�ҷ��=������,����9�[���4c#�
��6����^@�x��	�!�P�����ٰtO��և���Z����_y�^������ݵ�>|�~��O-Ӭ��c
6X��<�"�$J�,$��d��}�˯ۗ_~Œ��fs\Vjeʹ�վU�aΝ���q����Q���^�!��Ru�����t<І/9�D��Ѩ��
Ѱ���C�f�C��u�+X�wzy�r���6�yn��v��]��8oŬ5QO� ?K7%&Zg�J��x�0A�=�J"Z��v���у��{_��[�z�/��ꥻ7wnqy����}�3���I�Z���w��~���X�#ԡ�5��ߩ�#�����pP������9[�ٷ�s�������v��!������l��ڥ��X>W��'O���D��aPk��rJ4x:\�|<�1*b� ���[��4��!3V0�?�Z��R&�"�@�"�!�K�^�+��5ᤪ��@��;���d���.�d)x����jMHZ99�1���<��D;�%�mP���%�1m�p#`��,�>�Z�������g�`'��@���ґ>���Ă�:Mu�,�N
!�-!�B�yF �=ҡ��%��)��� ��}�_���u��Z�O�#�������Z&g�lN�B�q���N^~����o~�NM�x��|�g��o�쭛���K@��i1� ��>&���*U�� �J����4�5!�^<{����x��=�/Q�IG�s��8(`b�����nY��f�ם�9sCGh�SU�9�[�<ZR���P_�>#����hWSeT��Jm�!��A;��3v�̌�	(&�/���*~��%�Y��;�Tp�a�r՚t2yiSS�8F �f��OӒl�fi��.�tmY��B���=>% ���y�={W`7Y�0�!�@��|�It?�t� ��<vLr����P0���I%��W_�ހ���t���o���as��R7C&��K�t��yu�w�L��ތcz���~I	������o
�nY(���YAPv�`A	�FH�����\b���w�֜"�nF�K2����a��TwZA���Y͜�}����+�}I'��{�����w�PnE"�@�E�&/��!uU��;-h���/~EA�`��bpA�ټ;���z���Y�磂G���+~$C��~�����fvNv��x�}t���a��GE}�3�W��!�CN]����(h4���>?�`̈́ז,�k[,$n1E�$O)f���,�5,G%\oi=$bkWꖶ�����{_���O=���}�򝛿{���	*��~�&�[�U���N������>zL�`�8�BG����0͢�}.�lj&���g[ْ�jf�����W�ԉ)��Z����~�W�J��ɗ����9sV�wUU�}�ȃl�e'�G���D�1` ���k��d�	����8�
P�Z�����72�Fk���T^�!�bӡ[T/���*B�ZT���l�0߯���Ʋ-gw,����� K�O��kB��y.*5�hc0_����r� ��@��ׄ���C(7���VsY�>�;����yU��2f�1_��?t�t�#�Ñ��{���v��.C�v��)�#�e*o*\�����Ύ��@~��Z�����cD`9c�p�����B̃���lsc�^{���׾.IA2m�7������[v��=6Z��}��5
��� $N�u�?S�,�B�	Zyl�@Kh^��#l!��c`M�ø��R�tg��1)��n�*'��9���a�`� ߑ�A�o6���������<dk�붛��^.+A	�X֟�Z_�J۱3�������a\���m�ú�  Q���ܴͭ����]�m*QNX9|��+�"W�J�PQ	�:�+��4ZjK��4sGT���I��j���J7~jzZ^�T�w��)��c U.�`K@�J�9�f bO��\��`|Be4<0h/��j�����oh`��	��G}h�_�Ю\���θ�
�D_�3u���.��D����L���C>�V>_����{֍��I�gJ�QCf4�}��E{��9�	�PI�zzm���~�e��$�x�k��_�����ܜ}p���Ϳ��zY� �<r`����E��*4A�.�|��/�f_x�e�t1y*ʚ��S�Ӌ���]�~�Em���4�?��ǿ;�w�ꄠ���y���	��n���*�GE���$��
��-v��Se�W|ڥ V��dZw8oזl��{̭'kd�g�@_��7a%���jK�w�����~�;N�����/�������z����{�h�$T��>���cᶭ,/�_~�/$[9>8dgO����N�� Q%ж�2Ug�ɡ
E��ڢ]��oK�{�_�Z�ܲ�_���gO��h�iK�쯿�=�3{�bє}����le|d�,h��`Zr��������H	Z��VH,}l ���^p��Dq��Ǩi�j�H0������\��5) �dӏ��VK�b,� ph.�n�G�l~oݶ+N�G!ւ�B���!q#��3
�-	��8R�v�-��m��m+m攽%��m�z-���'�!x�UA�K:�]&�22p����c�ܰN1z���+�
C:��w�jMGܦ X�(p��!�����E����e�`�,�p^�♇�����Oqk��9 k�\-�5�K|�s/���{�Wu}�̞��?�;�n�r o�͉�_ɘ�WT��Q��uC�\q�1]�x�O �3��̮�}O_�*Ԁ����Z�T̡04����3뢣���Ea<� #�L�Z�{�>�.-�yp��9w��^|�����[Z�;swlcc�Q���,���1IL<nc�����q;~괍O��.�Ҽ�ԇ�y�n�n)��_�/ܱ@�S�1����-�+��t )˺��DL뙟ת.Y 
��K���)�����Sglj���&l��]	��"��x ������- k�D;V��0C�޹�hf�k`j���^��gft�"�jt<"<�w�{��x�-�t���7�-�g,��BHF��U'�vx�:��D�&?qCx�
�g��r�7oж�4�wT5�#YY�q#�� N�C�~t/��0)�����TŌ��7��u��k�i=?x�h�]�h�w?��j�Z���p�NO�ׅ������\ޞ;^̿��U��V�ͥݟR�Ut�)�:1��Z�P��w���.H.$�����tgB!��0�0$e�s���J���H�G�����m�T�Ę`ׁ+�p�e;��;[e� �:_Yߜ����.�k2ޗKm~&���"����?x��?�����?w�.�����k����ʌ�Y/|^B�X��w6�G?����)?u�>0)�d�C�h��fMU��}ͺ�_\���nٕ{wlu/o�r��2e;s���9*�x�i�ˋ�W����;o�`¾�_�D������j��=A��� `����)�T���*����F�Æ�[#2!W[��c���H,���!͡�D@�G�p�.�AQ�(�� �e<���/�����1�*�2IF�W콻��a~G�y*Ḩ9h��֩(Ua�GGY�=�	Ph�j_*6*{�[\����ś!��Z$��1j��3+ּ�-d7ǎ����i	�Y3-�F�v����= $B���RD#�f��2$��f7��ZiG�ʥC�����h��y�MKPl70��,�4�->�9��LA�<m� �RMN68�0��«��9��l�O�S[]^�̉�"\Z�t ����z�"$��A��MpH�v&���q�����$��2X�z��G2�H�(��t\F�|���٨����� $TqT��x�]0sdf�AXn.���^�<������L/޸l�~𾭬�*��dCk��E1�{mt���:3c��A����b������@6��zM�LX 82�L��Zy?g�\���u\�!&p��o�(��.K},��d_	�r86����kǎ����Ӗ�첥�U�;7o�����G�-�j��3)YS�ϻYI1�T�u)�7K�HZg,eӇ������˥#����˲�%�j��w>x��z�m	�E`�i�p^ϴ��ԭK��U%Mt�|�o$c�Qr@�3na?�O�k�L���1�3�1�=�o����hع�9^?��u��A��bQ�;��׾� �z]Z^E���7
:����p(�x�ɉiH5d0�(Ul���Ɔ�l��ϒ��L"�(Vu-0å3��\���t$? ?/��$��LQ�{��R��Q�c�
ߝ��ءS���!a�q�P�U�;��_ݫz~��Wr�k=q��|�JH�Vs�_�(w�*ш�^�YN��Z�[Π(6��� �g��9���?���t����Z�o��wV)$<q��1K�:��3xg.����rs����;vg��kVn�l?W�S'g���<oSG'-�������S�w��a���_�gv��sʊ�H&�ֵ��()�B�v���5�
C�G�<QC�W-f����c�;ަC���/F�W�l��Ӈ�Y��P���wՎ����%e��
L�R��
�}o��2���~�,틯�֍K���m9����������d� ��z�(����jy[@���e�.�[}+gi�X:W�꜅���T�\> �J�-hF�\�_�:��R��kCG<�A�*��pH�Fy���D�/W�1^��4 `c�M��I� �����g�В�A�@M�۬6ĝ�uhR�\@`uS
G�9d�F�b�^�ݭm��Q)b5�sN/���S��-���<F�������JK���҂�o�8��,��	�T�PQ�� �!���N�/��K�5ь��f��h4p� �,(��Y:-��g����]��ao����,ïm\��L?��4����\��M*��T��`NM2K�o&�>&xz�^��Zqg�j���5̓Q�b���	\|O��܋�
�� U?�F���ѩi���Pe������x'��jr�Z�1� �%f�$�$5	ǜ�C�'�h3(vo��Dr'Z[^�5�b�<�|�}��E�t���c� �k2�U j;�	�u*2�t�p�b7��W���Rg�p�;^<���`$ V�O"f��"Rѫ�CACE�9X�c�v]X�>��N������BJ4.\�b�7m�弅RI'��@�/�'�)]�m��

XP���"�b$`-3\�sb�����FV����&*�{�o%��㽶�F���H��J�a�vC"3�Ξ��@e$3����_�%�$���`j�x��]�VC2�/��uG;dO�A�]��I)E�n\4$'��P�����o����}�S������O_�u�����cE%L��CV*f��ޱJ1/�сa�T�/fpN���) +E[\[��+K6��l����!E���3��s�m�Фu�h�l���?��nZ$����߶��3q�s���O��G�U�B��A�ꊮE@��D=�.-���n��Sq�}%��{�#�B$���	�~L�p�M��v�m��C���V����ԏx��#�:@Eb[)����h�';l`h����-��W?����Q��ʢF��T�U�Z(\���τ��P�̦�;�y�f���������l�����o�*C�&s ,��wJ�9���Ϯ;�x���t�ZD|V��_�c{-*e��E����4�v43`cn�+�w���Ц��"��4�X4w��6t�\S%���Ցhy9�Ӿ��d5#���m2*��WXy �ki�+�֔�(Px�y{L!�8��a�豽lƖ�V����Fl��a�3� `5e{c[*#��i����Zo��	wt�8�Oba?8�y�����ܼ*�N�A�I�h>d�F��|��C��g�ˠ��<���p@Q!>rԆ�����!��Z~�*m�:48ZN|�Y�[	0����Ѵ�^���᭪�y��BI0 $�HX	��.�A�����G���P�:$Ź
�c"�J�bI(oTԎc
�Vҕ	V�HMZo��b�� �1���ĺڮ�Һ�5�����#���-d4��V����U6�̍ <��H�moMSI 6^������j������N�i�؂�VP�u�N5 V�BbQ�x"�0+7����[G(f�GI#h�]Lr:24l=йBf��v��U�����rRI+�E�2�=I}�hm�� �A�%Hk, �k$3ҝ�>N�>~͟����'����j���<*��:��� ���qw��i�<=m��ٯ^�����"�F5IS�?9��h�����OtC��G7�N!�U�EG\End�~���I�;,�hx�����#���~���|�A���w�ڝ;<;w�*�/�����Y4�͝u{睷���W�����>�M���
�i�#Ps�2���m��
P�L�v�5�GϴR��g��W^��M�hFG������z������_�S�NYG"fW/_���yî~����T2!C2Mf�����"R�:~���?#��`<H��d�JE--GMqU"т����xԆ&'D��4�g��jcC*]T&(�����yQB-J�6Y0�����İB��Y��f/ۭ�e�o�ew�����dV!6�`��iƨ}�DDX�l ZI����V6m�����-RA�%f!��2�pmѶ�ɑ�.Aח�Tu�3���>��A��8��h<ꂸxپ�X�u���v)%I7�fp����C6�/1`~A��8*V ��e+�
BD�y��ɬ	�f��>
S,d��BX칄PmF�̓֕L�`U��SBG���?{ �.1!�����{J,wr#�GL��3�%�P�5����OM�� C+��h ;     IDATmk��T�:I���̜;`v��Iݿ��E�tᢵKUw���X"��B׋/�d�+��Ï.�����I�J�� %�aZ��*dJ%?�(q�CAqj��h	�x�y�7mh0 hJ��źC�����'s:�I`iG{*F�{ѧ�l��[��2s[�4a���D���a[U�u�2`"��(zNe��>sW��8�p�D��q0�@5>>j�������>N�������� @⿄��W���ޡ�S��e4_(���C � ̙"�=����f�������?2)1��6�6�|�z���
(1▐�	q�c�{��9�mm8t�o{ż���I� o�K�/l>ɀ��Ǩ�P�����c
�����J<%�ޘL�':nrz�2��E�f��yRlY8� �T܎��L��/;ߪ�#f�o	�0'e��ģOQ��&���
���u۪قU�Y��B�xh<B��3e]C�nVlm��֠�;�!�@8��z������߾�ῼ����w���;�󟛚>i�>��t�9H7v������L�U�(��%y���#��1��z��M�q3���
�i�i��v~�}��svxd\�,�?��mv��2�_��/�铧��3e���ù����f#Ãd c�f��0��޼�>hG=uzFAx`tX׳�����U�W����<^7�G�RQ��z�v�ښ� u��������!��!�Ws�"6#@��ݬ�����ĸ�N�X�*6��HA���e�u+��֒{���ʠQ�!��ޣ%�܄���{Ô�������7E�O[�"�x(DHZ^{��\U��&���9|���������tGqld�:���-@ә N5��u�A�����Y�'˩���;��������70�9RЩ
N������3\�b�u��vt��I����uZVf�uA�Q�kM�Li�zj��Cxr��s@2Ao�X���+�����lykUm],��=vhj�U�M.��?&U!Ѹ(Q�@�9z��AP��*	Mf�'PU�ݓ*���js@��������r���ns{K���ͻ�C�$5H����+�יp���q��5Pu3m_O��J�^iu�Ƽ�G���!kK7�b<!u%�d��H�ũ�^�#ǎ)�#@��@.�4\�P₨#�$I�t�{�����_�=#
�؀!�w�tO�{�9�'c�Vc�.�	 �%]#��¬+鳇]�@G+SUU�!�9�f�%�Z;��gNw܆�o���-�<��d��� ���G�^�YJ�2�!3W���%��`_�"�t�E$�.[�D�3p��n�s��< ��%�1!TдyI
@�W���tư��ѝ��y�>Tmd��� ț��Ȭ��Z���3e�Μ��6��=���^�k@+�B�g��oC|%;�	���"kdrf���f������#T�fn_m�����`$wP��G$�)�p-h���������G	�߻���kw����{s/� 80&���֪]�v����[����5��^�F�����J�D�bj��M�$b�,ڹ�g�;6qHY,�6o���-,>��/!p~�D�WPq�X�n��#��V�L��*ts}Ӯ~|U(Q����3�k�Jb!����ҌP���,bi$�M�C�bf��&$�R�Ж��Y�U�U3���R���2���� ����C)J6y�;}�:��,��ۃ�e{��%[���>�TЎh� �IP�H`,�Ӛ�z3���V�����`���ֲ�]�#A��O��6���1!>���Ƨs�lߵcE��ޠ:�mEg  ��;�:�?�>P��T��Ħ��ku� ��y� �n�P@�J��<㖂1|`�,`��B(�D�j�y/όM)�hȺ��֝�ZT~Y3.0d��#o�Tň��S/h�Zӵ�&��Kn��3�Bs֣A�u��{p�BH�R-'�@����Զ <���%u�c��	p�=�M9b�[�%��}G~�,�ӝI;:y��y�h�G�RIk�� L�T�� �BA.��>�deM�h�?�b8���$�R �`$h�h� L[Se�K�\A����M@��%PN����5��-'�a����{T���Z�#�%mP�ۄC�"�9GZ�x�RY�)f��έ�4#��L�ì�ψ��������s�I�X+�uI*�,��=!|9����,���_�"��djy�-�)�^�_Z�`SP{��Ʊ:�oW���<;�O{4��K�%�^k��dqu��ڃ�GJT�P}Pl��`)8���լkh~b3���"����tJ��%�cl������)ºT���3�7<ʦ�}}xY�R֓���vh�"�G�lT�	�f>cۥ�m��C�#&	�?fsx���u(ԩ��-�[c�*��lמ;��li�|�m[��0�G,��+���)y�����e8\�����������.�����w�x��q��˯J7s���U�q몭����ڪE1V��j�7J5���J�	4����'�twZ(��j����I{��Sv��őj��U&GE�����ã�Nu����ڲp�i�&ɥ��*#׋��{O�F���(n��:E	h{sS�E�-��1{�z���F))����uxH,��l�n�U��m������D<mC�c���-�hKp���S�NX�U��̪�w㒭e�-[Et� �:���2T�6Ί0zSo�w� �\FJ�GήnZym�b��%����e��h�U^귎$��D@@	�E�,@��_��v;�d߂L~�I�Р�fc�Sy���W;� Y���k����Ek�Ϛ��}�~cx�rm��ة�/9�w�PP ��ǧ����74~j?��9 ����!��ݹ5kk���R4�D̞9t�me� ����O����P!�,ִ�����<�v"��Y��G@(�t�zA���{��'�B~��`���c�Ц��ǎY%_���e��A~`{�����@�>+Z�J,������FBU����=P�/��|1z��%H"%K��q���a���ZM��P��OP�!b��Z�a�x��������K۟�Nz;�S&�w >*J*@��'�@���Ǻ�[{�h{�0�(�:	y!��Y$�I8�T�^���>3c���%�=�����Ċ�\����]�r��PԞX�?�P�Ev�B͖�@ͮEU�Z��
^�J�o�|����O�c}��3������+\��y��z:�&?ia�)D�Q���������tB�=�g(�.�"W��=Zc2]g�$K�ϛ�@x�=ɍ�yѸ�N{mo񿱍�+�j:f<O�D�"��e��e�̫����=�Z���l���Z"lt@NK��1G���\�#h�Y:�V�(�{_"%w- ��]�P#%��@"�������G�,�G,�hYo0v������s�q�����MQ�����7o�э;w�v��q��&������a��^�G�����.�d��T�C�q�ҨDA��'�
/�#a�XX3��c�v���L��h8d;�;v��%���T���3�ڡ���D���۶��vv��ꖊ��\�qf�i�܈�h����' �CiUP&�.$iȡT�2���<��c�Ѱb�j�Hܒ���4����B�(N�^~_t%�n�����E�#�i�x�b���T`�:|�N�<n��+Fk����ms�
���[��`n��7� Ԃe��x�J���59� �g�K5��ܱ�Gk�[Y�P�n�@Dҁ���P�^P���~ˉ���9$9��������
��� ���j	ˑ�Yr�\{��}��d)
����{����9����Dϙ��A�����%A�j�Ҵ�@�#���O���3�Q-P����Lg�#��C�^Xxd�}�U+��&��k�K���z�v����>���0�=�kx��%z:-�ե�6��F����94 t�u��EĂVÙ�޲��a;y��=}zFZ���v��[ZY�Ÿ�DR]!��If0����M��P��/ ''��l^��T�ܮN�P�|�2�eHO����3T�o��8M8���ѧ�ц�+���n��X'�����ĚB)��+sdڵ$�$�B���փRX_�S�j:)G�aUV�g�Qoi�0��h�c��*F�R�x؇Lx3Z�9�
���e�
Њ 瑌���%��$�����5[:�d����%]x]'Uyʒ1���;9������ɀ��%¬�_����i}^�E�c �A{7\#�Ͱ	R���Ҿ]��M��Ob\��p�Lymj���Б��P����^��0	���hDi�Z�_���}���m��;�Z�A0���Ϸ�*�Bf�./���ΚeCM+�LjZ�0��B�{���@��9�{�I�f�.;<qPIt��rA�s��g�\/�,�!�����u�7���������_�2p���߿y�M���=��M4���}p�]{pN�Ն�Qɗ-���6�,0�ghl�z�,�j�V�j9�+;1u��?mgO�(e{o����[�\��s�<m��5���y�ݻg,0	K��\������q	2���.���km�J���������e�N%�q`!���UmK��K%ThE�Jym6���}pᢕ+lR7Q��&&�r��Q�>y�����,���#���E��ߑ.n@sD���2	��tP�2�.-��c�t�2���J�(��(��-��²�<\�v�l�&iSӒ�`��$`�'��S�W/�%�{
I�y4:n��eNˬ�1�	�W"�3�y�Х�N�9�֢��}�g��V˚��y�HHk*��p�EH^�N�	�3s>�N���|h�PF��1
�5s�d-,9�`/�G܁�����bթ��[���͚�f5S��r
¹f�"])��v���9diWv��d8�5IT���//>���U��{�b��}vv�=7��sE{����W�7u���kޕH %�fɐ��c�H�iA�sBM��T��Z��N��9��=��N� ���}>����'ڦ�:�J���!ϝK�&�G�D�}�� g�٤�`�|ˀh�5���t�:E�?��`8�Y%���ѝQG5c,�Mص�ᜣ.�H�������_�3��$�S�Sk�_O52nQ-W�=9��W��*`9M���i�{��0�6p���q�.�	c��gN �[H�	���6@��]�\_E�G]����n������(����_BGN�A�]��'nf2ˁU������j�g�����~��v��X
���S2��4���х��_
��Y����vec�2���"�I��u�ydfa5D%��gj4�3�yH������f�d��4�θ��_��2ˇ]@RTo�ƞ������~�b��裾k7���{�<u|�>s���i��]�p�{�`�ʹ������R5jT�e!����<n��C�����6~��m򶰿m�F��M=nϞ��3�'��w����wmimI��8ć��v����׵�V��X� O�#���a���������u޿�XĆ��V,���,��S�W���N"4'c�`�WQ K0j�Ŭ�T�p�AKj�Z�?��67w,��[GG�8(�ܟ�>sƎ����C�-����#�[���̮\b���l[��b��8v�mٖ�K�Y�����f����/��I<�ְ���YX�V�dI�d����H{Ź� �Q���F�а-�" Qu��#��p�A_|���e�������C�)e�q���ţ��0��V�'a�6� ��ô�\($���X����T�� 'W�A��0ɕf���f�R����_��B���d�yED���s���9@Z�s�7�C&�L9gk�]!7U	3#OD�CPR"a��8dG���~Z{;���m�χ����Mi���֟�S����3OYi/k����͛7-Sv�c����CR^��Mno�x:���̛ۻ���b��#�gP׃���=�p��s�}:��
�6J�9	��h���<��Z2�z\I�2s�{ȸ�T�ݫ-��]�u����[Y�l]��<w���T�	�
鵋�U�Mt��]�|Q%���m��p�	���9o�#��Е���灳T�;c 7��j��IZ���p��4��7?�'g��x%N�O��r~.
���0�BZ�U*E�����+��{���F[����*>�&u}jg��ϓ�F"�$ʛ�!W�H÷��(���w�m�z�up�v�	��37������K���e��S9!y��$��O��*Dr��=,�ڻs7��E���V��E�˧$�|:Mā���s@{h���VJ�:(� Z��9�.�&�0 S�|��b͖�FwN�����w.>y�!����z���[w���콹_<>}�^y��6:<����ݷ˗?��G���V%���%� �*��L���i������){��e�7�hZ�V�Ƀ��矵��O������G��åG���g_x�&��F<�u��޶{W�Yng�
{-L��y�̈�%��F�Ri�UF
��#�� `�	o�Q�~�1njV�K�R�d2-�t�1M�";�`Go��$�q�=ܹs��®o����`$��]>82`��M��E&p�����5p3<�8!�F3`�
�����S��1K�X�#jŨY1زF�U�p7��7EU
�B�A�!���0sk8^0_�9yU����: WP��v��y8\��fV����_�w=@U4� D�?W�xT(o.	Z�S�~eP�T��2��#s��3��N�������_�n[WGJ��iO�S�F>�U@B�Q:\/_�Ci���b�N0��⋙�ڝ^&�&��+a	�[t�0�K�,=�o�g���"��={Ξ>}��;�V*l~i������F6�$����?���!L����A���sV��m��=�y�me���<qlJ����݌���JD@asPvB� L�M:ܾ3�4��
ר ��?��T)�mf�3U�g�$���LdU��\�}�n�O��C0CA7����� γV���G���u�l�n�{�f��R9C�����s�����~��F�N�7Tx8�nd����N�����o�k�k-�5�J�Z�D���<���ˠ�$8w6G⋫���P��s�؅�+�KWѱ)�D�u$8�ԡ��!�g����}*��C�����mb��L�s�4�h��q�s bO��#���r����9�Ɯu�}�XU��iE+(#!�}ٵ��@M�~�n�g����5��(�1>:�I��E ζ�I�YJ��k��Aq�ޙ�iW��-3+�Ú	�$*���u%Oy������*�����*�liћY/�wh�G#����[�8�0��~n��?��?18�[���w>���'_�s��^yg���7�h�޽_8q���K�0��ٶ��X���;��p�J٢5�u�9�i+r3iÍ��� ������l�J�K��>xȞ=s�NNW����mo}�����^�����؄u��6?{�n\��ޚ�r&�P��d���:�s����(+%ب<Ģ648�kwc�J�a�z,|�!�;҅���ba��NZ�Zr-NT��szx,���.�Lu���m"��ٷɉ1��C���,/�鼉�q��m7���kv��Az5�*�
�^�[]���=[�fm?д����z���NY|���}��"p��������f�V��,��!��H̊uO�O��U�>7��Is(�Tu�a跒@��=�b,��0��G=P���kR)gE�D$��p�:�D_�h6@���jC�`�[+9 �'y��C�$���2��^����ż�!�� D��: ��+����*a�d��c�l-}-Z&�Y;0��,	���m�N.eՎ��8+J2�*��瞶gff�U��=����~������d���i�b�1�=h�'��s��Ze?��~���$8��:{%/H�:��- � W�d���^>+
Z�3���hFº6Q��u}�/g�k�$U����:D#�ٙ��4)q^=�Qw��\�T^�i��Pϊ@)%:O�=�{��g��;R60<�%f��� �ǣ�WRdC_��Q>5�d    IDAT�̏�����(PS�� *Q��j���:k����d��JU�'�d\�V�ɵ�֭�������Ob�p����K<D�7�g�PҸ�'v_YM�C��3��Y��
.T�b)|r��fኣJaL����ą����{z]����z��Δ�d(�[��R�]ZZǝ �s���X��(Ja��Jֿ~���P~rO"���
�(��I��T5���P��GG���P	�w콇��ޣ9��$�	Z�V�LٍIܽ��5�J�ٻ.�f���č�~�K�|A����p�H䲻{��'��O�d��������Ư���a*�k�n�������<�Ͼl�M�����.��B[�R���Q@�EӇ��V�Z���'����H����I�,S.�
���8vTg���lys]=��^xQA�y��{w��ŏ�Ү�� & t(=�|ffΨMԨ�,��5�����ʚU�9U��1�F9����<�!��\P%Ò�+ʢBe��:�ɠ$F����f��M4jv�������^�=Y�T�
����$���C�	Q��x"e�H��͠�f����kk��jT�Z=�P_��>f}�-�B�n�+:��#	K#V��-�����a���*5d��/W��7�r�!�*<5�:�&p Ti�Zu��|�Z<#�g�a��P2������@z��T��W���_�C�[Z���8I��H�V�Rɤ<�G������ݼX�Me��N�r]O?���������W�&4+WE�E�Ń=f�e�> *�<�s�i�JѶr۫-��m=Ã���u'x履zƞ=}ƒ���sr�fneo[Hw��4pkj�{�w�N<���sq�=���LfO�o��rU�*j�Z��TR�~"GKs_�1��@� �¾`�c�]7 |�0A1!	��Swt5�D�!U��f� �bфC���z-C��ހd�;�_w'�v)�,(�R^S���{����x�AO�գ)1w�-2�란�5�����ۢDěk�cy7�t���O:�l�gwձ����ꗵ��4bB��{�Z�/�0��y�z������%��{O�# �嵫2{Ba��5$K�U�<su9h��c
�C#Ú�S	�� �9�����H>��ڊ��������}x��RE��W�KM�N�� O���xq����p�Ft����K)Tw�.��X/|�@����PؒhHh�3g�(q�B��?��r��W�K�}��t�>\��r*�p�oCx�`���;�O2�%Ѭ;� �[��Aj{��]
��HBϚ}�yR/;8�tL�ӭ�����?��o��S���ƻ=7����nޝ���S���ӟW��hgg�>|�}�׃4}��̧�s��Ӫ653P�~��	�Zz���c��LJ2���	{j�Zm���M{��mekC�g�~֎��ގ�-ܟ��.�ͫ�,�횤%i�V��9�6v8вAh)����hW��3�\�����B+�I_:O\f� (]��BQ���\A�N h�b ���4ԙ�bfǚ��%#;21j�i8}Q��ٗbk._��R^D&�m���࣡c݁Bª*�m�em�X��p�]�F2� |��6~jں��ā�l�����+u%+�xl���/����#Un���t��f[�`i�x��j��9�
��Tb��94�c�ɱ��YT��3� $���k�}���t��x�d$W����mon�"&X�)|$��pKzGV.�ܹ����a+�e�s�قj��R��8xi�1��e2Z����'pnt8�/�C�~�N�ª�@�ڢ5lf�-ۨX�;e�c#C�� Gy��9;7}�ҁ�|iWv��?���-�[�^u�M���m�o؎�N���g������ma�r��C��V3����ͮ��cQ+�JBa��p�8y`:ޏEAأ˸`��GO��=�8	*S�9�9���LIL�n_WT���ۑ{�ڝNŭ��3��:+�3�Q<�4�]Ã�=�o]��j���'Bׄ�F f��{��)���!�����sb��ͯ�� u�3��$~�g~�@h�셖*��UR�bL �G�����ԸG��R�=V��t��DA�iG�q��rk��)��B�]��D\I�ǟ���I����ú�{���������#r��􄟿��bo���}�!Q�_7�w֋�8�&[�>����"�&��eN�wE�
�gý�iPn$���T�ǎQv]��@�O=��t�ֶ��]\�k>�k٘Y&�g�Ź��I��om����\{���5��{B������:8 ��4e�w��E��1l�m�l�����O~��ڴ?���ݎ���,��_����w�G��^8��M�.������'���#}�Z�Z�unX ̆����6���uvX�����{$Op����x�1z�م�licM?���Y;sdJ&	�؍������Z�T���� ���#�Y
�]�.��щ���r�{BFSi!0�6���.Q&�x�;Z6�E�]�J�ʥ�T��X7t��.;4<h�f�zQ�IŬ'�f�,@s�]x�+U�5���HC���*�u�,L��s�*�h6�6)k�0J���6q������ʚ-=\��֮g}�L�6�֕���&�̥ ꣓=^���K������%ҡ��� a����[R#�(s�|�k	�z���AnX>5�
K�HܢB�Z���a�kC�\t8ӎ�gjl`Z���;���t�C�o:Su�Q��^����4�M�P ��ߡ���U�K����=�o8d���6��8iI͡�3{B�ӎ��X2�J���C�mfz�R�t�يW	?�^�Ij�*��=�vx�0��������m)�q�e1����I�xsH0G��{!�Nɱ
�	F��P�M��B��0����s�3QF�����,��:��� L5GNE��#���
�Q�xO B~���z�`��P� ���I^���=�tʆ�G-��%��R�bZ��Ui�6�:���?�~Dbh?�2yI�6�%}��x���$hZk���|�?�I����j�����U(,7�p�8$q�"�� mf:����r�7�}��%���	�*v�n��y��:%��h���j�{B��3T�Я��������	;=3�{���Y���{pA�$��5����<77�mxɦ�n�{���S���&|"� �}�t�]���XS�y3���P0(Eħ��R=�ֈ�l���+��ң��O�a�T1+�����FD�BJ��t3��p	.�Hi��	��Z��ך���mM*a�!���������7�{�& ������p�Rǥ���+�f��ġ��+���?6%�����������c�Ri���C���WMm_��!7�A4��H_�|S���<l/�y��;�m�o\�PA���K��'�n[ZX���Y�3wWm�l./�(d� 0>��a\�[G8bcvxhL^���J͵�%_�K���&D��s,	�1yA{L�[l����K%b�ۙ����v'�'�a�=i��LYG$h�bIp��E�X+�jV�4-_��YQ8��L�Y��V��9 �O��-�R�-ttlx������C�����Ҋ�R�7�%推;HY��R�"�]�Il�X�,ڡ@]�/@�ِ)`hN�y}1��؄NѰN�⚂�KJ�9�L�#��vh`H�yÛ-SY3�e.�f����>�:��x}��d�i�&��pT*Kz]�m��H0ƛ��q���i�Z�z�����A7�θ�X�*	�'?Hі�3��5$�Ќ8,$"R*���f��Y,��do�Ei�vt���6<u�%�f�r�V�7���}ۖv7=��Zfr����6u��}���ݜ��.Z&��(.��8�h��s���V��=e:]긂~�9O�X�Vo�}dT@B�Q@޵⅐������U�֦�cG�*�v��?|��戮v	K��D��<ɍ@@H}zjM��q���x��D��kQ*�2Wٹ�C����;��ŬԬZY.Q��dqc᨞c9_�(�/��`6ͶuF�+�ֵW�� �(J2\t���
́��C��ଙ-�$f��6�yU(�VA�V� ?Qg�V�l�;���RU&:�ks;�J�Ni^&���d������'hd/8?N���jMv�X�N�ͽ=�626*~�ݻw���?�;���VmhC����^N�ʡ�y�$����RW��*hVM�F%�#���K8uN���Z|�6�L<�>'@=T�>s�&��[�;�����y���`����tۍ���a���V#AV��^c$�p�.N�x~\�P�tAK�����m�"W[t�x�,���9�/�����/>�J�ͅ7��]Y�חo���c�=���:1� ���!�T�r��AGX/*����kOϓ���q���Qsnߒ<qtʎ����=8��o}��-m��=uf�N9��+�����>���ei��KV�4`Ɇc�sk�,�,�hJA�7��v�q�w����sb�bq�&GȠ��&s��%�i�ұ�%�aK&�֙NX_w�F�l��Sx��Ӻ!$��v6�����py�ֶ�V(֭ܠ��u(e�������v�b�`S��H�a��TLݣ#6|��9dA�0����Qk
"�\^�+�c>�D	��NX�O����PO�^��ղյ"I%�^�K����.����� �͖u��m|tԆ�-�L�#��[�j��.w"!ʛ�ohE�ګ�eV�����Ʉ~��:��Db����(8T�f���|�jǽ���:��_���u%lFG���l��L��TJZ���}��E~�a�����X��:�]&��d4��pdhКͲ�x+�jG3����몦 AH�ډCG�_|]�A�.������-z�d��M1�;�E������4 &�I��D�>�vf��v5��G��ha��C�&��> C7$��.���꺒(��ylӶ�x�Ҭ���t�e��*�>�kw~2�u�Z�B�.����c�1(�fq�Hcʨa?�6/]_x��t��D=�I�S�s�K������'��#N4�_Ry��k�kv��1�%	CG�	� Rì�.
~�$o�坑̰�R���R�z�,�k��:R^�g%��7�&s]~{ׯ��� �U�q>׍��+�߷(�u`cR)=�G�����:�����grhe��pؓ�z"eO)K���<K�s?P�8�y�?Lq*��S�{�3s���Q�V�XG$���`o��B-�֭@���C�U�~��-5����F��._7sV��)ΤT�U��ZӲ[;
´��<��Z�n�W���W��O��S���;;}0�_^�q��8�:w|��͜QX����¢� ��dz�phU�umJ
(t"���R<n\��p��1yR6�?`c]}��Z�^�l�ho�-��*� /7up�z��mmmU�� �!i8x�ea6B$��ζ���V�۳f�dHvD���n�X!W�H�	�|#�T$�P���a�P�:�XXEl�Ö�ۓ������lh���{R֝JX7��R�ʙ��wˏ�mv��-�gm;S�J� �e��b���i�ctQi�sY�Z��ښT�\�$��>y�&Μ��c�m�Z�m�-�lZ"ݭ6?`}}C%0�r-,|�u��`�,ݑ�b��c���^F�Mk��x�'��"�!P\J~@����%jU=]���'$t-���є*mQ��n\�� ,:�?��7U��RE��^��eɴ5��J��T(��H�O�ǀ~"n�FK���W�;�ܾu�fo�t�]S.D�� L#���A�$5���^1KvvY�����ɩ���P�kR�)�**p�x������ۏ~�whU��י Ը��m�]�2���o|K
t7�ܰ��xC����N�C�fT� It����؈S����nmo��'8�� LU�SF�<'q�确�qmS?����ёUр���r�l݉P(ك��
g���͡���φ�J-� �Qm�ݩJ�F�]m��`#��}��Ʉ�0t��8=zP�{����{�,�A�,G������}���	�~����y�����N�'U�R"s .��ĵ0�m��sH����\�>�u�% ��2�����*��,t{ֵo%r�N{��m�l���n�L�T�r�adz�� Dk���Gb�x�*4��t̐���S��P ���T�Q�Q'D�w�y�k��<:�<q�=�XȔ�.<��PHcA�bkU�_�΁Q�	�@��C=�����\, _v�:S2�P&���}�̚�ٰ>�q>J�� �3�hsT/T-�nE@A��]>u`�_���+��ԃ�o��0��?\�5�o�&v��:iO����&��e�t I�AKn��y���$��=���d�S�p��]IKXF���0+7*������ʒ��3g�ԑcB7c�v��{��f���vk��p����d-��M�l�Ƞ�/�m�p�o�l�[v7�f�T� G͹�T���N$,�xg�����H������h�����;M&V�%��b�j;[�_���meiݖV�l'S�|C��E��H�'��� �Ył�%+�K�8�">-$6 B���'�sl�zN�v�b��Y�ް��?`�ccV(�ʕ+v��E�9 *-e�ڈ�yŵ
�F�� L������,�U���hA?ªhZj�0��L�A4��o�]����H�2�	������]Vjv��1����gm��=�Xd���Қ��
�IH�%J�0��E%��h��~֙�ˣ5�����agW�~��~CH�����29��!��&] >�z�Ƭg%�!w��9S�HF����	;�̳6}��x�� �@4 .e�a�@�6�{������?HoW��=�b����i����+:��n���y�e�y%v�z߾����������lR�LQ�%Y�D{$�@&H`�LL#^�1xl$��1�d�$�x$Y�$RII&)���}����W�����{�9�{�;F�X@�Iv�����}�w���������ޔ��^l�p3㓈G*��RńW$bA�:quc����>Tѕ� e�T�n�!�H�`�w��$��ڈ'Ff��<�闹�����b/Ґ��xp��L���3o\���v��94U���f�
2��FW�,���v�T�E�VךAn}��ds��F6�~>5�]?�X�d�ڰ���=�S�y��<`�K����q�5F2�3�/�O�aD�A�p�Fݰ�{.���L��le���3��j&MK;E��_���rO�g�xI�2�VZe�q�ޟ��m8.���@�Ū	B1-B�f�R,��\g_'L�31�V:�晭C>��{����c��AD���0s����k'�TƟ��Slh��R7�'�Eޣa��gˤ����	�H� �(j�v�%"�.#O�>\v�f����M�"2ed'�����tNb�i��T�Ґ�Q'w[KO��'�◿���ѿ��=���?����&���Ǐ���#O mE�8(FS�M�'=����ٔ�c�pM.��.t�{���(�غ�A��mcuk������
��'���# ٨\�9ܸw�܃������"�Ш�M-��hUj(헙+_ۥ.g ��'<�i���j�������]I�b~��i��cht ����.3��-UQ�-"������`}m�{%*M��|�~�=d.F���Po����sY�?�@�Q,E$N�j!I|h7��{Q�C��G��� ������H�s�!kg{K���n��e���Y�4<P�M~`��)�Lc>�EB�dTk
0�>��@�~�L���������^w0��m$E�,����L��߸�+��C��`?n߼�ٻw��Y�6��S��F�R,�C�2e�
j��e�Å� Z�z@�%9��ĳH�ݍXqk�˫Қ�{���k�y��b6>$��6ӱ��uv��@H�a$Á�q��������Y���	�����K�&W��ƛ?5�n����/#/�'��ٓ���(��[7n��w���ܼ�Č�G��>�tNR���e~�,���+�kذ�.i����M0x(�XE�7��D��͉�$y�q~-Z	E��j$?1|����urA�By��AG?�O    IDAT "ߑ�i�u�2�S��:+���Af)D�8�0��^T?Lh"��Bj�	� �����U8� bh h>_��<��+�疚({%�Ɓ�?kM�������?WS+#�����;D���-�='iH�?�e�]��G�1��iLL���m~��N�[�lP����mxvSe������h�c�0i����j�!O�8�����`{�hV:|_�\�P��Á���BG
(�� .@ѿ�R����@�4l�)����L�Ō���sa�SG+�+�;��#;������繣���L�4J+k�O�良@�kT<�jK��DMy^��F�ʤ?�|lp���~����'a~����o.ݽ�Ͻ�@v��!1���C ;e���bl�=�v�9��Љ1���q��G�؊��:�>�ܬj^YYӎ�ږ�G����L�jo��[���2���=��]'�����ֵT�GH�BÆR�0����i�Mvr�
����c�_���B��F2D<�8w~�-LF��e��k�U.�������ͭacm������ڠD���W4��*5�<��71;Bn�XX6n�hXd(����4��Z~�R�.w ��-!B��� R�H���=��y�..b}su�������+)oHAn��v���9QУ�,�4F�l+OYI:��y����L��f܁�2pw�d��a�^�1֑d��:\"�G�04Ї�7oj�}+�L#�H�eQ�41�`^^˞�e'G��B��P��qjKR8y�0�D���U���fҢ��ċ�~Y�.�3�#���΃G�>jX��+A�%7� �����Cةo<q��hH�R�g�<	 d��h���_ZY�G_s��	Y����r7>40�3'Oዿ�E%�ܹ~��3�//Ir���˒�{g�:��s7V�F�ncB2�.]A����%X�6r[�ɭ`��4����ȃJ���97��ܽ�^��_+wj�u���I��$���'������EXM�}����@E�òF�x6ݶy�M�CCLcNOmN�*���d��`�ec��y��u�ٽ��5�u�(�b��� J�rރġ��.��t��^E�����]�_��X�Z�Z'b�/]?�V�ۓ+?S4�gfZ��"��	Pn8/�V��`&P;��.̂�9�W��~�J�7?A�W��� Q �8�T�Lm�D�fZ]�������r�[��v��q9�����C�Y8)jl���RqYdǆAg�\��F���0Fp��wO�
��1���9!#���dخg,O��K$�G���2��Ǌ���ql+׎����ғ��Gg�ړ�sG����wfG����|���έ?nt��^й�5!)��89P|/��er$�d |���|�l;�A�;��	P�ώ���z��v�zYlgR�}^�x�ƹ�#xbhJ�`�mrvlc��b�<L�j�=Xt$щA ��m�A�
%�z=�E
Zw��jT��6Ѭ�V�G�V`+"A/�ɨ�f2��i���}h�	�屳�"��{��`ua�k�D��x�M�o@E�I�{|��-ྒྷ���"4�ُ�a$+����Z������=p��F���Ȍ�`h|SSSr�!C���p��a�d!��"�o���XQ�B��e+-&�_u��Õ��$ev�$ݐ���b�o�'U�i5��ԟjU�G}�'q�����Inp�ׯ^�N�1��>���I��w?�H��� u��C	�9�b�:�!����=��M����=2eە��0'�N���ۋ�l��m$k,T��I��w�8x�z9�a"����14:"��X<i�ݲ04�0��^qO����EM�|]�ܦ�-,�p��=��d���翤�J��������
0M�GL�� ��HT��^~_��N�Q��5;L>�|o��`�-lmoŢ�^�d{2t�NDj��P#������0�yp+��2іN.���A7��	�ϱ&f{:�t�!.C6�"���2E�mg8;�����Si�	�����Ƅlug�lX���g1T�`�s���A϶?TCeQM�6��iz�
J�����!iu�B�Y���r�p*�F�>��)��f�ip��o���&��I��u�i2���^�)y=�ܱ,{���%���u�/���
�������sϛf��߫u�L�`,ou�ѫ�ps�T���~6,���v�����P6W���!FJ�}�3}�"M���XV��0z��1�xͰ��߃��D���`�����$N)י�ym�]�	Ż�*���pvu�"��;:�nȎ���o�Ӌ;����{�?x�?�������n�<��x��IE�Ad�J�Ё�����K��V~�O�	,��>Ī�EIE<~BЕnC��:;o.��:�0�9�xr�0.LƱ���͎I�	(.��m2�"������R�Lm�!�&�zA:l����Z.�v7*hsZ/�U+i�|H���H!����J�7onF�m氽����l-���W��n	�j]o m��D�2ݝ��M���H��l�k�CpG}K�Z�����\�cae;�j.�����va��D���ءx��I�>}Z�Uժ��=����J%aA��R��G�44�X����@0uxB>:F������{7N>���!$3���ʸ%|J͟􀭮}�`ѩ�ב(xp@)A4}�C;15�Gcdr\��?{������O��/d���q�K�7�� ۚ�d$�P���(��=&!��Pk(uj���&��B:����݄g�?%����1���D��f�Fq��N�,���O*"=��B�	i�i�et�����|�RU���/�����E�~�ɐ8	��?g� �b%�L2+$�e�~�PM�H��ǵ#H6#a�MMn/o=(ómP��u�l�D6wcC�R<�-�(���v�|>��g�E�Dۑ�l0f*3��,"b��)n٤,B�2�`���	5�����eT��N�&�+Ru�0�?cB���Cܙz�lr��(�@��>�f����⫟eLj4h��qM��n�q��&g½��~w�(�Iڄ0�����%p�g�e	Y�y-��M��3�ƶٕ���]�0��9��oas�X����N7-s��}��6k 51^�~gL::�y�s��%��+����U�x���̛�iұ(�r��j��(�EX׮V7)|U#��D�rK���ky��a�%Ѣ���b��Vد�\�g���aTn���&�ȭ��4���p�0�U֕@�����9���ә���^�P�9���߫��+��o\�;����Q�]���
�&�% =��O㞕I>�l�qB�c�Ǘ���s��=a���zY�H�oM~-�R1��ϩ��i���cxj�0�����O�;���������v_�Td;���n(Z��U���)�U)���mBp�z�\�
<=j\�H�CH�"�&Bpq���Y��J>���
6�����Ge�����]/��z�j7{ܽR��F�U�n�7+!f
�pX% =�KM�*$#T� 2
	[�ܨV��&鈾�L�aQ`�9ܠ�wdf�y�y|�S��aI!6ED+6�r���5,l�`s'/�������0��7���RT���r�^cw�f�B���vK�ŉ@g�Ӫ�?�Ӗ$"��Oڐ�i�R(�����	�����
#2��DvpH9�\��]���rY�N��t��>�LΈ�D��"�d,��4	?<4���l��ɝ�T+汿��'r@�6�
C4�i���������z�,v�I<�'��S�̪���E��(�!�$9���$��w�@��|��X]]Uc��/U��{_y�,-��s`f�>+^��Id�IA��tM��4ҙ�^7��~\/��;�����٬P���u��T��<i �=�x$L2��_;uN�+�*�DIX�8�U�T$�w�2�0d,����N���[f'(�#��f6EA�Ǧ=��v
��GQ�,��	fߨ0Dֳ��3�;E�;v5L��y�fp����D�U3՚�)z���}y�;Z�]��)���#�|L;�{��2?~��ִj���$�YSH���M���u��S�V,�%SP�}���5,f#)r�z��ku�xa�՜N��S���S�h�j�	��/���>� Hff��BjĆ&��"�J��_�$��M8\ȁm=�5��AEr�P�jY�] A"�����QHD�d(��m4�wwP{�
Yh|���Ӹ��*�R���p�J$뒋V�n��TLs�3bS�{V���˿?�����ك���/^d�����*¿��_|����?Y�^���j��H-w�v��3x��B��F��B���Z(JF�Vfno�2�$�p/����p��Ut�^춪��@��#����8�?���a��P�?,�q��.����_ԞR�|W�߃�E˷� S�]�H��Ь�Q/ᦜ��o��0ZyzHF��&0З����m!���.�,c��]l�_E!��n����At=,�*�6���y�z��k�z�}*�������q&��,�NW�:j58���g�9�^O ^;�U���2&�{�PgΟ����x�駑N�ǰaQ�|��m\�w��n��w~�J�.XD~��v��!��Kr��,��ӕY�z�&Bn/I���S�@*%����Y�y@����.�~?¡4Ig�2~Q��׋��	L�L!�׏z��wn����5������A4=s ��8��G�K��"��v�,^"�hgg`G�lL�Aܣ�L����ۚ��Ǝ�C^/����I�iX�<�+=���;T���$\F3��: H�kʭ!�h��;�����)���_}�UE�����/E�'���G�0�C�H���n� t�[{=�n��P��~�ŝ�c����6M�2��vw���'�������v5�ΟGr$5�ԣ����h@��X���6a���
�~YTe�(,�M����*���%�F�;|�(����;_B���n_,&�\�(������g�R͟+p"F(hc3��F����*�Ho���F��~p"��VD(�8'&�ި>���ܘ����y��fڛ����l��h�jyD>U�ӝ�9��*I��V����ò&���"\���ȵSv�iN>���b>Sl�����&�Fd�A�6N؉]vv��v^�u5�'�ƩOM�mZ�3OS�}��=���05��XL<���aË�|�h�}� ˍ�R�ʖ-�ʜ�u5��2K{�v"�i2#���?�)����X���.b�}������ϼ���+��w��^}���ҿ���pb�QCl0+�f��F��Ԯ��Ѷ)O��"���{�W+_]�����5F/H�B� �C8���Fa+<�lU�Q+�L8&�(%�6�6��LË�TV�":(ED����#4�Q���p�X[Z���"v�WѮ��*���6qa�4�"A.���VB��T��bn�|�*i�����$v�U���ѥu~��B�}A�<$y#��
�m� ����B	�e]�v����֒�41s���o0�[.Zt�#@��� ���x�3���C��P�A�F�^jT�oVq{��ݺ���%lR�ͦ��@�������@�6Ƅ��2��Tq?�N��D�
arhON�`0�A6�.т�u�.��tV���⢊-�R��ӟSNE8�E�����a�iS��1����b-�*� 'N��ɓ'q��1[�e��|X�6%�b`�v%;��<"�Uj���M�*Jn�޸��Ak��x�I*c{\���Ȥ�}�y��bdܐ�2�s��;pJ>��3h��y{���"�`_�&h��^{MF4<����2�_ZYV^�{ ��&��Zm1}yh� 3)H�����h!	,r���)e��^a_"?�KX����i�a��d�<%C���1���:�..i��vhrz���pg''�3g�	�ʿ�05�/�u�jNf)=�R����_vLb8M��<̋�z��[0���8�-�#f��j�T����l3�t�ӎ�W6;�6��zlm�%�4��-	�ѕ����P�c�bB���㖠��y�;�W5z�<*r�������122�喜M�;s�KLa�+F����Up��(�z�@�|�Z�Ab���(��pRN���LCÁj`�f�0>>�T"���aC��5b��4�Uz��YO��p"D�y�(���mxE�#/��'��D�Ȧ112�ϊ�yw,�}p%��R��}��Y	0^�H̨�
��g��)�3Z���ohE ��kt�L�Y�)�>鄽��d߿?5z��~��7>�"�g7�yjn{�_][����&�})�Ը�4�T��(&�R�#��!��8� �rY�u��:5w$���R�@u��N�L�tW;�
w�Pb�K�������m"�H��Ŕ�J[ʾx�4"^���a�����V���~+�g�b�o���_��Mm!��$��k�H��jqOW�ۏ��v�s���T��Mƕ��C"[,B8�)8�ˇͭ��_���*ַ��_��+cڸä�,�pOŹNRW�!�4�7�u=�%���G�/���sHg3��(a@��{ɮ����yܺ���WK(2��Z���T�왉��X�����g�}�C��ZM��829�c��L�@���Uln�iO�&$�I+���ܼ�cN }}A���k����a`�K- Q|�ooaqs�;ۚ�I$�!��S�e:?=9�״KwB�]�K9��)4A��hl��?y��<hTj�����&m����.�b��<h�;Ib��l2O�;PK�9'�h2�h<!��P�w���J��v��R������b{��-�o���+R�"�蕕%��X���R���܊(��(?�vr
 C��j�.r����ƹ�%�b�񇃸sKkk��+��4#0U�I�������#)O����եe�'g���z�w&�ܪ�ܢ|��h���kg���2�[=�v4!�m��%n�!�f��͘k`UN��g$��&a�jQE׎V���"�a`�c#C�{�Zk����m=�%��l�o�P(�~��jBFX�Et���UP�n�{fju��Pe?��U|�"�����2��XSS�7�a���=�ys�ʵ��ʺ���r��[ϿM�li��3+�e��
��)�p�ц��|r+�!���V���Џ<�ɩq$bчtA�JS�i\XX�@�N����i�����l�m$E����3�"l�c�$�L���>erA/��.�V9O�����O�#�'�;5�6b���xv
��lH6%�ȥ"��p��p�yk�����������V>�"�Vn����g7W���[B�
8Hp�� �ª�����*T�+��!�_ y���<4��t<"i���#�T��zQ���{�:��y�06�p����XF���@,�G����E��P����c��ټ��#e�J>���7p�㏱�������L�C�^A�YQ�s�V���k�A�=���:�C��좢��.-�zmD�)D�I�NObxlDQv�X ��j�Q]ݯb~a_����K�*�2�:1	J!����_�:w'm4���ͤ�~-�J!�?������p��L>q�l��t1�:�&
�26���za�C�.�����;$�7�}��u}o>��G��h?L��:?;v���l�0OcrhǦ�152��ۃ�7o�NA�sفxAܹKHհع�d�'2�
Ţ
G8�T\�+H]tG��v����M]g�h��8~
�ΜC&�U*���wѪ�PN�#ݚ���Y4E�ٟL������XCN�*�<�zQ� �~���IS���i���Ј��I�V
��y��]ޅy�(&�G%���P�{w�?���C�t�|������ה1��_����V�V���~K���Tkf��x����4RѤ��غ��U��ln��E��v��TV$�щq��B�(��`e	ۻy��`����Y�ү?�E&�Ԯ��L(bCc�\�[�f:��:Cf���#��>z*
��&gD�-c �Lg:�).�bro��}8��c�K,Ԇ����nBT��c6>��x�FBf�94Я	����ϲ��D�8i�*�m�ml���l�)2"\I�������"�L���~��w�^���DW    IDAT��:��ɦ����JA�Z������op0����2`a��]�ݻ��%�cG:;ua�i6���h׫��fKE�^5Iaj�ms��Ƌ@~^�#d@����(��(։��p��AĢD��|fSb�eF*2tn�K�e�axw�d���8f���@����H�Z������8N��y�6���jU��n��"^�c~t�,���ڦQ&�����u��A��jή����4�0S�H��N��C��o���|z��?��S������c�����s�������-aQ��(dp6<���J�����!��N0I�:�MQT��:R 2W{^��m<+�A9�TȜnvt ��P��e>��6�"Q�e�pr� �R��a�	O@�	��q�Z,�����.ܺ���e��X.��nJ�&*���VU�f��B���eWI��X(�DY��6|����76���1���H��S�g0�JE4�Pl尼����:f�ֱ�SB$}�F�X��#	�ŗi�nNB,c��TZ҉*���ظ�fϞ���Au�4��Β�/�Fy�n�ɍ��1O(�ˋ�57�{�KX�\�Va_1'{v��;�'7:?�LU��J�_���DS�#xbb
���-�6%�D�Z� �ߏx_��>Pq��A�MR�,hO^�|���9��#m5��}e��"��6&c���8�)Iz��6"�;�L51�tQnT,�$mq�<83���!i�	�2��4�6ޗ�`Qpl���&.6\��,*9�S1p��}ܺ{�K�2A�����I�N��#c����k�}�B%`������n���W��ʧ]������=ܽ}S��ןLځ�>�c	�����f�9��W��#�/_ӽ�v���H&q��gl�D�g�ɝ.�"l1��~0�X���B> �y�E��;�ƢF�eCξ��G46�
�<�Il�,��H�dM2��D�t��w{���i���H�j�;����1��P���"����btlP	mcc#�ǲa�}#�%�u������=}�����&�H���S�eT-ڷ��.MUn��p
y�V}����DrP��A�E��3�h��h���~�|TD�χ��}���oi�%�M��?'tF��#w(~��B�iT�V����tR�$oc����c2�)K劇�=cbl�N���I>��N�.y�s��lj|��}��8	5�� I����NVN��s��f8E�� �`@�hO9,U �Y��y�5�ȹ(��(G}hD|h}f���/����l3��ღ;)�gm":C� ��:���*R���7G���<7s�w~����?�"���}�Ե��wcu��j� R�ʈ?�Pσ(�H����D��B�o����{٩�+�-�i�p�+Lq��!|�P�w��d8�lZ�%,�P�U�s����1������ax���B�
#F��kU�lnb}cUZԥ�y�VDS�[Z�t@%	Pnt�54�x[-��,��1v��ei�����H6�h&���rz�k�,[)��k�E�Wװ���͕�\ۻ5��ĉ�pYA�a�8
:��'*v�<P���	�k���H�pT��#cc���ఁn�Y=R�-�����5�fF���KM"9�w�2n/.`a��xj�Edcb|:�ёJ�nO&M�	L�`��Q��3�7�e�;*���>�}}�f2�ԣ+�1uʄ��;��h*!/�ͽ<�67�W�(Qk�{8�%(o��ϝ����_PQ�w�&3��pg��JB��b��v�͓��y��1}�����	���I�a�Bx�a(�c�J<�k���h<�X:)B֭{w�Ə��.}�?�T_�&g���TV�G�cc����r���$�b��~ 8���k��5}��܆&��s���^�}��A��|݄��îHI^cp<.A��s�$n�!Ǧ���<0�@4�+7�cuc���:��5I��ćD�ZSnBR$ԛ��s��S΄��@�i�uL:�l_ZE�DDG���C�[�lB��1yr��$�qU;��q��m�'ኑ'9EF�О�59j���E�!_�̦��p��)���(ؠa�U)�da�*���Y��>�'�)�>��cv�I��bu��d���e!��{��!�i���%9	�a	�/T���Ko�s���ȡ����E�0EQ�R����ʕkX][S�3[daۘ�F�u��o��?�X�<�A��z]E�v��9(nRf8^��v�p�a���¹���ɣG&	}�M;X����q�nݹ�B��������$Hj��(iI�-�^[&,D�d�i�1����C019�H*���r�
�v��v��0��^t�����*�v<���xb=+~���%͝p�,+^fy3���l�����<=s����g�>�"��n�������ۻ�K��"B�(�0R�w���Ç�˯�4s�u�S&�;����ŚH$u�e�������3��-_�/�Mzt�lk�;X�m�)��l"b�����0K �P^�B�
c$�9m�q�p����Ϊ����D�X�����/Y�2���Lk�wt��.�#�����cuâ�U�d�'F085��@
��ш��"��_����߼��[w�zoŽ*X����Zh8�� Z��@"���";YG,HB\��a����db�h\���	�T�uM���v˱d�O����{N�SBO� 4�Bܟ���������9��1M(�%-���]��p���!ң�m�Cau�9���蓴�s��[]�NnSל�jfxX;iDLOO
��}�6���S�013-쥭uܜ{��JQ�|�n_�鲷!���ᩳ�����Μ�q7/_<��DЗM� kq��v��̴v��pDS'�Pܹ�ɉ_N�:s�w^��IV��"�oBKX�H�#�K2���2�~�]���{�1'�i誴w�Иd}}�F��*v���$Kq�������:��"�SngKE�����3t��aM�������~Qfl��s�ϝw�L|"/_.��nG�N<���)��oa���n��,�����2 �lr���+��b�!��f������A��î����<�,��.Jt������u�K>�,�^�J�2���H�loz;���q~|��sCr����ԉα�g���CS�T�����cƤ�e�h�B��w��>��MǺ�o˨H��ШDǎW���5E��<~߿}O�ɳ����fX�"���B;>��g�Yg�q�d���ʰΫ���.]�s��5����eַM.�w�"e�(����F�ar,߭-�����Z�RJ~��Nd��#8w�N{R+G�6=3�a�\�|W�_�$,�O;:Uar"s���0ƝFX�o��Id�z�P��������C��7*��Q���F��rЍFȏV����M�3ϰ����0�٬/�(F�(���A��Q���%J4xb�p�mu&���yz����'��~�E��������z~{}��Y���PN#��R�^��Q��)�O���f�#�!�f۸�D�������)E�t |�9��M�;@�TJ���ҶwwP����K��l8�C�I\*T�Qf�B��Ji�ۛX[3f;;�������P!���;f"{�� ��,��.H@�,D,7�3����2���$ID�	R�h�m���ͅU��/cu~QN]�T�hR������v�C�R/� �|+�����4*2 =u8F���(�?�d�W*�պ�_@�w��'���L��$|��Y�8�$�GG�����s?�t�&�s���7�����U��!�$h�-BSANC4@!���0�FK��@2����F2���cgc9�yK���"�����6����|���c�d��081���-5{��&{l�Z2{���'�h��}��}�ݾ�����HS�H�5���A�R�ufjR)@�x\���"k�˲��{�LY���*���Qs���#�<bDd�G0;7�b�އ!_(�Mؖ��ܵ��"2� V�J�#<y����lZE��k��j��~�T
���v���Π�/�*rrlpX�4#>ז��N]#?>��PP,���U,o����l���uM�/��簙߶rc��L���2�-�y`�U��),��dg��
��S���60 K���q�<tpj(��܎��[�o�̺����^�D���"�9��C�q K�ސ���ȶ]�l��WH&����҇F��q��!�<~L�`(`��eXB�/�L�;E�σHEԟ*��;'�L��D!`���H����&w�W�>6`&c�pe�51>��~�p��A�Qt�5�Ih��b��*~���2t�����X_:)B|�*>nc��0������J� ��&V93A�(k���H�p��i<u�4�=fǝ������v�,�|t	�/_�fn�V)0���儌M���-�AR����SG�50:���)����������z%�Y^�-�=T�e�I�y��/'EN0�m`"F�\�\��^�a/<�xU}�ׯ��x�g����t��[�x��7���W��t��3��/H��ƑD����B��A�X�(�`�kX�s�i��I-M02�����5�}�׃D:�=��2�P]fx��"�0䞇�����Э7050��?��B6<�YfZ�fn�ul�sb52�m�<;���F�+i})��ni���3�v��H�1�MbrjSG ;֏P:�6�ը!��wP������5�H��vd#H��	��#��B��qОNͣ�u��j�EX_^���i��Éx#��M�4���%���ɘ5ᛱ�)�;�f&5� ���.o�����i�Zx���\ƍ�Yl��s�P'�C"wBπ����;���s�O�c80<���!����SgЫհ����{wM^m8~�H0z(:aj����S��dE��ەK��hY	+��CX�S��q��I�}A,ߟǝ�ױ��(�eH�p�d\�rm���'K�B�B�M~kK���w��!���Z�y�������p PA��������{�kz����%�p+��.�������� �>uJ6H?z�u\���`����We����V�{��&�p ,�MʔM�(S�����w�:vjrh �"L����.��y��PC�H���O�}�<ʢ�-.bk;�	Z�׫�H֤l��M��SH�z�v�7��̡G��߯�Z�Y���u�8p Ǐ����^���*��dM���el����]��Mi�Qkv�a��.Nv6���)���nOt,�j��O&K�e�����IT
3LOL����x��)��@�4��ŉ�\��1�^�&�s�]S4�mӜ)+���m;ʶ�d���M�3��I`���e?K���>��<�.A�G�8��^z	��B��ƴ9�G|l
H�{��wp��Ui�%ݲ#�8%+F�LЯ�1�1���)U�k��*�}���������я����_ʆ�}'N���:�_ӻ��f������K�%A\\^7ӮMܢ��?���x�^�t�O��%��>F�1r`
�3�(3K���V����>�~��������Gy�ԩk�k��G_�&`S읾]�i��0������^I���@�����y��'^�����ח����NٞdFD�����B���n�Q,kyM��}�\L�`�}d�Z���a���]l�,�d"f�8�,�TZ{7�zyC/�����*\�&�fZS��.�{���]lnn`ys;�]9{�+�1;.u�z��K�:1�a��C�V�6�7h"N�#��ġ�����)��Qj\(nJ�����]�a��V�/csi�bCŗ+g/��ii�	�P�t�#7@�g�����uX!�#q�KG�fCE���>�H���:Vs9�5�H�rk�����V�-��x�����?�C��TL�����(����.ݾ����������n�1�=�k�Mຓ���%c~rz/<����Vq��\�q]�9O�<!V4��E�.dO��Z�_��L�r�}�F���=��Y{��;�����*�BQ�[�c�H�;qi�\^{�3�O�(� ��t��^��CڰUm �~pTf�х-N����@`zK+kx����;響
�c��\��aww.��d
�dF?��'�\�>�Μ9���ڏ_S&Q��گ�Y����;��kܹsK�u�|n�VO�=��I�7�M���i�D�ذ јE��^�����٧D*#����]��M�Xmr�--Fjv��dK:��{���:��7U�IxS�m m���i��̅g00<���erlżu��صp�V�E b�<u�tu�3���C��^��a- �v��?�����K>�ԣ��*$��o w�=�,8q��y�<N�<.� ?e����[X��λrt�^T�5ga$�ɍ���p�|*XAE�2&��Iޙ�U�m�
��5	�����?{�4^|�E���a�7�N��4�]Y�����p��e����s{,��N�V��4��e���0ҍ���|:��,�b�s╆ڋp����������3i�7��T�8�%����%�K&l����6�� ~)����v��4���M����A��(�S�(�z�w�j��Q/��w��C[Kˏ.mOiڡU���x8۞�N����$�F�����2�g
!�Y_��������~��O���O���ks��t-�3�����X��8�� b!�W�y~'gL8���k���o�H}_7�ݞq�O�I�Z�
�,��Y&��ER��!�+EMΜ\P�"��a$����T�6���I�Y�ma}'��ZQ}�V)����ͬ4!��T��)����w�b�4����5=6�c����K �E���.��,��xp��kۨ�VQ�4�������Ӽ�Xk��i�	���h�������A����Y!Xޠ�V��$��ew�����=H\`�s�~�������v�jMZe"$\�b	�{��}��$�eK�2FN�����x��U��wVӮ٤�x�d���R�Dv'�"�<_ޤ���#	�=v'������x睷��G*��?ӥ�%,//c����q�앋�|��&5�|�[���Y6\'t�x��i<��y��z��<�q{�-5b^"1��F�I��d� �p��y��e �sc�{�uݗa�������L	�2���H:b�S�''T�>���~�]�������	��^��5�Nr��!��Y��Pp�y�ǯ��+(W���_�5�������/���+�����f�#*�$f�ll�ޝ;�3&�"&� �F�y��ӡ$�T*�'O�oxP��;s�p~�{��H����
>��`� �jFU��)����m���U6=Q�������O=��{�9;��v�����za{�o������Q7�l�}l�Qm�Ԑ9E�Ϯ&;6�6d�v<lНՁ�wͿ�x3{��b��}q��<��gq���#q����m"ރ�9���{x��7���L�r]ڻ�K]�_�S���f:�7)ir\�%;Hs^g�@�q���!C}0I�/|ҵ�T ��z� Þ�f�.]�ի���sV`��R�z@֠fv������yV+����y`17�H�G(�������_�2fL#��)���&��4"^�y ���G��_T���D4�o����DR�ڸl�9Q+ͶBV�De��Gl$����|��"�hú�6�=������8Y;�f���4U�\�d�J���eݞ�Mt�k�_��*/��Н�c�����?�ċ���/�vi��n
��V�X#�,Cq�[��.�l-�EM*�hX{|��th
�k�q�X�L�Ӎ�	��;K}>�����I#5��ha_������Y�����P��v~��]�K�+WɈ):�#�gx������d�Y��.�;m$�>�%��dЗ�`x �h��&*͚L@�
�6rhr<��N�����C�7@��A��D�זg3	���X6,����Ѽ�\�� ��F�XE�RC�Q�{`����=^�
%
n���Xk�F�$#3�=D#x�#ڣ�U����j"��#=2��Ǎ���3��:^�D1��IBW�XBf�¸C'a�:<�	]�$?��V2�œ�p��qd�1��ӟ�o��,�� ��H:E;;NǱhO;"F/�ue�    IDAT��ł�Q6-�m���(HJ~^8��	<{�F���q�2�������'y��C<�Ȃ%�ǝc:���e������?����ð�q����W�u���i�R��UM$��\l$}A�mn��vB�!��&�ɖڜ9sJ��/��Y!z��_~�e��������kW>RAv�}dӞ;sV�.'ҹ�����S���3 �u�R�~�"d������"�]�uU�\[��m��W)?�TH��Ra���L� +@ԿXTnc�v�Zt7j(j�2��Y�1���g�K��EC�	��G��ljrm4��ߝō+W����BW,T�f#���;#K4!毶{����b�WӦ͐v4���2�Ф�����>�O�ۨ�Rc�OgoJ�������
�7��n�\IL4�K'5�p�~�/�pɖ�a�kՆ�_�s|�l����E�����'��ً���ŋH�b&/���N�ٻ�i(�K*ro���]�a�05�.5��bg$Uz��xhmI��f�!����mw�����5�Ĥ)�� 	�Q���ֽ�Sѽz�*���ܻ{u��L��=s��#�����C0��4_~>����<f��&ыPrw�ݪc�[G��B�<�^�~���$�@�I"��"SE�q�"�ms]:�
R����*�Vr���f���'���g_�ċ����_�:{�_��+��2}��U�3� �t#i��ϡv����܇�|E��,�BQ�:�8aq�R����[�來��:��r*��dJD+2�<�;� c�AX�3u����/a����¤$Z2��!�DL�@�W��_��hR�0��W���~/R� R����7���q�[E��J%`w���pB�^�|���N��d;5�5J�1�D�.�3�h�eI<!���^۹=llnc7_��4���fM0t�2���������a�PF�Vq���h�l-7�OB%��������Y�ehj���C������be{[��*	ETO�z�#�l�љ8�ahtx�dBv�^ʅ��M�H�<rs����^�G�/c��Jjj����Çu/l�T���.��ܻ�]���Ϝ×^z3cc�~�c��?RQ '���9�����Ζy��r�>� �����;ylon	�q܁Bf�1�hJֿL���`F����2�߼%"
<B���2���
�ff�v�RO�>��������?ԡ�?��W�*f1�o}���}�:6��up����RnE�isc�[����l��O;v�b���+��ˈ�G�:�C�2=�?���2�p,!�<��cnU K�h�R�;��\]��:�k��W��H�D�C����_�/��sl.�>pZ���UFm^���_��z�bY(�i�K��	�m�${�2;a���5�����2F)���\(A��Sm<Ĺ�x��������������gے���\�v�������.���&���cճHڡ"u[z=2��G�H�i�M|mNlnY"�Q��g/�>��!G)c�i$Z#��S�/_����ks����VD?���ai70�4�����R�)|~}�m�av�r*T4���R:533��~�+������vȊ�T)��_�w61��>���=����eO�j*�Yo�r���P����gB�hT�f8��+B��3��^Ef���*�ݠO;�1���+��G5���9&l0�_�o���� ]��Wc��B2��g(���������������/�����^����ܘ�h,���B�;�j�F[��eպz�Ʉ�u#�B2���׻Vn�O&j�>6ZG{��F�3�G����_:��j�t[x\�d,\�"Hl{+���M��՛h�(�w�M�C���4�p��|�(W��,�
�3���7��<o�v�r4�E�:-1���rB����� �ޒl���Yl�Q��!\�����M}٬�GjG3��8��R&hn#���e,-�aeu��:]�ܦ���$<D�$�`Ba�BA��qk��b�Z$4M�-�VDN���NX�_�K�4�I�?#�<�w.�"��s�D)�!��!�=�!�{�������Т���~.�����	���������4����d���:x��������"c�� 1��S���=~�l�>}�"~�K_������;��_W��d�Ӑ�E�ؓO����I@��80=-�!"�c���$��L�NΔ��n:���"L�I�|n�#�$iq'LM�۷m�˃���&
6�V)�$�ϟ�W~�<󌒯Hv�$�XG~>_��������7�3nߺ���EA�z^!5q,�;��(����Z�OS7�ϲ�#���A$���C"M�fL#C=�#^�m*�X�Q#2��Y7�p7{BB�Ѹ��|�hO�j�T�-o�dJ�N|�3�x��TL�x6f�v�0�����q������X_�B��t��	Lb��+$E�y1�l�t��k�a���b�y���@~5g���U��vf5ߋS�ںq�����4���M�,}z��^a��39;�f�3�%6l4�q�ht�0��=��t���<��y\�pAnTlM�50��q]���dO.},āω�t�$����`�]��v��4+r����ux���5��D�����"�˿��*�1�]XT{Ҙ˜�6����ˆ|����Ѓ��"���G����v�A5�d���)U�e���υB��=4E�jҦ2T!fnr��u��c��&�s���r����"�g�7r_:��lwټSQ��*#�D�>+2?�?��'.��W_s�������)J��빫��w�������^���4bfl��8�]/b]7z<���"�C��B�Y��aR���M�_�}q_�g���/q�ף-dL�^)c{u^�K�2���S]�	C5h�A?�k�=��T�j��Pj�P#�C8�ٹ�@ah�n����o��BAB$��T��(+�G�X���uX�I������aAdCDk�2RN��c��v��B�(�&���K�/��^��@��ɟMG���=X��{����`�fQx�K.�-��S:k14��A��M�W�6.Th�FV��'�^`l{�D�u��T��,�D�n^�:}h�,~&�,Q�1L�R6�1�x�3�/�������l�܈[��<D6xX2ʐ��(�?f$��h4������$���<�iP඄����l�.^�/}��'�7o����lo������&�g�"���q�����BN�t��ye��줟�H�;�fk���o�UT}g��VX����ʪ�r9�qb��I�S	k�o�L�LZ$+�9!��.`|b?|�5a^���: ���o�Ƶ+XZZ���EM��a��D�.s����i1H~4"X:����HO�̈%M�3�09���� ��E��	h�� �A�o�D���ʚ��<]��𚦀�<<8�?q����p���&�������bH�kkaׯ\Ǜ?y+����/����Ҥ�(����C[���:Eٰؑ��c��a����AF"t��܋��3�\D��4��P��xX��� �������?�ll�t�Z��y3oX�]���4"��t�<$N���� �ɏ�����xY�Y��
��V�f�=-'O�}�I8E�7ƻE`���	�X(��������B8,��|�),l|��Xғ�u�m��mG��GM��=�����cV��D�s�b\��OĬ/|�8tx��>��춈���������᭷���ڦ�e��+��s�1�К�C4�nd���7�/te�����"oi��k�����d�x�H ݐ_C� ,�����N3щDU������{�+R�zv�t�����jMx*M������#�}23�=j>�����U�+���׷���B��HĒ802��pB�t��P#��"��Y���#�Mj{��=A�H�+��&��)�@�{r#H��f�2�0� �~s�h��ww��<��"c�Z]�s8W�]��(�*��F�u��\�[d��i,��5����I�C{8ހ�
:�:z���8=��)�A�pY��Ё��E��{���"}e�����#=8��0%1��A��Qk3% {;�o�h/���"*�с��'B0�D(�p��
`���/S�s
$�O�%�(�����mQ�	I����a���ᾄ<�irk�v+�w��N�}9�:>u��^��d��s�ZWv3� 	+ݮn��XX�����nX�c}̮M7��}�5p
�*��;@����v��>�/��ұ(���x�W�|%����|~[/5�J�QJMD:WM����J�$�J䌤�'�UT[g��kX�5Ή��C~�{�s�6���4a�u�2�^����0¡�+����Դ��s��Q�ko�.&)��|�+������˿�6�]���C�}���u��C &)��(Ж����~�%��H���5�M�9�1�G��y��~-./�Gf)?c;��#��w��Q�sG�������1�JFmr��g�ן�S�N������'��$�TÿU�s��z�*~�ڏ�������cA�co�zES8�c7h�^���񽳸�>Ra;X����"O���=0=3��|�Ӹx�i5
z�9�׃����0;aa;W�E���#����#�t�i6h��=���'�p�f�Yِ��,��l�����?��tF�afP������WG_�|E+��~$�C$,��/�L^�x�H�c��GGu�:�=�p(�4D.f�����|}�x���q��A9��M��7]�<z}~p	?}�4X4rH�7�g�#i��W����PQ&JC�7&��W���;a��p��*��xH��,�<#6��=[zx�������b��<%~�����P����吐��5Pp�$���V���ֳ�3��&�����;a~��~�������t�RL2]b�o���Rio��[:4�T�V��h�RQ�O���~ƅ�7�7h�j��ڕ12�N���̯t�Q��5s$y�ۂ�t��Z���~^�(c�^U1�6��%�U�����̂d,u�^K���!�}C� و7x�MC���\���;����=���G�>��/�ofX���l�!dƆ�@���}qx|�t�'�Fy�����/�c��"�Vs���W$Y��|!�I)DRicI�����u����C�c�'�3��M���4�~&d��������JÐ��~7\A}C��#�^���͌�&ev*����Y�vp7�}g7lL h9G�)�P7�Zj'�}�U��W�L�9a�]�CȐ��Tr�w�)�vqWo��.�XA���������֏�W���(z\5ЩHNDѨ���)M��ZM�I>���"��H� �i<����e^�q����@[M^�߯u�T	[J�TLb��������{��r�����h������/����w��||�#��wp��#�y�� �!�_<8Ȭ�{�;)j�i��k����a�M��L�+��_�*�j�$[�%[�˵�C� !��'@!f:�&���6�IH�TL���Nf�$�L � �i @(������V�7ɖdm�������9���J����y�>O��Ⱥ�������=�yρ��0�@�ӻw3�x�	y��cr��%���u�Ra�	Y�}�ml3+a����x*	+J��l�a���[n�W�������
NY�a/Q��2m��E�/��U��_? +:G$D%b�>H���^q��������ܠ�hV����zt�I�w@:$��T��ǈ���9rZ"�G%��O|B����ת�R#;xB]7$�������oT�H� ׋�����%^[-3hAi�햛r]@�#s�.�^?���=��I��׾&�?q��S��f����Y�G��Alxp����p=XH
�~2z�x�+�D�V�����ˡ����cc�Tu�k����ۑf�.{T�q��d~a��H� ��A��o튅j�Z6Ќ��u��E&�8�X�;u�'/�@�8C}�#���]e�uOz�a�*�N}�-E��4m���S����l#1%�2b�����������zރ���w��p�?W����l���BI����7��0�A�o��*|d52oKaA �@%�����,�0�,<h9b�U���QV�&��&K�K�R2B��k������A]�&ҁ�Z]��Q��-)�j&�q	�@gYY*���8������\3�aH/�Pp;��$җ�J��Ȁ��^���f$�bFzK����,�R��MCb�'N:��mJe�"�s+2?� W/]�k��Ҭ�x���+N�W2�^q{�-�{��Q$ϣ<%`��1;�E�fr�|��!�� �(�2�pn��l6x8c�	�d-)����V�;WVe�Yc����j+�*�
$.���'�w-7����c)�|1��4��q!��Js���1���0�J�����+��l3�-VKB��j�?��W�%p�+��?�9q�鴄^��P�0�GI"�ӻ��S�Ƶ��O� �Z�G�J'��d�) �f�v��ՙ@ҽAx
� ��B���D�*�\����)H.\�@a�[o����Xр�V��^�:�mq`~������=Ġ;�c�<�u$��@H�~C������`%��5YV�U%m%+T����<� ����� M��`�羑���yp�L�DS@ ,W8�nv� �]��B��z����w}����d�Q�"�+bV����������/�>�k'�#n�@>@�i�-T�ZB� qW�[��G�AK��y`a�vO�oaa٨4��f���S^��C�}r�E�`���� b��sK\G���5*Ciέ�o9V{�Ng��9G��u����5�K��W,i�#8$kUV޵j����]�\��u`䀴
�Z��kw��ӧ��ѣ���Ӽ�b��Y��j�_1 mT�`u�@H����s��XW�S�U1�^�Ѫ�8>��Yב�u��	Ȗq�5ʆ`�:��D������#I���k�sި�UX@�\��Q8��mޓ�z��H��~GfV��ނd��.��6�hX��� �Rtf�(��I�R��p-H��`1���{1^h��K����nyס���|ރ���G�Փ�����Z�T��Q�(0��lQ���HוF�������q�2އ�z��e�΅!�i�;�*O96��D�'�t]�%���hT$naD������dq�m�����~$62��^���ȸ����ŗ���#�c ��R�P���A8HI&�[�"�cKy�I_1#�c2��lٹU������@pDTH++�t.^����ȕ+�R�0 S��E)a`0(�R�8�^	@���-�
w)K	�οa��lp��Joi@J��	"hCD��nK�ӖryUY��?H$�_�������ڊ\[[�J�)&�)�fr���&fI�`A���V�5pA#�	T5)R� �B@�K8��諩Q5��n=�_�?L�`�Z <vV����+�~���W� �Q�����!�Zo���dc�@��ò��6n��Y/^e`��\�PT��
�L�V�'�C�A��		{�L��%���Q��X��Ͼz�*��/}1gi�VFE� �p�0�t@�����ʃ>@q �o$�Lt��AP�X
K�w��S'T)xfx@� ��v�Y���ߒG�8!Ϝ?��D��!�!zrt����%��
��Z�E��tZ>�=�� Ÿ�y���N�~�!ʇ�*��7<�:���z�Iy�cr�cO��p�C%��Jr]w ��Q�\1�dbj���QaS"�ܐV�z�N���+5Y����I����n����%�_�0h�kՔr�Bb��������E�<T���7�4��V4m A��D+\#GB "܇x�9���5�x���'�F�(C&�Ң�Yc#���Ũ$a�'?�NWN�=�9��'� �	p4�0�@����f/#yo���3k3�CСXԹ��t.>u����{��w�)7߲_&'��D�㓉��*@}miQ~�ay��#�\���9�\��7�>㚍	W#b�@#��6��;J    IDAT���m[�ot�:觯\��ZY�R�G���)d���c�c����p�ԕV�)H^�J�B�;�CWLx�BN�e·���zWoٲ�?���7OL(�g�zNp�o���9s��*�j}�Y�?5-�vF�n�@Ŭ��!�-��a�_���V3	��s�d������t�@�E;�xP��t�ff*�X��
GQ�g����~S����D^G�x:m����yenAj`G�:��-����ӫFK�Xڀ�;�۬�������a1ef��D��q�c$�?kJ�Rl�g�c�둩�mr����"=�"C�j�&@�,/-1�._���k�2��$���4;���-`��K��+�B����t"��V�}�ѕ66�a����pm1�/�f�LNy�"�F/����ģV�J&�G����͒�Z4��U���a��l�.L���-�1�&�ꂖ~���;D��Z�?f��*}n�G^���]�9nD�1_exO6&]Δ���9s�6�)�0�T�W���_�jټiD�����׿�e��
 �% �u�ّ�C�,z�b�F��⽩Ċ}
-����A$:���~qʜ�c��6��yM�z��P�YtF�z'��!�~�w��~资����X02�*A㗿�ey�駨[��Z�����~�Ǎ�������#���}j�3ۏ�8.��x��8~6	9hÀp�D6���b/e+�s[F�@��B_�y�,����k�嵯y��-��@b��!����O3?t�C��R�L�(��l�����U��)��*���G��ZF��a(�1�[�$2��h��d�z��}$@톓��S��xݗ���s���:����*{�	`Z:e�R
��W뎤+"oJN�����2Y�+�o�.�#��p�q:$١��^�'�b0Q:��o}KN�>���|���K6�^��t�J��z��Nd����)5C$��,�2RȫF�!�F<��n;x��yQ��h�m�~��	��IH�¤�4�HcE.T$: i7��]��Мf�לB�[�t7:,�k�ryyAf�KC����z�M��?F� ��@��]#nJ)Q�"Iʂ�=���4I�~N���R�Lt���~�����jpY��z=� ��{?��S/�A�^�E_n��n:�aBפqd��Ut���xCgf��e��N3j��) Nv�	�Q���.�e�� s�$�>4��`���$����:�4R�����5�30����$�ۧ�_�&A�����識]�LU,uln_�+���%f��`H��X��Hш$'E)0�b����عU6m��/*��E'���ۻt���]�"��5�WZRE��s�W�B���Z±a��Vo�
�%���C=��]�^��o 5X\L�w�7i���v$�p���Cq�oErT�\���[5i������!	.4b�,f�<x��6N: ������%ͬh���"ц��u"TڇUU0�� 5g+�L�ʘ�R$��m�P��Ҙ�y�+erb�<����_�O��Y����r�RJ<�Ԫ�!��Q�橤��W���Pc�����7�����+�hQ�� V�$������NB��z��{� �讻H`�ܺM��巾%����~5���H�ʕYN�����D�(�,
�x���'��.T;�|��U#a}2�i�j_8�!+����*��ǽAr�ML[���9Ͼm�f�q G�'\ʳ��*����z�+�5��A��X6;��	q�B�����c��o��MY]�J��_z9�d"8�����W��:4U�c%ՓO��p��d`
�>�J �
����z@F�	����(�1�TD�O���JAx��Qt<3+(pqNX��ྥU.Зjm�p,*;$´r�ȴ��Q%�9�2�ρ�0{�X�a$�%2�wNNqL	Hu�i��T�H|z�MP��  �
j���հ4��iO��d�Zf��F�]Z*�u��"F=�DV&4�0�P�yٿou�'�mU��P�3� �!�g'��Z�L��`�ox$Z�gfe�� ���%�*w��#�7<�3kf��\X�� ���=҈|�]E��9�XP�VS�!�9��O�|�^�3$ꠝ��k�y �0Ȧ�Ȕa���7:�ǷN���7���<�����l�[�o|��������+7�=88���#��A�Ili�-QKs�X��ʖ�1.*��\����U%����۫Rx���l���Y>,:B� MaF�ݒ�+�Ҭ��,�de ��h�~W�pE��*�Wgeu~�Tr!�C�GF����
�֨KymM� ��[쩂,�4T��7��Ċ�#�&}h1�ԗ�K��0�
�U�<F�2�4T�ɉ�2�}�l�<*�����#�	���̌\xZ���i��tR�$=#����ߴ��,�U��� �knv8�>1��l�!���Eu�]�Vu�{9�z	��σ3��@,J��+�%��Q�Z�-!�Kͨ%Z���F�58x�!8R^U�q�E=�V��URdW�WXat�bW�
�#�!�恦*a����p G"Y�|A^v�]r��C�zZ.�{Z�����'�<!��$� ֚f���Ce�7������x���S��.� Z�^���9f�g0��Lb�_W�A�E?+e���*3d��'�@�:x�~�'G�|�	B�Wfg���[�����e1 'j{>�lUҀ{��@G�V�U�Ið�l����*M9��+- �o=p?�p:������g�
-�B�+d�4 ;��ț@%�D��^~?Hx`�c��Uw?Y���3�#$A]���*����Y~�ޯ�Z�.�b�K��@��&���h��X%b0i������,S���cֆ;+��*hsFݐ��ۨ}�o�.VTx�\)�ȩc�Y���g��*�S޺NV%����| �Mq��Wdye��� �MV���n�d%�^ɻ.�)��s;����,S���X��R.������f�t�l`ps���"<���8jr�.�R��t&ڎ�qc��$hs���uHP�=�l��;dzǤl�:�m�g�������������E��Ş�꥓<-�0�j�&��4>A���\����
�xH�'W�Krf������c5��MI�b��J-K�l�ܧ8�P<h�o�d�Q�'i���CA8F.�{F��r�ض_��&v�?۰�W�I�������3�/��r�^��XvN��M���\��b֦|����t��	><d@W�H�yG����U��|8F�0`̮�U������9��S��M�ٵA�puaAVg.Jcu�F����
}dh��DV��>�"T�]��Q��p����=��p�����ood��3@��D���H��H1��@_����@I2Yh��҅D�ߖz��B��J���qhI6�'��+��
E	����H*-��)7�� d�"\Qr�Lq�C�#G�� #F����#t�Ƹ�jY�^���+}�}$n�`�w3Ʃ��CC{��@+'Y"+�	z��,��
�X>�`��B�$1\��p}�7����Z�k��B��H&0*�W*��J�0�����!(`9�[o��_rHn?xu�1G{����47�BZ��N�~ ��<�s����q)A�L^-��n�(T,Ӵ�ş���H�#�Ԃ��POB%��t0��Bf.���)����³�g�!4��dH�u,s
C i�zux6�/G�p/(r�U%3��|$z��7��������9G� �+5<+-����oߺ�����N0C�9y3��y���8��}/y����Ioo��/�g���ZBU��w��%9����}]ʕ�Z��#�;n�R$Jr�v���29+&?<�q��ύ�� Ǒ Cy��b;&?�a�zT�\��� cX�u|��/Pޔ*o);zC%��>�}��EY*UeyɖI�Z��&��E^#� }}��,B�3�yշ޾u��J�����H{�QB��'OS���Y��u^d�U�W3��5��x&at/�~TR��z|�^O5ң�
�@ ���˖�����m[&������!�l�����/\�!�{g?ʔsVʉ4���y��� ���D�?�g@v`82�iX�^[fW婙���Hio��8��LX�VMF�:�փ.n�`
�%�������$�ML�A7��́-;~�m�S��o��#��K�~g��(��PF7���歲�X�f�%$RLZ١7�c�vj�"KE�Cc8?��$*�&���H�&�""{uaaN.\|F��:�80b!�ѭ�e�3đlBVY�M��< ���UY�vM�����pEǲ(h���>�ApR���M�}���E0wu� !M���<67�([���*���ltۄ 1��H$�g@�l������o͏�
��V[�����M%��͊ED�M@�j~U- h���W} *cs�}U� ���Ijs�C�*&'�a��E���A��Kg��Y ?+���`��(��T�}^�'�����bI�Gt�cG���s'���"� �WJU|OV��{ހ]!�D޿��ɫ��n��ҩ7����2;s�kOU�*��X�v�y
A��7�c~S�Nu�M�%*1 �UY��hEHM����z��i�>���� Z�
&��S������y�}��S�<M�2ƙ���P4����K6?�/�#��1*6��5d����K�Z�;"�R\�:M� Y�v����?������$�z$�$�V1��j�E&�6��90E�x�K�C6QJc`�V��*�����|�|�[��j�Α;��W�\�뜕��� 2���ϐ< ���8%֡(U�><�p�����b5���3==��A�"-�:�ˀ �����5��c����G�D�T�Fr�� ~hp6Wϑ��@B�� �vT_8CcV�@�rY�[�,��6q$(O��4�R�#؟9���}�i�2;'v.#\��sY��Q��ӦQ
�v��#�:SZ�k+��pO�҄=���2�
���ϋyٳsZv��� ��ʢ��\�W�r��S��y�?�{���_T���'D�4i��W2��+���&�(�BeU./���ks�E[���>?���r`{Մ��
n^��D�y�ga|���>� ��-����.$���vzl�z��=��� Ŭ���/]~�b��kD�̝��mhT�՚8^$v�g�x|`H��e��������ua�7*SL��Y
g�Y;}hV* .�K�Z��k�+c�7���(I�%�JY�^�>Ӑm�r�A0W!H��H�RU�	�+L�|��3�rռbu��@�"6= f�8@�{M �����2\�H>c����z]�p�MV��%��H ��!�Q�LOI;+u?��zKV������Rmu��=H"^�׋5:ל�8�X�O�s�
�U)��Sz�
�I\�A�MB�g�������Re�9n�,�|tN٢i%��Q9^�n�}#�V�.�cիTN(�NqyPZ�e��;C��u�=���c6,����eS�_u���W�R��%�P5�P'!;�ٲ�G��h\��|fz�D-5��z�i5�$1���ͬ*a���5S�
1*)� ��)H4�d����������]"�f��׎~���[�n�t�8\�[d�Hv GS�LLP����ʗ�C͜f �i<��B�ZW�xv���1��ejw1��Tp� mt� ��qn��x죣r
`�ޕf��*3���=r���r��e��1�ύf��5iV�v��<��r���Z�EV���J2��,�<܃�.j�Z���h5�0	���	+b���H��9"�	fn�	tƱej�$+�];�$��-������p�v��~����ߥ7�JL5c]��q��<aX�c�z!�s?c�~˚������nE�_w�`^� �^!�1#u�]��������+�j �'[��X�XHP�Nk&A��,`B�!X�7�K�0�	ԅ�� $���$���~���d�OMNR ���XJ��i�y���䙳�R�����Q6$�tqR^� �*�K��P1;J����[���̵y���(�ՊDYE��ș�=z1SZSBL亁+^�5�{$�)MR�1��k,�E�-�S������7���yL>i����/��4�k�z���vd��&��3�H�N(/ <=���P���0������Q�q�i���Ք�å�	| d���j�n4+k+���$�{�O�%Ԋ�5)D�L��ȶR����d�D�����t��т5~h�����/����a�&|``�r.� �4H"q�{
x��,<@�k��� � ���Q*I�W ��`P沜��D��h�M�,��!�Z	"�qM2[�jӢ`$����tS�>��i��"5_p��V�:��^U	�=;"3Tګi�H�UX�Q 	{gZ��b8:�g��wR�)�lNt�D���� t�5L�Ϡ���	FT����h�`�#CW��J���>TZ��a��3�W���ԏ>�k��LG	�lp�I�͔�(��]kaS��ٔN[ap���*�T���;�{<r��Iq�;�g8t�~aj萣ʁ!:������0�H�� ���W��Sg؛��+G�T�UUZu�TJsʃ}X(�1	�NaD.to��o�c�Ki_h,"��f�����E"�����$�vL��9bP0����*uv1���������Ėq�DI��1���;{iV}��<��q�a�=[$/u�e�������+�	�Z@��H�
P�z��c%
�@?ۆ^���~�`��t`���=-=`�C���J��?�A�ر�i,���d�,F�"؊�*�Cc����A�\��O��E5R��7�<���^�c��аLm�*w�~�l۬��|&��I��� ��~��I9s�izCc����:#�sj)�B��Ң(e)cM��y�jU<F�0I��P�jئN�K�Sn9x��ܱ�#}��l���钠��#����S2�{W.��F������PgT"K*�hE�2>���6hQ`���nJ&48c���q�ƸF���H�ғ�)�	Xx.L��S�-�#��K�x�Н��!EӁPUes��Ϧz����������|��O]����z��5��0�+�v �0��b?��3��)�,p�i�B%�DBe��A��#���XB#��K����e��c� ��O��I&e���d_���CPoJ{�*^�M�mT8��`��NJ��K���AHh�*�A0�q�!ӄ
��$$p� �̊�p*e��,X�h����� /9��V`[҅~j�-kݎTڰ��
ܨ�H  �Ǩ��5��(9�@���P��"ԕ$gr53�8�2z�Ȁ!��*e�^Pݚ"m;�L6k�&D�%X�8|�W��D\�����-���p��*T��rA�F�����fP��I����{`��D\?L0(�	�h����,��Ƿ�In޳O�MM�-���UT���8�������A��!�s�'|E�Qp�� �{�,aq-F�lZ_�o
�C;b/�q�
��
��h^mY�K�|�DhB�N@J��6Ǟ����9j�O�sc掃�k?`�sz�|��lC�.��A��`��<�WJ�1����<�d$5��쬌o�}�v+�ɪ�d�ZY�V�Nq�RO��z�ٿk���m����X!�z��K���G�z�C�Q;��b��u��Ġ��Mb��^�PGá��t�b
C�j�������{�0�z�A9x`��z{h��A� �bq����1���Y��W���k�2��Y(H6���,./&��8����d�����s�/���w� �ͩ��;�b�>:iM0$b�Ԕ��%�VSN>yV=���=��4�'�H��h(�>�_�����|�p�N�� �kù��q G3������9j3����q��r� QQ��la� �D�s�'��0F����۔0�3K�����K*�A�c�@�V7���ז�6iJB��T���>��6�"f���Q�SO{����3	ׁ��1@D:jH��;=f��L�]?�����m �y��|3����/x�tb���,uZ�V�m�y��������&��$��: 6�Y�    IDAT�x�YY[2�<+�RQ��#�=f��w�X=�}gݾYjey���2��H���+�c,�<�KS���d���bחb7�Ֆ�ِ~�AH"R,j8ZYk�ey�%�NH��+`=�������/23-��IOĨА�����%F7����+�C����Ƒ,�k��Z�5D0ZFDMS*�p;��4ɀ8�������d\E*B_�R�jS�`�nH4VaZGc@h�+�4�ܕ���@�-<�R"f�� �Tg�i��yKX�E��7�)�٦� ~@��B-A����2�P�hM���sڑ�3��"�(���W��X������&(�4�TAϊ٩Ƭ 7#ت�[�|����t`M�R�փ.�HT��е~p�B�8�*)����j���o�?c_,w�?,��a�H�	��R0!�p2���N���g�!�ĥY�+ L&���V|*��/����� r���=�)�L�;��/�X�J�%;�z򐮄���@?Ek ����/�j�)Gff��c�?!{T�eJ��z���p�`�#i �ι�n�ɋ�gfٿ�duЩ^&��ɨ���)�p��.���[��n��c1XXKvb�Ѵ)���O�W��5��M%��;U�:�l�d����H��ΕV]�ol���'�5�R�@U:��}%�z�LMMI��H4NoE̲�Y�'?��3��1(C����+[$����Y�,�S���z�^��w�����S� m\���^^ i���̴4G�I�	�HB�|v~A���0qa�Y�.IT���\�����5���F]9��-O�q$�`]cv-Z���վHQ-a��H�ya���������4��c״'��nl��b�r��nA���=�� �|}�A=�����]��E��Y��m6+#�z�!/�ER�c)�"�ZK
�3π�Č�'����X�=P�*Wm�]A�8�8cR%�ڲ�mȕ��,����: ����ϰdߦq�Y�Bۗb�+n�+YT���ݎ4;M�)T�k�TY�%`���P=0�].Lm�%ʨ��ze��F�(�=��6!#E� �V$dH�fH���Z-)C>�ِ�v��m8� Nr�W��n��+�� "�n]CE�*��F2�kx�kЂ��Db{��k�E@W���<HVOQ��P1X��[��
��nDQ±��¬�e�K� ��Y��J�沯�f�UN��*��A8(���s�>2vm��|�H�4�X^7���66T��խ�f��S(�C��}� �^��
׼~p�kf�)�]9H�#R�<(��m&Q���~�B 8A4�e���P49����i���"h�$4T>��� �d��P��(���4p#p�׍�VA,f/>g�2�Wb�q�p���3��pɰХ��[o����"���IL�/5����ȥ˳�У��7xH�VY�!1����ډ(esӃ�3�Z\CW,�5#Y�+u��Z���X��ic���r���:8�'p���{b��ܜ�:}���h��_ H�B�04���m.${ZZ���p�p_��3�Ԭ�le��Q�A� s�/���ܾUJ�>1�6��;�:�8��e9��Sr�Ҍb�#xQ�D��������� �G�ք�I`�@P��p�P�R&���N�d��I�D�z�h��L �_�Td�PK�я�gT�'��ty�(�z�d3L� �@����8��I�
X�V9��RM�8L��s|�0�b[]�0=1L�4ͮi�m˲�b�P�P�X���-�l��+q�����җ>k���s�Y��m���_���ً���r�+��(�n�a���ё)�0�R�H����? ��N��h�	[��A�؇h4��XBd3=y��h(p�Q�K��+	9��=�-��#�n�.S��b�k�Ԛ��z�L�jK�U��ZY�W���>s�F%-�7%�Q&χ���6�U��G�s:��C7�E��1p��G/k` �J���4dcQ�2��&GV�
ʷb	S)\i�,N�E\5j�7� ����_�NK��X�M��I?)�[M{LX�j3�t_n�|�A'y*5����d�����Bt��u��^_(i�4�QL���ՙ'�:��_ϼكՕ5�A'��ԇ'��8:9"&.��ŧ���V�^>��4� ��@�V�J�T)H!�H����)�͘�U-�`i��<��{���*���L/�}),�3vݍ	/�NM���[W����lثׁ��e���<���}�����������~�t��8��Ĩ���
y��ѾADH`c�lR��G���-�һ^$�6�S�TB<'�Q�0d22{eN�=v\x�QYXU�%���5A�����p*'4����p(B0��w �1���A8m��s��{Ӿ���>)��Rꅢ�����-� ]�|EI��,St#5�7�Ɂ@�S�;E7�r`R�EE(�B+Uh���+�<)Z�u��r�YxXk�~�Ͳ}\��額u$//�	��\����/1S���H&��K!b�mi囎�qAK���RZ=r�(gl��ЪS-:L���:���;��z�Kh;\ge/U+����V`�W���g�&[)��q.y�q�8w�(�3+��)Ɩ� ᇑ�E�4lӎaĞiY]C�iX׵�f,]1��'k�i�MC���D,߲�Xvm��$��ˊ�@`�v���(���r6�y�+T�x���{��W>�oO\��׺�BՈ�>��<GE0��g��c����P�/q�K�gdǩ�N��j�P �f��
��1&�s�a�Rn7d�Q�7/z1A�+n7��lQn�>)�=}bU��6Z��)�&�W���܌�\���ZEÒR��/ȫQ),b0��z�lw��~�+u��A��<t�A������ ���r���@60'2u�a��q8b�(��=	]��ޯ�\�1�&&���?���\�V��m���d;e�*e&�� �E�͝Zu���=�9:�di�x}�A�Vl�TY��5����蓫5�wZ)�}��n���!�8\? �j([}��������t��)EI���Bz<�@Nkj^ξ��G)4Mt��v�+���y����H�E���dH���[_9���$+8�lx����?µ������­©�nj^O]k]����P^:��,#a �I�וt�`h����PB���J��ID�)$�轻�� ������$��.��Ӕ7�:>�9\��0�)�X,����S�屓��X�၍�`mw�6��7��D�4�����ڱ�� ��	!	��ϲ��>1���#��y��Q	�A�_�x�V��O�תf�J� Q &!�ӧl��t�12��z���T�1���i`KH@��o�s��d`��I8+Q�32�/^�"/^��/#�B�6)���$)���iR��ϴ
f�V����-""��2)e�}�f*fad	�LڒQք1���ʪ,,��}��Wl�rs��f�q���ܕEQ�q'�����ZEu��۶a��ql���g'��EQ+q��i���FbZk�Dkb��m7L��l���ذ�ؑ$r�$��,�;#��[�l�E�o��9�_����Փ���b��[�}�0�˲�d������Ȁ�J10$$���`¡��`L #�������*�
H�!M�+�c�o�[������n�Z�m�Ɔ��3�Y�J��R�b��])���eY����ʒ�kel���<\>��H3H��8�@$T�0o����6lF?־^�� ~��A��(*���!h�\B72Q��V�?�8 �B��iy4n��C���=y`Ce�1)Vz
�S0�
�)�"5(@��Щ��s�dA��K�!+e�����C/���W�ER@OE�H�3�4�z@�I��F�L�u+=eU�)���҃)�M�i]�]��1{=+F�Q��H��t?��^i��U�f������!l��CK�aT<����@��\'f��d��	piO����(:�hZ����AO__g*�������������[��� �&�!n��AW���8��]�R�E')�*��F�AXM��C%E�`����#qѐ0�֫$�7'�7����v�<2J(:�� <?8�Z,�Z�&O]�$�N���!��� ��B�q�/�����U	�gC�M��H�H��a��eA�{�n�(�1�i���}}
�`F�n8��o�%X�6��5����G��{W�P��I�C^c
���{�pו�6��g��8��<�`�Ax��V���g�2`r�<�.]�� �2{u���c��#qg�2��0��i��i��a����0�8���$1����U�#K(
8o��bA�2��|!�X(fAh#�j�+��}py �tuy�J�CA�gF���b��6�B0���$Y��h6��k��sF!��|N(���׶o'ۏ�Q�$ΗJ�J�������\�ޘ��Y��_����r�ʅ?^���5	���:8M����ۋ$%R��t.1$�I-��2�t)�eW�� �z���}#a/�h4�fG\ϔldI^�><${G�eK�G���U�|iV.>#�W�H�w�����߯���+C��u�VVde�"�F�f�p\"�be؋-�Uo��6G�u�tpDi�R�"����6�>�]���I�O���y0�����INM���@+��S�H5J��gu�T��l�ཱ�LE�XGUw)��h(��*��ϑ=a�B!� ��=Ĵ���;z��`��4��s�K\����v��%%1�>�V)K�֫2�5A(�P���ji�z[	c`���@���}��6�%`�þU���f�J��:Q�J:`T���J�9�E�M!8��WC�@nF*(s��Y@&Ԥ0K�{�d�c]�P�H&��u/�_�(�d;g��������F��X�*'3K?3]��t�RY��{��d�!~���J��� 	��l�^ed��O&�F�!����fl&��#�,!�L��tIx�Qa$°��h�^o�mF%�N�ـ��ϊ�_ʍ��	�h��l��@x�w��KC�u�'��a>6�v�I������ |��.�U�f��9M(6G�`b��Q�xa5�(�DQDn۱I��5�j9�a��i�͐�Ү�!��XI����z�PL�6��As��$�IL��@p=aF.�?�_/����$��İ�b#�l{�rl7�� �-�q۶�cYa�~ 
SA�4-�F,Y�!Q�$θ���q\�0�n�S�8����-�o���~ ��BA"m�u��V��$a��&K++�R��g�'{��>�Y�w���5'k�f7��}��ް��Fލ��*�{��9y��W}o�m&�8��-jX�{�93�I�+�X��Q�X$b�a�AfA��� G2"�=��x ^�uo�'����A�Qd��$$}�q"c}%�=6.���2 ÂZU.?yZ:�I:-)�s���_�z�����do�Κ�\mб#¡n9$����4D����A�W��^�ГZ�)�����U��i��6��ɾp���W�U�@ "�z~�}��0��a걉
ZWE hQ�P)��T�
��J׉6�ᜒqt$D浖gCU�yE�<tc�R�* �]�k��q���x����������u���LBT*c��1�������z`O+bt��윣6�����U�5��@������6>O�����8l�����*g-?Ib�%RAW1/��0�"h�Z��*tB�� g��c�\���]�8���?�|���6֯W��~�^�1��{O�nM�K+�t�x��i^�4�%;A�P5�˪[�z*b���L�lz��q��F�����,���d���>B�[�a��H\X�I��qBy�!�Οg%\i�9��`.�H TC�!+5qH��F�>�� L(_W��b�z;�Q�3��g3�0*a|�V��G�r�7X����Sg�[��}���A�t��3s(��>4C3��0�G�_��p���Nd۱�Nl�Nb��$2�v�,��7,k�4���#�&��؎�M�8c$Q.�Ɍ���o����^$8���$�0Ƶ�=u�}����=�V.t:�hxx�Yq�0�ضm�[(7�QǶ�|���F!������g[�e��iők�nd�A`Ʈk؆���Y�k�<3�ǵ&6�~d��]�nj�6�dikc�͆R�Z�փ�J���K�~�K��Ե������)��K��'g�d-�lC܂��F�`��$� ����Xp)�#K��i�`���I�d�+YXj>VhV x�����d�����۾�>�JI�ٮ�{d2t���ui/-I�ۮ##���
��QH7���2�C�W�Rm�ă|!�T�nNJ��J��K�h4�E�}_@�Уi7<}��.�$���HhanM�:` l��!��1 �Z��9��7V\�`��W����(�� �g�)���د� �����&
!���� 6��CXgL"
 �f�	�W��@��ΐ���:L|=��}t ��}�+eUE�0o
w�
j���_'g�s�N��i���d�(��J5�#k�I�(�-����:�7�<A�W'i%�����(�^��N+̍�iʦƟ�
Z����n�@%�"�� C��	��f���*ɹل��b�>�����j��N7F r�؟	�a��a�I!�3����@T�f�P�4"��8��(�#�l��@n qB	^2�ˊ*�@�cC���N��iu[k��_�-�)I�Cɹno)_�7\�����m�9�B��p��"��~�iy��R㌫)�a���1�u306Ϋ���+����9���I�J��!Fմ�eY�r�v��RO���-c�ݻw��P�:��ksb�pty��:w�O����B߅��?p\����ÇI�8r�@{���o��w�0�;���q3�<ǈ�m���m|�w����;��B[:��}"�j�g�^=u�����<���9R{��������ã�}?}`���2�m{	�|�T.�ݐ��ީ֚�����WZ��~�#)����{�?� �����g?�������r�d��=��R��(�&C�$%�(L&:Ծ嬟r���jV/
���#�Jb���bu���{,[
`Cz��x�5�<�'�2 �G�"�5[^]�P��>Q�W�lN
��
-��{Q���Zi��(R�b�~56:-�:I�"檮H3W8=�1P� ��ԕJ
��?�aZ��h8�a92}m��5�b�	�+`�t�Uy:���Y!��3��(0�!=ͲNGuTE{��<=����l��(��t>sc KG�p�i��tvr�^��F�����u�x;�d�T�KdԪ��\��p�DqlYVdF�A�q�Fkr�?���l4�E^��>�|����o�fbFlFb�f�D��8�L3f�db�u#�2#ׅ����@5,P�݌�0�?�</�汉�o[60�$�f�.b�q�	L�B��yA7J?���:�vXO���d,ò�l�qr��i;�'DV�@(�mB+2���nl�~DÈ�$��8�-�N�c*��#�.*K#ä��FM��z�O,+,t�q��/��@M���;��~a���?�oz7�,��
�U��2�ku9yF�=vB�����ja5��*^Ek2�}> �b��W��R]KZ�i\�S'gC?��Ī��c�0
��7��a���oڽ{����#��C�� ���ry�k���O>�;����?r��ܫ_����C?q�]w�{��d	�J襧I�M1�Zp�[>�ē�;y�����/�u#��k_��ޭSC��gz������� @�	׃ ��	�yҺ~�Z�|pq~�7��г�����F��s
����l��T�?���<xd��Rjc)�O 6L(�vzVQ�")d3�u���1l���!_͢��Vߣ
���y5���`�%f�#��%��K2��+#�W���P���[�g� ���+�|���g������v�ZoH���  �79��##���@��JqE��`�"<���ɍ02�۴Z[g��9Q�}U�6m��k
s�S�B@ F�r���.]`g�$�کt3�B���@�I)�D��p�}ɺ�@�@�Ң!<��E�*0��[    IDAT�G%���b�fP�R	z�6�ㄭ'T�`�n|Eq�a���0�"?Toj�)b�h&��Ab$�e��i��m�!�`��{!P��D�a�Q�N��n5ڡv�(�"?l�nP*�z�8v� ������Z�U_nךK��[��^a�ŠrF�*iA N�Ȋ#H�Ȋ+�]�1���&�c��0I";�c��e&��QB����^'LZF�v�0��4�r�'�s��-�&#+#�B��1559rd����>N���;t�P�����5���N�t�=���h��B!/�vG._����|@.���r����7�(B��� 	���#�	�����hEQ�D������y��x��G�2��#���|�7Ƕl��]��i��}���џ� TR� �1�����Ǟx����W��#G���E�߇����s�y���7�v����ΝS����Y僘E��Nb!�an~n���ӿ��Z�ώ~��j�>ϯ׿��=�v�|�];����pH'$Eq��VE�:;��W��?�8��>��/=ϗ�]��S��O�s��"�_�v��(��T@<�i������Ԕ ֻ{I�95g�#$�*@���Y�xp�d��y3f@ajb]��1�����I�����Q;AW,TǍ�4kU�9���*�K���ĖC(�Ro	�`�C٥5/$ hܹ�t�:+��c@��R�EP�D�<}�Z�h������eUդ��C��!�_j���< ��.�a�v̶���H�0L E�����d�|>oerY�qh� :��$�M�NȁL�������f�^��~��~P1��9�����u3�i0!���U=�	P�8��0P�u:�4L��P�-�5���՜�gE�����j�ڝ���h�	
�.C�8F,}��Ac	p�3~�N̸�b��a��[��fԣ�LT��8t�؉3q��b7
�����n�f�I�ٌg��dde�l���ˋ?��Dg�	垿3U�]�ɿ�.��ٟ��ݻs���NO�R6���6����љ�yy�أ���Krm��X溕���>LV���S���V3ʭ*���$��y�:��='z��ѣ���t��wۛ6�izώ_ݿ�-����7��&��8�`\��n~nq��S'���j�72�y�[���7�r��عsr��1�'�h��--ז�Ν{�=�f�Ф��{���?ݳ}���w���3c�Fa��@� b+���w)/+յ�̮,�ڧ?�����ھ��s
��@�O�f�ȋ^�TF��X�bf�$�DAd����ߧ�=��Z$�A7Є-l�m�RG@��P�9E�A����-Lь���k�q��mw �w'��d|�_��[�]��o�9��E�2V�V��~I����JjYP�Egws���B#�c(�qǉ���0�01�@��|? ��e��u,+�ضoZv`���A��i��i����� ��@��P~�q�*��iZ��8�l�0\˵m׵|ov���r���y'���;�2-È��"\��q�~�����N�_	�Cq?0����f�~^&�8��fb�mbҾ�I;��Ј��ءaU�����������v�b>oD���^���wu�2++�\.�l�t���ğ�*0�G�>�����om�������;�`��}����Hb d�( A��h���Uy���ev~�Z�ڬ�a'I2�1��hy��w��2���=yB F������֑�����G�~[q����?�c�ԯؿ�GFȎnCq/T�&�0*�k�K�Μ�͑���s�=Ǽ�ׇ��?����}2�}r'*a�0!����n�,./-�=w�߬��4e?�&"���n�����?�yt~aU	+8��n�V��?_^l��8��d���O��7v�=�L'�9b怑�Q��q���V;q��Q^<f�B�!��"�C}�c0����%v8��J���6 t�~�L�^��t;�V��w��$�H{�|q����knݷg�h	J^����$ݶ��$�.��`@S�#Q��5�	6[��6�Ql��3������l۩5��z��Vkt;+�c4��Œ�)v-1�GI=
��$�r���q�%��Vێٶ�@R'vP�Y ҤmY��yqӶ��HP�6r�8�hĮ�&�2�1�[N����M>�@D�==�`�?~<�Ç��WV���9�;<l�{� 0а+v"���Sv��H-�����?bi��O_�����-o��=;����NnU�"L�`�ĩX���:/�=~�:wm��f�uΰ��(���p�e���Y��%A�� �<j3��v��ۭO�ڝO���/}���Ѽ�o�mjr�?���[Fǆh9	�cX"����k�dy��|�ܙ{��G��F�7��-/޻��&&6�U�{;��Q	�_[X9}��{����|��u���,�G4?>��v����[7�;��Ƹ������ ��x~�������>��>�������s%��?�=_��]�z5�K�l�� p� �jݮ��zq�����4�q"C�:ɣ+]�+���u"�ۅ�Zd8�cDQdt"�:�ԍ��;����`S�"��:ݮ�8�U(�m~��7�����@_l�f�:�	6�ﱑ	64��AU�)Wk��v����r#��ӞE�,�-'�3�X�J��n��u��h4�NOO��y����Z�����{�|�;��Ç`�����[���l��c(a�sV��R�+�Kr��مٹ�O���o&��o&���$z�H2���8��>��/�_�:7����ڝ��z��9��~�s�?G·{��G�4�s��o�t��w�oanwથ�-�9C�\Y�����|#����÷��3���ͣ{��+v���UU&��gΜ�_��/��7�g��׾632:���;'���։,f�Q��d���;^P�T>��^��#:�1�_�q���x��n�s��|�`!'�Q�%&��N[Z�Mie���jˍv�b��<��}+:�DV��v�Q��{�B:��/�v��^�7�>|�Ўɭ|��7�l��F����臲��*�N��p�����{-��-y�%�����7��4l,m[\U��9n�0����V�h����/}���Aw�7��c['����}�96>l@���GP�
C���m�W��S�N��������{�U��7���7��֩��eb|/�h�ѤNT��!��_[X;{��=Q���"fa�j��ݿ�cz��S۶0�f9��:��l�9o4[�ry����g��?���X;�,o��]{o�7[��߾i�o��Y�c\�լ�߳5��4����p��v��y'�(��逸*��|�?ˇ{�M_�ߣw�o=|h���?9�w����!�-��GC�WM��Պ<���sK��R�~��8fd��-�zu�u�2Ms�v�dQ���n��Vo�m�[�
���k>�l%�l�w޳w��it���)p�3� g�r��j����3�����9r�y������w����m�&�MLLh8Z)�9�\�#TK��s��}��s���g?��0����~���~���aǎ��Ln��e�4{��4�sɳV�E�����:��G����x��՟�OG�ހ�{�ύ~lxp��\�����u����2���z~qu�t��|�.2��bL~�~���;�z�����lzz�O޴��Ѐ䳮֧V؅�I��Ғ<��#�\�t�=���Q���ձ�C�i�K�d�m�%�2]S,t�a.x��������=��>����������ʦM�x��G�����ë\�t�<u��3�μ�ß�̷%z�S?�Ç����mٹsj�h�U&�:�ߴ��C$0�������Qs� ���[��Ν��~g���~h�ÀBM�(��C��j����gf~��G?z��>}/���A��o{�������=I�H.�*�ˍf����4^��KK��k�^�o���ڵ�Oطl�_r��(�+3)����~��c=u��wO��g�~�H|��a�S�n�'ŀ�e%Ih؆&Q\�h!̚W����s�O�T�������������`��?���Z)W�O�<��3O_��ȑ#@�n��mo{ۋ�m��Ў��{FF�HF���f�C?��R��/^������w}�c[�!'"oy�[������75�m ���ѥ�s*�j(��Z5^\\�����#/��|^x���w��; ?�S�����5�'�<�otS�d]a�+� ��f"R�T�~��ٳ������/߈[H�ҥ�~��}��i�p_��W�	�J.µZ�s�̙?�4;�������&?<�mb��Ѐ������X�-�^��h���|��ճ���|���B��O����?�}	tU�����������.����(� ��Q�Y\gZeAQ������eDQdHI'�wUw���n>�o�
���[��$�Jݷ�[�S���h�dJ�fM���h�ز�����4
�#zUu��=��~�����ۺ�F����*��.�@}D H��sZ�;�ݹ�
�=H�`¼} 	C�/ D���ۿ�z��ǖ�|c=)���~C۵m7��A����؞�":n}��f,W������~����޽{_԰Q�כ5i�
H؞�n{�`W��c��z������OҾ�}��۴i��͚6·9�x����lx�c@µ�ڷ�.M�Ѥ�l�E�"@@�}�ݗ�ݺ���k��\�9�r�����7�c�m�_~�s�#�_}�R�����޶mΙҰa����\[���u��4d\Ւ?��������+'>�~��-

�4mڴ]AA&�'�q�A�0�(���UTT�_���l�}�hڴ�ԦM 	� [�K���A�5�@�X�C�������I�m]\�z�uqW�M��b������g��{����� �ˉ�Fc��L�+�.���~���;w�[�Ҋ�� �{�w���Y6h $lK �*oЃ�c�j��w�=?���/���ٳg����U�7��A�,���=��L�5�д�G��~�Сq$_���ׯ��xF�F�=^WF4�2	�I���fF��*+�Ö,�����$\o���8E��A�O�>͚�j>��λ��(��@� .�ׁΒ�_~���]ߎ��h�R���sG�sZ��BQq��99���	)*6	��	��}����.~e�R���ѣIAA����E.((���pbp�<N8`�zEE����c/^LL ����WXX8�Q��B�ǉI�r�0�'�)��'>>ZQ=rɒ�ߒ¯.�CI�.�
��"�_����^Բy�gο�>� '�tK�2WV>�C�0ڽ��������ٳ�B
���{�Ժe˹E�����eO$a�7�ط�?�8t��y�'e[�>}�y��7��
�����ghce:�C0�
�����tE��U�~h�Ćax�=���S6(*�A'X��<�
kI�g�I&S[����_xa3)���:����P�(���~���7�|�EjX� ��L�=�ʴL������B���~��-_<Kj<䐁ojР��7l$��L#�۴=�X<��Vݺw��a�g����v<����z� ?��u�A�Ԗo�Gb��c�V��w`I9r�}�sR^^^>�k��Z Z��l�Jx�4wUW���5k�ۤ��P���Bm��#0h� �ϓ;���֠� �0L��"��P���O�c{�7#�Oy��牌�1t�u���4,l$���3��`�7�	UU�>|�r���7�ڮ1cƜ�p8V���ր����X^��j�( 	G�q=�����4i1O��G�:��pL�x]��B`�Դ�i�Ў	g$k�#�k-���X׹>�����{���<��ߕ�g=}�Y͆�qY�>����U�<�U�:;x���`d¬Y�@���w���z5� ��]q�S��*��!MM�����Ǫ��|�I"=�p�O<����$�v��EB�W�1�2���I8�В�Pxu\�F?��c�r�O>9��,I3�Ng��%�.8��S)he��&��4-�X���mq�zxP���No�"�{"���e�&����
Y�0�e����C��$*��?O~��_��N�=�����-��������'Q�D��ސaY��D55�﫪k�=����:O=�T;�g�t(Jk a<�Ĳ庱�!c�z��F*�����1�>�(1��	&�&�����!��9�9>NHԨ ,�	I�,~�ǣ�<x�`ȩ�%�z����)�����������=��e��吅IH&f��-��WhG�Ϋ��ybƌqVO���:]��9��?@u4x冩#+*OS�T��_QQ���?���]�ƤI����FQ�s��!�� P��Y��_UUWEc��dIxz�����KJ�b��-L�IM�hc"��a�'��j��̤��dס$|�H��(�ӆ��)���<�$���f-{v4�L�{�.��UVW'�ˏ.JT{t��iDԀ&O��tJ��99�K=�M�@f1����L�B��Б�Oܾ}��7�xč��1mڴV@���VQd��RHׁ�lO��v.�3TU}3�&G�5�XNxҤg��,�Pq)��'�	�C^��� �����c$Ѹ�Y��	���$\O7��6E��D`���JE�����܎�$H���ͨUUU�W�/9V~����*Q�S��ɓ����jn��J��k�p:��K��탖�`(r��f�۷�YREc�&�j�9Л�|!����4�:6�}�$g�[sP��N(��C��<y��k8�Iq:��$��v�H���</�i��4}l2�z§����)��o@`֬ٝx�� 7���R��0�'�v۞�����#K����Hx	�\�����*'?�8	�킗�8a(��"�X�CG��ݫM�5k4���g�}������N�%�,�X$|<��pR&a��E��G��!�F������t�ԙ� �yMR���%����|k�X�q��0�#�i=�iu�)�LO�P(��瞛{1ˡ��\Oh��x�	@��	 b8j�k�C��,)��ԩ�߸�I��T����P^��|rs}�HpkMFf�aָ��9�(�?9v�X"��S�6�Ei��(���b�����h�eRL��x��Ph��ѣw�ԍ���&N�xÊoȲ�Wo�|��E�ݮd�φ~L7��9�\<b�"�g��O�%h8��CJ/H��s�,:״ҫ�s=�Bu�,��`ǴL��|b��Ƭ(/5�=��#��ŝ���%�������<p���xL�@D"r��za<~�?v,����3g6��uI�Dc�M�m]�d�IX�4�5z������O?=��c_Wd�B(��3�f� 䫧�d��ìJ�ƤX̵����.��%���v��K�/@`޼e�S[�s�.�A�I�'*�)Lr�C�R(FG++_�	E��3&@��'N��Pd��^��kN��x��c��$��j�XU`�cՏ���	�fM��0ť��ۑl�$�i{�'�0��@cs"�
E�<����H�k�'On����,^�G�fH^�cO8�F�aT�>!�,�$Lj��:� E !�dɒ�dJ_��^��ٞ���0��7��XUVV�E�<���D�N���"�e_���n�p4xtY��,	�a"���<x5�{�ᇉ�ʧM�V���%�t�[���|��h�M��1 aUU�F"�q�G� 6�k��\)Iq� &�G�"dvXi�z2�����"Gӏ� E�"@��K�$��b�anv:;g�Na�<a �D\E�TT�7n\%	ǌS�u9���ͽ���0��4��h�O�4��X�����0R�����Ҟ�x���6	�H�mOX����a���I��&o�*�|{�<`{t�te�#ܲ{��z��0�G���tb�'��A�P2,XP�PxϠТE<pX���$��E��h�;G��HxԨQ�>�{B^n�}yy9<Tg�<�� �d2i�<�:8<d�?�P��������s� Q�Z	�
������Ǎ�৤��S���L�N$��T/ a��"-�pJ7ƻ��*:1���u(� B	ƚ    IDAThٲerJ7�#ɂZ��S2!�)`yC  ����5��`RC'ƍ�v+��rss�5hP �W$�s�!�>UU5�Uլ
��C}��;�?37bŞ�X�(�b6ך���2-J@v��m��ՇG���#��'>ۀA����ތ��p��ǒ�^q�3�kZ�XYޣ$Lj��:� E����lqq��,kM�9��q%Ӳ�V����A������p\�o���$�5j�R\�?�������Q�����±�q\| Z�R�p���ꚱS�L!R�=�?�1c#Y�'I��:��A�����/��5M�.O<����!��1iҤ�`��y�� �pV���RD;8��1�����S%R;DסP(/~�&�Jm{uXT]ۯ4#5t�0����%�tȀHIw�1t�tw�Ѓ ݥ��04�p��{���������[����|�LKp�C���e10�+a��Pi��KB��)C�%8T�23X�՗�ˠ<z|,bP�Ϭs��C�M��ni�?w����_�^Ex�S9�c�H���ʌ��}�&����[/��h����6s�涘��1}۸�AiC�CX AA˄�|V"o*ʰ�3�J�?�6��)}m�l���8�$�������W��Ep�݄��L�cn�E�F��ږ��S����Z�Jց��u|�ȸb_�@�	�,�����]��븩{�+��b҆�E�|�.����Ƃ��>�����2��������I�,�q3AļsE�eM�3���yő���C�c�4��I׭��t��w'�pƚ�y�fz�6�"���oJ�Ԩ眝�G��.mq�P�l<&'��ɸ��y����K��#����k|�A����M��:��|��M��{7�{x�ߣ}-��kc)�J���2���&�L�=�x�29�
%��Ւ�ѓO^K%�I8�w�;D�_a�W^X���4�a�߰��N������;S�u�&m��iP�����h�U�>H�-&^>��f$"��o���z�K ��5/�U{����[����.�s�پ&�d�!C���B�#��^'��K�d��bi�Q2�����Zd�ú-�
���X�)��v��l�uP���B|?��m!�U�x�?�y����K=� ����?S���<^��(�$g3�p����X����
�f��NL�P>�c��ri/�B��y$ԺJ&�� �Z)�H����!��2&�ӆ�Ѝ"7������"F����(�pYAYl�:ĳ|�~��5���/����,{>J�]�R�ԡu��,4W��llߛ�9r$�@�2M�a��;⾴�~��+��F�ڷ��^�T�aY"�x���'�;ϸ�������2�Xtgn�I�*o��K:|o�f��`���	��>��uA+�^p�:N��flk˩��D/�9w�'_9E�o!7�j	̭��bS�8B��ZR`R�O9�I�ޥ�i�|�Cm�g�/��2��cI�BT��E]2� �
�.����u�����	���P�
�#�3 A�����hO�TqX��ƹ`��ۭ��(�<�!+c�04M�����E�>�8:M2��TH5���p⊖9�L��={��h\<���/��o�U�Ԡ��lK�w����-����(/!�n������f���s��w��Y
3�O�hL9��z�e.��l:�bh\60N	�}����	Ș*5�RNJ8qI櫓�v��dQ��4���ɂ�EE}�jR�͊]Ɔ�ĩ�����$��������/���V"��iW�}}��ǁ@�vO� �Lo��7}��U8�=��ޟ�C�Ⱥ�Y�.�h�ŧ{Oǥ��/:v=����>/�.�2����B�k�O51��å΀����\\;�P�M~���A�-Țn�	�q��,��v�B*A��;�JCF�r/=��.�Yś� 4Э	>��f'��˂<�t���l%2����G�;³Ѳ]�8�tn������Ǳ���}zJ��θӖK��I��b�f���&���1�N#E4��C�ۺ��IBQC:k�)���b
О����e���Hq�'��Fo���%���A)�"0�X� a?Nr���,�	;wtz%�U�����_�Xr�>��|6�hKhm�6|����)�� �/h��~�+2�q�Zs�]��O�H%Ԭ�Ȕ`��!���Rd[��T����������5���d0�4�i��fK�������aK�S[�VB�������1Swd��`���[">�T�������s����
�ɒ�W��g�L�e"�^� Z��'�Q�O�uSe}%͚��p��Ȁ�N��k��&��ߞ=�.�RT��t��/��մ,�ˡ火�(Vi�UK�=Q�ɐ�ETI�gL��Ao@½Ǆ��%)))E����&W:�q�o(QZ���R�H�:�$�㶮���d+�3(pч�<T�Ǘ^�E %�`�I��P���%��4���Ms5P:ʊ���E�+�LQ'C���jW�0���a�8a�-Y�7�H�n��.�m��و=_�'/{�	S`�+���`�1���VuD�ˢu�?a %�o~�0�-�T@ԡ��+G�Q6�Q�i��5���ž쪦�X��������Aܘ��f���b^��9h��n���U��_�ig�y�����.دi�`c��}d�u�{Zj)�u�#�xoME�p��g/�]�j��X3�Z]� K؉�'_�<y��{?�J����9!����_7���s��7��V�q�����hOnj�3a2��M�G�)Vה/ȶ/ZP/,���.b�_��w�׳�h�$����&�	|1�M�L�v�W=��BJ+�J�����dG�nA���ŧס�* �4,�"�W*E��N��gGky�L���jKt ������|~���F�ܘ��O��s4��{0?�Z�(l@� 	�&��M�Z*d��w�y�R��tF�}�W�������6�����e�[������.��\u>����X�֯�yI]�aV3�z�I?F�$}�"��R5�a܆��.�ԊA��e�'�l��;e�fu*j���x*df�n�K�Y�r�I����=�)�NB9""l��(�?gS"�A��Վ��#r���d�ǂ	��4�>���T�.���T\����}�y���&�
���[r`H���]�������w��J�!2���PS��Ȭ
�m�i���NK��ǎ�클e�ڒ\���z�}�K����(xu������CpF��7�gIr�͡bPm;�N9�0�/X�)�q{x��x?�cNĿ���ݹ�Ta�����VN����}��{�/*�~��?��7�0�c.�w��|,&�� ������MzX�S>���T�<��:;� 7����rX��%�A�U������p��:;�4dA��m˔���+5�s.�����Y^�>%�aW�I`S�'Z�����3q������ӏS0�=QJ�
!2a��;�y�-�~��L��o�����9��F�l�#�'h�k�J�A�G�W�5�׺l��^QdPl�U}�聥MN�g���"ǋ_S˷?R��x5?t�\0^'���;[�<o���������朥�W�J�����Ҩ�Ϙ�x�V��5N��k ��AƳ��J��l(�)��j�8�|D>� |s,Z�)bgzs�]�&ȣ�2�}�� os��Q���ݦ�����e$R��#�r�ߡ���^��{����+��	�$`g%盝 ����8M杫���_]��6T��3�E�W,��G}��j����LGƀ�J-NE	YN�3�>oϗǳx>QT+�qn#v�V�`�/�Yc]�v�
�0���MM@'��eČ4��^*hy�M�n�М�C����|j#�?��Ë"C�G���BL�L��"w��y��ñf�<�y�%�ɶb!:		-�p�]8�u���	0/�M�V�����G���b�1�o3���܏��	z^Ї'�+�D�f�������l��i tQl[<>�_� 1x�F��~��6�<�y�9�5M馋'�%�0��a����P��¬�V�� ;�5�}���]�W�Vv�q!������9;�F��ҽu�����
�x쫿	�����<Ol.��|kT2� ª�R���m�ܣ-��]���� 
�###�!���]bY��k!�1n��H�)m��'�kʉζ�x�Et�`F��w��� 
ٵ���-�Bgk�ޚ�v_����#}�`O��~�j*_X���U{��6�2w�ޚr����M,��|��'����:��toW��!���w#S�93+d�����R7?�_���������?�o��  j`u���<<n��ex���@���u+�j��w}�C�l7�{ȝ"tp���N�y��|��qh��Xz��3~J����S�_���ӣ��gO.5�a��moæ���긑d����,9ɾ���5����FY!:�t�bGܓ���n_�05Rd��GN�Э�Q�li8�WP��G$�]1 ?��#M(���l�_[؟��=VT��zE�g���9C<z	��������w�]���.xH�:ۇ(0��H��|N"|����nS����*��El&q	X�7��?�2��\.��$.�f���]@X��{c�/xh�!�2p5�ht^��iE�5`؁%��';�B\ T�1�^�3a{
ܒT���[_��P�������~x���V�1D� �w'X�h�� jM<.�֖Zj�t���-?kX��$O�ŸtK�L���E;��v���U'J+����3"�o�}��<��h��4�bR��h��SW�<\�����Jdޘ�\aFV��չ#"��i=�oR����/�����ya����sc=��}F�?���4_1�����d
w@#���xP�k�ep{���R{��V>���g9�;�.xPw�s��E�a�)w��r�kfcK�/��d�?z���<�� ��B)!"���O�M�P@1� ���j�I���TT�y�	Ɯ����_��3�b>��~�;K�WN
USS{��3�=��H�%����4zzL�&�,�S)f���R##�WQ�J�C��B��*4%�Ƈ 3�l��X�f�o�	^>'�w�����1�Q0G���ת��eQ/�m9���sT�P�*�2��:0�嘓9$�V��;Ttv��h&���K���*�\��m���M� �*Q�ؚ��f��ϥ(�S�1�b����G�ht���3_@�]贮Φ�V�"E�P�C_�5�+��h����uS����T^^{�¨�sێ�5N�����I�ns��rĽ�N��׍��0��+c$e���S���'(���|��� m�zh?���XZ���=X�@2��B�A5?���j%�T!oN���4ʊ��yt8�ȝ���-����m��.����U������8�C�6�3�#�p��
���X�s��^P��.�ꝺ�j���&'�j�tg��K:�PH3�B��*$�,S��MQ��	O�:~�s���;��Z5���-��T�ms\��*�X�Y���7�\*���Z�o�Н���U��<�kPR��UI(]C���L�o�YM�+X%SG;�ĹUz��h��x�����^��W�$K����
qJ�Ž����YY��W�r�����ۚ�X7ښX��e$�HՄ��T`!}���L��͞���j�E}�rYF_UƄ3��x�|8ӑ>;�=C����sC�I����5�
�����W����9�ҫ��;���Xd��i�d	�b�%Sϐ���W|�+'5��enw�7\ST���F�	[��b��DW������|�`��*��u�2)L�^���Ŷ�!r�	5��XZ4ɌGW)XU�w{�Eߌ��i�hs�%�)B�D�&J��J@$�_�}Qnv̑[QW���~��͢���Ή ���ѺpmNů�6�>�oU �P��?�����|=�45=�x5`�����-{��oN�i�}�c���\�`o�h���^\�0���~��Ųۀ[dE�k0�
>�+\Ʒ`}�',C�<[�v�ؾ�[�F�K� 0n�ο �y2�T��4�"q�l=]Sq\�9dƀF���w&�!��%}9v �Ʊپ�`SZOg�1�ȡFo�x�}fzZ�QE�-#���'#��g����Y��d���~U{Av�[IU����� ���V���y���d��i�N|\���Nu������u���ȑ����s�^������a.P8!�&˗8�� T��0�ҶrL<\�w�'�:F��dtb2�q�<+�c��P���3ӱT��Zt�b��K3n\ y��vX�͑�`L��kL{c%!i��T<Fq�kwd�3��{i��[5���W�#EP,�蚞����9��`�G��U�\ d��I�ıj0��q%�[6WX����N�Bȇ�4������׼ѓ��+U��1�g������j?6��+ߘ�O��N��f�2�`��e����T�,��;,_�x4�Q7
;�		��"k~��
^xwr7��D��v��;S����.f*TXC�@�&�r��^C|,�:q��y�����S�����flL4T�L�B4���0��Hn=�.x:㊣�f1,��N^��Цh2�c:\T9�P
�qLs��IRZ�)�~:ZG�~��G������^O+�4��u2{���"�vyƺ�ݼ�H�ObK��ku�-���L��򯽥U4G������})�%�E	�G��ǆ�����Χ򪛩K��tr޻��GMįq���3;X y1#*�"��dbCxP���b* �S�
�Y�ut������F)`Zu3}#h��Nti5y�R'��u����Y���{�H��[pPf�9:��2Iއo����.U}�3�����8p�����{B��u��5H�N�bAU��js܄w뎫�ł�����+�b�Ĝ�ƞ��|(����ք�]��O���t�dEǎ;����y��Fв��6�6B�=K�Z4f�L��Ɉ�_n�x�_�y�:�[�-t\�_(��VVV:����j�3 ���))����~�ν	�F{M�e��N�KѦ�|�O��э>L�	�~G�_��ҏ�2D�Jhw��e�Ww݌���I�ظ�g��o�k���<���0'�j����i�]Y��CI?F#s��u��P����S�'�B
��ӌ8}$����C���l�8_u�Dۧ���`�kG����4���X:a�[HV5���@Y��o�&��������5`R�I(��S��`��YT����Jx�D��&�N&��o���df<`����P+Y��
�I����^y����R���		FL�.fx6����Gf���[�bo�}RS�ћ����-�<�r�(%KBz���N���h:���C�C\��I�������/�&i�!�r�_"���g~5�j�����6X�`y5�b�i~b�sm��Ӳ�Y�Q�{��M=I��2i� q�Mg����Hr־�[�&,�����Gu��Ў�X�kl���k��IN��)�岎-��!)ԍ?���AW�e��^;��zc�ײ\3.d�:* �g��&�nB�p��@>K�`�Q|���"���'F��G��XЂD������>[=��p��X5W�,5wg����R��2��i�Q/q��M<|̐��XH��=um�3�cƎ�z4�[\5�@{��ZK�;�&��$!�z"�n�,���4tu�;zj����#]F���S�rR�GX��V�e�&c΁QJ��/�_#�xu���>,g[�e�qX�V����{�n�j&��jSh N�� �f�i_�Բg@��>P1̌�I��:��,�n�L����%)MC(I�A����j��W�����٠�ok!�^W��,��b�<���n=V����-k��-�����;�c$��O
RBY����L��T���a��G��/5zb��<� i�`m�QA�~���7��]b=�k�X#�v|���������ٗOc�	Nq��~���O�J`�qL�:;���js��3��?�ď@i|��8���!��R�5��(�B���ddg+�dE[W7�Z��4�o3������'>�D���ɔ�����?���>#g���p��pӼ�͵���U���B|e�oznm!��������������&t�Ii����+\�:��[�<=���䶹x�؛7�?n�*��xOɊ���/��Xpp�	qj���p05�쾱�Ba��I�^����s�1�j�d�8�V��y�����˅ɦPtz�RHƣ�����W�g���)�BL� ����������:��Іk����I�x$��v�U;����(/���(�aN�����ղa=�Hwi�݋-���sj�Wl���Lσ���2���R ?�\���.^�*�U���v7�'��R��k"��em�Xeu�[���@��o7��,F�����>GC��������.�<��
_f�CɄ�O���8���d�J��]:�sa����0��Ȧ�	�!��
�js�e���{J�>%��6�r�al�-��O��j|���	"��+�L��Ų: j�w�2���k��4��K�yzq�kߡ*'���΋b�
P�w���~�@߯���>��(�"ԕ��K�*�vY�������[d�@M�l�q 6�6��b��C#�Hɛ�r^�~���G�?P~#H�brtL��f'����/[f<:�r����s3G)�� 
�Ú�+��=5'�`" x�RD?O�
K~�<�U4�2�wrN�r�����5�m�U���s!=||�r>x"���:|�w����x+�TZxqØ�IH�;��iqY�ײ[n(WU�hK�)ff�!jC\�sZqNWVi�g�*����~;X$�j�F�L�@��2�[&�g��{�p8��wE=;��qefݦ_����+�:�J�Y����!*���:YYM���5JG�K]ٝ~�U�I�lQ#o���rp
;�\ܪ��K���!Y��U��*-U����r�i^a�]l��ny��D��m���ʻb��+��x3哥?����n��dʇ��V~D8#���)�"�w?��c��7g�W��wR0��w�x?͢',���-X��e�hAA�Q�D���5+���N��~��k��� ���5/1P<n�I%-p�l��W�-����[hR��9VJJJ�Y\�Ï���zK��f��[f&�6ڿ5��z����������;���F0,+��f��P�f��S��	�:_`�� -�65���Hsf`s���<�eP�]�T����R1P*����J7e̖h��A�+Z��۲�F.�
N��ó�oU�}�Fv�+m��Q�~G�:ߗs��Uq��~���<���n���,̠u�� ��%�mJ�r�rK�WwU��z�5�A��e�֣J�{��c�!"y�m�,��N7T�����Zwt���9��t�Ѵ=��k �`�^RR���|/W��v?�'k}-��J�t����F;
��R�7�7ٖ�?�ḿyN��G<�%�@�耄=��������'�c|���e��YA�vwU�4�q�*)KW��M�t0�����ϣ���29ӊ��ѳ�������^���8�b�=C1�D��P��Jg�����ސ�"T�~&�ǈ�|E��X8�����2O��s�
�d] 󶱸�)p
�6��i�m/N���_I�N�>�@"�>6������	�l�p�_7CU�����X�=L����m���N�G9��D�q�Lص��,j��-�r.���o�G7�*�G����U����:����++�훏f	���O`���L9��Ѻs��s��ݕ�Z�2r��	���z���9 s�����]䁏^�a#���n�����W�+��Jؤ�������P%g� PK   ��X�>�~�< �= /   images/ff8e3ab1-c379-43fa-8f3b-dd687c341a4e.png�zeW\��-Npw�w���4��{ и�[�Np�K�Mp�Kp��9�޿�lk�k֪��Q�j*�h���PPPh�rRPP���/�>�|7h7Y	��i�#((J(y)q-o�݈9��-�=*g7J�u��$P���?V���Su���c�07	��1��T�+ �!���@kȟ�?���>�����N�d�~�|����_s�3�;=?�g�".��/C�.B�
m5�lL�K�?�h �p��	/��K�<7�)��p,����O�j�p��\B��z9I���#�F��� �j 8PT?u���?B��/�od3��zr��ܜ����10��ǁq�����t�O?H��-0�Zp�P�.��9@ vU� 9�˻�	�4ʈ�)ޒ��W���Ý%Jj2��]T�� p�ֺ��;Ur���wAF������ؕ�R�D��d�
�*�����ۅ�����?R��r!e麗W����#^�������~�񩣧'oLDY����0=l��Gߊ��OU�w�*.����Ŀ����Z���2����}����D,�6V*"8��|����h�O�>]�|�8��&r�y����3�>n}��x�r]U[y�r��%�[���0^jt<�>[{��_�
��2+�%�*Ҏ��fq>bƤ�h��)�u<�&ee��F�Þ�;=�ed_�v	��^Uu�L�C�e�^d�T�T�ڛ�l��W`Y'��Sutظ{v��(���SZr�-\�d���w�ݝ���K�O�v��=���?��w߿����cggEi����U�%�5��v��&��8�+d�%
�qOi�����F�nd�YU-b3Ǝ��&.����M��,(g��]����ڻZ��ݿܝ��ooΖ��Q��Cg��4��x�s�S���k�oR�ovȯ߄D��T�9�?���ft|�C/����q}Dm�rǴc�����ZL�z8���I����dlqן9�\le�T�<Oj���QҘ��idq:2�U���Ȳ��n�.��@}��d�~�*�����]�OQ6��{�)�D�����������$Ly��ڮˤ~r0`m�E@a.���+���.�%�F��.i�<)I�qMcT�����_�0��խ|LGZ���jd��s1[W�;�+�	XN��t�n.��(��+P:�"p�6�}�8@��@�yk8#�+1��}~����
���]jnn?��g��ʇ��,����_9j�"� ���luzT�=�;�9*M+�AF|�R�Q�Ԋ9�9&�s��Z�QR��Q�v�L_֤J��6������,Ǽ^�맡w�#��.;2�e\d�QN2�p���h�Ө�;#O�u#
k>GN�y�C+�������ii]�*����W
z2t�Y['�z.��hO�X��"��U��x�Gd��5
0��<5ݤ�m�H��(R<�4��SYT$C������t���������9�����i�����H�ʐ?��� �#��?l����B��T]���zb�SN����k�����0^D�G#4r���q��`�g�K���6;�t�n�z����+����3�l��%�T�4-��T��Wa�ڕW� �K�l-M������v|��;����t�؛����cz�f ��G�U(��@�	�5��%�R��j���on�X��]X�C�h�T-,��)jl�V������"��4i���Ԩ�ٝ:o���+����t�L��,H���L�Ǽ)��p�[71'�v�TV)�Yf1kf�TQ�w<��ea ��鍧�U}���=��7��*IV����3������bȜ�7��5�h����f�� Q�r�ݟ�_��Z�ݎv�{����e9�lq���UMU�n�d*����'�*K�C�)��Gr�!mQ(;�M�8W����2���ihc����3eMy�H��q5v=��J5��r]���9��D\)�_� ��g�_�c���W:,����K�SbQ"۔���u�-�����J�:܇C�zE�V7�~/�7�nטo[^}ewd�����4Ȋ�Lc���R��������qV��������{ւ�4G��q�H
���#��d�p �k�0n�R#^�����?)S�R�5�=vgj�=��6�k6�͚�^����$c�F�l��P;̗_���1���d��w���"���N�D�N�Ʀ�Lĸ~������%��y���]9*�1*�/9�wmi�*����ց���n-rTa ���I��u�c�����Ff�~�x(Z����c����o���}����$�+��؎�M:A��>���ΘZ��,�tEP׷B�C�����p�c��>�,w(:��2�$�Q��oR�qS7��f3�~���U����~�*fdb���ℸ�}�N�6�|�_�`���U$Z|-�Ƞ��zp*+�5%E�u;��6���Ξ�(���_0t��q��]�4�{�z�5É,� m�
��)�5jh�����D�&���Q 2����N�,��y��z���e�B��'Ԃ�>P�q���z��<���O�4l��Ȧ���b�z��84�E2��ge�h���T#�nR4���!'��΋�E�	֒�<��v=l�c^Hrȹ����bFhi�P8Y�e��K��m2�e1��^P��]�'�����iӐ뇵,�[�d]Fa ���i�o�W���6��ZJ?�P���NѮ���2`оd�.��Pǵ����%�TZ
��6D�?eLV�p��YF����̞�k� �'NG�d��B�?Z�|-���,�%iuz�7a���M���M�d\�YI]?�i�
��JN��oUpb6\�Y	����:xF����LPL� 8��k�!�~y�W@�+��=j��<�A1���Jl�|��8ߗ_�B��*i�� (C�<���P�=U�t��|�j���lH<��K�?�VCܘ��h���)�NFKp��D�3��S�y�OMM,���?�Z�p&�e��Ͱ�&��0�)��5�L9hWR��2����j�O�{$���I+Ҧ�!�Uat��F�V�-�;Et� ՠϛ����^�4u~Ă(��Zy)w��Vh㒚
[����H��Ao,R�!ԟ�;��7Cw{�lr%����SѤΏ3�7�e2~�DԻ��+e:,�T!�iA?F߲�E�4�Ԁ�xH{)�U-I�P��i�0���>gk�-@yx�X�~tz�g�%��&U���zJ\�� H�r�$/o�p�����f�Y��榨8k��N�6�����֦��p�����K�?������[�u<B�t�3s��3�Bj��Jc��`�7Fƍ��A�6Z;���Y+ԢU��8l��g�c��| TX�������A�Vb(��5q��mp�9B�%���n�_��s14%P��+T�1�`��o6R�!��o8��FrS�Q����W||�F<�ݼ��ͺe]�T	�'��f\�f�����T�T�$L\M!Z�Z�im:�>�f���Bc9;�XĨ���^�o,D���������� ��D�����_�ܰ���:_�m�����:b�Б����,�
k��HNW���I����&�o�?�O�(�C�&Xx������<�D��9/���n��ѱ�tׁ�������L���H�B[��e8���b�&�N��\�Gk�<�m��}�/{��\.kq�ezAϵ�zI���WmY)�1�U�u�ʣ5mLԸ�������y��Vq�D�n$;�;�Mk�H�+C��K­O	K�����ʎ��4|����d�iO`���K��פha�V,qV������OW30��s���>�xX�J]þ�z�U�2OB6�:��0�/K4��k2�� ����"Ƣo3a���6���J>������	�[�q~���ַV�����pT{�<ه�	�cG�ΐe�oY�F���_N����s�����8'�1����8�wI��u����RI��xx�p1\Fz}b}��G,�Rߩ�g�N��&t�z�z3c:��>��!,˄�C�#��\�����<�]�U6����7�Kjp�8�W�x�ӳ���`�X"%�]���
�k7K�ow a,E[�/�P��|I$�wˇ�5�4�������!��EՖ{�P,��D�����;e�o�!����r���Fj�Ku�T�=dB�1C�V/;��	�8Rq�ܻ��/0?@VV� �c���o4����]�B-� �Ի鵢��������ĩS���U����S鼤�@ bȒ���'n����Ѩo~-4?¸ɸ��ŀ��}z�U��� $C�ɱh�m ����9%�������gֻl�+��CMC�"�+J�]��b�>�rؤX��>��,\��9��������X�Y%�R��J�r/Zw�!� �>��+g��0a���]gq_�dө��!�u!^�j�Z����_�5y�Xxq�]���Dd����w��k���~1����;3�5̴)�`!�z��7��nH�X��P��x��"�c;�����ύjb�u�S��,���i	$]�O�c��PhOXk7�\<{WSS�8�~[�#Ye��/@n�X����Ă��8�/G�����K��haeeU��x�_D�r�W��;8���2Ռ��)��0�&7S�n�%������-"�b�o"�)	2�N�qaU�������ƒ--Q/TM@Ε����6{MP���4e�V={4|R�/@��V
'�����b��[�,��������e����w�;���Di	���I�I����2!/�ؾ�-^M��V�v=L�Nx���ܞ� �=>���e�W���w�e�juY��́:k2��I��DD_�J�	ش�g#}~9�FB��.6;U��'�X�x�_��ʙ|0�֥{�q�e�j��<��I��(Rb
��Y�ll�a*Bo���9�`�����w~��h�J�o����N�QB����'X)��p}�[�Lx�Z3��7xw�c�d�nSR�����y+�m��J����$���M������v�W.��F�`��s�	Q��~��/�!���cXP�q�pߌO#���R��\�1h�v�O��j���1�SH4ɚ���"��brW�+��|��֮YIlW��_HAɗ��Tެ�yb�@�@>|� q܅Q oFeu�_���ǱA�Eqp�Ц�/�S�g/H�U��Ͽ����ɠ��_T�Y|�_�٢�q1�y%���T��^U��R��'/�G��r���%=(��$����#�#�I�z���x��x}wB��|��_�9�R�cNe�Z,�GuԤ�˽��ʉ�&k+2۷q�by;�@����j�{��]~�L
lЬpR�<�w�X85[TEMiz�������ĴP�Ʈ")H3�5_�s߾��k�{�5K���Ѹ{�L�-3�ڡd����/t%���1:8���|�f@G�q���$((r��k�Dq��ht�ǈH�N�!d}q%=�س&a�-���2�%�-���y4%�+#���Y����C�A�G5m�3GH�,K\���I7�����9e����G�_M.�7Zh�^��"~���a��w�P���7)��n�f9�����9&���uKL_ -9�u~�/��V`XpO�\�B�z�]3�&���F��Ut���A��Wk _>r/'B�����{̣��sAY�~����;R0�dF�,W]P��{��{r��c�!�
��ylSgأ"R�F�ʖ�{�M�r-Y/�Y҂|-�?�7R#�8��;`񿆲�h����}��"����17���)V��P����DŪx-� ��nVKEz��4:4Q����	��r�3��kUjPca��d]O�_1�,�N��V�/�����Qͽ�c�aLv9�����G3�l�ȴ���n�����xzL"�sV/�d����zT��I�GL���%y�
)K.����f�<�M|r9?w�8� %�JG��!lK��ݪzM�̻�����4�̯��:���'-L�1O��tȉ����M�g.'�ڝ�(�b}b�G�A�G\�9�:|B*�����G�{_�s/@�3�B\qR�ɶs� �~_�P(I}�C���ȓ����nc��)B��X�oOj���v�e���͠�XI/J7�ދ����#��|���*�2��!��[<�'�h!�w
�؂L�#�ܑ���/Q哗n��	j����(�tE��%#�D갚�r��*IO���/%6G̏9�6G3�a�v�y�˝,}/u�}�⸞~y�ڳ���57���)@� �D�I;�W �Y�W	Îo�ʹ'�1��&ı.h7��c�%n���P5�6�.���5}:�n<���T������:��#t�>�d~�f�
����Ӿ�;�fy|���b� L P�]�r���[���� ֳ�}����v���$p�g����1����;������s+��|Eq��ͯb'2�s�L���}=_H`���Q���7��'#`���\�����ŋ�w	"��$���y�ߴ:����z�@�-�X�ϼz?���� ދ��}@���� M9�`�ȟ�Ơ;�VI�f@���'��[��$��C�}�-ILQk�
>:��և�A{ߞTy[	�y�ۛ����p�O��	@���n�vIf+%��I>���AwwO���-�[�\��z��P��	>US®uE��M�$�T���r��o� |�3�1=nR��::b�B�>Zei6K�.UK[�L �z��ymier������Q&V�,�����fN]�����z��cGl��t�wǓ�ֻ��S�ِ�'@�(��G���;��ӗl�J�	�{��C��7J��Mce�۝�\��?f.2��S�s /�#A��B��O���Z�#]��_@�G,!��WE�����t��f,D�<�$Pۃ��9+o-J��ޏ�%�Ŝ��E�p��F,_Tm����)�g�fh+Ή�0f�D^Kv��
$���ZO��0�{Q[�g�lh�v�-X�s��r�ڲZ˂�X��nn����'�dW�	BD`�T/�%||Ė�!r�5��djp��v=>���fFͼ)��8Z�,}�#��D��b��7{ 	N1fc��5�O��Me\Ww[���'π�ڬvDBi�X8�����1h���V��E���\���<[�(�~���*�ʾ�6�veQ0��,�淥.S�\�U����~�k�Sd�B�> ��s��)�^)H?�^ϭ���B'�ֳ�?cn��/��h�'���,fS�<��Qꭣ�WRB�Qz[��ÿK`OU����,���G�F>>}����1S�����d9�a0t��d�5�
�m�l¯�#��f�Y�'Be��Y�~0���N:��mLtjŠ�^��H}�����I�뺪��t� S�,�����`DP�7�]9r���l֭ $׫����7!��,7]@�H���h��� ��_�� ��g��x���䞆�~�ċ� ί�Ʈf���'�۔V��Rc���p-�q���Uę��V�~�O����t�3,� �[c$��e"����dY�҆܇xɨ���	`i�(�}bӳx<��k�W]�uI�۞1R��d�,,���v`�L��c�`���Ez�ʷ1�(0	>�X}��*/�G�T�_}$=
b¾��^����i҆��+��� ����/z��3ʢ���к���\(��]g�O�z^d^᷅k���=��nT!=�w���d����O��J�!i��2�}����+Q=�W�N��z՟x;��
����Y�F�k�2�Z���IyA2~�H����Ӆ�*E�@���S��Z�&�1(&�eۺ��s��.��J�\�ס�ÀxDk�"��v�2e�8��W!_oy�$�d��Z�h�h~��"շ���6������İ)�d��R�c{�=�Xm!�b��e?����<uT�@���|}�cｄ#Aѭ��	��$��ucT�w�ͳJ?#qs������|�"��[���-�e�#)�����aΈ�L��%���u�"*7�R��7ژpڷ�����~���/+M��X�?6(��@�����S�l5v��E^ˍ�]?k�8#����@n׉�ܟc|��,�̇���:��6��۠��(�~��>��.�$��ah�wJ$�wݺ�"#�qo�!1�97!&�HGS~���gJ��8�W\��:��H���Qz` �m�M��B*�A�(�"�E?I��%����<�Vo���߾�B��ЉD�� n�]���B���aE�YvC��E� ����E�0&����i԰�i�R'��eN�^�Sg~�W/a���{u �������Z�哸�jL˪PW_��j@��;�I�i�F�M�uI�JA�<'y�w1�|���cx��.�(��ZG�`���π��w��{9�w����)�L굦M8znu�Z�XK�c6&%�������\D���?M��י�(�c#UL��4tm��ޡ�T�\~�7����}'�8��a����}8�L Җ�]�%b_д���h�d��鸫k�9�5d�>pv�AXBM]�%�����@2�	EB�`��P�PQ�&=���{څ"��A9q���jV��M2�����\t�X~��p���c���4J�� �(��Wn]ݍ}��pӿc�O�+��;`�V�bSfc3��-����PM���ʳ-@Ah�ӥ�����uO��,Zȫ�V�&��'O�krM�ӢE����X¥um���
%JC!�	ړ�Q��������<<s�*�����6Q�r��K���A1\����g�HY1��uo_yH��t7�wFq"゚��������.�s���W���ppΰ<�*v3����vss	�^���:�a}Ε@�$U�^pe3\���̏���<*�b�����q���s^��F/Q����u�GxĪ����H3\����%�2�5�oĚN���}m�j3���]C�GֆG4����%�F�N����[%ߘ�/r�=%z�)���b�5agy���_ �P=����1[���S��l@k#�>��X����+�F[x��
O\�X��J�>R�44�+�u��Yc��o��G$;�<���7��ȴ��q���]�n~S< ZaxZ�h�Vr䐪H��f�hH���x�$J��ǩ[���LJ���WK��
dܷ��?&+�mPɖ�{����r4w�7\n�+Z0�4w���eʷ��-.E�K�=��{,?r+*�@>h�<�G1��!H?D���Ϝ�h��yq�K�{��~T�9Mę:��T�e�tW#cƱE�~��t����\3�Ԋ�a=���X��G��ͻ��-�e�0S�~n� �NZ~���4A����"��I�O�������Wx[u���#��:�U�]�xgI"X����m�����$��>�I����b�ߕ���a ��<���Ѥ0�Jn.TT��u���	>ZS=�/w���Zy�(�-L�R҄���d|6����Q8 �}��N7��`���-�<�A[�=>z�߫!5�[���ۊ�x4�ɾ�L��-p���
�B0�xK��ݘ��P�_��"t��c���^���bW�
�/���W)��s������e�9�����[�q6ʍ�@�N�
�?�9|4%��D��4��Y\ԎkR.9[�$3�9��Ĭ�":Nh�@p��л�m�"���-�����=�|VnM}v���oR#a�Q�L�G���ه:-N�$�vth�6v��S�V�!H�M����w%$c�嚨0IgO*tC�"qh�r������?.�#6�m�Ύ�ݴ��Z��"a���<s���V8�]t��
�.w_N�?���Ϻ��x��p�������`"J�!��<ޗ��d�.@S��X��y�qG�_v��[���cC��`��f�����͎�\xW�6S"�1��W�����)��"�7���<R�	o?����b��8ޏ<��{����h�QI���xm ��6�C?ep�|�jQTjf��!��x�dSd�{����QK+����GJ�-C��(�<�,N����B*i{�&�,��|�4�*�
7�?��C�����ޭ��c ]$� �ˁ�Ϲ��G	�u�|g3�<d��R�������q쩁�4�1�ݾ�����|�^h��@�'%���w�r�q�ÿ],b:B�~�&�TA�VuZ+a��9�`
d�z6[���5]m0$	�CV�����..%�{�#K���h���4�V�����#t��C�}�ś�(��?|���e�K&Bd#�|�Q��GO���4���ހ�~%J����$ҋ�B�8�[��I"�Q�pP9z���k#n;;��?EW׀��ꀀ���֟��I��,I������`I	�O�$A[�_Ώ/�T�������r|���0ztU~���L�H�CU�l?� �s�7YR�Ņ5���cM\�t2r6�!���"dTT���Qdpw�qB��m�S9�ˆ=h���gf��-.�6��V5�r���s9�,0������9��	*�a��`V��І�����������>lzn_�󻜣��p�����zyǕ����l�v1�5$�uڮE�X>; [z�J�5Xz\�K�l};1p�E�K�4_8��e�����Zt^+�U�/�T4�M�$%�jH�M�56'׉V϶S�SZ~K��nN$�M���`��2`�B5��|"��qB&����� �S���4�� 9�X_nn���5B����\G��V�P���F�oey8�'���E*�eg�U���;�:9a6fa̺�5*���R��jg�τ�_!�΃����CGd�=r�jG�J�tRR۳x��3v��7������Uݷ}}:���u9�G*�lv����z���8z0}f���qf�R�5�'U�J(�:�80u��=�n�i�|@���ia8Q5~�.q�7�l��D
�-ʦ��>)���+��!�#��0�V��ܿ;�2c�È��dg�j9�'N^>�N�C�D��|�襉V/�yB!����(�p����g.���#+# ��fй� ��\u�)/�i�i�L{����[�TY�%.ȇ��aW��J;5�0�)K*}8�3�;��}Q�R�0�,?΋��� ������� S�^Kݘ�*�ܥ|���s�cI=��<��1�@7��:�o�~��հd �uK�o^�[�����8�5s�	����t?f��i�ؾZF[�H�`!������EM��L�%�G��:̚D��MS`�D[�,/��?ُ9n�����5��4Ld�庖t�T7TĈ���5`���@_N��rد9o��(����BǗVa-ߣ�0K�ǩ<�a-u�:���x�\e��B�sI޴��=S�����Mu�ٵ�&���O~��ܒQ���Ζ�4��i-�s+x޷~�:�w�0���=�i"�2�!Ǯ��mU�r�1�GN���2��O�_���Ftc��O��G�x_4��r��p����>�X��m�!��[ˏ���X�Aӥ���i9�r�n?Gi�#�;}7��=��5��.��;���B����N���(���S�a>��� o]M-c�6e���~]�.A����Y����:��H*��^��^E�1w��дy.���Q�;Z�>3�|�K�`�G����kv������Gw>�9�cLv��[ո����h���߽�2���ٽ��e&�pǅ�I�M�`S��8�ױu�������}=�d� �pv!���4�F1~vY�RM�� ����(�6�2�yek�0�Z��A,-͔l�@j��K�(�ˤ���rSv��)'A�zT�c�,���j�7=,M ;�zǩ�-;���Nص=	����֚d	�Ȃ��$?��>���Ɂ�y�����2�(�j��4}B&[��������T�:�U�����ɮ�+�4?��ʴ�G��Bk��)EIƧa��s�0�x8�/�۾ :V����C�8������{��::y���:�&��1[i�����Q0vf�kiK��6F!\M�����m���{�V��y8:9�ͯ�z�XF8��\?�M��+�V��#���S?;�0�vQ�0�/�֢�[ϧ���烯��1��C�*-#_�1#$KS����d7�*|����ڥ����ٍ���`A����8aC*�Q˯�����ơ@4�/�[���5�l��-�.ɯ���}�7��H���ݗR��W�<�	bWR�:��X1s��P��<��wa)W$�B���Ɣ][��5e��y��Б(��ӓWe�t^3il2����I�w^�U��U�̸�M��H�k�~�2�a�z��?���[gF�Q���F�K�aSxPJ���s9�W����܍���'-Z�	#5��9QG���+5�E�L�>$�	t��v���Tq�|�R��z��Hj��ۊ6_a��.�����!j^<W����0~`���f�A>���\n�b)�mN����AV��5k��M�Q��O(���MLUZ[�O�n��Xl�X��y��y�R]�����聦c>�)����H}�1G�)��T�p�=;�����L$/g��R�gjzZ±�ب�ܵ}
X�!���XS�oKEa8��YV��r~o�ѻ�E:¶V�j���n���8~`��=#����+��?UK��*wj}<Ճ�+���⏅
�d�2Y����K��1)�Gi	�`��I��b��
O-����D3=\�=������O��	|d�'�VǨ�%;�lu����0La!Z"����<����_�w�T��Pߧ�����D�hQ;���0䆮��y&n�YP�UNL�Ե+�@�X��{�����q��XNQ�k��h7E����壣�(�o}t��d�$<�\~���R*,w/x����f-�:��%ʩ(|�F�t0��s2��d�B��Hp��Wr'�FQ�AH��o�<<�����[�/��^�����\RLU�#�z�`��jD&�v���A���G�� U7�n�Y�L���2,�?r���s2v�.lc�Y��;#G?�6R/�W������Ph�w���PZY�v���	�`�{x� r�L%F\%�(�p��d�|;b<f�|����0n�.��+�����a^HFu׈H�m���~��0I�÷oyߗ�}SC����r��C�P�H.N�FK+?�Z�;�;oGR3c��N���B�f���T��R�;���$Dh1q��(ю$[�#"�g�80_.�����޺M{��9��w��>��k�+����}Fkc7����!ʝ��;�i��e�*T�;�b�V�@?E@*���36�2JB�h]Z��:$|F�
�h<��t��
E����᷸�k�1'_Nq��B��>\�@	Zlw!�!�lι�yc	�!�^b9�@XZ/d�$����:�{-p]S&�F�
�O�C�F�X-b��#B��p�|k-� �����<�Q&<�:�er��¶6���e�������E�n��?�!����D�:YO65���A&$
'"����2d�
K�e�,���v PcV��Yl�@۳@H�����Ϗ��n��n^�|���ѮV��c䆃���0���N���h oL�Z,&(��]jkhQ=�1�R?b�4E駿o"p�� Ռl0�m�Jye��d(���T������Ej�B���S�����J�sF��_2 �?��ՅR�>���%�Q�^؏��󭡝�
n~��3r~g,�߂�[����܋�h��,�:@M?b���=S������׃�{Q�μ��s<P:��M�WZ�u�H9 Cy56���Ǹ�d� 5#1/�<0�S9��'���F-��Lg?��VCˈ�+�*�*������LhWd��K�QN�%����Yj���;��!R�oU�����}st��C��&,j&�����я[U�|�ٱ	uU)�&S��)�!�77�J��(����Vd�X�E��%3��'����ꃃb!��״d�|�;\���F�/@�5��<��>=:l��ض�J�vr1�h�Bs��CW�[�x��L�_���З*��B�b
�D��Ϧ�_�7���UE�� ���ku�D�'Ow��P!L���e<��-���-��yЯ��	���U���R�z޼���W㒿�2y���[Σ�4���#��Ԉ�Z����*�a�×��<3�7��Ȃ�E��JX�.��c���ei�֌H�eG��=������j���,z�s���:B8Ǹ��ˬ�/�mY0-��b�f����
�qΡ؂I�[��htř��(q�$mE�S:�_O�}s:��Y\,6H�{����W�]&������3�6�>�ܕ�/C�.���6����Vä���G����.,t߫:������+g��x�`x�A�j�OPSS2P��ٕ���bs�-M��Qy��b�OS3�`kxs�8)34XJ���0�覒���1����,����$�JF[�B�v��� �����c~Œ��&��ݰ9*  ��"d��:�g?3~#��`)ee�Z��A����f�����5�E��`���r{/eXd��u�!��ȏ>��2h���U�QsH�L��]ZYFƖ���'�E�Ꭺo��S(hg8Ni���5T���pY1�b'�U1�~��{�-�����V�Rg-R��|�y���E, ��!��W	�;�Sc��P�2#%�b�7�ϓA�9c������B�LS쮅�g.����PV�������9���VF��p"*r9-x�o�`F�D@[B��Z��6��`��'RU�I�Xr�������y>.�����hĤE)[^�v�iR��F���9>;����R�[�P�)ez��߱U$�V�f���!�����xOs��ok��F$�
~�\|��k6���,%��1� A�v�x�5������ �|.U�J�j�Y�h*�K�%�Gw�:���-}��=+����Z����=S�ϛ-OW�m�/�`Q��Ad��L��٘�CU�m��!X�����-=�YM+�E�v͝����%Rҿ�H�E�{u��lt���||l�1��~���N����2,�t�V�ۺK�@~��NyZ�$B�1`^��C�����8���R�X<�k�sF�1�%��ג�5�����#��M�R� �H��|ђI����s��)� ����҆iӓ͔`�7�7N���2�7�*,Ǎ����,t�T�	Q�*�|T�_b�4h���(�J�]�+�q(}LQ�ݝ�u��R����/����W�JY�uS�mݽ�]�k^��8GZH��d�-j e�'|x�8a�~�[�xەWV�t����T��}v�������ˁ�<��r�A��{���n��Q���<<x�w���W7{��6s���ܿ<�m~�j�jxX�77��ШH��T1�|�)�чl'q���k�aA;ʖ�¿�� E'�s�%�>*�IK@�ݭ�|��@�����zo��]�]�^��O{��9U����t[(�q�E�������8ÿ�n%a0/�e#9�,����Wj���FP)��F������2���Y�0m�xֶ�v��+��2���}����� �$���[�%�l�A���#�3X������ދ�v*i�o��L/ۤ��;̹?��M��L��1�}��z=B�6��N��ND� �*7������O���?�آהGP5g���޴�q��(���
��M���_���;�~�����
��H�Ë	��	uniiq�J=Ea�t�9���{�pi�{{��Gi���O�u���s�:+mI��=�=tj�toK�_�\�p�O��������寗�_ܸ��<�I������İ�KX�ǶM�G��������|�M�^clUZ�����.��OG�X�9�DN�tcF��������$��D"+y�k���k�p0���'�J�>j,|z� 2��X���ӿD�5��v<8���z�Nٸᡊ��q���_ ��úR��)�E� }౛y�I��\�d� ,GۥٸWWơ
N�|^�����,f5����n��UU���xo���� ��D�z�>5v�����W]�D�Ķݪ�7N7hD����{���E	��{Xc�[,w�wL������t��j�r��'Ϣ^k)��^�|��Dv�9bac��o�u%�ozjj2�}k��6s�����^��G(
?���:p�����3Q-"8�5�<_"�/_~����^�e�W�����z���E��v�	trx���oL��'�jKwl4��rv�S�n�K]zx�d�V�zi������;0��i�>����;1�.tN�5�;��mZ}|g����:�(޸��}t����<H��j��8y�����Gެ��ǡ��.�ޖ�5g����i,����ҶC��X=E�+ό9Ǧ��TGbB#V��pEo؜�����}�3z�����K�ˡ�{Z|�W���e����O��pXH�x#د�ui!xNߐ��.��	s�]\\rR�gyAF�x��W���Qa�z�UU��i@��U_σ��auu,_��=����ߺy�y��L�i�����j�54k��ʹ����J�a7�t-�����+�Ϋ}I��5��E{����}֖e����wCCC�c�?U�Q�7^z�[���?ݍ�(@π�*��*�� ��n�<ʼ���b��X��i]�5�����16h���@3����T�q�D�����?9i֬��+�����O�Z��SB����p���i�@�>���wO���
!�f�W<����z0G��
,\#A��5��E����<cƌ�
�u]?� y�?���e˖́����b�(�&�+�dKE�Z�D�jQ���e��{Ҫ%�����Rz��m�q��!��U�A|Jg�=��yK���}�۶�;���n�Y�~֎����p@+���Ҽ�~������@��6�of��.�Z�K��.}�&��C�	0Fh%]��5����.��q��]��_��>������g>�`:�Y��%���57�$�%#�^p�ډ��$��^ (�B?��ߥfk�5��G�����-	�x=�&���D�>�̄�{?p�����~C���F��2id��/X� ��%U���=�FlRI�b��+d��8	�r}�.� ���:���P8\"�6|�Ka���w�C����c���ח^��?yJ��a0���!��l)���x���"�/������[/ �ړ" .?���=$OG ����*��S!���������U�|������o�ǶD<6nI��؂�g�4R��ΫY���{׵��5e��-�g1X�Rq�A�L:ͱ�D�u��k�v�׿~������߼pᓿٶu;Kx��7u��M�����!Oy����2 �'�&5��j^�F.<k�E`�H͚�:�d&�Ϛ5b]hJ2�Й�޿����k�7�x���&���ѻ��S����@ꝫ�4��������bs\ν���`�3ywG'�6��.#�R�@�F�����tD1S<���z��g��eRL��<6�N����J?�Ȓ��+T������^�6"߽&���1IZ�X������c��R^���Z�k��(�_���;��ݝ�d<ʇ �_C����bf�t���H����,o�
��jV�̻���W���Z��+��?�����C�)�k^__O����:��*��O~��%�֭=�g��س�>4i��~��\���ri%�R�W��kIɹ�oRXy����*!Pb��Z��+<1�V~u�5��(i'�w��_/(��W�������z�]<c�� ���0�}��4k/X{��*^3�V{R:�7��V�1�ɽ��x=�Q�1Κud����/P,���Q�ݥ�}��?��]����dq�7�"�}��ĝ���L��I�q�f�)�m�$w}f^�&�c�rg%?/kN#Ԕ��
��kh�H�9g�y����N���g���?��8����� �#�H�� �`-�T.6/����Y���2�9�����ݰ'�fs/�eW�56$�fg:�tޜc�Mh��_<���������'"�'� "���+�����kzW��w�J�%7��b�D�������Y��46u2!�|��ٿYZ�U�/�G`F���C���������ݝ��Pi���C�P	� Cb���f!l�T+d?�y�|Y��J.}���{�M��B�4)��`���� ֽ=]�%�5Hc� j�"x�k�������_����x������+�Lo ��=���J��Ր��WI� .��kiyy���n��� �\��_-cC""�TI��a�;w�����'y����\��F{�⅂�:�u	u(a�����q/��1�v�!�ϋ�bKB�/���tJ&ֈ�a��N=���'�&������ŋ~��{�5�@����q�4ǻO��OD\Eړ��d�\\��%�߫yz	��{7|�\��<�&���A�  ka���4O�13O�>s�C���i�{���������bSk�z�U�9XHI��o���� �]>�Id)t�BJ�.�/mv27�	`�^�>�Y}��c�㗖U���K>0�޷��w��mU�͍�݂��l�@�̘�����5��w�k���&�`-7�4��X
�~��=����3�]�5�#���X;Ƌ����3�>>a��)M�u���e��i�-.O����%e�TQY�||�f�S����Qj�r�K�ë�H�Q��W��o�s�`����S�
��.?��`�?���v�����[����h4Fm�Y�G � j�@[��4kI7)x��],��ڸWI�ſ"�mOߓ��k����9eW�y�����{�7�����:x�UWdW�^����CA�|��G�BX�"伽�R���/{���bC�,r�e�̿��A��3��|�Y����l�}������������
�y�}A�c��p�VQq	� E	�^3A�>�^��[��՞���I�X�5��f�0�7t���|�<�(�4��O����?�q7�����?�{�}WEqB��g��?f�ftN߃��{ZH/�Ia$YJki^K��r�H	� +4 k��rW�A���ҋ/�TYY�{��o~��+ދ O��/Fy� �TR�	�'�ƖV2�w,ҏ)7m1@I��w�k$@��{�Lqj���`r�f�|n�����Ea�>���㊋���՛�;�m	nٲ��\��+TU]Cu�Y	A�@`�1K���V'�Pfl��|.�X���d��{������Nd��f���J~�2eJ��'�.��{۶�����7a/��v�AE�0C��A���~^���Ei��ϼ�����KKP.k����H���q���0�^�sQCk<|�y���?��n�]�/~���;wng���.�ѣG��1���Z��`�B{��w�z1HοX�z1�����`��3�YW�-|�| z��NqG��o�^�l�۳P=Ƞl���JJ36�m��?¯+�0R��o��"�tvr�߽�X
����JГ&$�:�L3��䈊��Is��O����Fy��7��멇z����.�?�Me�`�رni�:z�v^�׻I?LC�j#ޅ���bi�~F��/� X�����lЮ1��H�w��8��9�����ܔ^�fU�96�!������K���>M���er)��y7���z��!��x���1��>��a%!O�T�2m�r|���/�����+l۲ɇX
> ְ"���5@,�a ����/���Q{ڠ���a��H�-�¼�ثqz��`��b�����FV�O��b]�<�H��?�������w�۶mì[�|�.���kиV!|�����@�лV^ͺXa����a������� i�aA�ď��ܟ>d��|,\��կ|����޽ڸu��뮿�����n�B�&L�@u����������W��ʈw�R1��y}Oں��"��Ь++���O<Y�/i��y��w	��������>>`��7���	R@��Ŗ����nD���^0*�h��h,i�b,�?�z�Ec"e������9R:~������k��_����������&3�W����MņX˪(	�LY㩌��e /p˿{5pI�]/X˿�M��f��L*]���}~���;n�ԧ>��yq7]������N��r�1J�KK�i̸�TZ"|�����R+�j��s����s���W��n�~z�n�ڌ�Ӕv]>��/T��;��c0��?�t�)���N���~���~b������Ω~p�#���P?� �CA?k�ȇ���vw��c������]X�B�f^0��8 �������ڔ�r�^�)��;n=��s�����<�{߽�Ŏ�NJ�2�po�k)�<�փ��R����
H����k����'W�x���xO`�
@h�xz�[��c��eмm۬�;��Y�r�g���#'�R��� k<�A�2[L�%��mN���'���,� ix���f�{X^/�7[c��U�5�5z�X��w��8z��ƽ���>�׬���o��ll�C�1N�UK^�e +���rrR�(/����M�]\�`���r,x>\ �h���R��S�c��C���wN�B�i��j��z`�{�<�E	����R�7��Ӹq�(=!�[���rǚ�[�&�.ǽ�j^&�Z�\p�Q��LC┶Z�Fy��͌<oh�,�0]xᅫ/���˂AMU-y���������D��(���V��C>*))��&PE9�����'��˱���fލ)5g��oV9�=i$��\�m�{`���u=,n��=Y���n�v��P��GqD(TS������yB�De-\>āP��..4�H#��w|�aU�T�L��yz�!�Zj�r�{랾�`���Ƽ�ʘ<e"4e���:�|^_�f�n@o6�B	@�K���/�xy�k���x���4L�^�dly����& k��! ��r�ht]*k>�/��d�v�����Bc>r ��	��X�tW����X!�����y�1�żZ<�U(ݢ6�\wA�9N��ĉ���u�'�8����>�`���__o�����n^������$�������6R�Gj�X(Hw	����${(_�j�R{��	�tvtS,!�Z�j��!�O���̙éa��?�R���҂ؔJ�l���p=#�`����1ɼ����)7{���y&E~P��. O�=oJ�����c�^��� �A{R���&���ѱ��Q��/������
�l�
���0f�?L�&M��QUTR���j����	�%��	��7�1��@5k���f*�f��ȩ�(�jQ��F�V@lƌL�P(�}��[��{���t�	16M�豼�K����r�$�~pw�nIW�w.�ږ\W�5�'�Dv�������`!�_�cm���'OfW	�7P�i�&Qc� ��pi�:�w$XKͺX(ɱ���S��Y<oA�ݫ�w�t�J��n6�?�� ���p�4��c7�U������FnJ�} lµ�\>XS\��1���ܯ֢������{�w����	�� �4����'L�D?��9{��{�}ޯY��/����ՁP�эj7ߔ�"��c_#.�D����J�/fp��4�=nh�V�1�u2�qs>8��� �(b�(���ӧsY+�:57��N�C1�(�w��1?~<|���:��`�Y�B)�VEe�r.�$M���k��J���`-�o�8k�2;s� ��A�!�S�N�R\>TKWiͪ�,��I�%�֠���n�a��� ��|��ܓvU�Ľ � ��@Os�=*�i����<����� �UWW"ӧ���͛7
WJ:�y�(`B�0��54���cGS$(5k��'ׯd��7 '����޹�mcKZa��A�����`����"��I�&�ĉ�34P����Z��$_B�A��`�{y�A����?�f)� ��=	-/���R�Z��A;�x�Z�cAG�� =�H���;2g���z! žFj.��G�1��	��{Nα�m����7��n,�%��R`��G�}Xc�������fϙ����xo��kַ~������HJ�pZ�XMр�ڐ�BS���.�	)5��e�b�ޓV�%(|���Ԭ� 
�5�U���EC3LI6DR����f͚E~�2��e�&jj���!�%R����~Ѡ��0X�I��2�w�	�	���]jP��l<8������a�h��;����.h��A�A�eǦ޲a=�1n}�8�}��i���4~t���h�"����7�LÏ��ns��U�߱]%@St�L*˚�,��� ��JK�3�Y[;�����X���2_�
Y> }S`!�;X��|J���Q���?w������b�.�T��^�ڜ^r����_F__��i1��k����ڲ4�[y���c���(f�w �M\�y�>ҏ�Bϓ�Q̫ȥ5-����usM��ו"�[�I�| ֲ�ɻ�����[󪪮`%B6F�-[��h"�",%c�1�ko/YU�����s���!���נ"��S�O�H�q����<*(8���/�h�<'��(�,sM�w�{oU��w��;g�����}�:u�����Z{�Wl��
��v�����糞(������S��c�C�u���t��/��p�9O�O������#���{�ّ{���Rc��-��C �0�h�k��&�5�����!Y۸8&�Z�8�0&�5��aO�=�x���(�j��(�Y��EK�H��U�/�7�Ѓ�w�O��N-6L@X�!f�@�����_jS��.�q���a��^U����[xm�/��3mc���01N����D
Q�����l�XcX���+�1��ۋ��u���[m�����X��Ȑ��F`�­��J^e&�35��Q��6PLN��n~6�UA��eZ�"W˖-M;��|���8�f �w�=6N�S
�ꂾ��^��9�0�m�u�K	ؚk��� *mU�#��F�뢧�x��:.�X�W�5�w������w�)6Q� Zȯ-�R �����Nȭ������[���_�u��� %1k� �w�F�Eޜ����;Z,�A���-��!�F�P�0��f��-|B_yq���s�rWf�q(A�H�y��u4U9�p!�u�Һ�OY;����~����U�.�������o�}{��,\�Ԋ��m���Q<��LuJ1:ۑ�Д��Xa1��Wl�L�YG����)��!�ۅY���˗�����S�k�t���ի�rFC�!5�|��A[����Q
�7L�%4�,ҩ �8E���n�$��Ĭ��g�r����������}|�C��j3D/|ы����Y�P�����8n�>�F��Ҳe[���픖l b*��+��s����k��uK�៚�F?���=U�W��я���ᡡ�ˮ����QS�i��mZ(��56`�(��5`�V̚<�~}�ª�����F��bW!� F�O� ��`�g*K�=��t�m��Zs���d3Ef]��(Pv�-��
�2�$s�.���VvË��������Rc��G��x�[m��N��Ҽ��n��������}��˗Xk��yg��آ��'Y���Q���^s)����;Sk�ߖ[n�^�W���Ozu|7���?��<v�M7-_�l�u���Z��e آ���9`x�\P4�j�R�H�Z516Y�r�z��\|�X$�eB�m�]��M�˅�S����w��b��m���{���k\,�AXp��P\&y�U��G�����:}/���\��1���^���=�%��(/����H��sO�ѕ���`M��i�����XZ��i�m���^J���-�T5��8�꟮�@I����Y�[-�o�_�Zr%�7�Ԩ����w������:�^V��c��2[r~�6[o��[���^\#�(ǴܥZ��~
�>G��uRjU�k��qW*c*��ƃyE=f�;8��|��'���+f��h��������E@Ӽ��aR�sH?��In��+>`+�٫�	�A���b�ɩBUoZ_���I�-��/�~����t)���²�r���q�5J	��6�ai���Ԥ��Pu��`8_��W\u�	�l�A!��X`<�C���+Wl��Vf��soa�,�(�o��/�7��UFe`�cޅ%eB����T敏�R0���իs8C� y�/�Cָɮ���=�5G�sE5��eK=k`��~*�R�y�{v0*�v7��R�"`E�~��T�:*��	�:�+*��!�7�E/�#���L�|��9���T8���30?�I`]5�1Fٙ=    IDAT%����Da����#d�]r&�F�}�}�P�0�;��wi}��jq���+�5c@y�S���y�qN���7���/���k�A 븰$�
Xì�>sX��h��f��o���A�c�Ŭ���e�c�U��:X�o�����	��N��sO ��5f\�!̑�a����',���IF��D2�E�#�8��d���ᱡ�Ĭy���W�b�{O=뼝���W,0��o�����]oAv�X��GǕ/M	z��E-����Fi ���%��*2kwy�ڵ,ܰ^�&a~�=�����4���}�����|Xo�������ד������iw{�GE��E�����vn���F�����ll���+�s�}0N�K�5}��`����[B�%�����~��O 5�, W�Z^D낡��C�ϢE	��*��Z1+W>a`��{\�bχ�SN�}���L���bV�EּF9�="�Ǳ�w4/<B b���yd��{0�k+�NO��6鯕\m�	�ُ�ų,�U�PH?��<G ������	d���D��Z�Xkƞy$�-�ZtX��kì\�}�ma�/y]bתHW��a�,����2Y0#��d¬y����g��}�W��`�wm�'��ۮ��]F��R�5g,ʳ-\��)��q��.���?�@�A��ߓ�ր�}��B]k;��F�'��� &f]����nc�˖�"#J���a�`�w ������k���c�W�k�u�|�%�_������j���Ra��/͋�^�E��I�\m��.e(TA �=�Q6E����I��?����e�<�-Ϋ���Lܟ�&f�mɪ�!�C�k���ڳJ��RW���9g��:V&W��SI�[�߀ޡ�Z�Zc%p�'L����;��BEړ%t#���B��$���1�V���,9��|�������LjC�d g��T"X�W��� =�Z����*�K`	��?z�Q'��?�8���x���'����%��۪�.�-y�l���Y��C������P��XtN�S�ՠ֔W��n�~��1�n�l��<�J?�yU6����v�D�f��Frֈ�OY!�A6֜6���5����a7��B^,,N~	�/T_¸)f"#�qֵS�����L`-f��*�_*��s=�ʤI����ȃе�XVd�Q�<����W����_�o�U��4�=�1X��z�wN�B������C���6e4akk�- ��~
YV�d�^P*��q��{�Y+�z�0߁%�E���b�Ĭր}�;�u饳q�\�LE}�z\%���w�}�Z�3:��#���_kڦ�+�/:6�A�`�g�0��.2k����<q͗�RϢ����7���Ա����P�:�v�.\�lٲ2G�Y�u�GvHkժU�w�G�k"�Y��k�K��I���a�E��F�Im�����3��&�B9�`-f�<pv7U�Z1k� ݮU�>3��5���=�_E�r�U��r�8��* ��gS`�g,��Y�k'Wp�=v+�ϣ&��\]Ƈk��d�"[���5`#�Z��Q��MT_�1s��Z��u�/�:��.���51k)��v{�HU2}X�cRDr,ս"I��F�12�v��[ -0��+kA`��zUfx&m�0���l�L��|��M"�0�P떆)�c)��v�(�<#��T�:�WC���o��Ÿ djG����/}�7OOZ��K%d#�f�Ŭ�y^�5/q�4�؏�d��(ge|����~��t���3�]��m-Z��Y`t�b��џ9��{lKj�8#�͹��QZR� ĭ�D	�P���#XK�u֠�}��81"~"��?��^����k�C�B��{�Ŭ���4u�z�E�F�Ԋ��"4����*��d�	�l3
�����R%��;�z�-��wA��G��.���0�[�x��5�{�Ff-�ќD!��{�y�ϑM
T$�DzOM�Y� �?�k�\RU`=4��煒��E���U)�xL<�s�=f�[c���T
���}������	X{�"[�=�u�������,����>2N��O�V�:�WF����Xr4�s͹�:�(q\�OS�̗h4�x�H��W󪃼��������3`-/B`����E2,��#�}��(`֜Fv-Cj<0�dj����/~�-~޼y��/���[m�����)�z���p�wS;���
r+�U��2Z	�
�&��?M��A-�.A�`�qI0P1"�XV����O�Q��`Ml����3��Y��qM���E���Dxb��ڪ�b�±�����a��I�$U�G\��RD��n��`��TfC���v��B�wD����`�g�-��e#��+7��/	r0��~̔l"�	���r6Hd�2� �Zm�ل��f��Ck����,vdW�"�ǹ-�K�:e��(V����������9ݰ�|���.�X#���K?�8#X��b�F��Аo����C����U�r$�>D����S��y���~��ݣ����~F�@�k��j6����`D�BrA���#e�(ߒ��]�Y�%� �O��<��(�(��׿��]��n�;� `}֩�<p�m�mױ�ʫ�Eʚ��^Y+�%�z_, �[�x_t��-��@����p)&k�M��-��Y��X�gMU7���o�c�>�y֩i�{\���bּ��ob%�	&b̿S�n]u����5R}'~W �3Ŭa��ڣ�VL�kYL�e��!�|��c��3[��}6���$��:���Q
 C,0��4*j4�q^{�l��~��Y�!�Gd���^J �����r%y����� �nC� ���/��_dP�E��D6�k]�,�G�b��/\�V��W����P����b+Zŋ�q-sjY>yAd��Ua|[�(�T^��Fn��[s[����TIT4dq�y_z�iU�W��t(l���4�2L�m��0f����紋������K�M�^ݷ�j|��?/�E|�<k�X3f��~ɒt����{���?X�N9��G��-Y`���Gn	<s�5��
�%�R�,�Q�cLT��NDf�6*�(�F�M�� k&�&u�s&��6~8�l��g��b`I�C�	H�c{kksN����"6���1��|)N�(T� =fx�^�]��23��u���(�@8���~`�VN��W������`�a�X�	�"��S`1�eς���Ն��vk��g���QZ���} �Fɥ�U�ڍ`�Ѥv�%���Er"����2�8�bh����m��˳�{(;%4�\���i;���	#(��G�՜����Fc�<='�BuSL�UKw�0=U�5�bڎ�Ģ�HzCȇ1�0�k�]`��4w�Z@sh|��2Yk����0��`�{�5i����6��
�駟������ `���[u�=�,�<B^�M'!���򀵪x	��u1����=�޶��qFB��F���w���u����M���� ���&4�������lk�'p,ڙAE�b��O�49b�Qad���T�O� Vo`ݺ�������~���I`���\�Ƭ�S.� �V�U��s!�YuN�);b%gU��̗��d���b*`�l� ��W�����-����U��`,�F�TU�j�����H#hpm\��o�Zi����#Byb�\G�V�Y=��r=�~o���M�̩���VD�_�E��agl ����1S�!�F8�A��{2��5�(�YƋ�z��<a�J^���qW����<�DQ��1���X��ƣ5ic����l���v�)�|p�W���������9������۟7E�c+QQ��
G�)�^lZLC«	��O9F݈h� �3�uF�+t�u5�Xcq�B	R^l��~OAs�ey̚g�J��E�B�.�l��-X���F򬣲�$�j�B@��Z�&@T_�Քy���3}��f	ּ������ms�sa��^�Es�
@��y���o,��{S̮+}b���UfL=d#B��0� ������}�2R�~�/r�B,3*u�h�5�b�.ÞS���.H޸��Oc{u�!�Z��6{J��5�X�H(N�>�>`����Is���g�i��\���37�Q_鏈���&�\c���gH�2&�A��W QFX�����g�r�Z�?�3����`Er���œr�XL��=b�x �����׽�=G�=[��弳o��^�ar�@�l�:m���T Yc�St�xf���^B_�n��&���b1��O=e�Զ�Ȭ���'Jh��pN�<��5;��hy�Ko���ɲ���I]��Ĭ���C�Ln�Q�&�������n7��h} �&f��5��W�Z,��cb�D��@�ei�g-U�O,D}�\r�]d��+;�4n�Sa�Xz�/ �0�b�J��R�ά�+/Wd�j��U@��:G" �hȪ��6Ű�\[�u����.�<�o8�
S5Dq_�"XL���_��ǹP6H�`U���Z�8qdH�W1���9gʾ3U���ԕEhC�K_�a��� �}���#�T�H�T�dH7���g!o�pg֏��=�Y�|Ŭ!
������o{�;�~s:^_0��>��^����t�.]�r�`������D`R�V�Z�"
MTM�)gN���X��j�>���))������� [սQ�>.����;����"ލ˲�V�M��Y�l	x�Be�V!'R��RU�5葉HH�c"��qQq#+'�k�J�fM?d`�`SWHAg1�
�rm����R��)XW��������y��V� ����Ȑ�3Șy�A�8k��`�qq��_�W�^�l���s��h��}�Q�P/��G]i���Ņ4����{�% �����S~x�Վ{˩�J}�N����
��nU� S���aH101>�3#fpOmv���S!�7��g~	k����S}U(0z	�l�>Dr��%�=ʁ����}e�a����d>v�'.y�����3Xs���w���_�k�o0���1�|r�hxOA��"XW�Hu��z�O�'���J�{O�Z�,i�� ���g�Y�v��PJtp�v?J)�la��)�5��	Z%�:Z`1�Ƞ��x^|�`�����U�.�]B��:i���$�Y�������m1'��b�qN4�o��d4��N��D�c}�`��hc�K�P��X>N���� k3i�|b<���֒�~�r$�/
ȫ�2�������c�=�+�9�����Z2�WX�1&2k��N8��<"�);C��2�}��Dp�s������FU�X�`T���6m R;t�.�#`TؒTL��EE6H��G<�g���F�W_���},	�W��u�Y��'{���Aa�����e�{����o]r�7���=W>��W]-��'Z��0H�Yk�#X+FOሓ�O��1Y�2��kŬ	��J�jG�v0��k�#f�`�y�E!'� �]a���<��L@�y���R�W�-� ��ޞ�X�*`;�y�:������S��p��%ϐx��,�X�2k�MǼYDLA�:������gd(�[dq��{�< ��on�F�ga������+�R6�����u�ъ5i�4V���4j{��ת�����^�ǵE�`�s!�v�s�9�;k���5�G̚����P��.@�?c$�_��(��I^�<�j�d2h\�uP<u�Xk|14�uN<�+\A���W������W�q�/ʬ�M}�)}7��ݓ�b
�|�ᇌ�?����������y��/��97��+_Ġ"Ό��na���( b:�~ ���)����$�|p�ȳFUu/�d�c̋	E��y}j� \�]w��Aٍ���s������V���o�v�	1y�"*fd)��Q�#C��ZU蹮������&��x�N2���T/	su��w�i,9����]&���xp/�� �ʀ�P3���ؑ��}������}E9�[��\غ'
@�,ZX��K6Ph��v<慻��h���غ�,�� ��`�y�8��U`���ڀNP�c^x�����^{�e�6�L*a6�辌�@��g��{ԠhZ,7��I~8a(�Y ����-�Q�xl]4�~{(���H�G�F�< ���}~*�T��=� ݦk��gE��GcAd̫`�I��K�$/�n�:�{��ן�ҷ���^���O>�K;�A��_�굿�կ�D�7��ʥR\P�)W��FpQ��TkYC}O���]U��-
���pq�kp�=�vsR��#�f�`�gN�ک6�r�M:��RTM�by��!�� R�M1 ��),�˳�/����2.c�.};���  &֦��ܨs	�N���P9s�藯*3��
q	�QN�!6-s���`mJ�7�`�|<��P�Ƅ�c~�`�3���p�YG�����~Gë�Gí��WX�ڬD��en�3! ���?`�!��x�&l�a��,!�g$+ע �6%=S;u=mі�7%�������7�u�.�vdY�+$u��J��}�"��UlY[��"�V�5Ő�0L}e�b&J��*9����,�4�zf��Ov*B�_��}לz��� `��o]�����{��b��~`���X��\���Ն�{��֨�Rl���{�Y[�N����	� �.�~By֪gX+��5��)$s1kkc 몫%����>��(�.���M��+4P]�����Ov$����5}�8�8��o��	:�,�.�P�b8jc�"C�s�O����%{ko�o����614�.���Ϊt�ߡ���+}J�'x_r9>��X�K��I���a?���122)�����pk�AH�?�h�l�sd��{ﵓ��F~IQ����K����y��:ϼ��jO4J�e�=~��{��韘��A�-���`�M/�$t�Ǥr�=  ��ac���ˠEf-�(Y��$����)bZu|$��(��3^d���ũ�͗�l��g�s�?X���O~��0 (B��e���q*1/)t��N��*�kr#��b
���Qe�����?Z`��@��>ְq
9�&�<kO�Z�]1w�f󁭸�=��75хΫ�Q�c�"X�;�)>`�D*mPh@a���"P�뮻
��y���ЯX�m���h,��
Vl���W�X�1�|k��%0?�&ՏYG0@>m���=��*%�Q�z�dXd�2,��(�\틔:����Oބ.�g<C�H����	 �e_=�@��-��"%�`SL�O�5�ʺ���%������^�f�<���gP%]X<���ZO@`�U
�cD�M��"�����T[�ELO�#�|��#?
̋?�0��Xr&���\���~F��Xz$����n9�|.�^��t��ٟ���_�Џ�z�����?���������X?��n�s������	W���8Ir�"�G��G���cl�#2k�AX`4 ˂m'���l��I'Bꞃ�-y�,J�)�� V�P�x�������l���1��U�QUp��w�[%&�����v0ZN����И�V�!�,,	����g��  �v��ř0U6���Ph�# �%�jOt	��Ga�1kO!t�H�@���%�f���r�uk_��+�����]�ѪTE1���:�Ȣ��RY�;*��Ic�<��֑i��c��[��XG]�Ƭk���fF^h.��ًs�>���]C�q|��R.9P�ul�^�Bѓc^Y`T�)�0N,��;���}�5{6֚G�1$&D��\r�T���Ё9��K�Gf-��=��E/zq����@�
�o&h`���r�?���?{7�bBX5��,wk���/����$f:D�Qj�����`F�P����R������YↃ5�n��+��P kb֖m �f��b�R��	��C"u�G��Ĭc_"{���C+�q5&�Y�D�_lT h.ΐ �|�/��; ���[��K��`]Ws��U`S�#�WAMlR��Q�Hs����Z������P(�/�4�#�F_����    IDATu
	c��	̯���)d�D."�VAK���F6*��/��?���bj��#� ��"0���F�q柘�$��Z��v�nm�*�����J�c$sɶ-?9�\d�`+3I��g�����W���16Ԡ�D�̶�3� �髌��'��؂g��]���~U5���H$%�v�֚-0�l �Z���.�ο�+[/_���!<�W����~��/����|�\����X��y�.G�\eW|�A��ud)Q��,~T���M1�lEX '���"X;�s&U�`L��t�A��&Y9�|ko��:����{Gk�� F@���|��=�72n��F���\�H1�xO���J��K�b���Y�R���Jy"PWe+�hl�Ɂc4��;k��Ĭ�BLX��R0�X/�jˢi|۔A3�""��w#�Ox@� ���b�܌��WdW�s��_6H<��ghq���Q�y~d�Z�;4wr����X#�u�'��:)�R�Xl�z,��رJ���Z�<G�06�~���rt:�����qq A���`-��m<�W�4��d�Xf<�� 	���HX(����i�����X{~���\�ˊ+�z8��L_�������������S�,�	�q��N:s�PE�Yg��U��d��G!:B+��K�(�`��n����^`=6�������/V�%���k)~Q�+O��c�eT'$*@A���C�g�0���*�֘���OL��s L�)�����v�mc���5̹����9�@�����\`M_1LxM�9��"
q��$���zj?�6���'�^kb��E�B-�Z� �W��P���Ϣ�P��ٰƧ:��K�$|�B��x��E��By���2���oNS�Ű�ȩ{x���6��GD�g�!�~�#�~�R����*n��̟�+�-t6�)��\��Mk��Q2AX�O-����Y�;��h,��Ŭ���p��Z����$�q�/�����@��/���vۧ�/��>o睯�'���/����ޗ/���Xۺٔ�P��F�e�pt_�x�,�2$��B�ùt��Gk���r�x�#�2aG%Ra�ܧ9�)K�˄A|"�䕇�(b���ބ�s�ˌ}q��0
�LBL�~�E��MƾE��<W�W.d9^�����K��7	;�{0k����])sL{X�X���=�sk�P��8��q}d6z�D���Kne(�<��*�}��x��@1����b�φ���^}�ѫ���a-�cS�k������qEGqN��h�5Nfx�ef��Dm�gI�I����*}+��8Kf��F�i��z�u�YD:eL�V7P�0��F^
�*l�w0�%/ �J~%Z���:QJ!aDI:��1���O=U�.��2�l���o ���;m�4Ł�44شEu�Xr ㄮp���-�6���N���F��Ccd:0��N�O�/�J��<��Vۤ3N;��җ��3�~�`��r�%��⊿��!��.�A�2�PY:IcĮ#S���NE`��@Pv)�>�@󓁍��	�j1�OP&��JD;���h��Pd��I��ޔJp6}�5��V[��@ .)�	he�CɰJ��9���G��i��,����G pP�(	,׋�L� Ġ�U�dp�|�R���]-�K��댅�c��� �b0�K��v4Κg�UE�EGa3���\gi�r�=~G���v�W���rҮ�!6NZ_U/Cccq��$�[�:;�0�� E��"����$�2��M��_�$ۚg���$�q�6vaT�\X�Yk,�0k�h�l�ČN��2��a�c	͋덯�����i�̂A��
q�@��G;�V�1䞾������2��3������� ��%�]鲰Cr�9�WU lX��щ����~o�2�`X��J$2h��ۢEK�	��w���՗<g���_|у<��k��ք&��A}k�Cy(���2����z1����
�$RJ&��F������%��x]��[��,X�p���<k6Ű��&���J���mws��3�t�L����C��b�NY��E-� v-��!��  
��Md <��r�/@�;0k��)����_�5�$��P�<�W�O "a�6�*�Ul�Y����kd��[d���2 ��@�v�v�����(�óF�G
��]�&��X���+���y���)P�
��6�8(�S�&�)0� _�Ɲg�OL/�1k�5`M�Z/�Â*mƻ��O �1�h$%G��<	D%7Z�YPc' ����	(~-y�'}��	'd� ̕��k94�yS�Z266��X�I���(g��)��ID"������ݨ���v��g~��W��566?y��{�o9�9��]�/g���_B��d��^(�2X����hQ���E�L5�s��tЬ��8~,���;�(�i�?�*�[�z�e�s���}l��}l�E�	�����<L����W�V@d�REM.2.��gkU�ZS�J	Y����,��$���/�{Hx>�M\B1 ��)�yalYI�76f?�&#��"�V��@;\# �9�ӽ�RL�WJ�@9�~�U荾���V��{��T̟{ ^���1?���a�82�
���J�js��:z��86U�Ƹh����\�焷`ʺ'Ͼ����$�)1n*�Mb�2�1�.SH.��b8G�v�3��Zٽ��:Oh�w�B.5E������S�������C���T�TvƓkeH���<Jn5_��ڬ�W_�gr�\zEį/��<f��|�w��]�{�`}�U�<�[����	-�ӈe����|��à�1 UlZ� ,6� 6RCJ�^ţĪ����)���!�A�ރ�.������㿷�z�����!c�,̑gM&!fMN��rba���L(b�B,[,)
���ݓ1T"A@�,��Lc��Z<�w�)V"����- c\�\�580P�5F�b��
�mL:�U��N����M�$ʀ�AL����H���hj�ca	��>�0�
!��M3Ɗ��3�9�lR@����\&Ηb��KU����>G�w��(]���K�7�xc�0�qY��I'y���F|nc��Vb��e�w�����O���<G%����R�=�*��=�ĵ#c�g�+�5m�:���[o5o��2�"s����h��H�
S��j�#������a@'_n��:�܂K˗o����������`��+~q�9�s@�p3''[�M���+�'��W�@B,�v7�<PTn��:�)u��J�RI�aּ��0-�Qd��VdF�a���t�Ŭ��b@���jzt���B���}2�M�mO��g��i��L�71Ml�HW�p��%*8B.⾬�cd�V��]�r<&�ޕ��$Y���X1�}�V��@5�&�EN��1l9�+a��o�y�A`'��
�7sC;�������"����.c�d� k����r1H��c�"�r_�'/N���Z�^�W޴���8��+�n�G�|it��TqW��Oc�}���)a^�}3��rk>�h��[�H��&��qN���Sm7�`�\��ج�D��k�|�9^`-�a�0`��0m��$C�]dFϐ�ƹ6��:!�\�/oK�z-a�������I�8F�~��x��;��=g���տ:�����,�1 �D��z´[�`1���V�s�j|�~vjb86,R0MH��s:aSI�E���`��}�FX��{��������,�|��k��H@J��*X�����KУ�քDA�J�x�b�Qx�wH����U�Sϧ�&]�M�k�1�E�q/YYw�s�R�(���` `xs�b���j6��8�U���R��Tޖ��H�G��җwީؑȸ�a~5V��
����l6\Q�B(e��1���jkDɆ\�x���y�~)~/#Âo�� ���ž��Y'/�;�P h���m�����^�&��l���ƵE�ܓ�=yqE�4��Е�X� ��W���p&��8Ǿ�?"��8Q�.��EC��m6��aa��\?˅p�C�╯|��t���`}���_��<�	�;]����:+��Q�5��� U]�bP��.��]wV������(7��F��P�m��&3_���[
VO̚�ق�e� ���b:�H��R�"&a��X��,�F�-`-�Pj2�{����"ȩ]&����(
;)f�gʊ����v�LM��g����2�⩩鼨R��(��O�K
���N���Xh�M���)v��V)�<7�V[m�u�_�=U��g���z�o�u�W�30B1#�)��t�*`K�grLV����2��iN�}�q���%a+�5�R�����q/� D��a��r?k[87Ѯ��4"و�@^�H���1$���N��F�V[����vK���F&46x�x�r�SP�yDY.=��e��4�[ɲ�J}R���-�F��=�d�����t�V[,X�^���λ�ϟ;X_{��O?��p���Z�֠S6WGi�����[��)����^>v��:(y�Z	�7jS/MĦ��_�nZ��I$�xP��ڽ�
Z�>�!��&��X�/�OƇIT_a~�qƾ�w륋���Lp_V���E�C���h���L,*�r:�R�g1��N��!�@_ڼ����ڱ��C��G��>�s˱ͅݥP\��@���R��ռPD���Ĥ���L|��]]�G�W��HGu�Ԃ~:M�]cǜjkK�0�k��i����ܯw�,�Kf�X;Fe-
�[a<<�(��{��7Á���-ث�2�z_���Q�T\ÒPP��j��S%�;^�Xs_2க� �ʻ��n&��
5ű�k����i��������=�3X_���}��_<�[�/+�AT�̪��Y�|�=�&����uL�*�:��w��_?�.��$�~!!�JT�}�,��0�>�h.��@�+�>����V�Y�c����]@�:���U��o=��"�ZMע\d��e��q�;���3Y����E	���D�T͕�m/됗�d�@1X&Q�_%&�I��5EJ^�}. $d���h~��T���?���F�kd�joIJ�y�1�s̽�;Ɛs~"��ˎ^Y�n��G�1��
��U��gh ۧ���o��(�p�(�y�%�1��@=�9�z�2����b�z�b���mW�O�KCRlr����	�9���`��g���w�+5 /7���a^m�����Ǐ\~�n��������-ǝp�`&�
����s�5f�+3P⟼�֪I�Ke�\�j�&E�:Nf�=Я�*��:��b��rvo�m����+\��~�̈́U���pԶ~`]ݮ[eB�����p�^)�/�z�}��+����D�5�7����i���U�g��,�|�%cT9�G�E1g
��*��������=.J��γ�7*���O- G(��Y�b|v�����:������Nc /M� #2��@m��w�I���e����|`�kg��;8���s��.�̚W;˗��ȡ�g�pd�[�M1k�sg��+�E���A�fPrD@�Sd}Ȩ��Y�_���~�����WW?����]��{̱?Ҧ�Z�{�%� �����ֲ40k�y���`���c�k�	Sу���T����9����IWLO+2�~�X�8XTd]_eőY^��X��������l)�%f�{2L}���?R�=0�~����<�
�6�y����P�P��i�;��b|QJ &��R+�V�[��
���~`R��2 �]�'7�0���V8����3羚S]�EYg���uJ��w�M��~1��Hg�hf�ֳ�`����X�[s��F�ŬE�z�u�m"���Yֶ�W�+疺@^�(0�W����z.=,� OW�-�WT��}/�Ɍ���d/=t�W���h?���]}�������(@Yڹ��0�u��u"Qt^u�g�<�d6{ۊY����'4�����:1h�C�2Dc" ����9��G�QW�b��g���Ge�x:��m�w!���z�-`V����7���/)G��sʲY�(�:0�``y^�w���Y�/g���GS�P�km��r�D&gP�ū��h�{��X���s)wk~7¢�?���#�����~�؏UW�TY�����je�İL��U�,90��fy�;�h�%k�#Pm�bU��ђ�g��2�)�Y�	��������I	��[���C��si��Y���'�.�6?8���;�7\{�^��Y�X_}�1_8�GĬ�5���<���)��� k�;�	��I,@1[kY���lX���h�ʾb��L �0H/�,,���O(a�E	��{2�b�ꗀ�*d1��ګ6��M��h�M�IJ`cA�9���z;2����=�X���BjU�9�q��,���,,y�z?mC���T"sf��1��g���D���唸����' �`-�^���Q�Kw���sb�C��?!�h��}�:.�
��Vu��=�s�(�c�{9�&���q�Q2��Jw4�ֶg�x�>�����}˱�8~�gx�Ⱥ���}-�����Wƈ�r.�ֹ�WW��f�m���X�~���w��?%eO�1F�d��Ȳl���.sl�3����-��� ��_q!է`ݡDjѧ
Îa)���O��1���`R������H�>d� 2)�"�;�������Gъ���Ǯ<W�aS�ZcT���W�'�Y����Ȁ���(�,02�_4<�_�^����+�$c`]��" � ?�Ns��D�Q�Gx^�*���:�U�T=��0frS�* �b��X�O_��>̪��|�_�)�;ږ�����a,#9�����t��>E9��Z��R�.��[c�Г�Q�}�z�Y+:3yXk�;9(:��	�}�j�d;9��X��qU��Z�0s����ӽv�}�6��K���[�9���I�X,��&Ƭ5yRX~6�Q�3�0�nO���rO����[�v���Q���F�
��!K]����c"�}��>!1Y^q�1��1
����Z����'��7V�^E�`ZY!R���~������/��%6'�	�����Hȉ�	��0'�ǟ�*b;"3R���[�r���2�.w�u86]m����
��8��*XW���)��q8^�ض��ͭ�c�Q�J�SI�<�G���\w�U��2_��s֜�{Q^ln)��q��\�dZ�)�".e˾�1hkKH=�6z�^���Q�5�Fm6�S� �*�lis �Pj{^����fm��ʅ_9�oxӏ�n��}^@�}�ݹ��?��_�4JsL���v��AJ"pgG�	W˫�ie�3���Ȼ�TO���e����Xe� (�&��ĳe	5�j� LQOǬu�� b{Է(��̈席 L}e�o��E�`!�
�QH�f�F�"��:yGb%��b�:XX�(T{�#E�W;��uj�⡸�aW5O�̢E�bl�~\ܦ^���Ac)��f��nZ1<���3��a�b�3#�����/��3�}?{��V�実і>���
�H��y�4�s7�O ��CL��<6����0'��q�F[��t�4+��S�s�h�
p�����Qa%�Y̺Nҡ�*w9�ω�(6�y!u&�����J���RP�n���q��|�;��O���{�G~=E��� Ĝg-�(�����{3S^�<�*��_I&%��[-jf��ƪh�\�B���/��JX��I���j��Fʔw(�9���p%d;fd�Z 3El���z����1��*`k)��Al3fNh<�����0�{�lήo���`ܼ �[���t���Û��:� 4�
�l6m<�ZJ[�B�dk�\Bc>88\x
��?XG���ī�n�;-0F���쑡J�8�ƭw��S�Mv��-F~2��W�|�a��O�iEx�_��w�[�o��Lyc��y���x�6�wXQ�i��v^e���O��u��7�����5�9��3��w���	�B�B    IDAT�W�\�����<�@�� ��s�ufF9�E���	�̴%D���a�L{
/�\��>���%�Q��}�:2����:Z�~@i�,���,�T�$Gea�b�n$i:oW��*E5 �`�W�'�k�PǸ��������3���̑��q�v�Ov�]OJ+%�6�R�;�F�v���צ����d�R����)Z/Q�F]#�W�٨]e�F���# 󐛗5(��\	��~̺�^\t��X�YG�察��l	�~*�%�����V��)k4,�ۭyt5�W�y�g�^�<����:ak�&�c"a"Z)�`�ϊ���[�<�f.�Ɣ�/��q��6�9F^]XX�/0k���3N��zժU+����衇��#�N�M��L�	WN�`m���S��9y�cL�Q��Ņ��/p�mF�v����k�@Eō.d�gJޟ+uϮ#=�vn�+���X�k�+\
��{նUYo�0�D��3h�+��_�;,�"���ʔ�IFX�Y]<��R?�6��[�7�5�����6��!�|k�SƩ�� ���H)j��q*�z�=�j�Ӂ��@���Ez���w��"9+�0o�a�2/��i#:50T�I�߲,��Ae����]}~o��DO��p��Y���l2�ٰt��!���w�_>w#�Ӗ��<��Y�(vq��lsǼ
���_k�c��{�����]�c����{���ȇVrx'VE\`�*���kt�-nf"45嵑S���dm�%(,��iM�2&��o�#J���vr�X1(}W`�t���@oI�Cؙ���
���Җ��V��
�s퀫2�*+��Z��h�X��Q�g��E)X^-��瘂��Ub�Ϛ���b�1kg's�b�ZlQIlK��:�6��PQH��X-��F�w�(z�˵��I"ʢ*HM���d��阹�/��Bj�IkN��W�:�T�o�7�!��ȏBZ5�jaӜW��r��T^���~	�i��^;p�S^h����^�on��E; k#'ug�8����WΧ/�Lށ���M�m�{�*c{�7�|�oz��^��g��=�`�z��E����]-�VySuDa�h��j���$�h;3���d�B�mչ,�#`���؍���)vd����{4,<�ʬ�h�5*U�~:�vw�!z"�]V� <W
=�)w V����41k}���Z¯1�0ֽlĕ��Ÿ���S�"N�[�G��x
����g�����y�﬎g?�`���A>���!+����J�����u����-���D6GQy�怵����5�O �q���ߍS$3萲�dx#w�Bj/X�����u3����0?s3�Yz��-�`]e�6g��ⰍQ[�^�?��Z��'�����J�vo�v��"�����W�dｯ�(�I�t�ݡ�z���x�G� �N�-@/���4��h0�~�$���p��:O��RVL���L ��ԑY���҂EV(f�L�Z�o�~���9h�� >9�)���1�=��Ȭgڽ�[�IT��	`40�X�P�y
Uȅ������i�)�D�7@��JY�v�!���Fa�� #X@�!z�1k�u4���2��[���º���L�&
���q�V�#�Xs�-�nT5�w��<�8��y���$�Yb?��z�o�߰� 'b�vM��%���N����t=-���g�*�]+Sq]��7�m��v�c��+��a=��Sf�T��@�3��o4���<�����g���x��Z�[��j�Yx�p��ʬ����Z-��_�`�v����u���z�ڇ~x`��?1Y5+'�c��qK�
�<�	&ݶ��Xw��P�H�52BV�O>J� Ի2�|O��\���F�ZF
,��4X�]�������p�ﴉ]�nL���y�RBF�r�&>�;����N	����Vz���gY��)����칖� �F��:V�}g����&/R��А��hi���Wq4_u�|#)�ؽ�ϔJ�.�nJ1h�)=F+d�}d�ҡJ� �G�*+s.c�sH�c�;��)KF�ۏB�+��T�rdeO��ndus+�N�C1iy'���,@ =8���e��)t>N�r-�b�Ԓ��|��i���I�@�g}$����	 ��R�����͆���=�_Û�4/#Z5�;����f�p��Xf�!f�W�f/�����,]�b�S�����IW@	����"��X����̤����p��4��k(s�F� �����պi�=��� r&�O��Sk oze. ���b�6�H��Y�x��"��pUr�o��lSO�Ɗ�F�t��6�7 bW��iz�����NO{>l7����߀��3�5�ԁ��M��Nɂ,ן������,��Y�?.e�h�dLx_�)�y�3"˾��yu���l��L���4<B.�ˈ�[��-~9���qkO����Z�KL��f۾@53ˡŽ��{ �^�猌�ٸR��`<gZ>�<����w��̥�P3��"G3�n����I�J&�b�m �6��{���EVڴh�"����V���5���[n�(
�{J�Ⱊ'��YҷxP��&dH�|�r+/ K/J�.�M�U���]3ƃ���r�U��V����X�2��3k%�(�fR�S��)5��y2���=?�|���2f��h}hs��X���P�o���a�4��&b����n�HX���v{67��P3-Y�(MNl0���E����[h�|jUb�.���LLΤɩvJu������Tox���ջ)cQ,Z6���n�j���f�va��n��7�~��Gׇ��:Գ��UB�0c�H�i�y��^sw�z���(c.Al�=�fff*-�b��k�8n{0M�fS�9��3ͤN�uo�`�gQ ��$z�u����?ED�JcX0�P�7�d���?6j�>5���G3FyC��,�M�U7�Lk*�sz6ML��� ��4
���i~�2���� ���S��!ע���@�p�(LS�WH��B?4�H��-���1�SZ�v���f������n �v�8X�<59m��"/�SO-�b+����ֲ��Ka��\	h�N���d�}�M���'�h����v��Ϥ��rd⤚3��A${P�����mz�X#��`#MONY�~j|*͛� �ON�VO��3��B��}��0��1���T2��7m2�!���ty�� W��F�C��Z{6���E楑�A��险|JO'��.��2�rj�e�\LM����T���Z��!#(����z��"��5G; Q0F������H3-�2N*�ŵ�M�_��g>�?���ϩ����il29��X�8�oX�F��S֏O���C��CÃirr܌��;�'�Z��ݡ41^�-�'��`�0��i�^o���GFj�>K����o_��C�!(���>�`���P榝RK;��t�}��Zޡ��Y�V��� ��fg�Җ˷�g�]3���R��H3�ņlo�o q�f��d1� # &�� �<�MSx�R��7�Ah�]I]so�<��w��ӒE���Eғ��4�6�4Ó�	���v�
8-�?�V=�:��0��9Zi֋]UK������y�3�����:%ت%�q�"���e� �NgV=߶�ߞ!g���.����jYZ��44<���Zi���x6aˠ���,�'ӊ힗V�|"m�H��8��S��#cK�hT�}BÓ�Y>~'Y�af��(B�WՇ�Ѐ��۞�[뤡&�Q����X�(-Z8/=�ԓv|X���]��l�n���Ǯ'��0���f�&��m�"���c����FyH��������Xlf��  zQe�'�:M��	�P�u=�Q���Ӗ[.K��
3"~�}�=�zIV��7����4o��oIk�np��i�Z}��?��,�
(����:�-s����Af<d�E���q�*�s�P��A�O�z�YK������4<��NK-N�i��49M%�z�����Ԛ�0�z����ϯ�*5ci��a�D%��$��B�'3ɘ0��V[����;n>�\�u��������-�N����q\�towmˢM�l{*��e��7������SO<��`�n�Q`��v���,�)�Ś��S�>�֬�L��U�,��� kgֽ�6ȗQ��Tv�aL4�MQ$/ ��:�`����z�|=5�iŶ[��w�)�z��'��Z�oxx� �X6m᳑��p�X��Ҫ�Sij�0	 �!�:3}���O������Q5���X���F��)���*�:�A /�th�is�|�����6ML�K����i�ؘ�&F��`b�@ɂ��i�����˖-K�����z�xjM��H-BS�Ēʪ�I؋�MBMys������b��2#gՔMc���RCQ�a�r����M ^���i��G���D>.m��؋�A˰P/a�̓�4����Mz����dk:ͦF�5c\��d���lE�ny�b��̰�/}�K100�Z�n���w߽�5k�fl�ڋ�^=�L��\`m@X��ѡz��;�%/�+��oN�9�v�44�HC�\Wd۩���Ng��E_�ZZ�ت4=�I�l0I�1]!�X�6P��ZS�2�{�����^���gf�k�V�y�o��G�(O�B�a�h ��Z:�4:2dH87�����K����[.K���p�B;k����J#6?��t"��������Ǟ�֭�J&1\)ͰI�?���1����E������~�`�������߾e�J E0��ìq�U\?28`����zZ�`4��{N��rc���J#�C��2�g���575�����@z�ɕ��[nO����P��nq�Y[uō��b��xl�6m��W	׼{����&M�坅���v����³���f�V����Jo9��i�Ȑ-F�d���>�v]��ٞI���Ӆ_�zz�ѵ  ,<�uvJ�K���EEr�/����0�+.,�sŞT�\��O��用�$<�2����t@o���������E/�-u�����8*�"��`��'V��N=#��o�Ok�O��5S��J=�xu.��}��G��ɥ)���`ϙ��,b�x�L�^��c�R���س �ɏ���^�G:��3��7ՙ!~9�,J'�d.���t�g��������x�ye]��Im�`��0gʄ^d�.�ģ��\r�_��Mo�?���\s�K_��W_���:��r�+�R'$�<�1����ҁ�1z����Ȱ{:���\������Cv���J�~��t�����l����M^3��󚔞�E@��)� U͘�O8�c��ϯ��{��7���?}���@�u t5��*���<^B�L�ѱ�4ol ����Nx�{Rs���ӭT����r5�:�\�]�W̤���t�]���|�дꩉԚ�����Ge�}l�6|9���N�}�{O:��c?��������а%1��R&c��qY�"�94�L˗-Ng�q���e[,�8��bflъ}��㫰\{�צ�=>=�rMZ����F���S�}8`��E�s�0O���N;�Y�}1��#&g�9����m�4'��X����i���>�яX��)��F��/�NLMz,�E6|g�0�J��z2}��G�w_���EBJ���R�E�%���/�e�̸��r�������cxx�3==�Ek'�p�/��������O�Ҋ�1�P��~¬gg����`Z�x~�c�]��'���.Y`-�{��3�0lY ^�41�Z=�ju:��s��yeZ�n�#����7׼G��Z��
�G��|�k_;pٲe�fk��4;��sGw��W�Q쫟R�@,��|�Z�N�72���}^���O86�LZ�Y_�֚�-V�\�N-�_��}���E_�$�^?a
���01����[���p�93y徜T����ݻ���K����/��c�=�k�V?6�y� �Ū�FžˤO��qd���I�����S�;����nM�n�JT�Ҍq�\�{�|�����OJ��rGg��U�)�!����Y����Z�Ǭ9���9g���o}�ۿ=�}���.��K�Vay��r�p�C�~t�p/�VV���@�?6���=�J���R�5�2��؎�fjM����=��䓫�G9<=���~|:MM�t��F���y���z�����g��h}��sء���7W]�r���\k1ո��UQ\�fd �Ӓ��Ӆ_>7m��V�AP�x3q)B*Eh)^��Ue��t��;��}2�Z�>�]G��u#�\y)T��aS$��16�'&_�T�+V���w��/�To��u''[����f��}��/�����H�v�]X��⥣i���>s�ixx0�NN��ݙkF��l��`��)ug���D��!���n{0M�XeG�-��]�
qU�Z8��CM�;3��;���>���-����C��w��ݿ���/� �9�= �SqO��R�v�zl����?{��SOI���g�!�d5���ɸ��̶Z���.�8���v"�7ϩ��#��	ۑUk;/����Ꭽ��z��s��^󪫫}�v�������?���=�\���
Y��S��/>k���#i��^�N<�Ԟ�4��P�TԜRj���aa�#�/�A:������8�Y����Ś��k��6v�#��)t�A�:ꨣ��)&v�a�8�?��g�	��G���{f����I^0 ���^���g�H�3�d,v�'|K�l��NJv��u��ϝ����ƴnÔ�%d����K
F.f�CH��{�@���/���7p٦���~�}��e���`�y�]7�e�s���K��P�h��!�`��z�[��G��4�H)u	ei4-�����p.�a�d:��O�;�y(�]�`M�Ck��[�R-��1�J�җ������˗o�T����⊟�漳���#�<�-�Z���Q��������7���P�b٢t��g��om��鴋j|��Hg+B7r��}������tz���R�=�V��L�4`�om0��J�kvu��r']�|�u��[��i���e�]���?7�	um]����H��y���pz��������-J��5@:��=�V�bc6�d��OzD����6���jYl ��X�j��Z`=0�L��ַ��w�}�i�>�o|��XkNi���(X?3X����4�zl�`��?ya:���m^[��vg:�<���$`4=�.���韾��4>9�ƧfM�1B"���	c���ڲF�1���>�����~?�T_���������+��V�5�KJY�)�;����x�����p�=��6D#/�wuC<0�~r�e��s��֎����t�n�ص���u��j��VL������-�w�y|:��}�#g\z饇��n(^�|�g�A׀;on��:i�y�����۞v{d�|}����([�HM#�J�~�d:��ү}]Z�aܲ}��xn�
�;g�X�����!�2Y��p�=����g��n�;p�����+���u
u���/�@R�LZ-���8}��Nzˁ�OG~�Ȕ�nf�̧�����-��9v���~�3���K㓝41	A!�5�@S=ؚ�g���_�G����+���jn��k���k֬Y�W�~�/�\�rKљ�*�~\h�����6q��'�`�H�v�-��g���/_b sQ
O�,�i2 (A���t�a�L>�Dj���L=m��5��a�e[����l+���+��L��vۻ���k�Z����;L_<���N;����4gs��I��ƗmQ�V�=��R������o:��-�۞1`ƨ�Pj�,4@臼L��������|>]}�i톙Ԛ��4/�Z��A�f����k���|��=�ɿ��%{��u�D>��O�����)N���^e�l�qfM�g4�d�=�y_>+�[�1<H���р��}�*J�tҷ��?��|��i�ډ49��t��&�H�,k�kS�e���g�k�n�b����|������>��~��/y�'�#�Z�2_�>�h�f�F-��6:���I����t�1G{z��+���d@y�������SO?;�^=�6L�S����p��,�v,+���`��-o��.��=�~���q0Q    IDAT������'��NB5��#��6�xHD!��4<��V[/�숓N>>ugIAlۂ8'�wg|�R�e�ߐ�7�M'�tj���I�6L��lײ}lIG;��̓c-��q��Җ[o��M7ܸ���1�a`������7߼�\A��!kgI_�n{j^���f���,��^��>�sGڼ��N²;�i��kYP�oX7�>��/�k��%�ư�F�u<?�Nqt�If�v+V�s�_����q���<q�������XCZ�FxW.+I�����I/hCۖ[m��:�Դ��I�XIı7q��7�Ji��KkV�L���ߧGy*�[7��n �-��0��L�\O���'�P,]�������G?�4��WT���i�A�K	�.��:��N��Cd���������Y�?�u�{��k�{����}��,|�P����s_�pj�`I��5�6�07g��n�uT"�ϛ}�NAekң��"`�^v"�̞�!q'����+���\�4�6��O��&�5��N�b���#���Y��p<zJ�����#��/�J����x�ѣ�:�>> ۀ�a;�h\�WTÚ*o>�k���Pc�3��]�����Z=Jl��{Il{hU��-��f&�4��w=�!R��-20hh�7��H}��5[w~Jz-`�>^H�\�J��� �&y�*s
�=/~t����,���u�ĺ5O^��X��R�v��V���YS��|:$m�b����^�
Ps���8(r�`�a��C�B[��w��w7R=*O�R	���jݫ�ӔhK��A�p���S
��祢����m3[u^r�V�恠�DV]�?����0�6	���]��"s��H~I���iQ��=6Y�k��ͪ��Wp�U�,���
��G�+ZmO*	H>�ȶd��K�Ca�UT��T������w��٭S��4ɓ��;ꋌ�m��6�կȸ�ig�l��<I?獵r���+�0?@��s����m�d;����j�d���D��c�`X�x�/�gc\��*ķK�Q>[^-�m�K�������!�]����*�(;�u��k��B��v�����"�Ō�q�|��M+��<�Q)�������Q�Y��ј�۸�$���_�r_0��>�9F�ْ�}�wk{ȼ���T����'���e�O�B��KWZ�I�@��I|����~[E��]�D���QyuK��G�)N_'mA�7g��Gޠ�T���y������N��z��
�f���*���l|�2�}m�m���ff���K��_YPt ���rI��]\��M���]���;4C�n��&/��^��[my�F��3h��&�h
yO����$v�����p�����q{�k�����^�ؤ���~�D�h�)\�+7��S���g�̳|��7��0�svkm����i��~x:H�����?��>����RS;�K�;!�)�n����mz8�_���؊?Y5��c�k�l�vjʹ�0+��=��@����(�f<��;-�ODWk'�����Kds�Ǯg�r���_�f"�]��h?�33��wێ}ֳ�]N=��hVlM��E��.Nar����n�������#o��]�<�y��e���e�'����o,�rg	@H�.*��ܳ�}MC�|�L�E�ӄ�+U�5����rX�	L�,��Tt�J2�^c����Te�&^^*O�:��v(�|�L��J���~h��OʊR�d	I�z�,w��.ɳ��e�]j�8�f��72�J���S�HQ��=�}��I����{�uc@��I�p�[�g+�󜸟�b�%�W����0�%e��Nʕ���$!X+c��h�%,��������8��I�#���4?�J%?�K.|S�u�K�١;��Z;��n�`�z���W)����N�2-�L�xd�[.��*��K��՗���2R����n`��C��	��Ԛ�]���Ă��4�V�:L��a�z���iɡ/��?� �x;K��ǈ72�Ĳ�
��d�:J� ��Cu[d��OX8h/����*$��'8O�_U��Vi4/�e��1���rVP;���j/.��fGE���+��b^�����ᯤ۸I�r2$�9�{vvƤ�s�.�7aÇ���HNAS��R�-ZsU%��u\��Q#<&F����Kf�wy?��	^�������_ޅ�X����c�z��z���#��{EN���4���{j���B����]�E���d�UR���7��x�uhL��ǋI�B�h9�{11��:�z5�w�/�/j����J�	)aE�{��|�w�h��M ��m>����l=��:�"#m�\��оi�&�*��v�M�l߬Z�b_!n+r1�$����w�t��U�r8� 9��I���J�v\�n3T�fe�nmk�W�tDqVN����xf55��A^T���v�/@���F��R���m���Ǐ
ɵ��%�E���v�H��y��U���.s",X�DQ�����G�T�fE��<
�C���41t�̪p=�l�u�c��� ���Il.s���Ruao��~�jh߯�g+��v��/M|��!�A:Lq���n
��w��ϸ}��Ww:�c���Yc�\g�>��yOl	){I��r`�&��7|W�>+kk� �%����������O�f�p�"M�Y�u5M������X�㭗��R�؍�s���c���5��I$~�o�9�ј��mu��M��q��~�H�c`TΤ��2 ���q~y�:�P�u3:�鱻�r��HN�t�v�Ĕ�T�SK�I'Ȼ�"U((Ȼy��%((/���ёs�S����42�-x-��P����QZ�X���N$3�1���ڪ5��M�ϓ7X����5���6��}ݐ�zb���77=Š��OSK��7T�v�
��|	��:W���w�%�xJ���p䗇S�8�:]\�>"�F���IA��Gx���q����Tz�{�os���u��j��Sg�7��p�a�⽫F^�ܼ���"�*�����K�����B��Y�K�k�;��J���
����"�I��:>�B.�c��\��_�N��r����w	�3WSf�aB_��X��:^�h!e�\W_?P���yꙙ�fi�QsnQ�8`b'�HC��g!8�1�LI��k�! mJDN>��	d�hpm���`����V'�KAh�b�3�i~dd�a�Jۮ����g�@�d�����%!O>��,�H���Q�5g�ؗ�>�#�P+�6�?B�N�<W?�2�ʕ۵?I���=ZM ��O��=�����<������=��MI�<v(��;I9b�i.�E�1-��,��������Kռ8O�ei�1�Ƿ��i:Ů�ᰟ��%�C�t�;�� B}�~��^������]gl�~������d��;��>����ѭ����� �Yy��R�X<sS}�F8���1��j,�!m�{����DCc�
��A�Ң�߃	�EB>%�hx����A-~~~�?==��jq�C&11�3444�z����
TTְF�yB�d��MD�af�o-�������G��{x/vw9$���,��`wo�g��ξDJ���ْ�x���j���#`������d|/v�S��Ďv���IS����IE�^���u�OT��Ĭ�֊S2+N������B��$�~��X�鱋Ѯ��U6�d�|6���5�c@5,A ��-p���w#|��%�h|qץq�/��_i1�嶅\�$����pt�R�d�:1��a=�@�����!+���Sz���Ŭ��_?~����x~�f����?o}��X*lY}���l�E\ت�`��Bɧq��O�d5G#D?	��H_�Iy�If�g;���O�c�g�%�띛��c�O�n���.H�q��S��� ��T�VV�U�.{"��1�/ot}g?z������h?t(�( �cFHS�����R��q�n�>�oJ��i��O4��P3j�?�v?���H\��}�q�<�=5�	�A����jk��3����Ur}���f�����˩X-��R��������։�-�����B!��Ȗ�2θr�Fb��;&��vx$�3a8�T��´��6�uk|�_����������w�x��xN�5�z��w�|>3��R�=��1ܦ����@�"d��tN�9���&ԆM%��\�m��{�#���~Qd�k؈D��4�����<��[���5b>��e,Z^rȳё���I���
��%��~n WAk�{��EC�Dz�,��QLP�g`A�~׬�}G���';���tw��\+��c!�/`w�n
��#;K���������W�k�z}���~�-m�������Q����:R��s7�;6\nj:1��E}���汫p_��{.M��~A��Jє_u �X��Oy��^Q�
ȿ���˃��͇V$��V�D�Qlh�{<.Z@-K�gQ�^H/��a<[�]�A�e��
�|�xv��6z����{�l�Uu�ԋ�,c�ީ&H�N����\OU@�%�#5��B}T��g+w����� �!XL�y�G�;׶���20�O�����0a�X��x̙��ׯr�cwkKC�,�-�j�6�?��h�K��}���T�XCk�u-�ǂQ�H�n�^UW9�Xe��wxX- @�.I��;2���/V�1Pϩ:��'�=$�5>zfF�^;I���ysZT�a��LCMH�C�jG��Y���\����������1dt��`�`��Ms���!�
%;�M���������*�h0_pO���Q2'�Β�2aGZ"�����P~v�:92���L��'y5 rֿ�X�e����,m�C�-l��(�܅���mWg�$2���tf�K�r^,#���$ļ�9�:f��hS tVP\���ԕ��ȑ�o��v���>S���Y�����R�ݮ̪�o@��Kgڰ�!!����/7`�/�;��x�˺�a��y=J�R�t;���π��|`hS����E��F	�@f�ð���>���36�?�����_vg�T���>����f(qd�pS���˚h[���!�:L������+l�*�R6�L��y�ɉk|Q$�s���^�q|�j�m�|S���ys���Q��U\ao"R	���S1k�h���G0C5[�W2�XX8n|$�Q�y��{fko{hRB�ŇDjڻ�%�BH��onn���Mݬ$�����ƹ-v�+��Y��P/�&E�M�s|GȈd�pK���ձ�Wͪ82���kPR��e��ntG� �Q�`��=#�ƱY�[�`X�fٹ�+n+ݶæ��ޯ���n���Y�G�G y�5�K��1�<k �g*�l�,�V�z�=�da�0���mh�ڢ�/���)��G�-�Ҷ���3�����Q�y|�?��τ`�xt��a����P<nb��5���^�E���!�������9��OA0�ZTW���x`~����_��[��zE䅆2n�V�oW��icq����V~�Ŕ~
׾Y6���<�L*�?.�I1H�c�@�T�6M�(�|L&L���=:��E��PO������70j˸��`n��+����7`�m����z��')�Ĉ}�B�a�J��jeAŠ0%�U�ƹ��T"��S���f/���C�20� J�s�1,�:|� 0�*��v�»����l�o/k�b%���m�?"�~˿w���l���������*TE�)��
��p�>�R�� ���\�e����+Rи��B�:V.֍w�/��si�C�o�^I�S�i�G��ZN���O�|o�����"y�QM�]u*d]_�;��P\a��l��۷m���sXo&" �VC�����3G(���� ��C����q�
�G%0����/#<z�"Fx���������HqKK����h�8dT�Uf!P�}���u�W��Q��̎��,=i󭸪$V �}�[����Еx�4�2Q��2U��A��C�??<O3�*&F�x�;�<�nj6�����ԫQ?���u��ﮫ_fF3���T̆5A�AR��أ���k�л?xe��g%���^�`6���
�Ď�:u4�7���*G�\�P���AEL���Q�oѽK4G���c�U7�Iے���{�h>	�y�泤]� �N;�%'Q���	+d��2���۞�CIit*�̓s?gZ���&3.��{]I�ߵG1���L�vUޠ��O@<�A.�n�eG!���k^\�Z���Z7��~�K��\����h������)�4�w�߶������B_Μn�d I�gaF��ejb/��>����8~g���1��C��8R5~\z�J5��~8�C���)��i��֮G2�2��|�(��Q��b|>F����<�B��ͤT�Qn$F����hw�E�K��t�v���,��+�jˮzK�\�������O���VH��Qv�\�!@���U�~!�'떕�i��P���3ŋ �4c_��Z�F��#?xJ��.90��_����R��#i�|(�=�?�����I	�n��ϰZ_ƻ���M����D��+ZXM�8MmyUD�+ف����f���2����#�P�k"�<-���>���%��-��z/ΨxZ9�F����Q��`���[��91h�1N\��������Q���g��I�Ϣ��f6^�(U.lY8���2a94��84��?	{H����"��4�=$��|�}>V  Ϣ����UIc|�~ ���,��H1��1B�����t_�[DL�/�s{��h��'uұ)�*$��W9YX���M�>*X�+�"��MϠ����s��w	9��妊h�%Y<�5:���wTH��R~��1 �#��t��rX����@ty�v�����!!��3Ĩ��UR"�F� �he���~O��L���-`=d��V�����]�i�Xd���ⅼs�*��r�X�^��T�<�|n��n�h��7}�����|a�t�蠭Ts�ս��T�V<��QP��X��np$τ#A�����>��x��2�`�v�+�k�?���y���:�h�nN�ӮIT�8�qV
�Ȩ�0��yUm�����$��{��}o�K���D�����*RR7.�����>Kġ��L�;^�S(!�~���xf{Ѧ'*�d�U'9��K�[Xp�Q��
`^'>���O_���l�ɩf8;�b��m�\��5��\�����T���i6P^��j��bקM4����� >� \u��Mҽ�	7���@C��|G��[�+\��h[�$oFu2��J�4�Y��S0�r����?�д�_�?i�[���Z&B����'e��}d|��2j��]���>������ފ�������/K���j�t �wtܕ!H�d�������2�_�ύ$5>��+�KL@���珟R�=kIDC-���|����E�{K,v?]�Jb}�nY��4<D8���Q�2�s9�D���.*�AJ~v���=�P���vaQ�B�v*I�
���#����R���b��ߣ��%�y2���
���n*�J�-�]כ�"}C��I�N����J�R�M�?��㷰u���l`�J?D#�����w�~�p��?8<U��G����RQ=���|w��-J���F�4��G�=ٟ�m
������p���/l���h�	�K�S���!� sv�I}����!��\∝o�& ���J#���-h��=�Y��G��(�(P�^�����f	�Xo{�ٗ������n'FV�t:��	��#נqh��ւE��l��y~�̡�'�O1���!���Kj��S�����s3=��*rY��2�L���!
$!�,���2�.(�I�=�˹����6w��8Z<�=��s������#h	�@a�C3 �`�g�(?!��R���Q�� ���%̖�鶿�Sq�,�>���d|:�5�uбH$�$��,��擯���)��GGP+�e�F~5�`�����ٕZ���O����=�����cC65����b��3�Y�*d��a�&葯C��TD8	$ɼ�� �hQ9>�����O(�ݧ$Wr$�x��7� ��fB��>+,��x|��t�&�9J>1͐�nQ�b ��e�~"��^o4Ή��K1��~�Xt��I�|S�" P�>}`������c�J�'p��G�&[&�����ن�@'Mc�<�u[���A�^�'��vz��,�5���������VAkC�Zb�e���5�: �ժ���Y�}b��_�5��39�b�z4��_�e=$	qoa��5|���y>|�>�G�:V&�>�����Ue�ZC�~)I3��lC��l�*�}�}�v���nG��|N�����)>iP�J�L�ma�k?���l��ʨ;g�HG7�c�gi�R<?��#H�X�DB�~O�T���&M��8��5��ռ8�C�A��?�gb���;[I�#��^����i��ժ԰�X�`��g�D�|�o]���	0��p�ˁ��Tq�0/� ?{&��+���wKD��[��v���8HNs�D�kB����hY>#��e�G�����~3l�1=!�+?���Y�Kg��X��WγS�4}����^-P�����������#rPt�U��nհ�R�p���v�l[�W��SRֺ>�W�|��l��qpY�/�x�ұ76�u�����V�6��g�t��ԝ���@���#�)�y\�Q���Cg/)Ioީ縡|����>g��
�$�n�d�(�vCB�[{��5/OZc��z���\}��PY/މ��㾯�����Y�j6N�ۅ�:��O�͍��֩KJZv�rr:�cy,I��Pt[�Ң�h���i˞(�V}O�Þ�\/Ml�{_�ܠA�F�{F1ɺ���	���=�2�$���G�� �jGU�J�:�;ƣ[}<A�W�ok�by��y���սq8��j܁��{���>��*8bp�t�˞�h�;�a`*�w�Çph]j�N����`�������s���j/ܮ�c7����Mi|~~ZlX��������J����\IM�5pk}!f�6D�	�|��<<������7n�F�L�U7>R�a���,��猀 ��]ák�?���5��o�Q�̪��H��s�����f��������N��@@�������L�G5�{��iB�JJ�j�މ�wP\��;4�������:N���3���pXM���4�R��~َ&���I���++{H,�I��d2��(8��g����݋��6����7&g��)�(�����d<��Yl��z�i��C����E��~��U�r2��Ki6[
�<�h�{n�g~��ӝ��{pr��Ua�����ޮ�I�����=T�3śr������pM=t��� �vV�8D���6��f��uS.7�u
y��d�n*���bj80�]�TڃK��9i�L&U�G{���� 㖳�����7����pݪ�~j&_�rx_�pB�ژ�-J�a��l[��=���&A�;�z(�\��&Ee�^��W��Zc6����]�vΊ��4�$��������K���}J����_�9f�f��>�h
��`�Ch����q�Pw2 9���� 	�׮g��Ih�G�J}���o��l̼�J.'�y!����0�rp���4�^�S�~zs�<���;�%n�k���OT<�aQFQ!����2?�<�Ѳ}�p{�үO!)��|�Z�`�z��NFy��Z�J�|��P�le(������l�ź�s�~�qJzvB�
,���:�]P̓��wܲ���
�o���N���V}�#��į��&,��?���cbA� ���W�͌����a0�).)��6޴k[5�m��|�gb^ �/��<sh�W�)��9~L�	�@(hD}<��5XNn}x�b�VxR�1i�8UOBbfM-j�nO��/>� ��Pc���GmJO��L�yϋ	���R�p��|T��\�2t�U^�-�@�R��.R �u�����!o���_�����9�=FUEb�ˁ6q�&:&���cM?Q%�j�3����l�&i��c�v���x�æ��dq:Οao`-�X%��yx�;(����yaoO<�3e�s�Ƿ�3�I���st�|G�� d %	d]�Ɇ�=:�Ut\�����V���^e�$;^�
`���Ƥ`�MY�!a�j���w�s窮	�|YBb�I'�3J��������J��ZҖ�|V��YcP��q=,�٫�Y��0޵,ܫ7Krr[r`c1�4���@Le`G䕠����t"���~��~\h��d p-�$�6ۑ��(����7~Hɡ��D��fO+����9w�⩔WOU�Q�#����q�"�=��M�$D4':�:(H��	b��Byf���*�䨽�vG�ąۛ�Ng	��fkx�=s������C��WG��jG���.��I�lhvZ)>)*bj��8[���G���AUv]L�Zre3A��8�/JlJ��$�.���͓і?��侀�Θ�`<��=/� �:��B�f+Z�[�D��°���X���a���~eu��I_�NE�Y�:1��n�q�$K�9aјW��썧w��K���6�{ѝ/��'<;F������8Q>��	�8��\��{��7��`���k�2S`4]���ܧ T$\:�!�4]Y�(��(Ľ'2�@h�-o�2�\�����_���*�����u\b�%�ka��o���8������Τ�D���K{��L9.��X���p1�^�g�g����SI!*��1��{v��)���x�L$���#�2e�!X���u>!��A��D#Y�A2��|�� ��isV<q�䀩^�� �"Ԃ���/�k'�g����\�inn��.

�^�R����TN���>s�9�m����v�@-����Te=����h�"��&y2�pj��4�%�{�}l�-Aꦓ�d&W�u���f��f�4�f({?���U�Xq(a�ӈ��J8�wJd�VMy���Y�a���X�����M!,�:�r%A�s���:�0HQg3�������w,,ZЪ����� 0`����Q�>��������L��Aa�b�B]f��b��)�f�Fy��t�t�����hUL�D(��X��t��B'��t��W��k�9��j_�^���C�̩۰��ݻ��}r�~0����Ĉ� ���Ƿ:Y�5a�w>�h�h���4$�p�I����Ύ���p��e�`���J/����f^���%�QS��z��f�������pT�����~�G�;���{����#xJ!mT,1�LF���J��F�%i@�|���-P��J�S�����;�0�VtP�����ۿ}A�6b�.�;ߴ����u�,B�/�F'l�e1p���S��F�t��N�Wc8k7��Z7c	�b����B��������
����F*@�2>#<��U�pB�KC-�:-5�IVӜ�H
}�Il �9��e��8��h�zL"l��ɍ/�Ǻ�i�30���9�m�㯈��3��S䨄��t���������Je��� tF����PZG�5��q��TUm@��r(}�*��G�ieꮀ���@��+%��̨6]��h�5
�;�Y�.Zz���2����p��;���_��Ԕ��є�K�ޅ��J�3vQq���TAtΙpR���b� �f�ƍ#�%��ڔ�!�,V���9�V�����T��$�U�6���ӷa/zrzH��!W�Av����8WUH6)-exUpt_��(��*C�4��|n�ض?�8�4x��O��Y�q��}=] �G�1Y�"���ڿ{k���Wen�<D!���Q���q"�Ӄ0��U�u�0��xN�7�a��mXA�F���I�ato�e|���;�gL�96Q xU�!֝�T���*�0�<�����	iS��n�ٛB��N���琩�YD�����m�UJ����l�Y��:�stzN0����|����%�W�I��<��t�OE��j�W4���	z]�l,���n�/X���b�c���,'��)�d�KT���^���f`f��J���D�VqQq��졀ć� p�W���s�� )s��O�1 ��5wRy��?�Z�o��`�T�r�+Wo��@?�^n\?�䍳oI�҃��p��7aX�x��������,��� �g�:����f{_��&u=�|���N<��?;\&����:��87�s�jW�����3/�&���[Ʊ�-���Gbkp��?\�,Lݥ(���<���rpm3��̕z����;��V_TF���dB���x��UI�8j+�v�Xp��!�D/t ��������CR�!��M��׳}%��K���\kiRH��y�î���O9����֏^��_~�5]]JH4��m��<5XcS�ě�P~GJƠ&��k�
�	�9�5���߹y����7�H8[��1��X7KS�c�'�c(��V<׀R\n��u>�fQ�R�m��yе��h�@�Kei��:��l,�hd��i�s{��d��!_�N�Z�W,��~���MC�Y9��\�Z�h���N�KQK�٪L���ZEY�ҍ����pq{ܤ\�<�62���=�l�ts�������!k��JȻX��ƊJ��oY�,�!�� �! ����	�G���� �L�o�Y����"��T��>"	�(G�e�!�m�}�M�q�
U"f:��*����"���Ue�
"��Z����u��1��VB�b������c���z���4;pwK�-5Ha
�%�m���.�)	tqRX����ݶW�PG`�_d>�BV�W�D��ѣ"�7�"T$!��	�Dӟ���*u?~��+��^�������Zk�}V?O��{P�ִ��AF��u'���\���6��}�o�� �U	jM�+}BW�=m*��^���w�CEo!!f�8
��t�UpU�f�+b�o�`$qv�/�@=O�h��p����7b�8Mv� o����� �<��T�iV�2������6&������J9���F?��-�F������6�=q�W	��7LE,㮯�C�7��̽�Ѷ�̠�3t�2��H����s��P*���e�4�T%/���hW��	��

��V�����F �/v��!�6Ԉ�
������Ez|��M2Ui1g���5�>9� �M"yw�I�F@�I@��2Y�$��&KER+D��v�����5���G�p�f�|�����e���A�am�Y3��0G7VYʌߋ�W)�ֆ�\�]i��)~ms��s��R�#��j�1��_>��c[h���+�h]��p�h�*��fOv��3��J�I@���K�CĈ)���&�:W�̂ǡ��ȷ��mpǉ[:h-���g��`]�<"���aن���x�6�M;���`i������R���1d��p���b��UT���+ug��	�J��)u���Zy���)b�7qRS�����BI|�/2
8u���O%�ې �k>5)��"I)bU�e3 ���m+,ᬺ����E�� �Y�+f���wY�I��S�ٜ}z�oz7���	�ϓ.��- ���BB �M�z���N�r6,��h���ZxO�*�u�,V�-�zs�$w�"��@'�1[(bp٠n��� �����k�~sd�=sUi�l��%~i0��%+;� B�
�X���Ov~1�HSmjl�R�6.fak-/3~��%�(�� �.H��}����	Og�_����<���!�ڱ����ZҢ��
LM@k}��\�~#��7���"�%�]��o��{x=��z�PhZBz�įwd���}�
8@�̓ӕ՛��F�s<{�L�o��� F?�� &����2EA�`�0�2��}���:{�n�Ͽ��	�ᓽȡfU�h&�T��S�K�YX���
��CC�W�s��_�0iĹ5d̤��¶�0M�y
�rj�s�����*�o.)����d����11F����GH��������:��9�95M@�WR���]��Э[%!8չ�z�|*}�62��LG�����䲳U����Tf�^"�9%d�I�YV�_|�������tq�Ѳo���������\�,s�5i�H��Z�� x-�{(rŌ���h�j�F�����I���	��E�"�x��_Hi�}ӄ���d��'}�!��
���!�ut��f��ҝ���.��N�߭:�+kZU]ӡ��7i����$���9nR_7v��������iqoF� ����՚"���30q�mwc��G�i�IҎ4�-���~���?�Oҫ�'�U��g�	D�;Vleڊ�*�ὐ����G׾�<pU����|w ��f¹������Z��n2~�>� ��~��%�U�\ci>���Sth���.fͅ�g�eoi��"���y'�����[�����71{���`/����?�
v͟�D��n
�ea�,,�wn���93
�54/��I����?��!������D���7?`�zN���zF�ī�{��=@3��+�Z��6S	�F��bCm�W=�:�m�}��S9���Ah�Ѹ Ǔ�1_�^����":GoQ�]W��������P�k?���?Y���Ƞ*� W^���-�x-�ֶ�yV�q_k`��J7� 6[S�b�WlBbd�$�j�d�{R�Q�1��Y��H
%��46�~i�hE��Z�*<\��I͈[Sq}���N��C���j.����:�xK5�7�;�˹��V���������t<�QA�]�R!@=]D��]fw�ځ-������`�r&Xԩ!����R��*��9n7���~,:���;�+�C~E�JٌԸ����J��jКMCF_�R��B�-���Si�os|)��`9�f�0SiF�mV(�����T��bNQ��"`��W���sAБ��;����JR��M��.<��-{�C���4�<��ؾ�0�Q0���n�;�i�OD@����U�L*��^ƍ�D�ΔF)U�������	���>�
���u����V��J���H�@#@	�i.0SF n͋q�-�H�sF���▘/_$"�9����nD~Q� �[��>�^V"gj(��E�rE��,��=����	Q�k�%ED�O]Q�p��zU*+*�(Qz���a���v�c�12��q��������G���m��z�h�]!��G�@*1$���d����8>'���	0H����7E���S�\�>65���r������jtHX������b.~�E��|(��V�G�w��� �pI�G@��/��k�äAz�.�D��/f���`Sif��y/�CIg����^�3� �py����7Q5u��ғ�K+ӣg/�R��t�	�d����q	�u�K�^J��,���e��o��ӑ+�R*L�����t{�XQDF�8Y%��?�/<f�Gx
�;�����bL0񉂘���rGe^�[6r�ݬ�y�6��2���vZ�g�E*>ѷ2"X_tqc�[�!��`F*��a*E�܆Rx���}����[�l���C2���Rf���@��\�b�~�+y��.��T_Y�j������{�PF,�e4!���!et���a�b������l���36V�M��ݘ8�����a'$��J;���0�����}�*���!����N�/tua|*5Ӌ�v��Q(�
�����݇��eO���1�|�_�|Ħ��o�E�a�����0�3�DI��F8n_�����8ח}|o��w�q��.������
j}�튋L� 8y��J���@Ӵ�T~@!7@{������=��hΧ����GwޢBn^��7t��2E�pi�UN��>�B^�E{Ƙff�,�:�;w`bt�o���FYy2�S��Ė��ڕ�Y�pZd�	-��Jbְc/i��׏�W������x�V������h��EceM��"�\4��i�OXʊ��MF��m1O��Q;��'�Wp����\:��Z���n�>+Y=r��^[�d��W7� � �vH�hit,�+�_
��	��D=o�S�)h�K����P��� N�I�O�$����[�&,՟N4���:��3�k���aD��iۑ��(���#m��wXt�
IHT澙������э��"c���g����:
��N�`�����Qd�QA=��������L�+������=~R�+�S�q.��R�W�ƛ����nG�Ǧ��=�WEB{d�K����a�)v�<O����L�
���Y���g)� ��/K�A3�*�����=r0����9�j;?vl߆H�Մ�2fwp ������I��'_
;�d�	t����w�����zMj�NE��W��$��&殡�84�
٦B5:�K�I��h��|���K��_��[Z�Z$�:��:f���5��o��p~��L�r�h��;̹=Q�4��~І�quB0�x'Zd4�E~a����;<��y���TH�*2�ݡ]n����A��c��('�]K�b.~��%��K���	{�z�HM�F�0Em��(1M��P�x"���g�v˔H������G_e]KHl�_5�JJ�E"'��q�|�1�;�nhSy9�5��Wi(�Pz.g�r��NC�R��B��1N~�B��[���ؚDw��K��B�oU��є�˥h��D����ƞ�>�4;���b����4K���W�YF��5[����$�{`pww'd���,�Cp���py�ۿf��ӫ�Ω���9MvL��:�T$��9�h��OH���\ۧk��U+z���2D}�����í��?�Kr�8w��V�T��t�@5o1IAt��s�!�%L\!0/fӵu%�����_��>N�s#��}�^gk�Z���~���g5���/ Zy4�RS��E��E����dY ��B�戦�/q)�Ҝ-~*�K��ڟ��ݪ�B�Ђ-aӉI���!5˜���Ǆ����e��K3���m9ױ#%�=�LC���Z��}��֯��M��L?� "�-�9�2U2�&;bo���Ӈ
S�>��=�`���uyFB� �x�<<��苩$[���?�>0�P�[����G�oy@�D�m�.�-87���}yD����ˡP���$.7�v:��,�	�v[{ؓ�7f�]<^ʍ��Sc����W��Y�b����t��5���##Iwm�ό��+9��&�;���͵x�&���0�F���@�=��==�hH|�Y~�֡b��榣),T&��H��� .� Ĵ�t6Nm�P��k����:M�R�i�k؁��kA7���{�y���@1�Qꩀ*,$I����}	:DZ�����Ӧ��4�@Ƶ �4
�h��'��ը��{�H{� f��Х��L�o]�b�&�$��|����C^�����o"���*gxt#
lg��/��cm��ڲ  ��( q���.��!r���嶭��(>�O�Cª�r��W�6��I�/[�!����T�~d:k��>�Q�eɣ�,���S1!�>�O=ξ��PC;ӧHT�t%	\�<���Yp�,������U���L���š|䪱�史_}1?����,bX�Vr�*��*م����m��PS;z����&�A]'���d�ssQ�EHy9�(q$1w�w��LY�H�`�x�<}9�H��B;/{.���o����iP�.�l����}�,���]fȾrH�ez�5��߹�W��-=�f6���},��SӢC�)=C��U�:���!��	p����~���I_��vFz��[���3hX�D�~O_E�K�$og�>�a�M؎��+�&�5����z��V\�����`��l/�7?�o��A�De��j:ѿ����{
@?�=}7���ǜ�!�_&Ԡ�ׇ$K`�[H��ap;C�(�n�f���(D�[3s�Mv�Z�1\Q���(�-G�����B �?�ے���K�9�a�������k�PhQ�Þ\c��
��fg\%�;�/z�*��W�|&B�}�1;$M5?g��UK� h9�ba�~A����C�o}r����a�*��>���zg��U���+�j;_�8<�t6�~�eӲ`��� ��,�L_�b9@L�䠘���C�A�U��~�����B��8���T�x����s@���_921Q!.a~SMa�x�dt�[�`���J^<%�S���&�īZ����,I�#����H��6�F��|༆o_�C"3e��ںIC:��D��\=s��	X������ȿ?{���N�6���ސ�O�8� +�~�D�`��ӄz6�Ai��2���i�v��P��5;m�U5KS�T�d��r�����9�L�ܻob��GELu[ω���5��D���p�z��� ��@0���x���D?n�m�s�~C�J���^;�hc�m�rɥ���ook�r$נ��5������.��{�In�:�JW}� ��R	��Х�3�%l_�b���B��ňt���ֹ�x�,[����.5��ى��d�Uu�lnN[o�vS0z>���_�j�f���"�L	��{���WX��8�B�Gɿ�'��EiN5��p������hkp+Q�B��	�7��N��!���W�{på���Ԙt�y��x��W�R�^=��K�i)�뉆�J���#�K��R|)�c��TT7<�s݉)�{]�wlڶ.)䒄�#� �1�Q�Z�c�@F�f�j ���.�=�tD�^T��yMMh�"�]ߞ���ƿz�5���3���hC-���vvJClL�U��H��l&Ɵ���An��ҳ��~)5�� �Hf)?���R�s��Rt8z�V�gee?���p�dJZu�CL-cM;�M�0Do�m���6B�_�i@���S���.b=�D�8|���F��{�W	��@��������6�?�=��\��5�
���WE�/���ڑ=�(1ȟ��~G�	<KQ_���/	�#�b���� g�^q<�L-�u�����'�|��
�+;bp�����jSqNw��IsO`�����II}	�����kU�cm(�&���3+�}�H���m����shP��[Ε1hA��8E!;�:@#ƕ3�J�p�5���N��AYd8��`\ZjMT>[� ���%Fko摆�(���h�ͳ��r�'��?m6���9X������<?����r���I�^��cI��sJ�q�~蹎�
Q���I��r���AF�Ex���}�_w�MN&�~��9R�3��ם��~���d��r��	�P�=���yLm.[�f6U��I��ޢfc�{���Z�pt5>&�j�}��/3���V:��hX1ۑ�4�-23�G��C�R���'d�У���H ���@�iEr���碖r����"Jt�Lh�i@0OW:hG��	�)n��-�$�thj���6m�iO_r��ܯ�O��ZecV�u���C��G��(C�|#N(�c�q0Q�m�GԄ����g�P8�'�m椷Q␽\��7���w �Nޭ��|S)Q�>�� ����6��J�g��@ 1���Ţ���X	py�[E�V��������C�h��]�W�]�e��p��sG� ����?�C
��9 ��:2�ڒ�.a����~qr(̃�!e�d4�����L���K��`uC\�35�ֺ���6�-���.���}|��� �Z�AK��ˋ��S����j�6���A`s���{�K�'��\+�ߧ'~�!x��/u�����U��a)7B�S�o:E��@�/r�w��QQ.�_p��Qt���Α��Ag�(�����(AH���vxl�:�geW�ԏ���z�P�m�A�|V�����`a�THK�Xb���ẓ�!�7N�}[�kQ��6�@���7����K��.���B�� w�Ӯ��������ǡ��1��jZ*qґ}�����=P͂!�J2�W�O��"����?{�$$�cIC-�9_aap�'}�0e��>��WZ@'i&�����Tyh�m��b�ejl���G���+�'b4����n~��7'y8nؔҺ���'�-ԣ�ˁ#���� ��+2�I{�?�E��fh���d�{>��#B8qI_j����г�.s8_��~{[T7'[pM�������r��.��a3�����O{n]�z�Rޯ�a���w8(DՐы�8�݈ؔj�cm�{P�x|}%J�_��S��cr�DX? ��\��j%�ʾ2i\���C5_D�\�Ԥ���6*N���hZ�P����J�p��B5?nb��-��,<��%��i��ݻ�g� ��(�Q�i���N���ƶ�}��w��8"XA�Տ��ܙ�0}��¨a���-��;4����E/��}p���\�/�i��B��&�Af���z6����s
�Rm��_7���5� /v�
<�z��sҪ��J�x��iW�ͣ�!���]峻{��I���s�-����#����ʠ��_b����8v��ѥ4T3��I��tF�ƶ���w8k�5�A� �u;w�E��>p�ު�Лr���� �N���z~`DlC7�:�������(?k�T����ߵk���H��\��<��]"�N��nL�X^9���l��ц\x���|t�Ht�7�ꪣ�c���o�7}��D��c�x	�rI<c7ui����`@�f`�4r��f~8TΌ!$ؐ����.��w(��/K�\�!PHQ�3����Z�=Ѫ`��7�
��p��^�QMcx�1C�&w|�'���"Yֆ|i�;�ہ��@��bY����J���-��%�A%^�/�d%��Z��%%b�'5Zn����P�Xx@��/U��Q���bc?�g�_�w��<�w>���$v\�&l�=HgR`:�>J�)�¨Nl�\�@}r���ܘY_w��Ý>�lW���9�ge��ֹ:kv����ýs+���u�4/"c���@p��'��j�5���i���YX������G�a���n�+�S����˹u�%�fy�"����7<jV���.�5+ s���OĎmv�!n�Nr���:���+��{i��R�K�>N���ٚ�xx@����v���x�!�K���t��E���c�	4Dv�\HfJ?�,�a�x �FC�5Y��s�%���\�0;��ιcD���K�r���w��B\�t���85�.������:�ܺg��3�'걖恉�jy�Uq,�Mk��R�iξ�j'�\�'�赼������T��c�{����"�L�5Nn�ԑ%Q�����2���}�6X��6F]�S����+e�`� ��I���B�t����a�BC�ONN����-߀�PIX�̓m
U�Oc��!D��oH�f���a��8ڸ���l���L:��r���u�{b]��l���]a�I�r����7S�vYXvM�9	�-mOk''��Eԧ���D�u�Xu݄�QӥDc3���T2���ׇ�t���f��6�OK~���(�txzl�*%��C�ͷUz�Φ�%C~;��Nq2훗J�ш�=	�D�ޔfӇ�NJ{�֓cj���C���0���	$~��J?�o�m��"!)�*l2��taR�`h<�RP����/�������}�[9�b�i���3΋91�Z�(����T�t�tO�j&H�?�
����:1������2��3�XYC֤GՕ�U+)�$��(�g��"�l�����vp��l�r �/*J�!��ŉ�2:O=�|c:A����u���� ����p��2[kJ���:w�����H��x��������dƟ���Ar��6|Yn��t%e��]ڜ��h��LI�+���ꀓ�s�Ժ:D<û���Τ��o��Wٕ=֬1��-(��/ȊB!R�K�l��=B�ٕ��-�������	���@��'6�$�$�8�~]���ydbg��o^�M��^c]�/:��>~����*l�d�,�&X�k3�ޕ�w^��|:8HX�H����f�Xl�D����T�5�z�p*���bA�y�5��1���o��B����3��=�E�ڛ�E3���$����xC�8m"�0�;�F�w�C,B�qBMO×������D�d�I�9Au���>=��rk8��ƿ�9���3��F����Iggo{��=+�M���>f�CS'm�{a8"�3ȸ�
Ht�3����}���	j�Se@�|��z����-�~�3��{R{ڮ��; �h9���+���_`8�Qe�7�/������k|K.�7r�j�!K��K�{����IJ3�����H�Fg�lA,Q_�Β�p��������&�n���}��9rLO�h�9�ܰ�Y���5\�|�	���m�m��/�-�d���ך�ڏ����d�
1
*���(�%ܕ9Z<a����-�A��'�������7ːh��VNԺ��?�rPy��4s��{K&|N�Y^?z���Ɵv��M�*S{�?X�R��[
3N�LO���o}���T�����c�f�_��B�ˏp۽&��P43�y���*�X�^�;P�]I��! cT1A*ي
���?�rL��?��1�:1��e
s��p����@8�	���;P_�V�������Mw�z���һ|;�']�	=.&�=�䐐�CC������f�G��D��t��$y�0�7tС���^��nu�OZU�ԚO����:ynܜ�5��˻�����OD��l%��Q��qR�F��;7�CA,��W-E�3�,�O-&8a!󘰵�j�Ϋ�>q(��J�τ��S>-X���u9�-6�	�j�kM�2�ߵ�D#����Ǳ���Q�\!���y��m�e6J�%�w�����Mj�<�O�;}\5�+���@�$HZ�-�I������N�9��m��&�	16N�P}���yN���-�-�ؿ RJ H���,y��ڢ��[�X������������ऺ��AM���f��^T19����4l)GP!	�M�<%�褑r���?��)^�S�Ra}�W�zV���qeӠi.�~#{Oׂ�KF�b;7�㦦�+P��B�V�I����X�YqNy����dK	�(u�U���Z�F�Ί)��ͱb�+0VZ��Hm
�<�+�G��B�E�|ĥ��%��RH�2Ubf-��^�A����d2�7b������(���u�^\B6=�"9n\~��L�y��=�[
���ο�K��՚g�hm��cC�Љ }D¯��fO'ȧu
�C}`'�<�̫H�"I����s�T,܊\��������Gh��Ώ���>�G
�S�!�)�����b#�B�����Ʀ��֎��
̾O�!��:��	��w��w���3�{���#)m`��Nۯ�'>��z;������{�-���u��K�B0������QM/�oRaᾸ��a�K�%@W1�?�Z:{�8����62�v5��N�u箥����4�����o�98�̓o7D�W���LU��jqh��eQaAAA�2^�^�T���S]�ڛY���"Q���a��4o����du�����x��p?(M�Y��Ma2#Z��'ؼ�pz���x�����O��A6W�����_�ƀ�#S�Yl�d�}��=E��&+�
����iPP�

��=�EMs��T���ΔV%�xՕ����j#&��]����τ�I����["�::�!Z�����z�笺i�iA�)����Eܰ�������W��/�!�.�@5���p��ے!��aQ����S'R���}��g���	ı/a]p����spT�gP���k~��p�n?FC==�p߁�� ���<��G�#��!~r�z�6�ɰ��Y��[�Dk��W�*�	u1S#c��R MiVL2�qM��K45���.p�R,_5X�.B�l/��+��u�7�������4������y��H�K�?鏒��{&@G?������� M�G-�ՙ��v��I��L��d>f(��7�;��F%���49ib^
���H��
;��6�Dy�IKoY�
�W�S�����o�?`I�]�9�abL:ݷ&0�y��Fd6\%�G�Z�'��ST�cc��z����C4wINo�/��-����a���M5/����!,���+�vg �"A�)���ho�W����"G��y�L���.�� [>�]$���\�7�3���{Ζ��
"b;D]�-s �-��ǧgg���f*�@�T��7�,Ļ=��b�֠X���;|;�u���I:U���EFFCC�5�z�e���^�c��)L9�ێ���T���Er�&��k1%K�<o̒32�1D������X-r��Q�<V#�m1��9�F����Ȏp�I��f`�D��o���;e7����(�7r/ҵ�
�B(\�{C6��Nt3� Zk�V� ݷ|<���vGe�i1��ʊ �(�����A��`a�����y�������e�a��� �G?�� �����cb��W����"�ڏ�{9��R�Y��<����~n�_3\��o�8Ȧ����*9��7cVD���_ӳyߐ eU�:��|��s���N�&��c���;���it�ɤ!A<��`�#hHXq�t�%�M\�c��nlNiq�kOXۨ����4P���b�a4"�ĂF �B]_�R��]��w��lmAmFtq!:r;X��{3��J�J�}�e<�%(mY�٢��[
�H�3��u7�I�t�/��&=�h�MK���y�L8��fֹ���t��XvɗO��H/����ԉ%���]^t��*�T�K��Y3�>�Rۃ�h5�m�r�o�Mfbk�2@��#	
� ��Ń�N䬼�J�J�� ��bi�A���۝~��T� 7�`rÏ�����uC,5����s,�$vQ"Q.*���0�6j�����`���h���1��U1mm����յ�
}c�%��j�F����NR��QF�������������3����MH^\��DB�a~X�좥o�1tDWt��E>`j���$>#�Nz��d��X(8e2���� ��Љ�N�� ͜�/*�}߻JhBFQN��)Tg���*nn� ��QG�J:i�o��.Ԟ��#b�+#���E�~� y,����}ZӺB�x���2`���%���u2�D��hկi"����n-«�ċ�PB%�,�o��30�	L��:U�� [���쮊������y�oa�Z�n��R������˴�ς��D���$Ʃ7@���אZl�j(����]ʐ� 4��ؙ��!k��|��|W:�q%')/�}Э�� �]M�F��~Ik��9@��	�	�!q�y�:���f='��t����<�m������2E75� d7!q[��ţ*��t��C���1��d����i�|��W)��n|���TDT)u㲼�!.0��:�"+�N��Ih���m5�� �66~H�O?���,'���B�߉+U�T�Y#^z�������kl*_o5BD���7��@r�P	�ش�w
�,��Pk����Uw������,�۰���/iJ݂�X���i�4*n������R��ށ��>�����b��VV������S%�o��+��X��BA���?�۸Z�Xbc֘�엹 �-�i@�Q*#�Y:%�	��&��%��gw�~�q�����8�@�v����x<�$Lt���Y��.��T[d�Ul�ƽ��ƹ#}r�o���坄g��V��r0WU��/�W���6�vM(Z�(�X��)�K|�If�r����U��H��K��������Mwk�f������q��1�R�c]�+w�|�X2��z�q�p��0���P��ӂ�Ղ����z��� ����+ZI1x�KL3�>mH�搒��3w�[k���y����ck������x�UgW��p<y�� 7]>��A~0�U)�b1L%���2V��B�E�asʶs@���J7�3Ͱ/�;���i�������D��R%�>%^`	T�X�F1�+��bx#�����������Xhrd_F�;)��vy�L�k)y�SJ�V�U��曢���fۚ�Km����{��D�$��.t!�WtT�� K/�$Uh0^#)=4[ޜ�0���c���{F�A��C� p���s�Ys�4TrC��
���ii3r�]6a>iG&a�JE����#�D��m�l�����H�t�@x��~�����B���xm��%�ur�Ǧ��ðh��~�\H��e�V�N+Ք�0^y�����ORƫ}�LC-���2X������jx>�x�w�wX�ywj�Υ+"����Aq�҅)*��ۥD�+Jt�a<yA�)~�++����싟��r�_1����3����u���`Q�C�6����Yn��|$3�N�P�p�P�45$\};L�ZSW/
����
����݆�3C���f�IH9�e��)���Ń�����E�kՍ�����tr/1j� k�-Qd�����"Jr��6��+Vm���A���̭aL>���Hù��6= eN�t���5-�\�z8��OI�kO܍A];wv\�S�m�L��DX�r��5���Іͷԁ��!�;N�م��y��D��Yĭ����S���]�|�d�p Je<�nζ1�q&������O`���N��'���������U�Ů���O��GCU+�p���i��{�Ҥ8�.C}�7wXGn�w�)�'x�$'o��u��l��WP'�#?b�e���W��'�E�B��2f�J����=KI��zlu��	kM����r8�	�i�Ց�v��ʻj���)=�Ƕ�5t*������c���(��w!T�
~��{��c� c��j�&:�?�B������9oh��/Zu�����F��w�� Z�`$�/:nDl�P�|�e�r�a�ۊ�=�+��L �hͦ�	[ѐހ��N��95
,����F�nn�s�n�.�]���z�؍8�;i+꽈6���]t��|�^�0B�r��w���b�����⭪iD����I��ܧ.@�oӰ���m'�:����,�
�:p�a���K�ؾHI�K\�8��iNd�J��67�m`t����Lp�a6?��Ż@[��\�.�Fc�&lY���S�LbU������~D������_iW���r^\˾�02R��\@�#ɭaʏ*��%��6���~.@��G]3<��ҷ��Bbr���)u����w�Ӭh�JZ)U}��	k ;&����"��h��G����:Lt'iA_���E�CK�@u2�C�Ƅ�k������i˰Q�^�� �"JT�]�q���ô���#���7V�@���}��e�a��`��4��:�ts[��e����6�|����Uæ܍Y�����=z"���.Yg1�jb������IbQ����`Ǵ�Ֆ�pNik�����2|D!bb�x4V�P�ssm�V.Q���7;���\�ؒ��e;pB%�
���Y�i��񛏝n7>Y�:��5f�CAh�:��.о:b�AfJ�������|�bi����V���x%s�[8*O4P� n�/v8�I��|�ŴI�'���W�/���	��f�����vg�K=�/���-cn�@�j�_A�<ۓ�/r�x)��� JF,��x�r����;Cv��J������n&�;W`̇;��&�q��~RŠ%���<N4�/�=�����B�z��Ñ6�Q}��*w����9
�>*6�󵠟?�b�׮����bJnHQ
�G�.×/+�3X���q��d8�k����z���G�ť��ڄ��
b�Q1�������y{� .�D�<����Ϟ( ���G6+ƿko�Ӫ&!'��E�gfԖ�xq���p�ۅԌ�~Vd�g��ot�o�.�����N|wձ���a�l�\\0#�_?ؔ!�?r{!�yUl�F!m�;!sYp �Oxa��m�2�Cz�<�ͳ���0b�O����'��4d-�^���_KKk��WȎ��!l�.f���!��$�A+�Ō�������ĔR�e�pX��xK�ϊ�"�ς����x1?2r�=��9�gq��/���������dJ�l���;�v��@$�"F��=������y ��x�E�b�J$���1[���7�E۷+�x�h��X��D�"m���B\?s������8�G�S�m|ϫ����V$f9��L,LdTy��ܽ{	b=͎Ј�(H��.bt|���5�h.�2?U����Yb�9p1@��mJ��S7#������|Q'6�� ��agz��!k�^QmXsU!L�N@O���{������5�~�8
E:��W�J�y!�6B�/F� ޕ���R
ݒ��!����+/��)`���u��guJ>6ȯ��6h���OEq`�v$��Q-�T����mn;�gS��r_����ѱ�(:�_��Ĥ�i�cO\�s8J�o�?���Nu��r��R��E��:9V�;����p}\�V��ǜ��M�*5���C�p�*�%H��_�֥�U%5�1=�೗62"�TyӘ��;s �"�����3�Ln�h�}�k��'����[ �����n��?n:����д����ҽdkү-��@J�x3�Н��r��d=�ͺw�r�6��]���'��T�yh��tک�}�d���b�Tj�VȤ[@N%� �-�o'���ӗ�¦b��M�n6Y�=)w-H���;���"��1�����w>�p�X��˙��"o5��m� rї��~i%+�j�&��/��瞗GX_R;�pgZ+������l�k�JA<�Fxؿ����6���AѪ�|�H SP3�
.���j����*o:]�L����&
�:S�~���X%USz�y*GTW��`�z���O��w���i-��Ao����:\�ZN���e�j�&(���ܸ�?͌,��&��M��˯C������!,���T����C�Y��	�Tr������tR�����o7XVQ^L�-���l^J������2Jaa境wI�~co:�)���Q�`�IE��d��è��a�&�i��H��K�OS�XG:�w��O��=�mN1��p��;�ٹ[�/$O�)$$"LW����d��>a>�n�S�e�K�@�ݛ� v����f��ׄJ�����l?R�
���\�%#�#��]�r�j�D���|�T�x.RF����WJ��S��_�l������h]��S�t�sy9-6㝫q�.���`�_Hz�c~^�Y >ҿU��d¶�r%�r�| [���o��,7���+d��o��89�;|6���ă�Dd%J1ު��n��[�]���𖢢���-���ٳb�a�K�?��Wa&�B�;��'7�6��������U?:�j��mRr��:D�-Y�P��j�X��AD9�;x�rԘ��ˎ���Aa6+O��:|D�d#��1�8�dC03֦�E�\��m�Г&����F(>������Z^0ꩆ�c��G3�Sd�|Md�.��}���?�����p��gUM�Ŵ	�	��̆�?�ԟ;�v�V�r��WV��˨Y�q�N˩����4,#s|�!��H�E"b/)�m���ѱ�����aXAhk��i��'n�F����"9��2'���(I}	��L�Ec���<C�ӥ��߿b&Ήg���;����B�5?#�7��Ʀ�֐�����ڜ���~��s�FE\ʜ䰕�3g�ؔ��1��N�q�?~~�#��-�{�� ���}XR��4,L_�**�hq�F��{����8G���-	œ*�1{��C�!�0/�i)S��;�*@�K�{-sDH�D�xTEI��A�4���F��C��� <����b	c'=�5���t�n~���p�t��'�V�F�!a,� ��hs�R+"���������K��r�����L��I����8q�x
^�p��$g7��b�t�:g�e���-9��E�%�S�-='�x���E2�#�W	�9<b�ZJB��)	��R�R������1�&��c�Ԥ�PW�-� ��li��d��f9�<k�QY��xl-Z���Í�vҸ��X��5MB���3� �ǴY3�=\n)�/�y�-�~l�1A<W�N���3:�vmK��|OM�4Rb�
F3�z���7�j��G��pfdQ�e3��-��-	q�
7N%:�� ��^yvC�$�̩�b�P�-�0��P���{NP�q�.Qz�3�^{Y�O[)b���)t��J���0�vV�0}P�ǝ�M�_ ��st�~5q���ڠs��b�|�;|j����~�K��F���'~�lO�� *����]R`���|�"�1H��rIA�v�-@"6��SRQ���E(��g)��	o��屢�aj�mbj���L��V��SF�<`��(:�(�A�98���D������b��Ɋ��'��T�Mo��(�[O[�TxW&FF	)�4�*��?�7I^>?{�{6����I��>TQ�X=BW�N�
"2p\�+��y5x�ظN�	h�滷�����G��e��+�'��#;��Q�b�ݎ��=���B�/��L��҃��r��͔s��[�ڬ4��a����:+���G�����nǑ�x	�`�l������:	���?�<0���ÓB�L'>�%#}l��.��n�Dr"Y	�[D"�u������v=*F��M��xqS��f?S5h$8�f��m�n��2	3&Mw��9C�N���Q�J�?����W� >��g��]V��L%i��RX�7TŇǰf��F��~�G��5x�-�%���Q��Ȗ�Ȳp"1Y`EbK��Q3a�8^^�.��_nv�;-_?<��Й����p�$��'0�a�	ވ���Y�P��x���P�ʏs��d��V* 3�Ig~�H�P 6;�S���V���� �M�q�n�m�����)NT|KTP��zrpOYŨ���p���^��e'�h��R��r��gﺧ������\cx����c9-̩,95N�v��֦�J�_����K�)���`�_�%���Ǒ8��a�ESߊ���.{_�����L����LT輹���0g��4G	�h�*𛗣}��R�u��f.tFJm�o$��B�;�5꿜\`'%��kk]ё����Y�#X�_��U~_l㙰�~����{j���0�pZ둹}���JĦ&�3~�%��vc����D���W(�����}�{�*�-������F��<i���fT��S�����'ǈn廆�v�gd�<EQG�)%d���Ƭ%ט0�U��������W��b":U�V����]�}
2�B�� 3w7
�F��j���S�ӏT	�z�ʡh?l��[�S�g�3ѧ�^�E��!^�����^���/���p�����S4�����]L0��Sy�[ʔU_,/P�S���*dy��]��h��c预�c2P��Q�#�&��_3�h�� <@^Hҗ��w�B�Y�	���o���#E�ӷ��0��!'�,Y-n�PK   I�XT;��'  58     jsons/user_defined.json�Z�n����F�%A�����4�x`�c��I�Zm½hz��c��s�Z��&�v�2|���Ūs�V�e��|���ǛUZ�S.�)�'�i�*s�AZ0�e��գ����|��絛U�����at�\(׋�s|#�uz�X~�7ƿ ����r2.#��Tp�
G�H�x���eC��lU���]-�i�~{;(6َ���z�Iw#<I��,�����6��2���I���D
c�g��NJ�O.��*����2,��/e/2�6`")!+�$:�$���ܾ4s�ҫ~���)�9�5��>�ݫr�r���_����\]M����gu,f�>�ۭ�ŧ�.��R\\��f^���o�����e��q����2�s9�^ԅ��Lt��
�\����_���)~z��EZ�ʹ����I�V� ���n�j���_/��sqͿO�W�+��\\���2��>�1*��M�@)g��$�H�9��'�J!x�c:4�$f,c$��DZ���.E�$ jlび�^V0�lӖ�M�0'A8�=�d��8��)Ɍ�6nT*=��V+���ơ�������t�x����e�y���\W$cD������A'�����i�i��&ЃjO$E�xj�9Z�`��Ӣ�1�,G�8:C3:`�t�Q�Ȟ�4���T����M�B(N�DQX�ts���l ���e���������������D{|�
/��YO���Vx�����'�$߲E?b��>�h�֑�fA��,��5�I�C��j���&-4�E_b#�F��SV����EN\J�B��Py�H��8Pel���P�#�Өm(ʆk�Q�w$j�FI�'o�bp]��޴��dG���	���ǽrb�+��^0K��jޢU"`1�	hzI�h���9r�:���H@HP.Kʽ��˸ �+Mt�����a=	�If�,X�dzA��эY
��g��b�j3F̈́k��N��&�ُ�?^�؎�f��N�AAd��k�=IvLP�i�%����b���;E�_w᫞�]��t=l]U��2�z8>����ѫ���vX�Ì���u���b�v�.M�]�ݎ�%h�W��Kͬ/>����l���v������A�����_`�Q���l�3�uH�.g3Xh'�ݡ����p���x]�f��;z}���O��_����w�]���m����v�����y�NX�%��	�Q;ay��{'1G��]��g�'�h7ҥ��|�����գ+�����MGoV��N�������%YPO$s���F[�O:7W�	�v�-V��@V<�(#A�������{ƫHXX�8���b �e�ʦ'W7]��BFh��E�+`�D�����>��x�c�����n�so�Ͻ���kg�������,��UO��џ0.4�v�b�  �P!��1��DCnka�CzY�����@�NP�X��F4�c�:��S"UF���$�*1`�~O��	J�p�.q���	��V�}x�i�
�))o7r���l��x@��
���9nlo'p-='NX[할�I �f�9t=��yܷ�܅I���o�J6�|���ɷL����5�Y��[��j��&b����4զ�����z9�+'䣛n�_�����/~�5.6�E´F��(�r�7|Ww}�]���f;�[6T�}c�n|w�v~��T������ӛ9��n��O�yZ^�j�������Dl_��7Ә�|x�\l���0����۫�75��Fȝ�b��ٮ��n���ʋ����#��>bg ǋͲD��:}��彝l�ud���m�o�;����j��ݍ������v1]��=�m����+���7�Nq'��s��Vܡ�6�)$Awo1�*�+n� ���X�Y*��|CB6������Qܵ�A\S���M������=(�ĚpU�2�å�|=(I�>����%C���r�/F��>A��1>St��E�0���*+@�,sR��mz�|/��"�uF%�W!V�A�䥧���ʸ�!	�n����:��kI�j���6&0�`��R	C\�C�怙�V����L��2N*cS�!�,5��@پ��!C��pw�.�����&q8��C��7������;�B7����)�î7����vy�����T��Wy���ʏ���^�~^��4���Va8rޓl$#��L\��ͭʞeo������a�2�1
&���z���+�X
�<?T��D�V��V��4T)�T�1!��O?V&0-h9z����p�@׏5x��`z"ma@�=�ʆ�<�{�n�]tu����Xh�?6�"����3K7_���z�R2K1�l	u*b�RhQ��(�Yu&�
�"�n Eq�q"���S$:�)�H�6�����j�䐁E�sU!�e�j�f���)���6	�Z��B�.&B\h��oų!0���f�;���O �I��I��Ǥ���6A�`�}$�=�s�7S��o��L�"�JTC����5q�`-���^��%�j�����AVG���7(��i�?�mA�{�u0��}5�]�i� UXʵ����@m�:�Dp��X.'�e���X���2��;�s �J`n���6�O�ކ���ث�7����p�k�`F.N�{�m/ߖ��`sn�eT�����z�L������`�� �};��Uq��e�.>ᠻ�i�O܋HP�S�1�qa�Q�)iB�Q0��j�@��s;�|@@G����XϮ��28� YȘ��t�{�1�g�t�8g}���<��W���B<��$8L�&�Dɡ[�dH��o+x�|�d���s�U�؞%����(��ܔ���y�T���KL�_�PK
   I�X\.ŋ  H&                  cirkitFile.jsonPK
   l�X,qJ؏� �� /             �  images/278ed6c5-ad12-4b42-b098-da68003ec988.pngPK
   F�X����7  �  /             � images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK
   '��X�l=�o  �o  /               images/2c21fad4-931a-4469-89eb-1a483abbb87a.pngPK
   F�X�0��^  �  /             %� images/3cc6de24-d07c-4ad6-96a2-959384ef4fe5.pngPK
   ��X�}�R��  ��  /             У images/3fe24426-b06c-40dd-b590-a579c31a1c4f.pngPK
   Ŧ�X���j_  `_  /             �) images/43e0edf9-5f24-49a3-b78d-83485af402b6.pngPK
   ���X��Y9-  �-  /             v� images/4fde46ef-4620-45fe-a6b4-d27a85e18129.pngPK
   F�X����+  J  /             �� images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ���X�j*�o5  �5  /             t� images/5ca6391a-909f-49c6-8bb0-8f0a302a1c0d.pngPK
   ��X7_DW�  |�  /             0� images/649de870-1a94-4537-ac6f-7e62814b65a9.pngPK
   Ŧ�X��~��K  yK  /             �� images/7ac84256-6e9c-40ba-9a9b-c812e48c1c94.pngPK
   %�X5�3$ �$ /             �, images/8251b1b7-c97c-4929-9682-a545aa133660.pngPK
   l�X��� � /             
Q	 images/8d01a3b7-0772-4c1d-bfe7-c89158596f47.pngPK
   ��Xq�q�  i�  /             7� images/963eb574-430e-4d09-a29d-074ae2ef552b.pngPK
   F�X�&�}[  y`  /             �~ images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK
   ﴣXSW'� �� /             �� images/aa6b1763-b16b-40d4-b079-865cc7d3b61a.pngPK
   ���X�V�4sE  iE  /             t images/b14b5b74-4377-48a9-90a5-00abeaecdcc5.pngPK
   ĺ�Xm.���  ?�  /             Ϲ images/b2b92e47-5c05-492f-ba01-c47f59068786.pngPK
   ĺ�Xq#Q��  Ț  /             s images/bb187b5d-1fc4-4a4e-a882-8dc83b4f659e.pngPK
   F�X�x�</�  �G /              images/d8843636-1db9-4a03-89e7-cf770aced3d6.pngPK
   ﴣX��\�  � /             �� images/d9fdc4f3-0336-4129-9adf-d1b56d6d3ad1.pngPK
   F�X~��a� ٮ /             � images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   F�X'�Y��  �  /             �b images/df4f81ad-bfea-4377-beb9-28b9cf54631d.pngPK
   '��X��*�  �  /             �f images/e8e17911-f8b6-4995-a3a7-245093d5e388.pngPK
   F�X
� E  8b  /             *� images/f891a845-194d-4c25-9fb6-ae7593a7f9e4.pngPK
   ���Xg�	�;  �;  /             �0  images/fb3f2d9c-813f-448c-93d4-6d887e4d49e7.pngPK
   %�X��%� V� /             �l  images/ff68aa71-01a6-4ae8-900b-bc3222580826.pngPK
   ��X�>�~�< �= /             !$ images/ff8e3ab1-c379-43fa-8f3b-dd687c341a4e.pngPK
   I�XT;��'  58               [S% jsons/user_defined.jsonPK      �
  �^%   